`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
74e74PpIO4gZbJBUimaB9+5QVZup7cbIpznjtjsi8ezAXo9puBW/gafhvAPQ5pXQ
2dGD6L2jK4Psi/kmLhkV8bMykUGP+Yk0JILtEzFlfTUiES2G3IOHo/qWAclTwbZ6
OjwqUHX3Iy7w3rC5wldY03dX4ZHkTe+8aEQ3lHjXDf4zmI/SRnnYvbMURJUL/Ahh
UeluemYUkXjekoWusWju4OFTDc024xW+wZ/ItHcIiYx2NA55Lna2Eu46HITf7RcA
+uZ9Z0XtsOYaQwrAKn5bUCSLcuk61+bpOnSTaXVmAKb6dJvTMaEsNm4H1X0TtOOm
qODHxIGSC+3dkgPgYz3H9Hq8y563sVUMOg8LgRt6kckCyrKe5GR/xh1a2XrY75gl
KW2XttjBw/zQAiXvP2xyEJKps5Hz1710CbIcBWdt5rqkAJl02/mdbvk5p+lA9JC/
8GPncOBchUQY1tIFW4U/rmUMLdQkgY5fMtpm5PThBKX2rlHuXhXreHt3884AWcBs
CpYLPLmbpuuP07jKtx4kfOPgOHRrD/131A1HDGzoTNekx6Ysu+Kqg1o6y/wJTM3x
S+nYi8lwtM+iUA+YnVrWEP4cOws+qwGVKEhxMl97ce9p0lDPdVpXxjEZqOo0K90n
2ok/OxFivx+g68tQuTeYRGM+JjxGk9FXfUxBSOqUAWD2i4IUJ9IdbKpOJ72EVH1p
mJDIcz7DzMEJD2pH+T1Wr2MMHu0i+lGfAKMd6CCGwHgWbYETlDe6PqDGdsS5tFgD
Qn8u5WhWGvYfDHrtYQ1Li+zlGz6lEoUzYD4sxppMbVeWF3IGZ0dfwgY0HOGpdtTk
8uuRqtzQC08aAh7B9XXDWD9f1pFHIWUAC2QP79hzqAhs4lzmsYPcVjU+IKjU5dFs
yl8xZ4acu7hTGwdRktEHmTPVVC2DVwI6PTRQ6pzJT4cprBf+WkMVfKbmynzMjP8p
KWhi19SK0u1hwfY9A2OmLHDw7CADiqlZIWdUbpwakGmRlfdhLXlDNDJdW6vRV5w+
wO5sTdqkXjE4VuH1hZb3m0joao1MYNmkmd4TNGbIGT+vW1zqHR9RCGQoV6Fa5JF5
hf8ws5PeU0NlCXZEOQGZ3TdX4RH42NdE0nAW68KxSsHuDrMG9a5FvVUaoE604Pee
9o2wODyPvoC1fAc/xmiSfc94d+A0H8qlu2ybmhu3l4YfpQRF0mO0tiMz6bfsySIe
W6ToOABaS5qgdKeudZbC+aI5WeiEhxarQUquKBPwJqWDbCSVVHEkIZ1c0xbeahNt
20RzTAXhHZS+j/Tt2RO7EfZrvXCM7RzaFYADjlSWX3MDC28jzmSHeZHcORXDAA+h
akQI1RqRaI9mF37azzpALQUoE3Tn/hRIbGYk9JCO4oZkuKQVyhm67UR/T33i+qBJ
OOhbhWxmVD2bGO1o6hMVGg/0ZCEojITGXDendcWaAKUakI1b76H4xeFGiKT7AI63
dKErHCQ6eDXCcGnGPvNQhEI3uwgfZjMeJh8jqUgodxM8YVghLaEQ0HkVKTOrOq5s
ezpB8BAbry2HS4TxVxnVvQnV7t+1yG/K8n0HokJyalnvos+RXfgmyljAVB2xgJHF
dj7JEk3A3BXpzIht0AHqaowlAY/hsRIfyRnry+geGR29I3mJ4OuAlPcniYLJEKwk
uH4feEl7D3Is1ekfgL4Z5pCG2Qg/jRrBBTVDiZGy4yHlohSgM+nMNKtMauFfout5
6kCNTh5Tmdt9uVBp04RUCuBaCFgCvbaU6VK9YKWIXDGCrCgwF7sLI1aQcDmDMyYB
92CP9QvCrbBYh/Ky17YetKNxFJjH1xIPn99EfX622Z4luj+a0GLFZW92oMMpo0Cy
f4nrer3GPDGyhmCe719kCP4cE/LXsqG11T2QxRtYptZLk3X3B+Dj3HYXcb84r+8I
URXIQQiLnjPFCA7AlHXhoGJ8lSIILVUUdAEelnKjHXe0+ZDY+oIxt6ngDuisGPQD
JiYWkGm5GaCGK2+tjApSmYVauyv8mAXY5eg3pmfv2/j2fS0Ub8iIUOwSXeJ6fCdH
SUIFzFpfoVny+DWIO+oV4zNv+OVBvaPevORxnkDyrVP/aeCZdbt2zaf3uJE6kSty
azAtv0QiiPHc9vBJWQH/Ryw1ljYoHtD2TaE7pTguCjN3tJ8x25I28lpyJUgntOAb
2OAPMJMF6MR7TYP0RnjmUoqm71pTCdyMFoF0XveKxJGMva9WaXs9iVRMAI7OEGP3
Dprm2j15exuQyDpepmzzMezOn5Lm8w1eESzlB4fwa9Vp3vDJDbMfcGV63kADGoj1
g0AhVqk0ID95IjqwMeZGCQPrB0AQ2JLflw9dHc7k2/Gzgn0whI5fFQT5RWvwiOmc
26ifXfxK/THRiU3zJzlLOi4qnQg164Ben69cS3zi3hPUJzx7OLh3HuRkZ/6olfho
MH7IuXSWoWmDe21QL0ErRAC1d0zQAk5XXzchRQkB78jD0ypoWPmYF+r00ISQ53//
3obSJzG+ktTGAiWZNcgaJ0o0QiQ0YKK6Xg3W0zOLfBwBVnjWx12F/vftO8UbzzWa
2pzi8tNq3hjo58ZpRI7r4JP8Cs9YaSp0vvL+wTO7PeQKgeShvFyUPFjH77lu/D/H
M41l8wDibfKXRIdWgxdC4pj78oaIp1zWjDzgRQQXohV3Lx8Ef7OHfF37176gDzgT
BsAOZ5SPKb2GA9VCdPRXP8flp1QLrnLy5LHoU+FwDZD/U+6Bx8QeQacR/yvQVKDq
fgGdETXYAO9QRKcfFd8/E5uHXEbpGG+CLkQjYMznGUUDWeEMzXpHiNdlwqwmMQ2U
0rKBe+fOFLbgn5td3ut1KquaN3qSyEuhdIwcnykoY13BFUolyQTQLVFMswk0c23a
z7P9H37ZYmGTOUbMXfvaRuzlCvV2JvqMLSg87Ymuom78OSkUjOFlMI669BAmsHMz
/uHpR2TH9H7vrkQAOSW1Rs2i2umoUVYoms1HvbZRwLN/r8ETXrUaR8d8nlhtJvrr
pGuUFYJ4kJvfyael2sEaDMataPjUmy5yle3LwOn8B40IoJ/9lA7o0zNVktQdPeF2
sEV/4wd2ehJOzX7Xo7TPM7yxMUiw7VOHCloyjwOn36tTJLviztui1pE1/gXWl13X
A/QZQEzlEsu0i4k2JQYfkIpb68+Ni2bDRDn5FXZHabhDUEWOVPZxmdSIdiIarNIs
VmAQgPi3uNyRRZjiz9lj7O27EA+FxyJE9I/y6QFEmSn6wWzqGm59nIq2hpcS9RTX
hTw1wcaQW4TFyZSC5R0xZScfBH2bpKPYzDTn1QKFv2sJ4WJRblbqLXTQBQ60rLQE
Yi9igU/5w3atzavcdNKwFvTV1TuLsqF16QkFsADmhwuCC8EEjDE/hkGLUu9WHjn7
RSDyEUlCSSTRJPpa0HMMV/PRRghgcnRfHLzVCCcoAhRXNZRPkozwz0qYuEceEpQG
E1C1TYG4N+jL98JHT+S/S49+sgAKzPzb7p69eO82/QXkHVgmatDSdVJnw6w6iCQy
8q6wOyZlEjsMCZtSskZkY1iovhzwjqPacO7jfoUVqy2VGcfZmbeic1xr0K7R7vCC
S/Uv9R/eVQFVCSK1yezG48wGoo5ra+5R12I5DVRVb1hHoxXHrXv+fw7dY9XGiNM4
W6W2W+yUwdO70ZLy+0STIWdg5aXAor3Bs6xDmggblVPBHL/iBdenyNAQxCQSUli2
X9pGIq/nSWSPVfqhPrdHJeokfS/vY3855Ard9cilPMjTZji2CY1di+od+kZkXL7K
LIQKY8yCWg0aI+2r+NN03eZQzHIKFfPCcFF9Tpu2EA9KSCHiWkQ4pE8MWOKQZMV6
Utv2JpvqOkZP3OL6qeXMRj7w2Jkh7+VKaPiw1WMVfWa1FkfWr50px4TJlDeCjGYJ
/EbX2FTaoaie8KhJUwaXr0sC5Oj9cDiJ/xuWoQxVEFbAd/M7QbJfvWL2URNKsTHQ
4zp28dJFyN4IRiSMCktm/RZc+zjkTLkjwjsLh4zbU0jqzBD/c8Jw2WLOVbT1d+MG
2HOoHjyhPGabgaHJGQ0bvSF2W1oKlP4twvC0QrHYfAiGOgaJ2I76LkcTkOVGsVDD
gW4AoHaUs1niFuQ3pGLqxZ1S2BTB/yggSKcOsqHx3GuTEIaNygBWtz9M32MEG18q
TS+4zTfjSaiUUQXwLGSK6bTxCSMB5dMTBnZ9FR9P5tT/Am2EvUN3F/FDQjZpnpg1
geuZMCpUEWrMtW2DO0WwLW7W3g41DnX66cstuFPic7tu/URPbJxIWJmb2JHl96yn
lUlTybsPwqSujQuwxgadxZGLaEFTucMCxhL9wCEgvmiQSaGQejqVztQTdWfzEsK4
658ldyzqg5driGYmVdM0cDoTWZuvGjloqwamSbKzdJXNX36lcJJdAv7RjdggTxqG
WQ5+T7G75mjNKwXix/UIEWMP7GBNP2fkQubkvuFrLNNXliSlp19fKV9Vwlc9swPa
HY46uV2b1enN4DacfMUsHZ2DtFLVMOd7DJnF2gSAPUGxv7Kv7U8bujp7+Wyoghjl
R7ImaslEjUE/J0IuBYTQKwmGxsGIPYpZEmAcD4UgyEZ1Ik+9cfJhaWLaRnca0TKZ
KZgRJCBBpvEKxatcvlSlX4E6vR00tKXncFozCsfZ4vYREneGe7xwOommfrvh9TVV
4eU8NqYpvXepy8ICUJkXrg2xc9HYjXOdKGOEZuOgnBZZHwE+B+bcGTfsQICRHDNa
VsMZsVxli5aziyp0VtaCePoMcj7Z27e9fw+ZmOkoIi2sZD4EW2P1GQbXTY2Y54Je
ruiguHZWefVH0RSHE4f/pBH/qlw2TG3wng+HUBZLmcDXzxsAE/I2ssSRyt8dn2Dp
NZzUrJw/B/lIA7AqaGUaw20C7eXGOk9rDZi4/4CJZ/Qi4SJy9R4tBxj+6rwDRQ/H
FwGQfBv/X7/cBk0jkQ3dJimg1qicZiUg3FLv99ENurJyN2RVVcLV7mK16REi5ebU
j2ex8L9e+7uuanwJQwJh1XiXZ8waM6Rlc+396yTfC4q6oFAYn2JXV1Q8Xhb7cnbp
wAsCQt8AWazByqwSFYQHdI+CLpm0OidqCXL+Hvdfd/5DKexPT0Xg/98SQ7400FoY
5cMbiNqHcDlTvfW9xethFZEvPyaVVJwYiaET3J+P4bVewVck4cHwr6wZVcdW0BGh
fjUcpeA/3CKHw1Kf9DRBoyJ9kn3APZWL96HS7T/4jD3cZ7qvLPeBRq++3SHod1S2
CnK6ubm/mXiB8N+yU8yWRNR5sAANDtAGu/th005z8yjSeG0Dp/VdatKiJPHkubIL
zk0j6UJqPeHSun+8dRvV3xeNvI16Ixtuj8JxlPUHGvaS1sSf4IHtj8KFUq9UrjYH
P1BrrmaH+qxy0MSJcB3welY+16yWKXmuwpRMvpYiFLm98fFMAidUCkHXjZQT6IWw
Q8S14TymV2BVZxSbVXABouTmUQfBkbTY0J+7YaZEP6TLSxMtDdnWee7OPJDgQbJx
+Bp7XD08ACV4GiwWzDCcQj8RKBl8rHsPZH68LH+GwA8tk5Wb82nO198h1adBjU6O
FL/a1w1Dc07+qtFBkkJb87DPf4SQt5amsss+9Z8T12Ffio7yzJHJOaMja4UwVA6F
XQdpWjCHDUfllzfifFJZ/+Q8BzGa1Eef90wEZRViqnKNRsllCfLGgRyLN0AvsTiW
dyEU1j6WWfz1/ZWqqWYCZ67Kr3kvsWKv3074JQZniWrGPDRK1lUbMRZUlHg9Cabs
VPDMNA0/WScDd0NUqEC2eY2APCaswOD7y0hbK674CMRQTQaBbOwsfJcdh/GN0VY5
Q/x06U2EFTyrj5K6RArKehguuG9FzPOX7+t1LGCzVLB1mCtM/QPCRRXZvHEDYS3z
RY0+iKk7skAeYlOTe7mJVvxF6xEMjOoBRfo0un21StA0XybO45YN0CZWkcIIeQRe
o0hQ47lkGBoVU5HsVWbCxcs3UppZNzZ1U+DRcRFAVMlRZoPlj7zX4jcT8N9qFDDV
5iBPw8nfPFNEl6BYjek/D2bO5WQS3QRIrG8MNyMg15G/KMaceckTJPumdm4Yc6Sr
DoSaNqDdFeG4ZPkThKI9AJbbUY1SB2yalJSKw5x1cJ8CG03PNDe8fumBUnv19mLV
NLardphgn096auWjjoTRaztH/F+WKfsZX9EWRBSnRAV2L9rKgBNyEQZxbHi21cW1
x1d0H6IDKrso7vVlbBH2qTR/o3aenjt9Y3bq5kZjgL2dzSylCMlOieTOM5bwMmHF
nUObgmkw2bBp8tmk8OKcyQJ+G8qzfsqn0p6FyD/1fvVMNkB0U9wVSz3gJL42yx9b
Nru2NLzgEpga/YQzKjGuepCH8EIR4vnl0y2IjKJVVml5zsdo0xrOvyYEsUEBd0qd
sOH8+J9KLtcjS8qnlwHkPqZBXhPmO73TO9J2MIUH9/s5nlPHV/P4NTOKQM5LgYgm
n0cpqpBON51s0xP162kacakfeKYdTa466BCLiPB0Blv5NWTyhvw3n4sgvUqFv2Kr
LfDcJhEvPBD3DyRpjoBk67ziC/cMnQAp+lVg3cuWnrDsaO2+HarDXBFmfclxLfdK
izfw4T4wayQbmoBjRbaPKADae2aR1smR9vztce1Gn8Q1imrTgjE79b27UTCgG5aA
e++LEUn+f26rRbtkfERkwDitEFhQGPOMqdTdDnxUd1b2bQtSiQ0Ixph6SxlUvOVh
dBlfQHp9LjKBOKB3HkvtWQ306ZYNUKPFijl6lWQ7I+g/Ss+xZ4z9mzD4ahi1riXP
kRao3XsVJ+2uVqIbvQqAnMPscn+GOychdCXkXK6bgTsu3Kbg1R53b6dBsIx8nlaN
tlPn9SZurOeWpynW5bBzaJuVi1cdGIHVaKGv8GjmPcc19JLpK3EVVAPFwivfTxYl
ObzT90ZB7rQPB6P2RWH9K23bH+6rz3ZeKL5rPhIyCUe3xuX+VRFgjZaVmwh00zms
7zd195Zoz0iZXEt3IakRRdKRQZcJtjRNB0i/sihlDD66Cq0fUVgSDbHr9pSOSCa7
6wLfL7H6RqFovxv5pgd8h2LnrMkyrEUl/hpUbdvQiFIKBwN8hIYCk5PoHh+gsFV4
7AvtZaIs444OzERi2G9iTfWkGM100tySwO49KeE3GruS19AOETT4Cvj6tv5xowUM
lB0y7iXNnoZ5p8ZEBr0Thi/Do5cG6sMO5mKuvhS7TWm7MpiI05yRvQ6kAoOxtwy5
/OtRQTyRM591Rj9JvPRmouu6+Q+Xn6BFeEdxllX3r14UEuDG1LuUHOhOhrfWENBP
UdMqaH4iH3kM6WFd3+CLpi4if8YHZ0tSnvGGEaBxhLxzLMZcGqYU3LveG3r48Di5
q+ZiJ7HKJKcimTsw3GWVV53/dEoMGr2O4WjO3DBfeH5RaD+5+0+sl2bef1ga/Cxt
YClfzEa6kjwlRTBenwdhfv4L9a0RxE74mQgQwX/7d+tO//8MecFz9qC8T8fRSyxL
oHahfuskwa9jZYNxRyjDoo51TLiO1lfLq9QFtrKnHbzyY5mvKxioZaecpIbjn6/Z
88vrkceKBFyZ+dRkSkLEP+D36g9vJhEBl15xmOTowjoq2fQg7FlerqVEsbwdrBxI
xn4uU+pLXHWX2bqDldFVO8CLlsIjlJAXc0BdrxV/QilSgp1X/4j/vHlpuuLoGo//
EUuPiJV2yNT8t3EbiHWz+mCvF/NcdPT/GeEOnzFDPnqtPGC/CYOw1ab9DfmBOFbc
B4WVW2cMPlOzrbK9egOXgX2qAbl4ukyAGeYnuI1p4U8odt61RsYNU9CL8He4Bg+H
idOqafRJnjyAD5P72bdzKdHjtBdKNZFuw5E83LFi1SbwU9b8iDWHBHdH+IW2DJ61
Oe54oJx+c7OyXv51PP1v2zUcbxSjY96M0bxmUMbO7YV0b8DRiOVFKlrss8DIYmXf
ZNHSj4mxjO4k3zl5AwHhtV25VzEwiE0KegWsSb75uavjXIz1hXixnUj4tTfNuW6O
TWx/3v73ZEZOMkN5y0Qj0RZC39xHJSK5WYeC/iN5+QmHvW9VzDFsKrTphOcvoFTA
nSyO2JSw6IbgtwaOLQlEREdOxLKoeWlhUwR8CW5rU/xF+aGtI/Fp5l4ZETNZ+/iU
YbI8FOdSuZaA6WKLQCfwgUaHH5RLWORERGzHCJu9S9Wz1vubNGu04couogFFpt8x
k+nee6HUdRGm/CGaccOinLU5S3u5poQOM08T0gy/AmiLB2C0WHPrqhD1HCE2Z6p8
sHxf4fs9qrABEZXcVIWyHaAuzkTILeNiv3jsc5icpFPzHgX1aGyujLwF1R50ZSMK
haZmcZdN342QiA2iKFBH/1GJGyTVLgnrQKIBr5bZ1taUYYiWF59Hj6pfgYAiqmMp
qDcmWZFy3I3LKgwTuvdGZ+B+VC2iFd9YZD5CtQhAzJwIQGrVRzGkFWb7Pr+nBDf4
9j+98GxdOwgMG9ZlS2FyPcZm4hAQG8ZQ3YzoVFAV4qQTpfeSPJw/nvEID+8dFCA7
cUneHutYUU6wZC0/8GrPaiLY+c1ZHiKKzh1zY63uABWemNg9v+k9ALWhrlt748gZ
OXhn23fD5DkwEZAXG3FRoASNy7+ZxXGuV+zpAIV5/2rl7N44Bjxg+EvNbQtb2Koo
ikCsQID1tRnzTL5E58E3ElIatJ/hx+9vV+G0cmkeekyFQbzmSUvAMYSFg7CV7qPq
Tqu31uWKRuvATJ+E71O7/S9AusRZZ25PZ3mVggmL4PDAJbygKWmpgUlYa1m2ohO/
2u5d0f/zB+pGljT06+IyimiZaNdySffRZrck7ulpq4sP+7iFA7TpbP+m67XpFhxm
uJ0a2Gdiy75Y3x80DvYTi7fEA6Yfw7SHNb0ufkDxcQaRmki2bhg4dxJ1bAahT6+R
sWKxb9Uc7DgtyOhMmryyjeT4yk1jcV+rGxb96/OtFRyY6om8v7XNJOmRVODG3/Ws
mvG5fhGylq5MjDXOrGbbzEHV3rLK2oVbmpGFwkdhfpfAUjhJtygdApBr3yn2a2vm
XozT45B/D2ki68OsCIDUIXMr6MM3vKBrRjy5IolSZIlGQjSksSFYER5oThTVYkX4
GHTdkAccUKgZjrlbMkQrY2qHQbmlmQfHAlhPtPc6t5b+eESIA519qJ6A2zf7n2uj
fqLnJ29nfUDOLPjs1OV1LM5d2brMm4WO6ei78Ls92k8qfU/PUrf2v63UH2lbCmR0
ufk6tLN7kPM48omPONwiQtmgJxeLukiUhdDd/heO/cixXeJo9lm6mAAqTKtMNJuC
2GU9nfXkT3hZKmGx3d/JOfzMgNrr9Ebua32Vm1UJBuwEry/9N1EP+FQ/T2eyd7Mr
ibF3IDuQwDMdXFgSBcjCmuIx9axDIl3ApmlVm5iTpMLPCnZ7mrg689SeokL+7qqI
9HAFxsg8ytZDZDKOxaD5qI4i6RR8bZ6AF6TcY+swluJQXw+TzTacvs1eKlDu3gNF
cIMRNQwqSvdFbr8weSmLpVyvL9PLd2qspgWqjjOSW/KxFA2cb3Bjyt6Ee/S/HEIb
hO76tB/jTyEx7vhKEv3+G74u9zPbQOETlEloPCYtTfNFgo406LJIqioq3NBWND3v
6jRDqmaXNTgcj1FcQqZvCYQAlPT5sXpVcGBFFD6tfLi5OgVkJ74xkRyA2tUwXwZQ
5sI8TUpwl1qDlfRQOumcwm6DafY6L2pSOkAiq/5wdTCsCCbkklZ2eqR8ZU4beNfr
0fTCarKLhnZwUd2P0af0u7xQAN4Wt15xGuQph4nKInSJplV7BHNE+7X6L8tFNbde
qkW1X9Zz1U2EzFt4EdqWu5cujoLsHM2JjScZ4LZ1PI8Qx3BkhVqtIiCR5k2EO0rz
879SOEcLj9mVETZP5v+Tp5CjaeG6x/DA2xOjoIYawYAD2sHqDx/s0WRWjxUjQtEO
8fBereNTqcBF0WQAmhQU8lVzKWsnAyZ+Fbqa9TRL6pYVaVlXe4jr6ud2KBfsLwtx
IeSy0/ETOCsmYc97ZH9rTej2K6v9PyQH3AR4upftDFr+KDILnY4HGeE2AP5L2wQc
Pug0k6fzR8ABWS25QVlypJOf9laBAgDnFo5RpLe218x39EB41VDPMtF4p8/Ncbpi
nIxadnjszX4S8SaHady0cXKOeis7sAnakZZCyKZsduSYDXtCltz1+pBIR1v9lThJ
kDTP8fh0bLwElY1P2ikuS91FTj3mlkoR78h0GBBvFzOct3MTMjnRMiQ2nJ9+gVRY
LRd8yjUbI1XlkUYgz8h4EDJgUGKpcG15cjmLy2Wodup/99NpvyDzUwffonSL98q2
CmoB9CcPeKkfQP8xdFJdfzXexEtkmGLp7+DlymbyXRTmNMaFzWHaTtG33KlflLZa
m9oAord2VoBE1Mweoc+p/IstS2hOYrer02Z25JxMCGPoBt4fcbCw0e754Hvd+gdI
Ga6lzpnjBWW+hw7o/5IdG9pJfIDNaagTDtc+eEpRLI66NLRnR4eguabChISbgOZH
iDWnwQleZgnG0Dywv76wljz2y6BBv5o4ZxPRKx0P+bx/fsmFhhMMeiByj20lV9ZD
tTMvLsQuzivqfk4WD+zDpE6VFKxPGN1KyEenZ35SogPJ8gQ15aZcmCWKJHuWkQNQ
XMg2rwOGWFiPtEz8KJyRk6AQY2ke0/JLVDFJ6d3K/+aSOZng5EWl9ps9UKRvLkH8
rm+ZlGzysQ0JZIFVhBE+HvMEn8V/AySQY/+WwbYHQX/KX3YQjKBw9rZDBDOJjazK
OZRYjCws89wHPOxCP419VC//Bx8T0Kic82ECzh6OPQxPK80DhWOQN3l4MkJthPbG
mlmfuHMJwi0EFghHVeFRvGpnGJzwpGFLXb55JBK33WplTU2yv/P75Zvn/tgSg8m1
VDofyzMr8UHrGJ0u6Wvx4qjlnNySQT6zMRUeO+DSrqhxwAG4aYS0Dr3sUMDr0AO3
qiTBPdavOI7MKcR5y2VSIyDX+uAwC865cyqFwh1lS1eiIgvRukd4yWoPeHma14Hf
bBTNVJEIdstdiBBFnHIpFFKHqM2T7aLEs5U+WnyQQ5VDWdlKazlFQjKvg0AXNjt8
nr2micz20dSITDRe3gA83F1xA5rO1SEktVJwB0KlOrwXe9WpP1lBiTSGXUqF1xUH
o6ANxqbvN05NcooMpwaWCVfMFn1ZY9cgMY6qC/OqeR3v++hKnN7647bNj3u3RkSn
q1zNDuIVs9J6+iI/Jcv6Wq6pGH3GSOdqu93v6tsYm/Vj0l5XPfHPTBMZBuk5fs0m
UhOT6QkVza5hlpnbDkUjX+0eO19dsrBY9L7z6Dr32ekcZjUk2rgCP1Uqb+0Z+DBJ
eDcUHThxHjt1b5vVbMwgYcMXeQCNEw6eNH9xvJNqsWC4n2/dVHP7v7T9yJeCDDDW
estq7dihSQ+mbHTqzWy59ZaHJhX4bYVHgBERONOgomn5w8knjIaP3Tmv3DfpdD2D
J1oQ1mz2qtymAutG119zxu3CV86+w4+6ZvTbKu28ziezf/yO/KnemxPwaL1BU5c3
bwYee+DUBDPH3PJsBFiKFj66kDRtdTxrKsvpMoqpMDkRgkILxgM2jcUX4QN8W8SJ
p103iNy5Utxm9n/nB84MJpV7g+sN2XBQlBsBYnwLJn4Jp9u4YO/JkSpTZcnYA0a0
0CHe5wlXKRDIxFSYRXvUnHWIcIUHLqe9/I3X+5Vxc/GEdw27lrw6Ma0vuAtwCzL+
FZc/6KptFQnQdBWUhkj4PpCu2dOhh9ZjGcWwSeFZCGFUZ1Axa8wFD3mJTCPBpwye
Ucu3P/v1nyBUK0ngJDvUvMGPi+uRkBNd47QHRQqquFj9d13BuoGdo7/8kQ2Vv+kn
qT2rFdUR7XwWG2revGYyLo8ZESIj4MlUDdm1G7n8m+2x4hN+BefGzPOOaNigwX3a
Fs/XgDjV5gv6Zc/jvMm1hbrFztK/ND9fQXNlwWwufdLU5kJCcplyGXiy0aNKxxuk
AKcYT4/Aj+FFUrckR/2UXIMmSEHe11fKx4HrLV9JsAU/86AXADbER3lxCH4D3/jH
9y6CTqaBMOsTtcOdlc6roieS9pjhKd4DVfy78bSrrr9QW9jKHIt4XX40S3Kc2xUW
OYDstktHiXX5rTzWHiudQJo7YgHMuM/wgPqd9SCz8GY/m6F2KE6gpwh0wZsFqZLU
DoVUJfsqYK3dYZ+wgnUa2qmxN0/D1OmvLm5/kvkYU9CqLwCI1IIiHbwd7pfLY0+e
Suw3To3+ORuKQpOTVc8Vv0v4FUxKIJMfcZDN18MmWTmGTK0YlYTF5pRuB31Iso92
ohhSLbisDJeMRtRHy3uWG4YpjIkmOv757F+zRDezAKLbH9iTO+Gjl6Hkc55Dkjk5
NXmql4i4PZfX4UIVsBo4dLprFxiS4QLgCUOmbGGLHVKNiKYW1KVk2n/bbmYuOmNs
ZKfILBl0C6VSlIZGyR65UyaTbsPVMzBJIXVeKhqRrzYiQ0a5xHGCvJlANhJqj/v1
lmIH2ymuBCn5od4j2306vX3hM93x+t39+9zh1s9at5ksFQlTT2D7tBdWTKiQc6XL
6x3/YaX1oqBh0mMDquYLsg04M2MyH7oLcZiTiLLyE5EfGFhQk8y3kYFc8k0ug57b
+8BLHffk+KBIK6fVUoEtU+N09CZ0qBQeBpFOr3DLyZNGoXeq33+I4uQmtnNboDK4
nso3NM1tAJBQYJpw/rZP5gcOqyC9YzSVFRvdxTnt3QqgFqWNJIAd6i244AH7Zuoj
L+KCJuj1xTJqoTKc1SN1bD6MuW+s5bfcn+yRE1EjKPdn5wDa/f0kfRO+TJxagJr8
V1pPphtN6IbjPVIa42WCbf1+DdA5nn06q9NoW8Ddaym0GoJQFYmQK0MibXfrKrN1
JBAAeQ+Qirevb6FjqhmTY/W4pCLYf2fIV2NW+pDkTs1SakbY4L3ILK4POx6Et3/Z
0/JpIOcoZ/UXE1BzkavGm0yVslQFml3y5IiA5aIvd9769PQ4Gb8FMxy73s5YodlH
gBW65gliZkUYyCICzd6yCAT4pUrh4aH7qEOTViRo7E063fwZCiJgaCsy0ZCRctNH
ln85jQbxs4jhex50QZLh67QfR2BNKwQOUlmZcOAGYRV0K2p/LL3wdJvmyp+D1FSy
YLcF1eGSmixswBkQ5QApHH7QPPfOPy6Csfra9jFyLMpUeVGxBAWXfBHMMByU+01F
PWxOYcADc8sSLmldiW9yr1fVr1um7KjeL1IQD947y5kgIJkCJknQCXe1EL/yCg4t
iuiL9O8MKxmuVgzzmZACWX/flYiM+cT7rtPPNBboezOKnoJgkD/4LVcFaBryjxiN
omm8w0r+kG7K/MFLzOj8oHO2mB0wa9gTzvYRqief26NVjyp88PXcH0dBga5tm6Ut
Hc3bcuCM+XtcfuiEUmgNu/xCicDBDaVKraxdjXxF+S8qeIQBlkrIaflWE5DUvn7p
JONOl6SY5oMQ05sW5XcsE3VmtCk0WIwVhsyF1jK6zH7a2bTm3Awhc1PbfZrGzx5b
aHibQMN0hNhL0Oe2YtPlfEDTuosfeu+hT8Kt7t4TJAblUEb++/1CEltK2EBbT9Rr
IZYBPEx3YxVqx/RjJZR44DaEjbicI4mDpNriwQZ0zlUltflW/8YNYHe2ymmD4IxG
n6AS1J5TByGeOLf4oxZctvWhW5NQ420YUaI9aKiyHQdn2wuCrRXZtu5uI7l09bzN
EfXk42XfHFcxmwOSzmgRRCKwUV1uNFectjKQdmhk3Y/ZR84xeSe3bHhWMPBNKEed
6ccCafezgGp/3I6PGo486FVfsNX0pBOYrwZFfrddO2c4d4hYSTTgda2S7U0QUDW3
xa+32O1LZctAe5rBzhnEy5K4E10gTsS2+15Mf4WnSYs3F7BjFqXi83yZJnj/+ik0
0qedaYcklB0cynbYpTHFj0LvDs9gjeXKLKAfyskOODD7n5VktovwJ2+gi71Jtitg
EaHRVW/iP43MJ8XENJ/lvVeut8xZOmilPZN+LylP0FiH9Mf+jpCdZRU3zZaJY44K
/m+aK1waB8kP3tTg3xnZU1BzQ02aAT5VO97wIHd2CrOqygxYfSYGUw9czY6pEJdt
Tk369nix3UHbYorO9y7FX+VFAmjWQPdw7tYG/jkFIWqMFxuaDkdlB3mhRaO1tCL0
0aItjTfjrhFZ5DHPnV2YrCNvcpz71F6C6+hHCojo8kohEHFvlesLq2xACb2VimoP
vj4Z+HHF9Q8SKBFswLI3kCymsRTLy8ApZ7oIdw2gBQiXHwr1G9kvTM94nEUTb7Cn
TdqX2I5M5cvO8T09jSFVmQYXgtLXNpQRQQeTW/SFPETzFHPPd7Fkn/dnlg8oXbcy
4dcMKXe4Ezzbnvb++0280EWoIhR9wsdfoVTZfj4F31PBcrj8NtTL1LFGG5KllH2g
Lls8NhkKJ0WAv0vIc1sPOmTOshEhEzbZFWVT55pSUdR6ORpPr52Wtujf7pG3Hzm9
+2HpaQGNM00haLif3Qqz0bPr1O4lBe7EgQXpZYunlSy69OUHoqVCd4QqPc4MJcJ1
+sL8v5bl27iASnIAPRdD8F/1lXF5LX9O/Zvd5UZGOP1e/vnkwc9sdzM/HUUyT4NX
0hUor5e6hfLSzoMW+O9zrEoW2Dvlh8LWimdovr3Wh+JOhFDHiLQzE8g8EPELewBh
cUTFRuR4QMdaOIUpsxTTzqJMWE2WPRwtwbX9r1QyQgi4HkoL3vUUYtvGK3fUBFXa
jIRjenRBqOMlrdTUsA1Qo/SS7s5eW3pmCAzk5u4XPwOQc2js8YSpDvXbv/paXS1H
7/NrVAlDjLtiZIfnLiH8dd7eJ6cV3bIoHIuKhObXxrQIJLffibUPeUtQ27UMq48X
HvP5goLZeiaiPpKrJbHfD9kLauu3t3q5Q0SVPQoZzz9rWQNOy1ZTS6IDSueGXiFM
9Gy/2d85AcOHuao655lKRIvFd5IMSGjWNpTrrlJlmDgbP2MI9MIkGKvAH2gqHQ2V
ghWGqitlAVKkznbVx08AYLpXaQjHeG0r43l3PfBYL7sM8+6n9kPPK20y0iWIF/8l
DVS7YQmQ5Gwvq0MnOLahEBlqs/v6Ux9Q5Yr67CLLqSOa8Fu9EZcf2cjiogu1zjzN
MoAyaF/NyH/CLB4EIUk1Qg+GrGECtcIaR+5cfW/h3xrtADjHEUxk1yw88e+W/Y8Q
kiBYvbWeIG939S23/l6prpcskh+Rs6oATANs0a05wRz2jTXl+17qGfekAUz13Nbt
wmiidGv9QIrepS4GYbFN5dUKdKb+KuTyUXF1+Ube3oiLzmn/XBY23x1XkQ6I+Vob
LBbKwE4t7KPVT5WMkV3DSRIFuygakUc2DLwMxcjTUhW0WFQQU/14V/WnCir7vDAE
N86lvumIt42jOzp3KF/rvV41ArzC72E0LKdlxmCca3mJTjQarUuxVTvUuy12XBiJ
jNHX03/YXRtWNpvjzHHxCr2FOV35Hs11bmNgLrzamXTsxTt7xa9iIKmds2p14wa5
qsZl4kF4tQk9hR46PYQrl1XHPGKSPkdSdzwGlO6iZYJ2bWC3MY1G5lq4291zwJQu
44DJKnu4lsG+VriPx83Sf2dlipW023cnZ3izMv5ksL5sMCE7KjwI6SaG8dSbrna1
Ndn2CCUOF4kqysrqleYBqaPk0KBRYXfjEAy+69tgwb8oQo/ieSiOKDJc/Z92Vz5u
mFoFR2cosPKLH29Aiug+vjpDTg4yYeZ+jsB1/8HzchRLmnTeYVWA1LhTKhU9Bjsu
TonV2Cd1DFXHIiQJr5olYNQJUlwmrHwpg7qch+2/q7uiZ37/OwCkG9v4a/o4mJZ2
OsBwOOR/0urV8RNCG5QyM3Wg724y0Y5Z2tM00dbL8puV00CBLd4i9ucXZPRp4iAR
tkFrDBxj7f12RC6iO4OwW7RRTI/ItIeuln2l8fsqdF6GPIeEt0Ru7QSl6qM7ppxU
sLNAoKxOgJsIiB/Aawji7EJyEnh9ryg7C+8ZDIm0Zo3csMXRoYQVGMIcb4/G0Odg
ZAuFple4VeT3WLvuCBukdLMKxRgSlSOSBFaV0fS/fy54idzzgt5p7sq1wY5PgXUK
Msjxr8Agb6LNbojakrS2FmyhbW5OYyE/p5jVPToBPgy9M2l1YBfzbulhnOZ2B7Qb
iaazGcNmpEhC2/ZEFOTiwabRCmtKlVbAT/Ws/Nac9p4Wi9LK9YOVR7CcQeoNKir3
2eHzdlsCgQSFr7YxuUL4BE2lzwGkDatD0DRtzB5kxp101I2Rxfp4BIz/BX4O2NKM
D2j5d8RwvsPTGhwPOzLQlud3NzRFoqBq+CDkDc3w+qfiSqGdb11N2iWVwlis47lu
CsD7tv9dVCCCHR1ywCzeznyzwRE/Hg4atYSIuETH2uU5qHJinr42TDFTithX/NBC
rFgcWd0JRy4BXOtHZNvjNW1HBjkkxPih7oGK0fkbjRNE79ag/AYUgx8y53nbBUKG
U7t4G3H3yFNG+DXTjtICdeu318JWB8MZBwLTV/b/28jHjOmC5LCf1F/r17jIiT26
BLySAEykIcp8iuBWC1LiQeERq6ifdtHbYLuwMzAg6SWTkpEW+PPZcrGsygYzRPKP
UCvxZ0ySBrYvEUdi0Sfl/L4YeEjLnCccV0pfxk13pq+LSaqxwqyV9JLn3Exud53n
wJDxwKqJk6+S6aNY/Jw/J5DOP81BfDyz85VCm6WUlsiOfmt6uosKrbVQDjEFGHYR
ldMUcKPz5pfnt0w9hggr0Kb0sitnRWNKnonEmjPEJsI7kk4k+LsQ+gy4S03VUdON
knt1OoDvoeGQrel6cHgHRB7C8YtXUlwmbpdKUADavpztbFw2KqVY3bV8napJnYHk
xmx0TXY/5QyviasTkqBiKPAZobRzjZQJKoyPXn3hgmApYfXAjGcRD+6AWRKzmQn0
EGpiOHpL2QvxnNqpJGdNkcjZD5Gx0KZDWYq4Dkn6vOMzvGGD76ChFABlXtW6fBqI
dZ3C4BIkky+ZqNqxGGwlYAje0519r9P6jGzUPSldaSH81RCRX6bJzzUPnVEf/65j
Vup+0yCxQAMXQ6+sY6azAD16i6sb6WNQyHmj+suim8qDQHebAnbbs23PrqKljE1/
7Vh0HhpdXbP1cWYPbzABNC0liUhDoGR9InhDH+rns5ETC5gnED/NaTMyI3kTqD6L
x1YuZjyISXDLLVskkHsDKrCUhyHOAbG+V/mHyKBfd6FxY9hk/JYdPS4itWKExrkN
eNa9xeM+pHyS4hy6hdWfsYP11dq2cqZrYix4mYYaP/TTm1bk4AOiqaDd5l8sM/1w
PdbYCxsZEPHaKLtiIvz6aG12ash9UeJ26KH/sYwNP9Iad6KX2+VDPJpqhk4TEO1d
IkOTtjclFGpYGdGJsLMzLcO4K/xNtofkev/G70SESYKWqq8Qp/BtkeSOPtzGB6ss
K5Cv1TAGnEoW52VGDsizsJp0+5AezazRaZYC3wnKfVmMxddKmDo2eBRkNgrovuhF
4GMLTVCN2kKe5LBG+o8yasZP/xFfM+wNQUWdaS3V6HB4ExZ6SJPK1rzwNzvVDARP
V/Hk4FN8jKhSssFRG3RECM83/psVDSRTvXWY6w5iLSe1MrwcJAAyOPbpvwJX0EF1
4nz5VOadPRreJc0AFBl2n0EiASuK4mI86uZYO+kYOAjkEfg4/t46OY/Pyai83FFs
OgR12BWezO+rr92leQiAZP/w8pJgKJMC9elTPoopHUTrqnLj/aGkJ9csgAftHT46
MJ32djfWk6kdijf/O1R0kv4zLoOg0V8ay4slDUGHpfPTESzPFJF5OtCgJySwr/xq
gNknGRJrxJvGBPKJlclEXCF8LEHYEX7Gz+8nbnkXskkiEkeX1Do/cgALo4gMvJCQ
Oj6r9969OAwcVM9tQGPQGWRMBVv+wdi37cgl3GMpFakHtmPjP5H92vGUyjExMxtd
xGHd40LbjJlHP+O19R1xNOq6Rla/rfuTTLWavkfahcrGAm9R5eoGC0Ue/Y5ZXR7s
rtUTYqYRNSJIFpfPFO5bCnJ9uRZauDcifxFY80r6nelQesaclASaXGhsM37rske4
3//d73INDO4juva8l9V52T5SYp7AyRLwwLzwuvRIWDbKOyX2mvOrue8SaBBxj/Iz
EKN2kYXgEsNPX2dlkopPd4Evk7+AXDkmXRVVzrE9GsX62+ICVzpU8yzNVTvXo2Md
dmBzEsLDNlOtvQ1er97IdZYpG7/5poGVewBgKnAKPz6BjLLJAjFqF/ytdz4v9z5i
xGGM+IdstjabVYcjUiPEY7MASJcNdXCrxnMCISFuArnDywOUj4sZDha5UM3bmo96
2jIxH0wDF8jO4DFaXk+ps5zK+LYE9L8s8WYL9LdzHdeJW5iLoVyMxfdEHMcHnbox
ZpCg3kLTJ4l2ih592fuzg7t1PC3A711lJyU1rzb5G3fZGiJozlvrkXRiZgFYgV/P
KNlNGiYDIZr6bcpXVn0hASGuOdVKeWIS2BsbI1tK4BKeuVWZGdO2VvqT7h1nY68/
X97Of9kFtoQy+W8IKrrhCT1e2kGIPtPnmVMYvL0oPOPdYclbeHYJDiRQSi46qjTX
5XbtimwgYOJvKVaxOcGMxutbx+l2JUrxWSbuI2KnUNUxd4YCli/Crl7ZiUxPx9N1
IuTnVkXHXGJCVBZqO3z91dcaaeqlPvvW+ASOaPhnnpLvDXSy7rvNiCC7q7pxOCkj
gWBFDm+VP+FrvFz6YOqYt7vFc6Fiw4whtyHWixr6Ml/Yv0j32gLob12O2j5R3KKd
Mpbj53xgrDUf+YM0fHLaPqW6PDkiqvNW7TRVD2YK/1/ELHk5lDrmCG4CKoEoXH05
SVMW5dAjbk+vBY8ESgRwMwJ3jEVMNbBjPda/oYwzYZmzjaw0CFaZVlVQTNFH+fAU
S+WEj7K8CtPJj+SC+w97v6bpNmRNiWiQoyWgPT7gM9r99cxEDpNwl8YGMiAXbwhC
OPs9K6Mg1iDc5IMuX1kdsOrgo4AZ1HDkdHRvAl7pvEaHK7fzmXTjYhpjOUQRggvF
7wfN4DcNaOkjwI+jSL1LpKT9PpO3ji9AOLl6yJTG7u4IlBq3EILVfV4ywJDkvjQx
M5fqCywVT1oBYWe6jR9VHvMLkoYUvV5WZF40upwImR8v83GlAkaDeOGTiV68i+WF
HK6/+LwuoC0qjkXy/WHUWoI881r9Kc1I6lKm/fZSGYmUBMKAs8MmJsZns+5ND6VV
3JSeq5arnL2a0v+U7qNqdzXqjHEKdGdaq/He+mhyZnZJ+hZ7tiu3ddjQXOcHYqwq
2Pt+543JRtMkfUTXdm5mVb09Ci2lIwWyZoUYna1B86zVN2SBCT5xQYyBQfJ274RZ
v8Cj4fjcuoJcJ9/csDJAWPVG+U451lNJTT6L8d7maKBYeZDV0YCmesfzehbd1b2N
gKKLPZ77JPxwB1Eau0vOnynPcgJiLFokDYuChEY1HNHCXymx5jk+I0ppuMPviD5I
i9U1dSYRopvuxMeWWe26kAjfzgtjv5o0JU4tOUBmpP78K2EWUirEB//w15stI+uU
PfTu+qMxDPTY6tKQ52jFgxhv0eVOsXuKfNsnxjEbagFoiJ4X5nlwjWaq4agXTSdY
MZTVG0vXIrpBto3AR1vKyktFjh+J6+PPSDxPkjDPiLCmJ/H7AhPZ+jOgAMwG9k+A
OSuQDUik5O33WEKk1Y6rzGw1+3uyqLp6JGn4Xv6x0yvwcMZuEpPb7YP6g0t59tQe
bOI/wG/cmwwBESEaGkr/785CF3wAIL/Oe9nWHnNo7JaOkyEyGSEPXGbwhltVKQNU
IR6NRl20DTbAW/ezPWJJk3f+oAHAEdJcZN2nzQ2FG5DSs45xRXWyRFnpsa16Wy0Z
Fa4Jzp+4I2bcFZpsYTPZbrq4CPiInLyowZ8gPS4Qr60OT/E3nnVG6RkUzfhxpJye
8IWOCG5ikSG0JKu5ysZi1NE8OqDKwPPq4VVefstxBJwQfQ8WmVGOhCpGXnKo+XGy
J9KlDFaDfYgXGRHdyPDAJrr/UiA0F4aQPB0R9wpsW8AVfUX4YiQEhapRcRBjMGZn
JDOp68M8DCLxibU6TfNd/MEZxO/kuH2I0O6OYXoGxI6Bb2fvK8/uyHjSXdwQD3Mi
3/glm37CBMy2fNF7QXI0OUp05Z/dex7qng8WScxBuOSO7wmCzQE1LYww5pslokFm
vb4OKjWRf+G0a8b1jzgYvSSVgI69FkNl8MmCyD1h8SixFFg9+GQ45hpM2mV0Ifir
w40tESyrYBDtr/49/toUWxwQuzfdw0+zqVaGCkqAFDAkxNvGX7BxjnoogL2zEsry
n67cWgtJ6wEmWdrQ4rBnBp/GrCaoec0it8LJm1DXhQjrKVuw4ZBPv6UJHc9d3Wlm
eE9QsNY3Tjb77Iusfpk406ruIxacFwyGOtOIC+D9E1hR/kb7crPkPwXdm4f4lY0x
UFiBIDkJ8TLncJrgR9xb+0MylcnhWNw4QWhHa0pZ70AbooQlkMtGV29vrz2eMNC3
7qua0Cnykz3/N9gWTvk9w5CqwHQ55e8CIT1DZUBm0adI5Ke5rtYAhpPdSPJbcCCu
bBdmHT6qZDokORlaKLNF4utVSLCz4GyUtQqPjt48QjGzc7pJZavwjMJum1WQmL/M
MH3y/EWn3jPZe7PeGpv7pyuwA88HsB/j/cZkm6wkP1O+EkqcL5PmI1kf0VbtTJWC
gub8CYa9ciQvdRGCCzhGxKR2tsr0660rMoNnZNwkH7wCHxae3TIPAFmjBZQIjsbO
Dyb59L8bTrl7StJYh94CFDtNFcZKT6gbjOc8TXUC4NENpNGsO7UMUNqxufC2TXbq
yxsEdfATKTZWaUe3urVPK5Asux3G7ZTY1rYe2ZEYT44sRFreGh53Gw1PKtKRfUnS
8qv3pC82znIcDw7jqBikZQOEVtT9kUsLdDH0RblixBLWNthEv0Rb7BZalxCADSCf
m4zkSSSwgFBgInMBekXkzhc0fHiwtk1Bzc+PXrspzNsGDOIH+hcCwysTg24E+tni
KJ6RH6i0F9fZ1YcBmRtHyfqBpg/rU8E6c6Jsg5qGCdZ0b4nN/oi3ZTCgXYnxpBVW
FDofGq0v4agAqTRlFPhs4AuCmNNYDkdjw8YcNUmHc0CkF//nsR01COMsjC9oIt4u
hykIjRsavspYZtljeMRXrMnt6+Z2x4TSA8NF0AmWN7A76Mne4zPGq0NCu4gA+OUy
HTLNP4HPaAr/qqbOpnvfCy82fR+865BgvDPwyz/xPI85Oitma4qe59YKVTcGNdYT
fXpfe9tZ8GfyFaokDoePBwLmnQrzWWGQeSo4ClG/5LuVywoH6KRCuNszcbpJCg4h
BzW8vKyb3AZz4LKImFbng4JoUI7+Nax1RZvTjqshTcBgPQfuU5sTOlXDei5o6yOO
hYHtgPQ06tTMt70Fu/UcVf28Tg480UlUWjS3SwNez5dK5bmYh542q1hl7r/VQmP3
eqoNW5+UxBdvSxDNWA4B5O2borDBMZyfj5NzVbCasctJEseGyTdtLVuPwuWAIWBM
zp/z6BNRjx+5mDtZQ2jPW3PUT0YMep8ciIWx9SMbuAAIKg/Lz07cfed3zHrmJ54r
SsuSRxz9905+X0Xno2PghC5idf7/DhuW/w9mN1B8/EjsakHuOrlSShZCdvUd9Z5G
xa2LG0QK5c7+qSq2WYpX/4Qsb76dSzxvl8fcNHK7uNtfGzXOZ6/BGc83XGhbXsJP
dBt8v4UjJMGc0Y2RJYG5VZdJZI4LcdtHpBPq1r2rPYKP0vsLPRgW9pxECbn5Reek
0vQFigpNixf3SgruuqnGmsK2ZM2burrUViEC7m1YWZ5Cl/Ks+zVF4up6GexQCHMj
inTB0FWAHBLlGNFC83qIqWSN/9oEUXUZ0/yU/GktFb7PUrhWYIP9jfZeBLHHjgyt
Yg4w80Qlv9+RvMVOFKHPgsU5a7xHblmT+dKkqbXFAlHYPwu1hUKP/zpNkVKdMlgn
ZmZNi6DDEdoTnAqJWNhdRgTQzUhawG0/piTTt1My1MHruazkq7/PX8+5Z6XZ7u/i
bk3wuiKggEHqHuwOH2xRTsLW7Y8iRrKIIlllTIHkWa76IC6Pgw64is/TD/kvK/zF
ZpVzPMIxJ+A/0/u+YZHVGu9oOeGQOg8kDgIB8iy2JZV1TEBqkPgdtZW5bYpuwX6K
DINNzVyQh8m74a72o//kqm8816R+Q9NP876903b9F1Euar8n1AF2HcPWNtPQHgyE
iGE4z1JBNTCVpyCjEvqomAfjyhaf3tB8HVCsu2nx1qlHljOIJQWzGI86MZSP6EsH
N6hqqofVRl36V8P4gRGfRH/Kj0EU//D0GNKREqvclkrMwvv3bLroGwDYSCaFixiC
ZT5q5TokQLMxoibC8H15vkpEYHsT5C8IP5cSNu1AE+ALwhjBNa995NaMixRquEwK
El1EeFAnGCQ+QAEb0eska0RX9vgMHwDOWy/tZByPULMy8UVO5dfsM9gXTSL9RvvX
FeOMEU9vcL0Zd5MFcW1hzU6axF2vbPZZtt/l9uyJsVzP0ZtU+daEhKsWSc79h0pm
/hUkAilSrzFey834jO109Jmun96pGAYM6dXYoLnL/M21/mmeoI5Vk4Y3vNwX84DU
NajQ6CBs2yTS5EFvlhSthERLUu5u9JEANRB3Vq476KT19FGo6w+J6q1zYFMYidwO
FPn9Y7lDlsK/JSfZQQq80dng1RN5MkGZ0N5C0PismosujdJbbYb7l4MD6ktZKS0T
A3zWqZoEspIs5AArsHkNI/0+Ak35MI1rzJcKZTX3S1Lvi4RHMoTYf9MW+D4xV3sh
XIY3COnPzhXjfCmHDsoMxuhRLaQlZ+sY4JEU2tuKQXJuJjHhDUo1YnQCifZYRK2H
u6QH4kO4XTp7/dfq5vP4VnBvpaluwpPYOBzBmaJVMOWczSHqwyVqEf84L8aWQo8f
+Yye4nRj9uWbq3Na44kI6MCZQhAD/RAY0GOnMQp+BMyF6g6RAraCSdT4H58tgZ1B
zBuZu11o3Tn5Vn/mDrbF/jUqbK9hxi+jN1/kiaEF9se3ZnuHZEmo2RRfqlQgTMa3
aJ3WxS2BrkN1UOn58uC4BZJ5cji9zZ3m6XzfQ72YnS4KL++oGzbhsXS94vIhjmp7
QDTVWv6C6S+7Dic7TMsfCR+UTZYutsWfqyPLg6DG/3Qc7kXhEKvPAxAGkYOO5/KH
9mXJOQEDNgUoDnkD9w71OXW3duN0i9xKcrtcLEQwhJO1UYKf0p/Lomc5SyofHaQs
eMbF7JZMobGoSfBZMrUvIXkOcGaJG4KGwteEgmnmuY+ROivz4iXIraX2kMqjSPGg
UBg0u6D7Zi0sqoiJcHFQhprKITIHPchOr3D9s01rgPxvuIzo1FwZtKeDXTiNQ0yJ
iia3s+6s/SvFVdhkk4OPVkhhheRxdr1MZFfBNYz/18SPepA7haVtD6NKuA4KibJB
+qhIls+3GANuRA9sAJekVLJHMGLtaFyQIH2lvwQt+bV/lGL1bD3pJYhUKGQKoly6
cLGiZwXV46wLTMiNQpvrUIwbjRRBdMhMffUIKiqiBTwLvs4ig42ChES0G2pN/CRw
sDCfARVzF4KuEkoETFAMBVoJYGIpVVcKrdeos6gmwvhCQOmrhgrweW3zhPPSTLLE
AVFeONtUujblhtBlkW+pQRBbeQCvPQdM2hk/Y8ANnQGCl+zk6rrb1O+STMHvJa+H
Wmw7qOOeC+KnElODPoTtfrjp7VYeLwECkZwardVNxO/xbtqB6M/cmu9oo6k6p1Z1
8psQ9pecNXK+Y9Hg5w8AymSErsTTulJ30dwXU79DAiIKmZPpmwITL4Z25sbqsAPM
xHTZiD6cbWokyyfG2+IPiGUV4gomsHjBsDfNdScmgipsf/+eIAtE67yJqNV7ljn5
b78+t4cUCoYMJQID4EVxB/5f98C4hvDQeAnhFr2K+0OwEgBnRggxWzmgtuR9InnH
R+xAM1MG7gEfJ4liWSrenXzr7F5HGncLGAmj1IBtfyee7Lhklb+iypMxQScCcvJg
Jh/lf3m3hT3eDiVFOhaYrTgmIxJXbIHuLekk9OkjF8sCtzYFgieqaq6TRuMlzCOf
ZK9v/I6M/qG7GZARPaaWQFwGZReNVM3GOSlVd1xpGrIrrmN6SjMLVAVQJ/Enmr+8
KrtZDlCqP4IuOKX6VS+W+LzJ/cNYGbeUcqMMlXeTrQFRWeHNSEJS/C5eLwt7pHcU
6Pqw7SZgwHPlpziPcRwaiMFClSQQ3LutbvCDmjuLp0bKT3QMMLuR52yCGCz6NYuJ
ZPicrxJPtnzyENdC+LUtTQ0gmPRIJq8bdxPUdepcvP5GvGusGikn51d6BCF/GbFE
ymQnKaVvvpeLmELUBctUoq/HUHmESUWn4vbnGTfNs4ANTzZRLKA/nCRdTzI7M/xc
a5Od9C2T/UAg0BWXDOey8dp/BHt9BeYBVqICznrHgt0Ai5crWhmJPP8DG4G4ghWE
FNHawK9w/Jhw1NT60XhZrLmvETHnkfKtG36pWvH6bbmsWUsa3PhlzVr0lgDduuna
JFh/bSle49N79Z5Ra6txqJeRmEs7nIs78iVxDed1eICEvmo6S60G+BdU9ZR9HAte
zmY20Ge504XH+j3JxiHYMWJ/EmzEum6i6IMxp63IcSK/i8VpZa6xcWKDThcSeCwT
eI0Oewnrag6vTEgUTTh4DhDS8E0iL4wd6+kIq0o2NLNX737IPX1w4r9L7F3MJIeu
EdzLlHoHsNwGvJr6CzcLHMQqgYXmj7+HumL6XzypRDSn3ZphC9hphMZV4nfuPYkf
fFhOtmrCuMsNODe8p+Fzc7VB3n3RyAQDaLn61Wi/uVh+a84lY7cmn0wz2zklJCI/
whlU0YjOKudYIQ/Cjsr3JI4yehuUmP4+aYG5pz0UT4Og6Msuf6ha4AE1IMUz0I43
UjLna6FJ+YzKVzr/4fCLcZNyKYwNyXWeJoM3f4mdH/Ck57pY3VOHNwsSZUZXcpAn
dj/F92elpzaRp6LEA20257AJIBWTzTxPFSoIaeNc2EKBvCmDUY8PjpdwdI1Bv24p
prNx8w2S+gIFDIei2rPuwKk5/arn6uXIYx3RkhGCYyKHFJaKBADkQFRE1Dt4OrI/
mihuGCR1HiPxAeTxRfwzrEXRZDR25rvSj5pVF48IkmiWGv21qMvKkxHTqW0g3qQF
piIuvBGsJFSI2eZ1lIyv+A6WbXiNqPPXkxnCH4rMSDQbOH5oZcZA6R0ffFEs4BQs
3szCk7UdNcGFqqNalIbi9yJUPRxMTofvJNtSA3nzExmcmiWUZQzzEMyou78QOcb/
TAHvJcHHEGpTnK+NOeKw0K3DrhNz0hcJLuE7ctyanv1tuYbUW78N+TcwaRTHMdd5
fI1GSQ2si+CMkg6hk9mmrS4tgFqyUExyg+tSsDowBfK0EVgTE8DKl9LBiFNOWcKR
FeSsd0ISdIj4Cax6hYBiTW5y5kikai+B6NkeGuGI+uILKNMNHUwCMUaGpV44byjK
YfYaphf/XMRK0IoAZ6NZpoAzKHTWI1ECXdoNVIi/ACKRqru+Cllqza4qj+A/JmRK
ztZugFfDSKrwiNqY71iWHrAOJBlyLRPyqlJn4pUuRqLQfMg1nCH5LWhG4mUWCMZ2
vHX9Gq3gBSWsTH7qKeo3aIo31xAY2vMG3W0SnoDVORbkXS5V7Wr7lO+Yyzo02q15
R0QqdudMFN4mTlZWj6hfeEvRmtKgjV0CtLRLvdJU+Y08xnYXxOjLZPowUNkoGk82
R2l/dp6a8jOKrzJRE8OGB+r9ysWfCL6Kzsar8AUDBXAGNMhGjN1yzPFV9ZcwEnwm
de4IbTTQ3OvnZVKQTGKaBeLReHjqZvjnhmSzGoqZxYAJOOvY7aLKdc6JgX7UDWI7
OYJbHSRQud67S/dyjt3l3A7Gyk85tVYuEHOLQEHAwFVxVjl0ZNaYApBP4i/Vj/SG
7kDb6xnuDjsO8/As2jk3SBpcs16SIlFGSzLQ4HRATI+IYmPH4xL8D4F4gd/slKmX
zxT2Z4GT0T4bS9s32h35g7ai6vt599OGhyK+4wE9Iqw0FaKPea9nfKs1QO+Gefte
yJ+S3yZFjb8vmHMS98Dp/KazHjpB1MQLbRKKnvdpyzwFJfGm31Q5QlIEnHfHOsNb
cGwdSi7PoqRjQ+P3asmfU1ObHEJjWuau3hrrcvpTDzHmQ/m8g2sMmyLhDCLik4Bn
MmWkAVT322olcZreiPhHswMwKlbpSX2HKEqe88JjWwF3CQtvUwSUFQb8JNU2q5cw
5jMuP5qD8OE3kFPmI8wHodSGoVGsEzaUJQQirS9vF4pLeg9tvykMQMiba+E7UYPW
0tkWa2RTj4e9DoHcPhxFFNnSqWect7C2wYS8lJFJWJJAVhvrjlJfBHhygNlisAM9
d+2+2F0Tm52I137HlTbiO7JHEjDCE5/zyme2O0gMY8fuQm1t0Yb/dDooqvTWX0q+
L5oSVZIIzptIsgMAS2xd3+GQ67W/CyvRQ7Htq/qnwQIX/YfCh1YszJgsFDZ54s3i
Bn1nngjt/X3oEpCOC+Cv4Jspp6vbzH2cmr6uBSOFkKH4bDmMHgILU06TqksKDsGP
Y6NenQwhqIlte4MO4bV7Hwlf+hamT71ApG4Jf8gWMU06lBXk7Tnf6zJ9K5SpyWSF
H2MujleGqWGJ5wYJYFBLT4EjJtRzZp6MF5XzElfsrMydci+BtLgikRgDwubSC7UJ
qoJNmiNQxZFUQ465iGd7SJQY1hbNZyXr1Z9GWDpHHNWvBprdbU2Qzt4Zj6g1XWyu
pvudo/WiWtGuv6y0UVsi3LoRJvjCxdKSO/lQBxXlio+aRwaB4LYwUlOS8EZ53lNJ
xEJK1TbS43sBlic7YSRyzfyzllkDRMFcoo5tQkhtP7oWevBdQQuRrPBpMwLXRT9T
cL4FUMFNuB5Q3QliTNgomLJ0xSY7WlpvVVkQ238wBZilzQnylUlDHvywAH5ENaOx
UU6cbOxmT50qEgyzha/PQFOJYqyu+Qi7S3Es0VzbP019KylVg3+rqAF3UkwIorqc
ju+GuQJ+NIUsDySMtBZ3BcCMTJNf+wEOcrGQMzlhnW93mPJWDk9QLLYxRtxYQ0vH
YwVOoi0oBxweWfTchxTK8KxA0gfQaTVFFHNURkUrWLkjL34o+7gbSY8t5t7FkLZ7
K94O6to2PwdXG5pHtt9uYc6bz0Zhia05mDTh2KslSsr9LuaUAsm3/6VU3fK91IDX
EXVDL273HG5HtBQPsq+CqhB7A8athsRT5K/ZTdX6fREG8ucVYEo2qXy3bQRK4L1F
zCpqg+wa3EvFlFJmOBtLgd9/xHyH7KZYU35MJfBKLqm0HNBeddiPZKdhB3ighTdu
0eosFbAjKd18OnPW++1bYZYqR6tsd1Hpqui5ZPNr3nexCOGHfKBiJ9rsuWNaPxq2
cvFImODaO3SWVS7jqR9AByl9gAskf4V0rW7k/wgR5RfpCzVzF6rNrLy40902aycJ
G8XLmyjGFDfYFMp9QhOouneahftCI5vgEenL7Kru2DRm1fQfaVMdtuz1lyDpvUcM
+3IoYWXj+AMDgz1+1L13kGb8XfjPiCMyUI2yUdNctVKBSmPMII7Hkpx6wOVFp/jx
Vvx8gDcgrOncj7QoBhDbeT6QuXUjxtW+lucVOK252Xkbzy5eCCOO/w4yNRF2+OLm
TTjt3nmEbumEwykpqlC1e3IDv2cs2/NZn7RyWh8hEXeQmaawIoXzeoWKM3bYOepI
4M9MloN1Wf+smuCjY/LJvvKl71IZdxLLqiC7XwWYSQegDfgP7aI93193oAgWAxAB
NC9baCUeeCxwsTcYSkiRS3Q3dH5+N5MXm4sp9UqeHCBW5H6Ot9gE0e5AWjwcYT/W
L4mnfm20uV1I0nRv5x82O0Y9hO111rNRC80UWqD3gcEidv8PtVh+isMMyCnDzfzx
/t8qtVPsNaXd1pwIKt5JKjBTzEoQKJAK9a9HBUDwONhoEQ7BZcziKClpVmbDmK2u
NRc+YnV/XZbuTgVdpOFP/Rubq2oG6A4/jzWRF4uuzKIKeC+1/fxan8Ik9GeavbiC
3TGH+J2zs1CCNUkJy8H+IDDB3s/dvr8qLNyniVJV0lGQ+enDnV239LODgfotygx7
mRTn5z6Tt/FA7ePyaoMDQ+oFeksXYHPsIZhGGkwsleOT8zavLFJ52Q2YUryF+26K
gvxaigKPO7zp0CvHR0zk+Alu1l5Mi4bXHwm3QmNFCrNG+Net6gs97YPS8CkKtiea
52ukPg5cZVCev6LzqegTZeegqotRD3BnUZRqOmOCeft1s2fMFYOfMBypU77XrQM9
0Od8YAjCJGUwnVmx9nR0xvydT8SIfPMWwzU4S49lsLzmd9K1RAdcPvTsRsyVGmHI
PsPOkBWA/yaqzoyKStv6XbAymJsWioBB0eAz8Ls8pMyemKNoa/zpl3pMt96WsEgH
uhZT3NVqYYWdCpYBckvo7uN1WVe5I0T1wilf3+DtlYeC/qXRXFAnEZKqiF1Gpc2a
5/ACTFmoCtnxaprZKtzxHSQ6/fwYx+QSruo/n8BrDCF9kp4DTxKs3+qU1mBvYguB
/9RVWjOPzznaz4VJ4c5lPBpGNdsjiE5Ws5APMFX22xAGEqn2+ojWG1N0pa+YJ5dN
URgYkrKh6PRuQfS5weBD1U+Xj+KjNgv65JEErRcxwbB5dmNvR2JMzC/Qt2khmC14
4GrogR1hR/6p/uHLug5FMunURxde3a5cCOzR9Uqy6+2dkm8Mv9xApc/MFU5gtx5/
LIS14t5/5uwsYlfPF891EgrFFmAD7GGn+DBjThPkl1497ajaC+Cquli3lXNTW4we
Z3QcjIxZdp1fnaR2zMt5PxXk7Mp4X45XC7FGESUIF7igUeX2IfGzOuSGQ2Ll+8py
L/Ws+IyEi6mKtwPJkmnlm57XRxcDUEse/5Kp+euB4fotKjyaBsJlglj4/xmlwicX
0X9ozpZsa0w9TqPf1GaSBygoK/u4EK4J4vYSKLU+KDrTFXTlwEkqUP89i88vXQMc
jVbpc71c3ZsBT0spdeiqODHVDWoSu735Fsogkqo/nLoVqhVJhiBuLeJ87KCam9VY
mgYkezpYOWk/SFGlQ6s2+ZG40iqVRpJS4iw/BMiGCFxi2oMSM1xnFXb19EJUCoEL
Rqb/ZgRiKUYIzR2jbugiTT9MeY8UnJH9BvHiFcG2FvElFdoZmMQjgRE85hf2Hd8l
Le9Z/Yt3r78Nb7b4C0GFKzK0WcZpe/rv7gbTF6XM/FDmt7/S0G6UiRxLGlSRpOeU
/NxxZRDMH/mzMcyRqol6JyKZfaTJ0siiNdceVz8oyrtzYekkOGFgfkBgCB1dH36t
4Mj3N2FbdUsjRkk02vntZy78vxuQ0yHVEyAAm7EQ8RT/XnWw1cIIJmlqaOMbYhKj
rFbymBqrGKxkv85stg1ONzZxPVRlJ7w0tnEiZhRlxUHX+QN0SZAPz00hbp9wggeD
HZ1Hz0VnL/y7d2Tx0v4X5kzyYldF2UDt7PePUHvX5wXej1PlkDYEwXH7MNjtrp5g
bfaD9T6kjuJQSJwGqs6iHbBMNn2uQrkiEA0BQBk2c80TUBKv5HyiCPVUvfIgTgXi
xPInA+7rNlPDBR9AmCm1pdg+itpjyoZIFv0N46pii1TFoDYiHIhwYhuQAv5fJ3hO
QZSIt3FGM3UvuYv7XSICyMFnePXV3G8IdfZF1E70GN6XvPhcIrbOEA/QPKuywCNd
jw/ZaiLzgtCSK9NQiuZDNHRImluUiEMy/kLSMnAbY7CGLth0zaq7szg524z3L6nK
eN5OUvJvCDaS1AMhUktJ5rr2sBvZwwpvxYY6Ru7D5p748GinsMdSfI4AHqOv7yI4
STCBI4j0vA/oWNGwggv/m3TgM5MgkFnCOiTrP8Pd2FP02RVnptP7j4u2Tb7sAKpt
EWO9xUgr+g0OCQrdTKbsn+CAuj+YdD21kzOeN4IdtR8nSffT+4LK500Yuus0I5bn
VRuNXwkbPhyivT+FSYuEt6xVyqfjdnx/ouMXPqtayKuGt2wRsgTtY+gSJbg9G+PI
VlKOAbfNVgUpYvWJV+2oU86EC9Evi9ZWiuGyC96u72c6fA7dslZl88sGdzFup1X9
IdijrqdvTqao0XKXUX7nHNqWfOnXTScBHyqkLG+nfq3zo5D8wXP5wG9n4HAUX9Bt
+wrc+zZj+PCeTcV3y0AAfvXvUpRgb/Ysotub20+VFwENm4gvaIYhAifGoYLr9lI1
nz31wB+ZKDeLbK2ZW5rCA6f1235m7vF+EUJTc8KK09HGapXWDqDihrZqEmw9K+rL
vYKFZZDwkzPUyHOUojSN739J2YVxf9kzA4FBZCs/A48UcoFYSoeAOVItQdUPQUIG
PS6LUC1g+1JWJ1y3/rB0cSCFHoUdpM/xMTchIT2K1EaLl6eU2j3AJ9PA9RYJ0uls
ot2kwSyiuu7rt1Hawxl8bMPOUZq0gGMeIJBR4o+BvsKNMS5voXJubFk6uWgd56hh
1PxTf5IJtUTzzsHVVh/QX3EYvnRip1drFMcF/PWTYF9x/mqKcaQzPp7whz7Wr1Po
DycqI0L/+xMbgujczBjcT0EDqdAUtA9iCfdV3lMS0Ctl4seZks1Fapmq0vGX79OR
gpIJAwJs2Dvv9Jq/3cgwalhqm899jbNBXJLbtg8Y2G+JeSONNM2d/vIYXAABzKtY
8jvNHpMqNBH4Htlhin4dVKUd1lpecGlAgix5jBmUXwEjaHG3EtPULFZfiPwn/XTU
Xq0CS9l1MH/+radFA/pWBImz8W9zzM7V/Xz/vvPlcU+KCFoV8U39ZGnBS+F1yplx
nO7OM19MnK2kBQ5MksRDwjBeVWQzUYmzcPtX2+mv+1U4om4gkgz6PBDlMD0r5nrD
zlfEQ+zRMyJq0voeW7Blcfr3yS0W7xevPqQ/+aWixn5uvSli4v+5Zvm0Dn5/gicU
sfsKpTxRRGVz/OB99roce8ztqFLJLhSSDA36R5XwhblZS+mD9Hn+pkifIPvZHdf5
JKSghiWrgANNSRF6axXBaXnuB4p/hQ6OTjlbFiMhUohPxVyje5GY68LWr7W+5VIf
QEHnbWrH8WKIbfZNUbsxXd6ZjCI/CEogVLZnyM+TJlMDaXvGGoTx/yoqNTDTOgvu
95rBCeWwNwL+hPC+tp9c3HckN4HS17iKUfZMtBeu/Wt2xUJ2qoXaOZmHQ66Oz1hQ
EOlZiWkG+w8i8AVtlT6YcQutq+/74QuASJU+Dd6kYaYDYP6HezE6uta1Jkf/5MM/
W7FQaWsY8ZfZKocRvhyTr1gaHghgSJ9uAs0fIUfnJMxUgM53kcmPt+9SnavE7Cyp
C45Cn7uy0qDy1M46uzxs7svbgLpARHaGQgczFJ8fVX6HoEEvzu5xqgD+2QKVvxGx
w3nd+Tfx+2ra4bUt7/lEdz2sVF3mH08NxoJ63WGmI5DZQcqkZRPF6JcF5GvKURhH
RWe5U8B3FPdmSXB1Dcl2rfPHEOJ24H62Pu/H5In7m3JZAIfzLpLRXP2ATpfdrk7X
UBU/+Nr9/6/r3it2EkYr5hiCEnCtrVrvnk/SsgwsP762E1b1e13os9HrMLFM17+i
dq+Zhz4+4HhOKb3RyLDw8jvixwgVD4b4H1ue5T5oAu61PZflBsBwTCr7zfZSnI4u
D8Mi/FHT8QkjkDPRrtxdrryHUJT5u9HnwgV4iEAS6HzNv/eXFmIYfIF0uuM4iUuO
B4zpYO3qhu0uR4nWPZGujZazgVcqfSzup6KOg2cMrrK0VmkS/NJ5AcRrrJ9mzleC
G7mn4v8NPx0Jhkh5gRT0h2J0QaSL02hXWmbsVTR4cJhqfjwpry1WXuhD1rsdDuxb
VE3xQL7Yzf01xLxj+acz8P6yeIigj6rgR4n3fECPcPO7wBA8TIfbgIbkFMXSVpsP
JGOQq/6EZrt5N4tp5VToW5oVHWQ/Qu0BIyAkQGN8u2BitYRGM8cPwjp/C965ruDh
c/0zPStrvXLcVJEk4RUmv73HKe7t7FJfOR0qm8QpGVTyrIk73+IB6EGUAeD+GdvQ
z1Bf1xYbyuQNMCw21r1gRnYyK2O9KcNh/Ce/15y+ZEoJV4Lesxedf+ogQGunpT0W
4wGfp8GJ9id4ekx/Wr0ToyhOMrsADyvR28wTsenFTdCEw5KFNcfeTD9lnbak3ety
SBzdur4Oa2G9G9E7C/bFNC99X/vGulYHDJFAuOuoWwlNDqNiPMValYkvOm+9r5Yf
J3k+bt9ER8HlGwsvOKEOFDrPF7FY4fgpZo+uwiuP3G3ubXxHzRxoOUnflEr6RQfn
Aq34DDcT7M0aJK7ZYtBxmZ6NC/WC8BATeKMHEOPxyN7GnsaJrIUwhpqnSXjRPIFp
RTz6TjOwNGKYzDdpF0g017VyOk00HEMU4l/1nQyld73MoUmfLqQbcWYnmDTKIav+
9ikcxTE8A+uyIB0vjD1h24idX7Fij4GJdu9UOW4nt6mBPqcR0uVwt1v7qqKe5hbM
+D2vBffDr7YHGPA0q2OpTKOJJSvBJA0zxnIAd9wITCQJEVQZzwBteu5QlNNy8U41
HBnfRV8uorwXiHOAjdvUuQRLbCv+eQE22YfdffD37eA+cp+RKuyLRLkOBk5mZY+h
udztFSywvVlGQPZGgIWuXquwk6kVMexFxH+MQWW6bmd3CdiIZxEbrqK8J97BzI1s
BEeq1fZcOluFkL3NBeG0danY3m9frhVEeL13mqNXOTaivOrrdwWhmbKgkSq2YjrP
vUifwFdOX2hHf8WtUeryaRu8qHFy+REIgr3VauDsD1HWsLehGcyywcvDlaEYwpkc
Xy4s5JxbfjPREF9cq2WOvir8kO8Kt8LdT+Iu1FNdv4kObh+8fxK+xk3HloArNYlh
25RI3H0S0OBNgWyCZpFTom1d1BPy1h08Lfos2TZzLscmvbFWJM/Fk4xK7VIrQ6pO
7Vo/hd5fk33lPj5TCwsVzCaFxJyEtuFQhtq9ClIDuWGOTCVIqfYK4UD/v9hXSjl6
fx3/P6qF2tQHG88WaHNCLq0GjqvJVZAcQ3zOkWkNEAGUK3RmZUvsfKuRGYTpUE4U
lMR81K8jbXqEB0enSDM1BI8+FTyGo4Q/fwzG+hPWh5aCDhPHuRsoMDrPhTK3UFyK
WwehY1htPGkjIowLmifFO0uVEP/HgseGNnGLd4TyX5YiC9diRG1LrlBFuZ4456mS
cK9yXh5RBB4lIxqzgR4FvIum0PNR6CmZ8yRfMQq2/HZbJ1cBsZOj2Yn1IxzIJwV/
wlw1Kh0c5AtZdwf9IUADG9oyeoIy/c4k/Yx+fzhw0rw3HLsgVAirOIHtyHn+giZg
bv/PfMj40ptCR1JcsUzgy44XZyfTrNEFILFUjaJO+EJGm01/XezuKDsxT5krFUrH
QUSltCAasqkWdzYXWIKXgEbWCoMdZG6P8CbsC52RyKLtaWTWONtyjL1KbQssxtRm
DyJcbj7dxWxtsHZcd/RCJWl+jdHdPKG+k35TbDPSEa0wYR+UA+Qk/LvBzue+Iq8K
+NZ6TMrmcYfrw5efTSXymXBXUtK1gI3NZSK3i2/Kjj3ZKKugB6HMKg4ULhZE21nB
VksAIdWiDfWo3pT7qgqMoVnfbvPWHLv/ASPf2rR1lt2hzcHFIUo0h8gkbAzMNa0o
Wwb/8zsEsQZN/lx5im5sdcFO/Q+0ZaTvGgRhL58p8KHwkT0jRbogr+Iy0axtzNBP
nNhjrvf+8Jf9Tt50ZQ8lHGJx/UfGyoAKXrq3kvJIXG0e8yzYOf9Jx9aUH3Er1WCo
Qk4+PNcDKOkY1/R6vydf6tzY10vkNxkjNYB97O27ehBRkFjxd7XI947rfw4OY9mM
LBXe1z1iD0Qg/r9wn/q5pR5Cc0IPnLxb17L5SMIzzC9VGZodC9hxQf3w5/oO3gKG
4kcC3TS0p0+XHIyzKhukNzwhTx5+KCI1n/Vt0HMoefCGY5ZV2hW9A3ip6/fVLjKp
h8UY2sXdDir/XOTXs6F2fYMVrrXYaonUnIthX4cbtJYu3SMjEJPz/KHUteis7fCq
aFRR8YfqWRPNNuss5Cj5Zis19VMfFjrg6x4897x/lJVu41Jvm38fQHoHRb3xDYpO
+dUjvn8aBfhvIedKzM3nrva8vMmUQuE2rBfBmuxsUCI5oc8SpxiaQFrObb83tF+I
yKDs48V8koozJupu2ypLfjcPvpI9AFX2Agcs63odzu5AxQuu3I4WWkL/7dvClCVS
Xo8JKTmUYNcRm1hGdZNS3MIUiZqqRIxoKex6jfUQrz6iOf2TnPJwPK/Wlr5MXCbN
tyNxZ2sEBOnXuL+NCOfFHrPxthzTRSrAW2n2zk68gLuZKdBQhdKYSGo9GIGwtKfk
fppqMM5DeojSZKyLLk9VBTd7Csw31G22FpYvMgHdJ+xitTU+qvueMAG8msI/33/0
JFbpKH4zTKMw7HwLvRSbW+l1nF614ujwOhsTDrwSRbnmiGrE3P2lpBGDl6ne8mqi
hfm6rS6QZNGEagepRJnlcVBVustiIj27i/UfurENcGUMrkRhRbOlMD0JYEMxuAQO
1cFnKssiQ7hKIWPKVhxyxWpEyw196bqiIKo9eC3Xmtfp+lgdbGmdW2ZjZx3imvME
mHploMx/PTON81Ht5dIxYDEK3ffNo4Kld8tMUoJo13R7Aaao6vc1Ltj+5yjeCTtM
XpYKwF/4PM3cU0+Kp0QmtqK5C71yoPhbNoEJ0vR62Mj+xQu+tgxSesvA2XBm/8W2
K/r3u2bYtkLQ2DCZkhhNuw2IXwwxlupfyl2zP07ZpYMerP8BsTanQOuA/CSAvDAG
m+PFGk9kkbYCwQf8kHUm3TQjcx9PkYKmz5TVFBC63g3qFd6e1U6NLfYlwbO9Jr3i
WUXGLwpPD5LVMPFTASomaxLTu/BXSatiC7EQvVIqQUDNphdEqB8F0ijMVOVXUcy2
ShSIyhQWy52zmeG+QDJgy6YW3nhsdbW6kSr1rKgZN066M+goFODJLJVELBr79yo3
31phDRv9vloiPftzMgHTP6UeZ9852Im0nPOlW+5vOGdQSKra96E6yv92MC1hlGv+
w36cQg7O57N7Kc8hwyOiC2yO3/5qPwKK0dbacc12zVAbNoks27nPU3xB9gphD1tQ
zWQq2HzW61afQNM16qp1wHQlb/AEIVx1tqJ53mvHfLIEnnmAVE5491rDLUBXEnSl
Q+yqANBWamzqh0aGG+esAb8mv9ziu5EmzuRMOpq+0MEX4MhoBWwTMvUXaHCaE7V2
oiSD4lycY8u3ETEB0cZerdLXqwaVhcQUylFemGd6+DxdIYvFLLEO8r8ibHjvJHjN
NG15kHJJBFbQTfh0D6G/iv2Lf4oSN+Y02lQsk2X5eIu3OAK2/ogLX5/o0T/eCVuM
WtuWEHem+5cCiVIIPKHdpG6TbnlnSPgfgkksgGzXtjCYAWpZoApdmwxOO4Shc4Hk
U8mnBxT4ctR1OdC8Cots/egobkbDatlMJyRVjPIWKchSdxWjp01A+Pa7KvYVFsq4
9fABk5PG4swAXGKKUUFgUNKSqQcheC0rH0Szr8jJdvK1b1fjtg1tX9LUaEAUmFuh
x8XVgAMXAY6KE7eZXLDFpDWmEtvlbmkpXrmRm6BV1Rr9dOhwJaJ8PuyI6gkCM27N
zoIbIjgasf8O2ZfN0X+9edZqSv1sZWgcp65st5BRCpFX9YW3L47XjT9k/Ezig/az
tXG1g9bGXMT3hdz1KrjPHb7rZmZSQ8eCGexOMbmluF38mvZKo+YCqiSNRlbVT0QD
AfrvcvWXbPrV+evolDlvLCpO7pbrTNvN0jR40jUeBDW+SGu65FAIHaU+OegIF02N
hwPCXVZUSG/vNssTnGxi/SMz732PNDTqOBAmNJTZtXgRwJThRwwt6p+05BMxWlRZ
O4ZHfDwA7l1xvg643w5Yq2ga4Yv2LDePqT9p3g6lnXj2GeGX+zhwUy3GPrYhGrdr
8vC582ADR1xJPF8sK0NliyNggkVakxW02Ofnq1Iy19OvLxe1JyyXofmvAGSHY81J
V0JImHXpi+d0Tf2pMEjBmwjwwOUX+egST/3cfvL/+Mz06z5Ld0G/dRKX0x2/PRIw
9xm6geMHJ5U3hgHAO4ftEQGxlRWpQ5A3ZYZX3ipFmTxGQewd5w1/wmwLH6eTx/p8
1UUVt9DXCNsjleS8GPsimNVtQEyXNFV3uHFGD/h3lEP1UJgEjq5yrdEFdyJ4rum5
SWxGt9zgqbb8cav6GElZ28DQ2xawt/EIXeGSw0G3GytciczbEZcu+/YTZkdi4izc
bcNOo+IQQr+biaJQ0gHX6OvLuGrD71Wmb4410xafPiZvqmWgdVN/L0qbk4GGSG/5
hyMBVI1FZ88LqhxWem5lLCc1dT0/pMhYlJnxPFQKRaSqGyXBNy1mrkfTnlO3gBPd
boo/Hg81a8NVNQQTogaQdTCAuPsu8ooaBB3nDmhEZ2fWOhAQGikQnuxDHQw8sThQ
kE4FZ8ZvVSeG/Ltu5nIWjfvjrddmsb21huVxp+v4E2Dd3Ic068wK2biGMD54HGuZ
GZBA0UG6YdQ5z3jOr/EX0U474LaQ7WKCtv3qcRItLYEg5VR7Ec4ayZGRwhcZKR7J
bXFsm0txbGH/EN3+ziLTD2+pXf4MqkM6Qnyexj8eOud/rlG/zOW4eCX2KPQ9opVS
gfmoYjNq5OBeFKYs12KyHQwd8Yv3ON1F3t2Bff35UQF0nPNlgcDUjDSMErVVGnwl
gotMgjGRh4a6R9zgtXlPxQjbUud3b2XR5Ht86idNpL7sFBCWnecPepCJ10l4NPyW
HwNEc/M26DPK+x2F9mjGevYcmvJy7CAWlLMipadJv9zoG1uIRR4V9+Db4vdzx0Y0
Rz04KKkp4dlsd6KuPJPr0EwciQlNJqifH9RJucIqOhCUHK1IjHYUiL46r/DRvIGO
Z7I/iyJhaoKmNd0+vJZKxa6/FralqAFRgOAdKEuQcO6cf3o7HaYCUQCVGEYGXbXO
HRHKBhfwfOvXGROG2paKhEB3R50kfQFEjgs0lxPWWT/jsZ8OybBOACuEAI5UR1Dh
zNoH6BghHNCSi4IjgGFlK9iGh+V3YUbfj7MeZQPmRPkMjF/YEztuLKrmIpytCwhi
M2KBnkDTFLIxo6Xe3WhDbwiu1kjm0oElCR8acAb+jKFXoMyY/haOR7gZQJT22u75
PZDg9NEg7VR0h0HiFQl43rEWIKCyOt566VvFQFlu3nH9PkbcgW27SQp12Mxo7Xl2
a9pNtdBj6a86h4ppEU2Ul9wSe3vwrGbEwBAlgDG33zIkDXCCSkdBtpuaE7qrl/Za
13jTrJaEOfJvF0499hF1rQ6W14dqpUFYdi1Yre+fIKWcUzo2ujhHmMe6QLVvGN23
HayDy3bEdpihUmXGhV6u6CIkJqYirS+vKqisjlgwghIgwyKw830PsLqr49kfPfuZ
qexJNTps5P4JB8pZ1NDy+UA+7fZ3xtPHX6HgdD5JGVoR9muqliyNPznISxxXqSQ/
jcSdjlhAOJe/uAkqApS4BX/9GQH4prS+ne9B7CLnXfhlazmaPWhuA7fwZg9kd+YL
/gIC9ubPXmjbC9Ua8zsT94NKh5FymPEsFmwzOpOE5q+cJe8L0SCXRE2S6yCLy8Bt
eXxxcIBbApEs1ltlEHILCGO9jFYhfADzOuVvlzz9q8K5lfGCKsTvIUpu4qh4hKGH
1Opz8CVYa6/88NFQavDnLvTPX/pZSRENmtFPsxSIKdd/h6p3tLro1k+3b54G7k4m
UUZQ5v/KToxbDYdU/4nE8ovYeOJlNUKIhwUUI5lJe3scG+J255Bv0BIA4dKjqHhz
1kxlLXjhpEFc5u8Z1qTn2mlga77/0p1Nj9fUnzbWo9lYDJ5g4HTTxRD4Qmj1INNw
JiTb1nYnz4sPx1C00F6wE9Gx7cFAV6wtwC3U68QffhkLigWk/QNQSq6XRN38Thh/
aFGtVgqoZf4VXJtc/fwGdf/ne6Ia1l2Jos91GtDihQ7UtV+apBXwOyIBjpqVtvlr
WiT5A2sajikhpJUQwwZsVu+00qe8GzWwbvRf0gRpwSlqamDElurWaa9OHjnfSIpK
IxRwgyJYd71orhaYBXwE7xauQnjah8/nHB9a7kk1qqLvUZv1L+RDSqR0b8fAUZtD
ogIvvxq8+q0ntSBz/c87YGpeUX4RQUkmntb6t0BHl0ggAxZ9CTW8TFxhhqIZCkup
C+IEWpwEPFqpjZfXLSzjoa9hRF0jct0SRDYsxoAgH9EuHJUeaCAWQSWNMnsKoxrv
G7au92NJfIMkh63QNjUPF55Ttn9ZWFE7ZqjLG+HsyF4YUu+usf3jwE//nkywpIVL
/Rm2XqOJwOtu+9mIjBdYBBs9zRMiASfw8UmQ9a9hiB5bSJJRCY+eyI5De5dtO/KT
fvpgj0hWDu1l5mDFZoj6FFqY2y9573eqJ/0Rm4cz/sI4pO6hnbOqnycNvdmAA/HM
E9WctNURJZiTz47YwJrvSGBNSUDoPiGVD5gtO4aOCDUCc7gqU7BJiaGjeWabbGYE
TQR6RxV/sOelBvnnty624D1CN3BEP1t01bmPIJKbo60sHHnF6nlnSpWnZx1lFY2d
ffzOiwIfy6h3R8vGd2hXi/OoQVjg5QLpburmz69oiT8YtTYxpQG+sg/WkoW12zq+
OULIsMj11L3V6yt22qf1lyiKpG8n1Vd8/61b8Res5vyzh3cRlhcoqFLaIPcPuF/N
2qLvJidzIJidV7F4u/8lhW15x7kP4mC8guAoiklWVY6leirPVmG5Xt8g/KrLXrs3
YMI26HmQtkp/aTQNJ98kICnxNjwKrEdkqUHGUDnjbC8O5+eaqZ6e6KLd33ElOzHi
dK+m6eovaHYvciYV0FayO0rgjIQ30Fzeiw6Mglli8oddfJdFjFtn/n81/ob2dc9w
u2I/EHoYWL/tnynrzyP3BXp0deaItCs2/5j1apvVLeXiK9QK4bsgavZpj5kEw++r
yZar6yrlgOO4hva/+KA/YLnQs6uChJog0q80ygatAk1O+NyMod4hBhEFbPWpktuv
qSst6JvcI/wRZWvCttIQQMTkIKzpqzwHGX3Frz79n45mVmuBEV0uwJD+oJ7DSKGS
saX247ZYM2cx78BntwwpJRe6ElbPW+WtL3Zs8+O0r6kZmqfglpkjMKY7SxOEHj/a
LGn9LViSDVIQ5DhcxbEyQXVjGg4d/+YOMgOpLXo8aSyHLi8VXmGbjnbTIExP7C8b
25NYcJhgdzDM3P3D8IBm0gArERPhkJIaRH5GN80fi7Yuzm9XkoQGDoPMqCBg0gSF
FHMOqJ4qHmLsyWBGOkMG09OS0hz13cXXDlDksZS8fGJ0v9ixlzYCvalMRB+j3fUk
JFp8gGrrFNXyuH1mBJjzKNiRcvFJjSr3xPsF3pUil3NAU0xo06E9cRZ/h9jg/pQp
RD+lm8c9sjlh6NhjF7e7LQ6fo+4IRxgZp6nGi+DM/7/loJ/omB2YYohTcJDhfR2D
/HhRUh+7tMVuz3SLosmlO4TLfVll+naoxcmixBJ67AHO8gIGrz4WGHN4oXn2v/Tw
texY0WkEPc/B/JOu/mUXfYAniaqxIV1TkDnM4w65BvTlaeCKEhp1RA9NKz28l/qx
BIHM3TOouLXZyBoFWuKdLZM1RjeVhaUxZFryLfeQLx8fd6ozzu/yM/Wznorrz2JF
AyRBTTnDiyOJCTJ8Hu/TEz7HZqKTOLmSbEYQIsTzStlP2I+zGPlKMn8yu7WgKmx+
jnWK5oR8w8IUBryryJ68adWxAqr2/LxVdyVXLTnW6JDucst8r5mt2Zmj1FUU5T64
TGx71ZQp3drQia86Wr1dL6r0FQrW4HvUKOQH+NFwAxqAE2DTSVWAwtAM9U/vWQAw
hCipia3F6d6oidAa1Fn5f0wk924nk1OrIZUQiAaVwvzvePsMxZr1F+oCipBfrsS8
e6qV9gOsozjDvI2/8gMHIO+jygCs1x9wVQ24+xwiRQeJlIiW0L4lNiapGZykNLap
GIfZpgFLRdkRvR8dFdOk7rAGPUagCZwZz5GLCbjvJlyxAselb4IeeinGWQYNT3FO
vj5R2KyfHmI8WrVywOfb9pFWI+4BFPfJ9/SyqtGw3beTU3j8L7d5uFJNJ+AC3tjR
bFYcZj0Asp+wE/hwr+LIvPTD0pIcOtKq8RiDNFOIMs60OQKFBP6N3aHmMbC5Aud/
Lsg13qTbCcB7b4TavU+49BZ3C/dfmw5Ud3KXdznH0hsf+L3H1iUBAft1BbESpokv
QB/GP5eAWi5jV7k4dr1AG9qXJlPwYwr0wHjRhjO6Lib/W0UxG/qibKevomZS7bXN
Zb8NpkF5x6VozrBUQiaDZfEhQ/Unc03EkIdo2grM/fb38zNwz28De2bCCfnsEvks
/u1F7wqZSiPjfMzTBNPG3LJGwlE1B7AvUQRL/YswyQgOVklma2U3xlZjcM4f958K
4N2/3OtxIl0ByRwIw3hTKGP/cIRR73SktH5dRO3ULjo40dnz7l3CY4Fs6R9LkXsb
xX18Ilyq6ip0zYRM/SSj7oCP8Z5rHk7xc7TA+YgActBwGAklCmtOwpkm9iQUtcr+
TfBUsrwgIStFULYtvyWq4sriqGPm2vHtN0B6dqPWlCNjc/MDsiRoWu6gwWgEzsqG
Jp7xdMpUq3IbcyzeCVA1kH0hYiV1Evhphz+UFjCxGv6SGqohNXwE2/6wZDczDv62
uBM684W21UxQ8zYiSdIshTZXtcaQZWda8zKM05n45NyejEarTFmaqkg852938srg
MhCgvA8vkauktcWZ1+h/c3BqjuGp0na3txjtAWxiezXyLyCE/d/BPHhua25iDgja
C1mnKqSC2NJ5W6NGIcVNHAgAhK1I9DiyNBXynRHlAu4+qY9B30dcwea6F/WDZFOn
hH/owlwLOlbTm5jP8hFrAwARNL1/zs1P2v/l+my+2fFk2hgBPegjHMXWIfYYmsWZ
X3W0qlqBcik44wHhABXYw+19badhArz6Gd0LK1D8SfAde3VFyz7UKuICC6xbiGpR
ycHcYpSgrxJC7J7WmuuSvaH/dCg+BviVJwGL5tLGpKfOGClNTfymQjpiF1qMGV8u
Fo5ckeQQLnr7tsBqGpKGUM4ugYZmicEP4pf37el3d9/iN7mb3A1sPGyEIeuqYsSu
af9/5Mo4XrfCTZFlm3NTdWYpvBLra22YlRDABwz4k7978TPy66NPamd0g3UTOTew
s/BtLmssXuXQWlxgT2erLIs+qqkGyWQDm0Nq4/szlAlGd13hQJETEef9KM2q365g
8/iYB99tLZooARr5P9PNvHaWPuveAR8zsqs8HZoUI3z5uFC4JPTPy6w6uMOTbid3
Syn13jDv4yKLzl7YutGN061uFWA8c7gC1gyVfI+4WgU+7BS6+3pLvjIGIUxulwOd
go3TocxCLIdWuT8VlCVM/XeAxO/1v5fRjChMjKPa1w0g1Ki32Qp3Ydlco3rEE/vb
mj7QdKJTKl7aFry1Vnur6AzyDP5DBy0MZfWNiBe30ALX6qAE+m6eUXQ8GAlaaEjt
4bJlzIcN6dwxjJBNHQOfVoAwhhqXuqfaKJ7dlj3horg=
`protect END_PROTECTED
