`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94aMWaZO1YbE+HMjnwMM0yNKFF5bkmcUi6nepXFYEriR7aFwRIn61lvXzbha8h3k
KLmmZdEpy0d5No9zuy+4e1FkatHJOjmNPAl+skUueFYt6qBZubkHZMW2g5/JyuCN
cFEUPh/UP+VD2Ehjc3hNogyL0e3HAK+F/u8GOdIgToEoLcW2d1PJMcYVYhHb1bCm
kRsUWkKnumUvQ8nWTw7aMGrTZ2+CyzQWbvsGmxUM0ky3ql7+TaXt5nchR2acBhVq
6SdjxZSdGSQ5F49NdTidGWnrlow9PHxHSQ6yHbtKLJrLxim12uIDZE2FDhGlV9A6
n+iciLSoKAvcvv/5cr2zSsF9YJ/xrYrrjHSyRVMMkk9v492XsjLA1elvmEsVpr+W
a4vzc4CMAkQP5xwGanPn4QBR2bZ4XtiqxzEFyDGWZFVAyNIrGTqABZNi2PE0CYCB
C5YaIZr8ew32f7sPOY9hRGoUGKAQrWZdYqoQxsg/syOyxIwMFyFhYbcpiZVfjvr+
S1aqRDv5vk7YYbb7H5rFzbG+cqioS+yosru2S6eNmTUWmChRlvJ0n1J47ynyEdGe
xW+48z7rmLyObggd/8oTryqzZ3vUPDkV7hBskq/tP1U=
`protect END_PROTECTED
