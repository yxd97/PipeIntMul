`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J/+S7mNzxSTeVyBdBaWNkoBGoXNGr5Ct4i4vUNFR9eZuyko3IsHXAl2ZEDTOvc3A
R3tLKfYOS37WYEC/2mBXAlWeg35WYyWpG68FwdFF6oAmhuKdP9Crjtraxf8oWYwT
lrVSz1jzKM6QC4Xqvk3mzXDmwrBJWOXg1e/bMkPA2qI8gHMwCe0FEQIr0UoU9mmf
Q1YFgScE1h6TRRkzQdEc3U3DUNnAxiAKQEFWiYgpQarGMMjpkEPlINB0ngOfOdEt
b2k/7AjqRV+3JxqQPCGHrYqtdvPHqeiLqAarxLTnneE3TwACzCYXPc2GhkFoI+Da
iwLmWpn5OuY6Wm57Od0saTpBR2d2La0t/aPHjRq9P8zPpH2mA0eIka7JhJgvORNW
oorHrYYJHcOmhmW0d2bv5IRSqvfdZmOW9M39aWRfZGTFMljmcLquft88aFbGQ/xk
GVsAK370pt3UpwrsqacM8bFWnAJEcLRiTOPAOzS/0GJ0pQAyTrAH9QgSr1h0ZxAW
gG3vjXDCi8WTVKE0PQAbOT6KhZ/qdYAoqlAhul1jZlG/1PQ4a63mAwjSY6Eg9JHy
`protect END_PROTECTED
