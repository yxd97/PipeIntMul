`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYSjbpOH1cVE1pcbN8t7IKlWkuGVDZllwNj11KoOFdluAGR0vJBkneOdjHIQQHhg
o+E1ZU/GR5mRC8eqhLjIq2Ch5qF9qp9EJa7h9BWIzAQD43xjxN1Pq+bMTfAcXOnH
WTXHKQ1eWEDkIrjGbb6KyUMuwEbN5C690zONR6XkuzfXkGOp0cLnwFFcLpih0sKv
Ew4btbNIFB0SU59+TvusjFzOrTLGiQRw2JRQaixn46Jelns0319LHY4Qdg7luQrt
CbqULRczd6GPgA/06Dek/JWvNnE6Qqrnp3T14Lv6iZ3wqeckaGX5G+rjHgWT9A98
aA73juNZm15p1MG++dlexV9ib1WVJbTWi3cCu6hMOQkZQOxaP/eZk9l3OKnDikHb
jE+QFbBAVELOEKiq/Uu8bS9hzE0Zag/Ia7k0GpiMOYn3SE3LBmhtY/sJCiCydcv7
4jnoAw/HhYeGoiERBP1CNHn5duu+81Aidnc2yEUU8MCf+XcleTTU+AQdDnmXOy7h
KnG+CIaIcC20X6HDj2Q1YYbtSZnqhoAhhvNBTFERoKoxDgWoLDVBqIRm6Wb/vCZT
Uy+XNSV2UWPxYsidLf1c/WG7rRJyHUlAatEZ4ESqDbhO030AdEek0cl4/DM8k2wZ
VWTTIuqQ1reauVgQbV3pLElC6zBweDkyUKC2S1XVrCIwLVPEX0iSY0Dp+fxwnxNa
l5/LEuKJq9EiM7nMxUdH8sdHVCr0fnV0GadZxSKrFqJ3Qg/a2UhqAUdCf7NU7998
YuD1yB2vxEdUiUNjKYDzHeeYaqEa48cxl1AHNDBbQm6a+K6hgiepRJQNZTBOyJ7L
ob/+JCM9FHbfExIwJ71M7iMhxwPnS8wyeC0L/WbJuh/mDQsCmoxxF5+y4zR2XNS7
cQ7r/EAQS12kyoRoj2bot7deocARYFxQBC9ZRHIthN+UBc4P8+UPT9Tz811smLJz
eqxTcSZxWeZssuRRurX2e1cYniINErfbTvWtWEslvXmx3dsFjHEClD4Hq4pUMumz
VPPaG/vbn+jtKH1DtQfJw+UMtVJ5m/tXca1LJflkyf3NUGEqees3KwsuBcFNNLb1
2WrbRl+DzWugyuozo1CNfyUbawlpWSct4/v88iQnEOam2pFCPp2aeO3d9h5wCGSt
EmncTa7vx+nDRNfJwoNbdtHNbacke6Sp9pvX4JeLHPeudDwb7CNdnr54Cajk0kYT
ykXbO26CFcFiK7oPxRIQnJejJDJSrmSELe8b5zygUoWNfUhxKV3I5WNffFuHndQr
PWd5+BKL/b90OP1ovkf1hqZ61I0RyCSaaKgE9Gm5vYuj4ikpdfiMQqes6R62Cgtn
gbnZBODwRhSARvocusgKS7PdpE6wQ/idz8rGkVTw0E2VyM58YkPko1eKqJ256/bK
2LPgKzFw5IiRemMjwN17bVOttRu9hYZJT0vnJmC/EliWTpUyYAY0Ik3h6pM7YLcH
dJX3eWl8wpyGqIQuGcCqLoi6I5Nlq4LEGVnqvFhype7UhdlkPaRQ4GNVgyWYgeHS
9qlhct+27zJaXax43zsBHvBJjl+MUgv4ipzx6ygu8GYxSt3OyWhFuniMdrECe92U
`protect END_PROTECTED
