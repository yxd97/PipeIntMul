`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tCVBKjiVjeytiswuEsIleXGIeA6WS57KFy/ufpme1IWXOajNiuFWdYiwUmvcPZk
iWHoY/nYLR3z3CExdb8nGHnIMNVoT9af4oAjiikfoNJfVg/FGy0vQkn4Oh5uPqXu
CYWVm4xenTKFKxHRqVk/oEcHHb1rB4Jm2KAZ53FW68fIfMCpnqOOekVFC0Vjc1Bh
wZ1Mh4bF+bd5goam+kyjInsmm+i+LVmFsNxUTLY7aF/s4Ilj0pJ9CQCiIN2O1pcj
65c0eRBFHBiu+dUbwgUnNTw7TajgUT9SS81H0+mxie+JaSAGgAigG7O4mxZSltKv
Td7e8UJBgwp7J2raaoyFazBKS9Qcear56bVvIyWXlftt1c5nAC0z8gKuPS95AQg/
MzS5T2DIjrsm20QipLrOEGeNnJpeIE8LmSRF8dgO+4J3cqHu/AMxDgcE+tTZpR10
Qxb/QICw2B18WunsLbrJL9zqH9I5gls0yQsRXAYfHLw=
`protect END_PROTECTED
