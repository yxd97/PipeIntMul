`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RQRzuptb9OYiDqZhfXR8TTBRNAU9tU22kJh8zHKjLCycYNwh3rDdlLOIcwMn0puf
OKILjsmrmqrBq+9MxCHQ7rIZB4n3vMdrP9VmM2OzyvNfx+eeTtGV81orTde6M9+I
baULxAvfK1ClONipJ5CDERlprYR6oEwo0i6H23vwA7DhPo8TgFpl3mzFYpscoUjI
V6J37uE9GEUgisyEIxqsk5N+zhHGq1KoOkoc2tRZY/lUn7zxwt0nAdUf4pq/HTdl
dGYsDqRp8RtrbMshIQHWDe4wssnyFNTTh40ihbp1hlawy3n3rnlSdYy4OeuSW08Q
z5Y3iuCZm+9vuKJHVgFgtXBa/fEGbvVPLemD3kxFMg6VYk8RpUpWhD43SG4LXNsJ
wLOb8oVPciXLO2fxu8BxbVArPtJDrsrpRGhplysvLGykxuaQkRFyw1jLP1s687nc
tEJAydOLlY4VAYmL1vzpF45hdAiAqJoCaOHbPVYA7789kJYjaE2tDiFxdsKnXaIj
68qGUuqjZYdseMxJwqEBIHge4oMVud0U3E2YgvbX9ilwnQApETrFhF47LkBotWse
FOMslwloJMV7MtjvxmUhYA==
`protect END_PROTECTED
