`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Ns4zNr1G2hP025tYoGQfE85DnebtdTt/jKv7/KeTLyRTuQ8V9C8bhZK8iJQI1ap
oJ2g2TuKXh34IPleiBa28oLRC2qrtqcskETzfZye+cTHL5BOxMLlaqvrYFjx+7tY
ZEi+EUY0YBjg6d177oJtGAnFxRaFJXaSTWwKc3k9tQA3MlQOLSAni7dtB7zfY6Ea
NuKEtQ+ob6I22OEl8/tqvJ20WHkZabs1qoPp1SMsNAL25SiZmGcekRw6r8vW5K9l
pOCD7CEkKuy/6UMEi162OQLZF1AlLCh2vHPdTBvQxvmz1PCidvxBcXqPBGIub8Jt
LIHnflefNRwJ2r0zm5feNrH2Ly11Hz4XaIcji6hyObDLgCXsnzHtghYPQ/dBXzkv
aNYkOBa4xGZS1h9VKEA9c9Sco1ZW9WOzVj1Ui4TpZlCYTtuupKt2LATGyBqS5ujb
vgiEOJVBhx7kXflHzMroU1rkBltxFgAaaqyKqrn1/J2ypgvm4JonvjMmhGO4Q3OC
5YR+YxqpMOin952eVaLRlg==
`protect END_PROTECTED
