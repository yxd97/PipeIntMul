`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgBEQ0lTyJj8eW64d+0UNChVd1aDkat1sm4R9nfjIMxx1qPAXeagYWT6+ha4Yvko
AwCwP5yR1VQbcKaXB8g+24iuy+zauLPHS1DWwgNc2kW4F3VIcWPJNyXfOC1uk75A
LXTRT8o9jJBPjJ5jYJZW11pLhsi/bl9gco/UttbbVj+cho9qhAUW+qWBxxPObeES
I/ph1DqE7VzBWQ1q3ae9UggLLF7EWg+ctYndOImvGcbm/xBdKb6h8aMm6kLTdYKr
6y6c5c2na+Diuf5INo1s6NankaihG47++mrh03JlXvdAJ0QpQmyvw+0gpV+LTLVN
QDSBCycR/Mlh/ZNJRLVSQDGeGOvUJk49Pj+jrct97M/cApaujVQDbBRu92YQIRl5
GhhD1/QKgdQKrhqWowUfajatY5UGVvHtey7Q/jy0ouNtXPW/RhzmYxYK/uWpDco2
GpXionYScMIGatIL6FAkw/iduAJXrKkR9I6MEiDCjdfY/yjxKsZIrvWVm9dI12cP
hafpvUeyeSDlI/8dJfmh13aPKO/9tUz4cUGEi161zDJ94Tlwzs8JWver9ZFIPXgP
JUVQj9XUL2c4cCcGo2ALBnOM6P3mtldbMDTGoK9hLYnsY/vdBOyzA3Sw5rY7hdw4
lzvi3lBn2/AvSwxL3kSfSmWvV7UL/tu5tcCqJpaRAgOa7X7dhBcPBZBupi1AZeOR
VfolCUCoEbr1yjQ8RYXhv0g42y0XLeoyKwobHPCmx/icGoABq7PhxGVUdfigrC3C
KjT0eQw3CnLBeorsP8eeg+Gngtn8iEPuO0jtFSHqQqB3aFONINcGlADrgUGEhxV/
37hx13EQCEwXQFukvEwEEf4x3Re9BPejzZ/8poBtFO5LLFsKKvUcL94X5njRS3BI
MYNw9zraKKDEKexHN5zQB/D3ErVaC+g3vCPBMGIzZFkHZkNaciH7uyfDnbpwW1PZ
QtIMW/77bXR0j+3zk00wXe1iLjnv8CYB++a20YmOHhQP2laIxL2MH0N6ckkiGxFM
OvVfk9obTItJh7VYS/XTLUwHfBaYZU43ui7EdXBhSjq6HjUx/G9U9lpPNxisYaCX
8JBetyft+hRoBAjtfOaJZnildqpm6K3WqvbmWojasuv6FeURjz+WYKT5WH6TQEqr
mHCZXnjZJ/iPa+tCsD8Q5xvVVCxXRy6PX6pQ34OOF14=
`protect END_PROTECTED
