`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJVeuytXQwFsi3GgkRTIoNqnh9eftRg+smqpjAq+rsCUUds/MBuEAsAxPSIc0KjB
LsbSLz1FI74tS6AXufsn/jgeBuIlTs2ckk4VStrnXZVJc4Oz23om8nVyLiMIlNlX
bHycXqghSYXLHdmFgEjbc6EHS9XYaaVb6YFjfiNCvBUJny5juvzW9LK/TlQWS9yW
3PUAdHbfowd9Id7HlwFC8xwiqUiqMAIxV0zVut+TnQc/B9GH/eRy0UlA7YzNupaE
izIdrVyksh56r30ePiP6P0u9cmy8meRirXthfn+Ov14D8P7TZgaJESj/E8idp6MR
a3F39NXIc/6Tv02C1SAv7A==
`protect END_PROTECTED
