`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kntpnKjzg0Pvzkpr0nJ6uMwVbOwQsrFk5ov/s8nfsHhDnuTKrDYCUYOch5bwN9y1
sji1Ydx/Y0YjA3Ig0Vl28IBm4raDP3uvMuqPhf4Nhl/LwtsJlcQkxxy3DQkPcihY
L7KHq/EP7dNOAQQKy3/TJz0Ar3mawGId2RkEdlMTs6pq55SyS0YEqzPyUVHCVKXM
caEAkuetr4Uz80ga6Xw8eHgKHRJ/WNuUZG3Y1JhsVqlX6Ba6+mvpQL4DvghPXHZG
/0VqBFFNpNCrXnnQU93yFR/NRSY4T6mQwi8mYnQiRLLlQjBAQL2brIIByf15ljF+
5c+qHkouh9SOtoD3CHxP3Ues9KVwAZ2mhqCCmb2V0TkL8wTa9LVmUohfPzbneDQu
pgAo3Q8OnkyyI5xwSZE8fgQjYg1gnv0CYQ9jB8uVP6yX359DEpEFKFK0H7s+M5xN
OgY0ml52k8bIodXAFkbUogFxw08WAI8Gb6M3ZxDM1X1X0ZECr4uf7COto6ZXJXk8
SeugIa4LyjZQUoFi0tmbfZCjbole/6NIW+MXwOOxkcu4snnsukFf5ayplYt88OME
yQwTPu8tgRGIB1zQaJsBhdX5BfVwKCVvV13Gplg9uazPRS2WlTv8/sZbLaXvIkMa
mF/mrfKRfeQpk9KRfO7Mn0PQUQg+OA2ueZJ4b2QX54/saFRvpZiHmcWilKJbSDru
`protect END_PROTECTED
