`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXpEh9LUV53A5l+lKjNqB+EoWkzxx/oKSgiOBd6i70CGeR1zUpKa9WPSXQFAgykg
rLBSR56Jct9xRiFgQEMKzSfFQOpt3yZaq26hhI274B3vzF5ZswbTaIBL7dztkp1E
9E6iDlYShg3W0VWpdyZBk39Bo5Q2sxPBmzP/A8xDqhNsJ3klEwC3ANT9TYe7589U
zGAJakLkpYoU+utSCuYat7dL5LQUuj5mUx7TtS25gB9Xm1x1K8wdDzdM8GHOAgQg
dZiifAvY0MY5TUjiU407EeF9sXtJE0IRPujAawT9bbwuh3zWTstkqd8ojKnXMLV1
+UV7ZD1E+kAHD11/le9RKhBixC29h8cotznSra6nIYTqespvB+NY6WOGbznLGSJ7
9UgUmAiTPBOCzxGtRk1JhY09qxpkVk0gCSEsolecdJT4n216Um/SBc8CoZsp6EVf
BdrqanwtMnK6BDhfSdxpJoLn0pFuICubT5Mbt2zf5cZrEswKYXpW2R09AG5EvA6q
TLS9eQS8ZEUoiUyJ2gl4Vodxj78uRbDUfKsdPVqY6UsNrleEIBk+I68gkuXkif7M
`protect END_PROTECTED
