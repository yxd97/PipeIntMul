`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MtYMVZANpqtO7uU3/58be0izZfAjtbHj98HGJRgXGnx+Y7gFXMbhfDoufWtiXtbs
y1Ko6mb5BCfqDA3eDtpRj7d6Txkw0gG8f1GU0frHazprTM1hcaNwPQJvMp7dxy/a
QLOZm9kwoTwuRkBXhXbOJTR8ORNzVCx+Csyhzb7puUAy4lwRnYgP9pP8Sb3Veqza
mFJIsbPgo74GGk0vOA5b3QyBpHqEREx0i1aXejm/TCvjvmIodUVkw+UeOg9WUx1E
PZSrh3kz1Yxvo4DjJhAgjeAcETBSxGHcSoXkQkSUZH/9V81GhdPc15MrFNwCnB+L
TKDq5jZeCJC1SrJp6zvfDwWxjp19lYzBJag96CScUa5Qo5x6V8tHBfXJSyYpFjXW
L8/URkjTbwYsbdc2EGrqEMpK3TYd+KsOZJk3GpiMYReQjtyJPJYbvKC1BBgqTfvT
uCtKgiY1OohljgEJUoQJ6ZLqMgI/fHEk7R8aAjnIQeuokq9Y1PtafsmlworpDVG7
LSM8Uqzqsm9atfPy4d3qS4h9uqW7IcbEXfwzgCfRk9v2+8zKy9gecgGSX+P+9HgY
Upv95sxDIO0BR5YWxVPvwZbSfg3g8qrh7My1I669dXikge1AiCs2BQYWk5+w+V4G
Eqq0bdsxb1SoDEasNtueIXt7k8Swv1Id4mpR1lPq4lBHQsLvpGnRlCAizuTkf4sF
8X+I9C7e+29RF08Mz31JnMoZzDevLurpLcwGlRDJzEPAWXxnV/+fmJVY6DbDw03d
Dljv/pz+GxH3L5d1dCHEIo/8ifBSYVxXLXsQeLScOtc=
`protect END_PROTECTED
