`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHnfOhwLjqhjlbbdAyLdISXXLUXWsexv5tZDzb+PHhn75CgEx/BPqIJV2U9mcOkE
ToRQWNxoLVD4zs9Zc7Wc04oGUhrlhfl1lEJeFYkG9Fw9SH8XPKJUQ3xRz9k2uhGD
9F0MLEpq+Htj3G3Bsd/RdgwczwxMDCcSu+fnSzjtU/H7Au3uLtiQ/zFymMGElak1
3z334scUvDTO10TywSt7bvw368z8N02ksQlL7XjF2cEWG6VQfmQEXm44EEfFYXkK
fg105BCFnrwXXhKZVhgQCoDgeeKaha1jaXXyUDnBpx0k6FxAj7IdOrEdBmxN7WPx
+DoSo2TrJW9GLKmQskzno/Us73WdssPcygqu3EsL0Mb3fYY/nPQgOpMfjb89b1xJ
mtKh7EHBzI07h3HlyUGp/CPVaRN/tbgjL1aYyy5sFylNPBfzXHRmgVCZLMObV24V
6v9jcYdAPCHNTqKAu20i8693pQ35u0I1d9i/tEV0fLiyBGboct2m5c+u/OHCRlo0
PBoftq43A+GoUriNoa68k/fqACtpDPYhcijdMHDzNWWgoKndWXK0C3/30RiUIdUJ
ZnXJS81fr3GY9T3OGgvVUpeoufZHk6vM8T+da667Gix0U8XzSVLc0Dkzxvhggenl
48fzovD2cDYm9hm6smarBc3Kljf6lrmk34Fbm6oQhimWCzVrzXNMGW5XZgbvZkFe
3kS92U/zrte5yCrvJOPbmIWfI/ItJaMTUvnSJdfVy1933+zIE3RbBYHFJrSnVu0u
rXUk9t9yQxTx1+J/hgv0z3nrp+rXGhwa5msbBrt8v2vUDv8qyNLvhNdpQDi3wbjf
k3U9FS56gni4luI+fUXLUeNt2QuYZNooMm/msGLSSLgfppQvsx35GO04fQb4r7KY
Nk5lQ5gk9fE6Cbme5bGZZn6HEwyzrhbK0k7hsst4VCpim67nWXyp2eOsXfh3rEh/
sbat6TF3vsGzP1W+KIrbY/9bbXWF0t8t/8YN4ShjB/j3MiJxsL4h73RR++VRBPKo
C0e6qD277ZZoua2sm4iMiwYcqx0TZF6IfVAKKC3qQlwg9h8O9jlJFJ+DfaULIkNf
RrLi8569iaQ2QasQWSXMIPVwIsa4H27NiKDmfFkIaCM4PZgTAB1grStYAdSszXu4
sbnV5uZJawJqduKNY9GMjYzVMaibqeXXa4L0XLojoeFnJTAWo7LEMG/SqZrcovha
vBeVGwwxjULxEOGad7eUkhZPkixfXMWATaVjIAaHAggUJx4oKQMKlfwOV4ocYFWZ
21TB5myS+0AWntqsaRl8MRCBKSbZxxgeubd/qYthqn0OfkVdUwU5v+SOH6mwW60Q
TaDhjY8v3HfPiIRXObR+vdo2uAiYgTRAQaXVJIRI3nFIvKwtp+cffWEGQg+ekjBi
yG8ss48B12iH3tlDEi/mRSLGTuW6BHB5dqABm+huIbY4uiJn7Iuv7watH0qrABGr
NE7rzrVm+YCXAmID/CX6Fxp2NNP+9nW6sNIT5Z4q6BYA38cteAB606zqZQTl9mHe
ooC3Z5+Fy8a4p+F6qooxVuEUyHlmBvasM0eTdHZH6/9e8OvVOtscmGe1p0bOaplH
wrLzBh2x/XTSlcSLqUY+2qPn3nZPVU8rMi2cF5emciHNocJfK8NijlQ4SCsnyal8
4ATLZKDiN/zLpYUZH1XAxbwKmSR3Pz7veh0+tUNbQJt9QdiqV/8eyaclZXnGQ7Ch
oIA9j6+62mmPqi30zWrtSwEWcq15DFKALsO7OnMHWanMCM8JhQfro1DtaoBWyujg
oeufkAXA054Ziom2oLi93dujMMRTsp9s06Xcv5U13rKgaLQu+mN7yyI0zkHJvoFh
y/UH/IOnw+pZXxs7MbDelvzi6hBrrxLbz+B7n+bEbxDLpK7Ao8tE8enM19WJzWkF
l5/L2wV75SdSRd9C+ZKyLdEbUyDXNAbs2NaUPrB8Ef6TlHfKtWpv3UL52NYQUxxI
DevwQFC9OgMr5HIFunn0YaitEii7rSqzXVTGxQOekwNRgfxQKMpJG3xG/n2Ygi+s
PaSS2R9X/cc3rnmobQL+NHsdDQ6g9dstWzU3TdFs1rfLygA368wUfpRyxnwkYATZ
5MCqvK2fWMAceDBq4tPwYY4nXvO/GkZZS7p1QDKxf2Ufhtn2Bz1hig1/H07qKWzW
crtZ3aiaUo7c7hRQZ32srXi+p/18jeIRYzu+VtvZUu/+w53uAN1bo1jpmBydfy2e
nJLguvIwiILjXhnzVQACo0TKeAf4ybIDcTlpPCe14B8JZcT6iYo2EXJR81V9iIvz
Z1ersRr8NqDcFLeNKOC/+EzHkrWv73EqkC31zeHxEQD/sKZzuH95/Y9BOSUPPBOD
JaNlYPMwUltNeS86FCjW8hYYd+kkjqIee4pDlC51XZbstfn17rqCWoocAaEquOCO
mjGxZoGTqiQ5I6Ey11klc4tQocOB50fYa7gUcTMivLA8gp5Rkoe7DXAhDfbRLSVy
OyKCDBn2X4jrBVpeI28s5wp2hLyQuiK5LPE1wZqjPgesy0GszvCObn/zOct9HLRP
x85J1HYAntONCdQJZY8P0TmQFVYYASyX/ghqQWtwSKeSd5oVL3PTfQap685hGFqs
wRWXvCV7LzD5/0dwyX5yAzy5JGfQNcTk4RrZSVTMt5r6lWr8mDz2XJORKCdd5lpb
ms5Udvc4nW65jV5FEo7/3UiKp7DrtIdaJ6V0v8gtixtoqKlWPdPI8p9L8sdhm3xa
mS+BlPINlE7sQWOVHaeXOh8DbYWPjnrHIfv9D95hNaC4HUFM0dFinIpkrkkJ17Rr
twLYFBUzSJX4BXM0tFvWkw5uENG8FZYR6eMzcctAUZiDRHkIs8X/wM9IUztpJRth
q1Na0tbDcmNE/wGtvIdXxf0DfeTjndDS23cHFkv5+MIOSYQ9UHeNjB85tmUGwL/1
6HMHD6JxXy1o2FShLZJ7sg8aVF/pGK7ixVyu6MJf9Q9bb+SHVBahzlXj8Ibx+JVx
NLy8xglcYSl+fef4A+75UzgxirhhEeoNb86m5bo3lE782xwn/+WhRdU5MtE419tu
IxBf0qYiSALv4LUcjOXkhbMuDpn3ijsIa5OTF6+MUvQskYwbag2W4PyVpWrCBOBv
BPmVWkUkOozHytmi8l0Cmj30WarAAJ1NUlmO1nYkYdP6C2cr/wSTzydOECA98jvT
qbxUSEBU7utQ3EE8Q3vJDZ9loA+IOo6Dph0bLeibAwX+umukua3el0Nx2YgePsLp
7kvU0lvT+gQGYMhINxXZN1+qHg4H4xluuQXx9AOcv5BIpFUdlz8IGHWBczkZmqzo
aaolF5WK7xqGaMTmqZEErc3r8BWM9zexM3MgvCZvbIGkllAp39jKGqq/i5Mpilfh
ad4BAzazHRQMtjM4eluqOkRpgN31/Vdkmd61CmfJPwcr7UCPgaQRiACIfDz3gq3G
spDhiu4tSWqprdej4zLnz115Knr+c7FusZAVP9ngNHxsG2PKdezo7oBMByLJNseW
QWkE+aEI89P9ij0C1zCi8TqBi1cbd68j7uH1z6h3K10eVtneZB3HTSn3JClne87O
bFtj1GDTGZZt5O4Mdo3HHpmXXFqGsa7UPCVOV4HVfX7iEb2Wlxr+kwoRTxQaC2p9
tU69VfCPOL+r+iwH+EPfLDb3TvSUSpc1iAYhTI2X4d3rIw16IYG0z2gI86GG5z1e
7bltHj2OrNzCeH2iJ56+3uNKdxmk4MDwKpdjNM8nVbJkH2VQWvIE4gcmgT+g4bCj
eZ2g7Pz7yNg0zXv8O76bQ0w/Z77oVWaEgg3m2BmTQZH3/uNm8TmG3I/NMzamR3SW
VSprMR6zeZj9YKhvPJJafZgmTmb735iD+5qPV4D8Zrmo8OZhF5WCJ9ga0CGVArCd
VWROXMHaUi+5Yaos/6XFJkrZWlApBSSrQwlMYD2M3MH+Ynd0piD+/9QpFYaFYv6c
GmImQk+f27c3etl+dx4s1aUomYz+D5qQR0IIiGINJDezGVItmW3aseJTNG6lbEnY
VDBRaKSRfiaGGORVf2fPmEHgYJI8KHl2ST+AA07v+7Z6ukKbgKDSovkDefhm49d2
1iKmqtdn0pG33prKS0Q9xW2zcFj3FcXRTOkV6OstfxfAvH7yLI32bl78t+1/8Itq
+nUQOHjIOuvLuQc4u3BiNEFoZamxmCjT78GtTMqK79O7yfZSglYfF5/yETjdCJVJ
ICNQvPRgWxY18VOrmtqUDvpehVR8IqDt0yuhZ1zwzp6jQDsBOn6EdSNOUfODQMKv
ZlhLJ3ZlW6mUpq1sWjjzXWlUKLV4VxquSnc+erVkrBsNiWT0iVviP19H58UgwGkZ
BCvgwqbEAW9wqJkuF7BYpZxqw0QoN6Ob1tZtGXzSKK0UW103RWm5rnPcmZHli4fn
hjm3QzcCdQLKMBsQkG4eNbC2DxVtiJBYo1Vizj+WtRP4BV7taXHbEDKbKOJxExYB
/dojBMOMZlj2bvFBj3BMc6KJTC49ZsFNUFWIg7078naM9zHKDopZ4c1J+Z4INwS5
igIsE5d0G9q0MRjLiGUUEw6CP7x7FmX2r65nrAxqQYeDskLE4JLdl0okFAMMJ+PO
GQskEkXsFofefUHM78NBpLR3B69I10LaaZtwX0QG9cELvJxPnWPV1PW/h/8KWL7y
jNvGLY+0ez8cJSjfsIvClKaRxx88f094evZeWlvdskX1kN1WINLY/h0DRtOanhtx
ljp8IEr1/EyRVRj1L77rl2z3w2wdR4t9/qgxsKAe/mW8h2biUL3BiALbJexoU0P0
rqqQ5wB/KkBabXH2VArz8+25sf6DswdDKMCv5uRTu34Xxr7PBjvae9loxIhEYz3D
oKJqnLuWLx+GEuOoKURw8u6oLFN4NDQwUU8eumkAJUkSrWiNzZPX2KXx7mqN20JS
R9IWXgbsqWbLvkg2XBD2DY7dge4geM19JbOvX+vI7xkz+yVY2RE9mkxryOyrAiU6
1zNhzmV8SW2Xwk9LeDpNo1/xFdjzVnaaJBqRd/LFJtf2BlU45sbKLR0mfkbMUT5g
Ww+9nIPN8RXPFwq4WDp4pZSPvHzWXJYslxBN1x0nclRTQ2SZpDxDefg+Iob9HEgx
e+q35/7uvwhDZHRzyVzLvS3680agyRrlDRYlmVhTDcWz5mOXx6EQh9LNVu5Afm4s
wbBe55gWIgJnYpCPinkoZ9liQhISSIjwHm6cPoyCJLYcyokkRs4+adQpy0H3g9Rl
vXBz7kxDOlAQ369jDhRZ9w8pRg/wykS6KAoMFiraW2MgjNgjBZ4FWSKsAfzRGnii
weHfCQCZpwQ1rSp2fDfNgNvlNeKI6gmGVdwY1ioETa/SR+d3J8QAol3Zgdgn6ro9
xYp5B+87lOOsgX2KN7dinze5d3sk4h6ZzwA17NyyZ73zcjIsYoAoaccTolnRal3o
4FJV21J1eIfGLvo63X8XBHEhlcanq47pasapBumOUC+sMkMOd5McRvXmFB4+drS7
cN5zxhHFCxjqwhfpporEu7oC7hUxIsyRVgdcWQYgNGMcA6WP8HUXoyuORKmNkfS4
Fnl7ROXJFV24dFkkJVO+45dImpXZju95+UH2iy3QVX6urEXacN3o8UtdLT9QTMm0
hlVdihdOChMXZBfPUN9JcAz6oCxcV+YzKI3+Y0cV81FdpWtDsYi8rDA+oXLQ9Cvr
KIA7GF7CX7itG7l+r8H3NtOAFxM1JTrBR+m6V53DbDjXPRERFiN4YaVO+uuoJPWx
r2EqTGcYxdNWoXJ8i4JmMfUX29tR8Ne8QBsiPMalxKf+pvn6M4sI3h/ArRvpmYfD
dhMZe1KK5HvVOdqyXgMZgzhwfL+hZHMwt7OLaeH2JVdbjDCO/nuSkFl+XK7i79Xi
LbgMksIleDkHuFbW87Q4S7upPF665QKbkVPfHCqel1SEMLfZwa2temTtGYEbd1ay
9suokxMyU9jcxFQOVnFbYNeBs1+X1jNEUVb70GNebDZRMia9ELPo4t6iHPgUCYc2
csxklzbf7d9va+CiJZI2KJY2YGbJ+G+7Qgb0CmLQIK9zqTJHYyx2VZt38dWsbI+n
HborgBozu4PGPeH1W+Eapps3aICrVZ0SpB1UmlaFEjD2iY1gRjn4Lj40IEI2m5tT
kxlFDz7Wrogk63GQtpwJQM5aaFaT1fAXUwfrp1tDxsCuAvMUkA4zT3Htdm9JEwb+
MjyqquNKg0C1bSEN0edqPMx97bqHLYG7xszuGb+eufgiwNytkbEKKkcmqRra0HBa
IegyBgLefzM6r9z638wXwbXq2pNUuEWSz2SDPeRL2W0uAsu0TndnU6HLTPQz8Lce
cUV5cXTkginFnsO+uiftglqh1/3GW/h6HWjyeOwifLhhSJyoitprviMQf2LV4C99
ezsIxaTW1B/IVUDKwJfVao6ccP5unndOQKUOwMekt2Ai7v8Ab0YlBiIxoDPzF44x
SlkO+ROv7U//l2qFCloK8939/glfG9L3Pzvu4gCuggd6BogYg7Lw+J7ElffN7L51
YSYx2DKXf/U5FislrgE3F+B681deoqAU7qK85WYWnt8AfO+LKq7VKyjIsN1gayXZ
mQ8Nvoqoj0wCxZKG5/QJHVFW+eUifq+36p1mo164ytvVgtcTUo89kuNE0XGGdSgR
k/XesK9SVy+yc1wwdNAGfLVmlHSVBVjD1iRiYisEGl+7xWbvbJjwHItUB+LzZtqJ
PfLam9eoDgBPDkN1AJIs0TaWdjYsGqlR6jRNrc5rYn2rEVxWYQ2opYb1CIAwORv9
kNsxHgu6G+HlsROTFVJDAQXfGXUgz3E/aqNBUS7zYCt4KENE0QlZysrGZtbGIo+W
pq17iN7vpAb/IwoC24YN4BjVV5JtcKczqznGCuIp3+FQIS/5JuUd6tKrXsaFQsqs
MrLCsCU3PdTswndaLEDikvVQyA6Uc4Oq0pS1fxPdRrxntEYu6RUAnsVLXmkpopi7
hnidRqWRCOTVJfhfhRvxc0LlKE8hVSiK3m+HoNqGgkyGTLK10IZ79qNg1v/FLYON
AzHbsMA6XV6ShPR9x3IPXIl0GpC2RvmyOUsjJhgTQOugEBzKv0jE+KgysYBloK7W
FHBc4Jgvga+j+xWUYVA6Xd1r2gG05OqEiSZ8INXZ45a7VzxQYxch2dUvSvqpqatN
PDUiQhaweVDzVJ4gJrRQobpw8vcCex9oO1JijE+K9cs5NAVPiHMasqEA6D7hJKjy
+XN/IfwMn7XClEMYwgmcAa/4Bvs6JpQwGOtjp//4GlCU+qmbIMTvvs+QTy1TrGB9
aIAz/LprRSHSR2HWQh8XZilUtEUqAc7bvqGXDvUVIpojQ6liHragFkVTG6ahRebb
zQPCvOEqbV3NjJvx58y6f3f+NrCTzGIG7YHH1FcuIi239alfoaetOSig3sIHAH5I
g4If/flMvIrnZrAwb5Ill/NNtTTGVrGeSB0WGlfkJUc7Nf83SEPwSrZh8QMeHcle
C/tliOiczmvkL/pgoig7dqfibFSMSSLimrIpswM1XBwhYK2HS6y5wI6OdYRLXFcx
qH8chP644jEsFYbpdRCH9sbcR35vAXqeE3GO25vqkbznaOjW8bS1NEnV/99x9tIi
+EfIro6CrIjPm20+c+BG8/MgEUlshcXcbSPg8XxyrBna8yq/jTtHaA9xXYvyCDvk
k0ggSY2SKrl792PIuOQ8wslxX9HXENf7fTAkHXCB9ywE15Nf9kUj6Z2IwZGRD/fQ
1slK1BV9ujMwcrl3V2/QUy1hFgVFcVhMStbJ4deCWYgdz3tl7zx4idk62UmLttCA
mfp1qfNqye9O0HiossY2KVW/p6jcskqCx7SFr7ReYp+gyRVO/gSifd3cIRWbHFYs
Ro748CzfPu9nvxmzrlua7fyyyJDofoCU6R64GU1bqRva4onhQ292kGCq21+IBAFj
cPMBUtMdxFJtJwI3mYrNqmMn0Hyyg4t73snYMqRWZWepm8qPvXyhfRDpyQrsjqyH
4myYW/EBNCE0zWXJcOzCJ/ans4bWiFzMMBlvmxG4DrXj21h6mhuUiBrMLPKpmdF2
T6uvru5AhahtTJKWQloDiEgKtLFRiS8TmEyrJR/g1U1yHrDczaUBqvouCpG+mDGn
bSNTpa1jIT2v99JTptur4ughAntP93lh66gyBn6Ygzlv+xf9h0ZhB8V4SEymKTcH
nzIB7VQ/8jLDuwhRmv7TfWF66oUftF4zF8Oi5KtOzAETU7urshVTJ4GpvEPlS4Ml
bC678oFeCOJnMUwfiuYHqyipOZJ3S/1UwuHhOQADaQQUWOdHknuPKi162bDHqA/r
0AsRzm0qnjwpXSCSnyyT5MJPB8KgGI9otGvlBK7CNMWG8xcnkPIPZApqg8AMgpX7
Ex1ASezTBXWp6xwcP81LzXIDrdr8r4ugbRFhctaFwhYgPMxhu47utNmiwsqiSILH
n0L8UbkXDKktAmPp9GptPfFUnAldyS1QI3A8A2dPiRxvpUjtvf6vjasZE6nIeQzx
34PGtgx+WIax38LRB4TT2avu+Nq9/tivja9SqI4hyYlgSzOe7zH+tHug6HfOZCTR
AkKNsb5J0NGqRm6rwbjOQvdhwMS/7aC2laIpqzb6b+4xbqVrAPyBAoseu2BQD9JO
K8jrMbarFGTaeizLL9LyoLU1auYFR7d0pjsR20L3Ttl4+I/qOat30plTVA3LoKfD
nIhMr87/L8dfVnBxiDR0nYzSJFYwiD1CzSD+gmaoVm7DrFbXoAkKjEEqND3OpPbb
pLrEpkHKnukNjyJtjySjcUDJw21zDVCV8rW68SMmeKdM/UJDIMWg8ChnmudnRCk2
JlXHHJy9sMXX/w5q442wo8F2q98KDQ2jMdxvwMbIOqgwwSEDvxObKuTbfnVsAOJm
gzl7DcRk6i1BtgD6H6PtuTT07nGDM6uoZY/6UnfZSJwcWDFhnwUwChmnOO5LX3TW
LlMBArhaMr0857VcSHs/86rR0TNyaEaTjk3O+sTGj4XFiiIPus3UOh5LRsbvG9+O
dIo+BNLTHRNx2Nfg732BLt0cfwU8SfvdNGG0lfFHGfp93kVof1Dt74qiJeBzBx2S
kaB7AoPTKMnUvFeFsmNnXUXn0Kb4krQk9fzoh077yCg1iXx/MoIDwT5PuyWuBB8h
FeAvtL0DI/GBRgf4FgLi5I1vfgt7zjNlLv5Vkk8dbyn7S72IuS26OEiw/IfPxuAP
pQd79ErINWMKTFp1XGEoP9m56S/0mrJF4LuOhA0bEcgGyfiyltMBfFc6X1Yo1Wrd
ApPobiWc5QjfElppCswVjm4JH6iBoklXdlpgPI9frCN5iXD1TnkN8zpABLyWtXx3
ndyOVeJVFG0BzXLlcw3Thf7DSVWFvDojxe41Zmh2TZ+xBl+ih/X5kR32D3D7IlhD
IA3SIykP6KzcXVYq6oaAOquyQVyTQfxONFNKQhMVcAeWDASYPYpQJ7MyYt/ouOEX
EG5wQHkunuhKNidjJiKqVFVUGOqXjUJ/d4Q+dhDT+sV2P6ERGrOFSsjJKb14k8YI
eDCjmtv3coqT8DpC8adTJBH3lX7P4njaL2NxFdMdtqw9eZ8SctkJG6psOPbROnvS
Rwx9mhyfwgkzkC1JHXBx9t0m/JUr/33KjbgynVT+7+9ShpWjS9vYEkOtWrqbJO6X
Uk1XzbyIJzpWfvlAe27O3zIM31ZE3EyTXcvM7ARbkbKcv8pqDr5Nw+VSUW8hNWnG
LxCj5rWZbOHL09CqQuwXPBgig7D2hpi5ws2vRq54w3E2xc2d+G1Xmy9ZdHOUwWXZ
FeWBd1NTUVpFh/oCLdrILrGQBtB9jOtelopI9GZj4sW6Cjtz/U2nOdUEys5ZLU2s
a6+rmxkOmyPDErPbWxjQISvtND0s1lwBjXMiPQtA0KK8VQuKr9w6evKaErhoMd1d
H+irvySVRV+sO1UuLRy3SHY02vnh7mfOlPPFllOH9ygs0gvC4mAijH/9PLeb7Cqe
qXp03uu/alh7kEl/n2EPa6df98S7OFVcX6jrCJscVaUoPFlmKkhnpeH2T9R3oVjX
QnXxoMMMOvs6N3gLKIKhwoz5QbWssUgLjBAfSIXG4OLi8WNSrerODUakDPOzve7n
c60YTuT0NybayqszP27HCRXyNpSPBYm/iw+DwGEPcxxgb0Hf57p/glneKOLb/vVf
Gn1BqeJtBkG48S1W/mpaiwYu7S5QB0+8r2UbsRH9iLxKvv0XWfe2xmAPToi3bvaT
sexf0J5ICED5mRkU/9HP+KFI16mnVyPym11N0P8UW9loIbFkg7ExY36co4yRFkKH
Cnr8YPb0/LZDSjbvkloh8eWCboovzcHbjQy79Yaj7RcLNhPTSBC+YSknWosYeeTm
2aO7IP+HIoUPvGHwYUwPfsj5oQvzoPwvxA4FcIlaFs/3TjijaLc+buBAj3hdbxFE
XUL+i/pdBIN8RkSFdSABSYcpuDBHK6hfc1EdSRkfVnyRlrXlvZcXfYpqSJomlc1k
ieLfNKAvdqaduIYc5jhRAtrGw5umPd0d9Wx5rEB/mZyrNCnpUQs0tzfQMbTCP8Ak
HYqcv+5sU6v0DkRcxdrRyjHG0nIPHb/W3oiF+/1SeF3jirve2g7+TVgKxn/4TV90
lzLZ8ExzZfev+SQ6dOmVecc2bXRR1GRzf6HyYiLpm1mDJRLd23nCCELTC655m8i9
n7HiylOCe6Ses/de06x71ZDnBMyfrJr1cgSYgbu0gpCHNfyCoIhtjlgD3m2xhwXq
hRoTfYOd3pDjaXtX2WNVvbGx3/wHiyEJN+GPks2gurfvwW41CmyVLDKfIIyJLQYR
5Q3wqLE3I0KBbIKse43o9q9L3Gx2hoKOWlDy0p7TTyM6TwJFfkz0nUw1Q+Llrs57
RgSHaZdXHQ4RwEgPxejDuRWNcWDjHQLN/x6iHK+68cpa3AcJGvsKs5oypVb7ezHJ
sXSY1v7Htp5sFTPTuD8oEDFUqBgxiiYJm+CAMaLM/wdUmGfJ8kNBL3cU8iTXY5pl
b8AmixZFI0x4JI3bcjnmLYg2dehB27x/7gT/TVgvSxuX8KlrJG9yzckuveSkZV6B
ceUzdFR4XQMMTkpbzbQd99EnM0uHTepGpb5pmTATvjkuAT6BAGWv0Q6IF0H+3d+V
6HXGvOBNT0ZMlbtpjZiwec6tjLx1Xco4/KNbWVauummfbZ+D6lZt1f03KMz4ew+J
cB7PkikcUWMsBFcwKyR25+aE000j/O+dEraTy1Uk2sQebo/qtIto9Pgzgcu9f/XA
0UV9NFJXuOm6IIadJFBTNLghjIoOGF2vLDoF/NkjEcET/5a5/gJTmS5brH/TRAqO
a4gu9nLKt0SXw7H3MvFFtMTUw/HwLAJV64X4nCXvQTCciMvnVMJMgC0W3MSbImSY
3wgH0NBz3DbVyj+jghyjIFaeQX2jLC3tV+4puVu2EDx/eJ321pwsV3SX4dIuny7F
vP3Mk6f65lrhx74fd5TYRmuuAEaqMHOKwX1qEyTyjIr5uHULVB/udRCFHJh0ZNyS
SUqb+fm2FE4u9pP8FH965vba2hrKjemGcZuucvQ9nQZWCyEGg1YGPbKVl/sJ+1ui
k4WaXGmBO/5yw4tEGTA7kiKktp75EOvqDeq9IeH7RnRTa5s7risroj1O4uaIHSuM
zGcdgAwfup9gAJ90/FPfdsOMZQcSa9PWSnU1MgAk+KlmY99fXQ7/aEV+JZgw6HPL
meXM4/SUZIvJw90+3+IaJXO/stfXgg6+97ZQu35Pc2YPDkboaBpB7FwcW1Xf5NDD
tcMY5q4N4nHLtfo/29PEleTUTftg0t5soNbCFR2UUKUcH7CvdxRKwfW0GP2+k2Gx
3qVfxrBZhM2DA+ifb88Xoh8I9VmBxVncUQS8fOcjWsgnikDVCZEhN1zQBizS2gVG
kEX92ajEaDJeWn2vmBuUqHJQ7c1vBNYwPvrjsJWT/MaL325tAZG/28w3fT0Y6kIx
NgROaSdecUxktF6k+7JNXz337USxxEmpCf2+0q7xhuhxX0JC9RXEzSKMlVdBEgK1
8eQ5E5fSlM5qtupQf3c6cskX2rrHu0m6AslLxacY4gvqqgTFvsHcysdnAlC4v0F8
adsx6eM0uIDwmfAjSr/S3b/qvMZ5d4BN1PMFd6ziIRJaREbc15JhRwR09YQmM3iQ
hCMbGbdfqUEtt1tgcLW8/Ft2hzM7UTqPOSwNmG5tNZzJegwulmEt7wlSPtlxCc3S
bN2BjYpb3be1xeuKIsGtffYSD/v8XRSPPT9kI3CE6b3r5pQ3I7t1iwKeCtQn0NHN
W7JtQ/kWPF8mo3/RomFbr7AnI9riy+QBU0UOWZFoc/fHUTFOyDhy5NTelnQQ6mVm
V066XcCgD+gpf+DfciDGstx8a0a45MEI9ayzclYgA4lSk7515TKmUepN1iD5AP4f
uv0lJ9wKcYpjmuGP5YKPo2bJ1vYpICqVjXuh+nZyoLC6e6/bg2WEe5S067JYWR27
749Xz1ayqKegvN7qU4qEkz/7EWhDqu+FA0kA+4JTyOLVZaqOmTsP6r0Xw/JksEHZ
6SXnX2bOCcdvPR0FERMkQqLovlNmDLbQ+3O6heVFLwnCR8agcJCzJnrg/aR0TgXv
PqTT+IBOBiWF7APlUA3jgCR5yeWPVwZxyAbTtFKmQvZlhwgAy3fsN+6malqyX7hl
Djcy+uq12CzwXf/zjlMjF2h33HPdFpuM/XiCPc0szyFgFUEU02a45gwIwF8TvZ36
w/4CQDjSDQjgNlqGeFtnTawGNBggBbg6EAqMw9kGELH+YC8ssmxw0gZ0ttEnd+dS
moCXataSyuRWbhDx/vfjEcM+EgUmsIWLDxL1RQTc0RYePcZNihyoCc5h8ybmD7Zc
c4VpKJxkVHDx+2OwjQDzvYjmvvttES1L+31Tsdw1m3pYbljY4NeO8xkgFm0EqlUH
P6/QRIzrATv/oOoVFuNgj3DkxxecnjBIf/liSWjwiulrdTlIiP0JloLOJlChg3Og
LPfzzW70NZ8z411sp7qooSLz5zUusfgPCGbxuaXni0v4NveE6I4hh9/8PA4sYxkQ
GyruYhdXYX7JWOHl03wc6uAPS+O62Nc6R0+myI81mt8l5xtwDNN5Dlgj0ZTbB2vE
fslv6ELOB/wKT8n99Vf+g2C8V45977QIrvLS01Re5QGTqP/GPjQiKu9XEB/CLUhK
2UAPlSy91FvESnMRprPsdqWABXe3KT+IE1PLTWoSzgn2S/k/+4aTTxZ+uPvbKGhu
Ds1HtM9gMiDizeHW8fSb8HHSi4RGz7kNWwe6LAXkm24cHy8B9GvtpoNsLlLRkvT5
gDJVZAUYeKmh2GItMQm1kQdB6Ix0ZB8/Nbi/xnIjnJ2/uLIjw0gFm4BkdIydoA/0
ucRguie71/J81T2VTQCNhUHcTf3tBB90LsOPuvINQH6Thn2dPZDQFSgunsAJIKdM
3VhqfSoBQ14a0rqgEB9WxrXLdNZbk2dpYEMYJPtvDDmlMFarZxqeMMlysyTfJGpA
jMLAFOeQEG2xjWLAf9582WzTn6cJ/rbfayLumfsJQkDG9lCPTxrKBchWuuW+TPPw
0YAow5dMBIYbFd4YaXxrnYYUEqTy3Vcs9Wc2mqWQmFPCheyeNA0/kEqgNbYDuEOA
kH+/Or7P5sE5Y7kY3KEkQcADCJpuKB4rx6h1X1YGv14eQqAz87yHaTrzvCXuV68c
ZqVP92F31rhc9/UMDmA5H+wZGGQ/Fh0mZxLwnKNLPmBfn6h4J3Ce6OoT4icG4krt
bsCJSyEX1z9C3iBp3OyCyBwRTyy15jpMhRPjxhb/6IK4p20p4b7s2e3UDiYnrrdq
3IqQOgxuORLKTT6xC1EbKAe9mfm5vhJOQ98TPhwrfEE1PKmumNNoMGy3HddWJFcp
uzkop1U4MiqSVz4Zv+ZeR6FMNnLHxCeRbP3hU/Eq5lNjJ2xEs80ctwkwUyGqCwss
/lFh/yRHSIeOcqelR+/q4LlqxYrVQ2CcoeMngZbAhl8bVpyZpVKpTLi7kErNQatA
t8O0AtLu0TbqICnvnNhPCkKaJO0Pg4cwgVW2dMpznqj0T6/PYtR6YkFZjMiZlYWU
wBl28fLq+9DL4upQBc0EccLcPVKEkQTvu/s74QtGlbhuOEcoijCZNuextaH8Ko/0
vEiPrRYh9G++Cj1MNHbkayrxbRck07yaItIvYVkvVpg7OYWKhP1FF2658bATvGxt
exYeMWdaq5WlaX608UoO7Jg8v1njez3RhcpRzRcPQeRx1CrnTonZYXDSyjj5wEih
YU9adW+y6dWi+z2yoRYKaNaDULdmczK68iAx7DmUJrg3YXNHemDpK1E+yqT/mqOF
CmUDqT9ld3fvx3uw9ksjDPcIE4Rb/PEqkj0ArUOkWZefl285n3dworEN97708r1V
p3u0UnBHjJrv7OttFV1+vrqDqJcP/4NjBZ4zoDwmGg/okIn0U1NRskF6gRDCtlFc
MFqKAVf2z+E0EH/FMp2wrO9XwUJKBc/ibl9dW06Sgj+GHsWEr1mLZSiAoYSyOq9c
c9Tk8OHaMdN1cMVP1kMV1Aj7XhAhrXykNg1bF44TQQAssPWtlSI/zHF4zZNmc5EW
I3L44ghohQPbZ8vN7PyFYsZLem68u+efSMGKyQ3hLP5Phd2E63aS3b627sC342Rp
vgFR5G6/D9kX6KHjHXLUp5V9TNsICNb+v6IJHeFRutnvx8EjFCa6k4LgJCkFBCUq
RIEZTddXuWjpbXzBU7QTSEO1lOLev+5HQxrdrFtRQUFUuipO+JmdxDVs64QcdFxW
6hXkDE3Msyie7uaDiXexFgA44cH6KboxQInIAKtf0XGyVB/sHNNDDfPpqemGWvE2
RTVJqquFji7vaRVcoCVO0d3nDs0QEVRr0O+/ylHJn8QtfPzBR3y9Lg4CTaNNKrUO
QwDcP6WgwcOp+XqavI4gGtJwXrIIaRfh/22LZAQJqtfNJ3WQMGYuzj1cEaXhNTrs
7EthaXSlBBLiN+uzF/6zAe8hVxpMDpAsoXkgdlBB1VKNe68bDi6LvXa/VRl6XCfd
ghVHwhh9pRcaCpPa6LGp3cRy3Q7Hqi2+0wZyZb86OOwmhMtUBq4+9uSsQs82eH13
J/62dprEU6UyFr/Vji5are6CyKwCvznMOCsY10G2t5qwOoKfw+IrqE+l9i8BXtkN
cZ9o1N9V9xU1jmhUVwpIaOiO4Hte9hGPAHdHXyLYeWYrsML8fL2jNqcIvLxnqSdq
x3GiagG1mvypV1gZ9XWCjFUSj2G1W7xzxYN/Ogjc/1kW/NaQLkyTN4UC3TQHFLsq
bvVRfPmIoREalqx8iCVSsehnIqKqVs8qPzgZFtp2IYCh4NlGa5bDLBYX7WzZ1lhF
koCoOupOqMZ14aPlcLQs25bhxruutXWYVHr5S5xvMp4wyZJxYlaDE3ck/K/3i8st
9uVHYPebM4+K1TGU8l6dF3gyPbdneRiOG6uUKxJkYJQK47KqkPOC3SOIbPjug4fj
3n0lGzii0UnuxAZo9rd6PF8hopISPYOpt6F6mtEl/mPLGqoJulCE+u4NqcOkKU2Z
oOvCLN+CEbxe32u9e2DK8bhInFBk/Ub8fhXqZ4SSkDVeq6zAZ3pF2kT/UFwjSn9N
tFGMJupC/Er///PMsW6LUUssh7JnWzc8USE5QM2M6KLjqWwUyE4UrsgxYXMGZi/M
bnpcAq4WHdUm86SiuJG2pKlM/JN76RKnALLBgbX4Xim6M9gdIIlqdLWhucuqoRau
EDfkY2zQOamr2iNPEMdmC2Dca7DSBxGdGR/pvqmd0IJVWZmwKvkYM+mxpdACN2ui
dXhpDl4ofQJSqOgHltieAN7z1lcnUZ1tNQUSCiJ8sJOMe113o0DoJ8TVY6y/x/4i
/bkvgjAx5JCe4SIbvVfjRRx8rRRR80pf3wtZD9pn3acOYayjKVCZOAfy3q9vwkrf
lIX0IjsoOu+iZoaFDfQ7+Cw41tfYAmbR6s/yw7ONProvOWi1P2QmuPlJHDdmxQaW
j2yaXuyhT+LDO53TPRDWdZPbqYwewLsAM/ecZTahlit61Ddwn6A234voS3C894ck
e9uiN8H8QW0i05NctFN/Za85ZYy0AY5l+A6+AM6LFsEzgaVLM642dVh9H2SyrQ+z
3Ppmgm3uxhQXZwQDt9z7wQt6dOnPJW1DETR/fzIn48+olVw/PeHm9LrxTAwpyxIm
/xPncRqLeSeQgypsgoR2izVKIyIYS9hoYadBbf4noz1S+5h3ZCJuMqvqGtCTZdss
AniFoxXUIr4cV8Cv74olMnMRG8qKlh7aO5Fyt6Gch2MQK7ht+Q6qv4fY2a2mU10p
fZwL1DL2hcnDlLgD8cyzC2xNOi4osghXfTv3vRHRyggfIL995kfU/AVmLXam2aJ4
vZjTqmDtXSMRbfsqDy0O2gJzpaAhd5REYDaM/dTRIr2W//BEBNz2+IEtTQ9EMCx0
AyjAzLUtd1AK82X22/T65fZvJIv48n1bM+kZCujoFyNb4q4jYFkJGXyu3YyjXtRr
06La5rs82d87qAJBodfYd0IYeyN1P68fhaEFmyL9z0wF6oirYrq6Bhy5xbbA3DVR
NXyrB6wpaoLxE5IIYk7FqWxqeVMH1wJ94nHeJB8dgO6C1/a00FqHaoNETqOw9rhM
NdILJZjynEPkiCfkPWT+Xd50uy2crhXrHUMJnvOJPvRgLxrgsKAsgn0HVk8fL/ZZ
gYS5a7WNp0Bx2XFgeHwqS5uYPvgYtI7SW6zUa4OJmsKamf1KjBTzqwQn9fQp2dJq
/f2p4RIpBu3IPGtsYOvxgdRQ15XhZ/EQWeH+jMLX0JgcYGRmlwpZlE6/YVezmGIo
/Z4UlQltDNISR/0J76vavG5jrl/weLS0hxfuAmN1WTkpYfEglpgLnmQTROlJI/LB
+MqZEop2XQi3IEdeMJto7QD0H2XErI4o/9B0cM9igeauFVQ29KUBtpNnxTJcZFUu
t0VGyMa9K+CXvxHJFaG8+TxjlEXWnR/KxevEGYzi0tStqMVASTmLish+NYAJByLR
LD+bHIGLjSBE3wX+oL6/Gjwc/vkLO7KvoR8cLZQ2kDqceRm6+cgFh6GJtXEnGg1U
9UfadEDmUq8D4bK0lSrKMaZ4mfo0B4nZGOhJdEp3USJ22qWzK3+pdK3FDqw5JnjG
l2oD0hqr4/XgA6IIkkoW7A+svucVkI6YxnfqZCCZSagJ0qu0D5FPJ14FC7aqm1ok
GAfUfwLPAuk4qAXCEWp9IXsKbD2LbIiqXvgBwKFYCJnS/KYbR4DYkEVkjHIT+Zb5
SExqIaUgbh2nWEgjmLiFvaS0CdFDKDXD30qq0qhmVU0ubmEBRPWOm45zd0iQS8eK
kEWOpGK+sGZoTPDXGECZUj1BO8CVm3EllQTPtBRyWaqS3hTANzRP+TW65opPBhSe
yAbt3D7rGILKzBhgq2MyLxCfCEyCoKaXFRUVZOJ/yAwXEKVwvAb5CFYPafVFOB6n
mxiQrubYsMw3LrsWGUN/0223SY44Oj+FDnfIsup3MSME3R9AaQOlU10uUJEZ/1Lo
GJ9eKoUeACzkbnGiXDjgSMASRPLov50V30zfiSXt+6dq0MZa+uQqJlkhyXkxHLew
pC78SPDExzx2xCUI2zPm6CqIcORNT/hPz789zJfpcJKMkZH9JiqviqL1CFuCU5AA
6jj3ezCrjv9AmqsbuDWoNB8ZMHi+4DEkEJ1ivubhzL8jvxwrcmKdCToF1RvFJo9v
3yGlZFDLqa32iijIJWibDloiB1qYWSLjc2raN658Um9wwJEuAHukCpyxw/2HcUa8
bTj5pj2lFXhJIXIT9MW6dOvqM4QcyU1GP1BwZpiICsXbloybWO+IkISBQZeaGgtz
+QinrpJNiVTG8tpT7vVXCoq1Skt/sbbYWJ7Eny6vXF9FYEOcIGhCFZf9uFMeZSEx
bTKMRNP/TI1F6HamenbA0vbjq4QKRs8Sl4GffSZ/1xjnmfApwpw7u6I7NjDmGM1o
tnIHHgdB6ogQGMQ9xVxcTpW8hl2qKPRpMNXS84tb+QcNl3X8s1+FK3jOEMP6+lnz
tQAHDl7rsCYG0XpvZNRkdveBa2yrg1+nCHMVYFR3JigVaE8kLMWltq1tzjeqBAmq
tt7WPpbxOUrS5aHP68DvlZ5ZXbwb6XcPsmDfxMvfPTmHk+ssDGUNHTvcqG/npvv3
5Crb59/Cfpzikr4GOYXXidlSOwArpIR2wAmOhkfcxoIgwSHrEXUttY/+pV8Aq3KZ
ugwldlBUcBlJGdo+j50ae7O5SYvKRwzj5jrn27RkZxoPFUjF1fz84j8D12V5Y/B3
8yu5+ejBLX7WF9kgbOPapFoAxhpd9B520e2qKLNYG5SlP0AqgrAsArxK9YRyWSqN
TQNkICjS4HUoq1Dg9kd3klEmva8dIpEteZo/G/bKXeGbRm+SX5CglCz+doVTUy2h
78KFpGgqHTkAhpJTz3rCcw8GP9defCJL1fGIkzM7kHd+EvMWCrrJA0cZsYaqrMsv
91g2knQtCn47eDJKuGrTC7UoZKUeYRQ3Ve25xEglXQi4CsUBI6+ix7gX9bMAXv8q
KSggpuUMUWGO93ho25ry7tXN8WJFblQ49bX2odERX+jC1xAsWpvfwVHJ8UW0poMQ
YGwxEWEajE3HL83LH06ByJACPB8yyODg5crWvrPeFQf13/qdUr9RwnURDMklX+t6
6Q5s2YB+iHuTW5Hg0N2cKACOlt08OejunZDhZVb9P4m+18Ety+92tIl0shgxWvFf
RM2thZfOUWH8O7FGW5V+7YY8BtmyrmK3hQbdNOh73+iIzNlFvH+d9JIDdTeciej9
mMkm2y5Cw0EwY/1H6oqTJGRukyl4nhBVLaDvTy6cnAujZtHoHIg4vfSCYjzZW3hu
CvN5fBoeIO21yZO/W+EA2b+/hmG2wx4hjL/B+FSSdVLvP8C8xxB7O/dm5k2hPBmx
QrnVm3eOkjsgg0DyRL5EI/pqsXzblC+zEFqP8OMQxuWW9CEnkM82yXVlxtGy/4rc
fz4Juy33CAz5ewNuZjoedwiIkdJSyBizqVty6OPfSLtm5SHSWp18hKrvcTcKU3NK
nFGwQ796yfRfi7wlRsmMjZPvSIOkXeh2wtb3xq2m9OyhzbzY7K2wbgIwOfqwDMn2
WoP7VPXH9ExKXf5UPz3pQcguRfbLj9ndmz/CB+JWF8d2mUFnNPsbqb+8IjBet35/
keXY2Sr8KMGypmg1ccdtu4WrwVD4dwEicHAeIyKm8RK0XV1/jjLe342+TyJeBfFk
g7EEaI/pIcgqLVSj73pvHVeuiGGX2HsBBaJzOF+SdlaMFDoHmd7CZLO7Gaw70pkN
x3FokUyHyY8+1ZUDGhZ2bnvhJDP9mtr7cR230WpAOIj3jd0CFBooN8z0zboSHIze
gKTdr/AiAdRPakxd5WOgVOKt0FtE0x2CA2ZxXZqwQgma1mgeL2Kr3TL5ahwQy8MN
a+MTjPLOFuejNWISzBEkrZVsokvTTVrUkXj/EC5eI75g/PM+XKkSgv9jtlynCCBU
mQ9hsXvbbnmlEfB11whb+v4Dr+khJcG25C2AgCu5MRe4TZZkgqW4j6oaQJqXRIMz
TYluQ1uV3yBlYDZg2wFBTZY+pE7bIvLUZSvVZ4FmCoOzercSBrE5G0RQTSMUCeQ5
HhLQvi1eVnaD0xwaKxqx+/h9WgKq1NbRdcnNw0m7C3pT7ekLOlaYwgNbcrDTQzUl
wwoTVTM3cRalMjtHDS84KmGSjj6lJ6GVuDtIj6uu59BcWC6spUJhLMQAyXxYPaQe
Hg6av0PGIl5qdWL5y7dAv5o1DG/t3ezN+S9c6TBADq7zzGcxXoMSuM156NkRXFTH
BFP3xmOMJZssIgOMSwVjlBtoCpVcnT+eGkm2v1nc+scGBoIPi5tDuALGIHz6QGVf
lB63jeVguX0AxcTlKE5IToMnm8ZAAywScyFhlif9EjfZe+/nSCN/ZwirVhXKZPJN
DgGkWUrwvaDaCsbrfz751+BtCuPbn4xpRjjbSFZDPt+kWVShrHtesLuXgKc+YerY
imHTHrPhbEQPFuYgD8m76kX5lu2K2RMr78ypH1axAHeBR2O7GhQ/BzovTBz8rjD8
DA2lIpbBTNw7Nvm5XeR+2fibg7mnyO0/XoHcyl3Dy2QcHzfze8/vyyFbXR2j1y4M
r1HEYUoWkBwzNHUi0S+zCaMyCiQR6zL7x639yWVH16JFmS2I+qp16RsoAANzAnyy
k1KHm66zwsiOyECNsNv9mGw+dQ8+yC0gPnJQljwyTTpqTxjCRBHyXaZr1lvJPS13
9WphNlQBevpdlY1vSuuBXEYsY19A8IEK8u6bJGUoA7hM1zwAQpAMHyo/n6q0+72J
jRKUbldiE1SLY6EIvzIlEUorbSgJUT5jfZL7rLLcUDjPCUeW4VRn6oU1pysQKZPm
ZOtVqq0cYHqWo5jUMpsl++KSiwxLuc1N5K6u7U3+zXB0drqORm0VMoUj+LM9XgUN
+ewVlAeGKa8XhtOXIjsHB7rEJQklsL1gVydoHqvbEVdVm+z/vug2aOikApIZstGJ
6/LIfpD36+29JiNWuEh39pJ5IfFA0IlZfLqh3tIt8AuX2KeWyhP7UZ/O38aZ+fng
2NG56l5OYIC3B9Dc4SEjIGFgVWLEkDZ4W2GZiMlJQxi0J98IoHR+8RGz2CL1f+My
pXngZV63rzL00IbVbxW9xwcgRVTXQUc8GEdW+RZ6AY7py6ghbRlN5ctQcDn2zJpw
zC8jIaTFrw/y3GIr2JFOy0ezdMsa2WOTouUgUVH5JbfFGTEen9VCvDhrxUmiVq7N
D02Ctud5Zu9p9L7/8k8sPsaNjrv0aiy4bLD9ePDtMKrbFcYgFJ5OGvYAvMxoBZ5k
enEA8jCI36a18bYHvfJXBe7HCZEmHMBpsIyxZchcPZdKp7nUxAlCkziWFv0Swwb2
IJckz/kfLInw/6GQeLCFcRue66vIyU1WciZ0svkUmLYh0aLmTKQBIJUd2YG3dW/7
vCWTgVmhgUK9Z+kdo2cFNb8yjLaBSz++sPnrnO3WYQ2d4rED9uBfWWpxwQVfmfXh
mnY5UXxBnYAxCYJwouhdA2/W18vCO3OCllMP32Z2fLTouHr1meyk4F37gKCcQfq4
soqNP01PxqfpGPo7/rjvvIhdaJKKJTQSYhgck7JVSv4+gnoAgMAji6CcQcXCiR02
4aqZxTVG/kNGwg7McgpGi5XHXwWFUHeMw8xsnXqk1/7wVtnKRmuJLTc7KLuWxhym
Kj8kp6OY1ye8lktpDHZH/lth00k7DVBwLXFZ5B8Tju8bMSoNswrZ70Zsp0iXgq1d
Jz9aqBhBup+wt4AZMRHLlUdMjn+OYeDPytJo2VcvXSNI4+nHX15ssDjoGMK1XbfT
7YN3IErLvaXDO3z9ttM5aqjn5GVNNvkI5Eo3DY1jpG8ylg+Y/9k7qblyeN7G3ECN
jKQy6xjXFxoYaFOSx4WAVXpSAJwfNkT6cENE/thjtCFRTgcv1H/sI+oWJcuPxaJa
70sRKWYdwYDQc6mENDeCQQDpyQOHJ0NFXN4i2hGE1tCl3EG1/WxW3wKAELLknikC
zLKtU0v55bfi1QuNj2DQP3YvAzUyu8cFvHIgWEcDTOz749u6K6Jz+pRsUw7QK9r+
5QRCeiVWcPSGkVdPLHCDk7eBBHydx+nUj4F/FSO0xoBQXydOk2DS4ZKPz/cmvTxF
kaLKK75uukEAn4BuNjsE0qixeEZGsxYa/2OQOVSVCIakVOMFSH3hc9dq7GN+YFYW
qv1BD/Z7/sKdPGX4cTlDMCIfv8o5gt64XMR9aVTYllnRsWDQYjLdgzFmuvhnono1
IUxNL0qyXP1gnjWSFx1kgAB1awPtnfSXroa+Sz3jPakt4kxFBOjOfVMwhrwhq699
9XBZu+s4vPD+uyHA15Xy2orh4thPxINLCvieHIj3KkxWQW3u2zFSqslEkIqYfm/W
R3RjohpohsGuNChBeFzVaxtZpxnUoT4nn/bbwcpOFSBQjJ53a1OTMNuF9MNvtE9Z
LGM6ybXBlG0pMQuC/5RchJ+cOuIGc2ItvJv44uh1lFyOP4karZPA9OK3lv+Ws46W
HkaQ2gTFxpL5LGzxs4IvnS1SPtRwq28/1vL4KOz4qm3vcFqp87Hgz7ZNEVDrztIP
800THjpxOHtg4b2ApmJ+/CYH3OKA1J6924WI0ZUq5LYAdsJZTFjRltizj56NJoZ2
4xyUClEBxBEvbuoBJvn2DGS0hA3pZy7LuI3cLC82HzlzoVhNlBqEu0SvrcFLXDQO
2VgFKkSIQKFf/KyPCe+XRyMbib+pm7q+SBhq0xgOByDMqSRXKiqCaWvkWCWLQZFA
tRRxia3UtSWY5qIQwjjd2hPe7zJK/aWy1dKiMKayWuJLKiw2pE1hdam2WZbTHhwQ
20xA2QJjRTJ4t5hhRsKy68quKWxrRsgUBEBzISrXcCgbQH7SwuV1Qs0FQLRlpPDd
ojoqEa56/PowzI84Ny8o6L4lFz+kYVzKfv2z+874WxUj2+ovKR2oCU84XiEAEab3
56Nr+hfHe4IiYYr/+V4RsMvqxeUbVFKu6ed8tKTA3sfywb5PIDJ0kgMDHOqLNr4a
tHI8MmvZWSQRgK00+ZOwDfbncnJ7hxXGhKEusIyYIqR9rV70VuFVS9aqA78eg9La
hzjnZi69X+wRcaqzmQOoeINN4Kay4TVrTHFYptQYdxfY6rmFSkrAXdbXmRw7Udgo
F/B0v+zTQG/12dZphFrGBLvtHgc4Vz1sxEr5IrudUbY99zSPx3HmYhbZ+gBzp1jL
cVESPOfwQ/TMPwRqKmC5od5u9kkfEO7Hv71dLxAvtezvs87hthEGmEF6TNR1xM7q
TCFaA4Ni7Duf5v4tQW/OAeRktio7MyIKh7rnNgHbZ7pFV63oa4TJwt4OImg8YCaX
FXbHQyX003ADlN44yg7bYzGiPfyzGzytTmsp8Ay7GyPqiRi4S/LymaO33Eluysp+
eu4mf01FvBrks+jniPEC/9HcJdjiI1nF6qiMvMmRMbQ+hUXPeLaJ+t7dG6+bjJHJ
C7wPohiZShw1LBQZQfCcqL1huFinpoOT+GlOTBLyo5LDA6W+Z92Lcmysnmdnl/Ow
zmS4hzf98v1sS9aXL4BeI3LeY1edjgKLtlTdH/IwMTxN4mxv7lA7zm+fBxwXfrkD
AyQnd/4/RzHD5Qz+3jTORooGB/c793GoyMbuhScF7Z/jziyAMaNvKur1ZxEIIP5N
Uxo/18JXIrpzjZ4HekGgOehZaGlISAlJgb0hiZDW3OBZjqJuQlNmfGbaWsem6Ucz
qB1AUityLbSGqKhb30LN2ap5LRZ33/91bBcZJlXT707f63aAGkTEWTPhFltuphVg
ZY7FCwrxmqyaYKhwZ31IfrZ5PdUmFY36HvQ7RwBZCRIlSZzCi06659VVyK74m5Wv
lOAsz+JbvYvGWwLySW3KMDXGaCfXfBAwSFLrkjT8NGTDhDMRFgaPakyESFHKLz7G
ih+6MB0wVjaqzPyDMC/T8sUvNDEtTIyy15SZVrJBphkOGSgMsM7uMl/QVUq4ASmV
zLM0nlPydWOWQGdjWs9mY+wQfe/y2KHDpUc1ZS/WswZ5T5kIvvf2kUeIkHtI7P8m
Ej3C6aP7vs0J8AXvlZY2t3p+lAgDVpCMGdhdNhNgUB6fiRUpPouIcal0eVHL0CUk
J+gQBJdReHVo9sL/61wV6hQqA3BJBIfE0b/oouV7cIbmVN9Z2j2hMhFVtRwF8r4t
woYOkaiVHL5D+MEiBj5opT3wtPvx7qlKOY7EJ0APIc2RS0cDw72ezv6wRFOiJsRq
mdJLbbnTUvrMu4vhiI2aCqNUl9SpHs3AZ2UFBJigp8xNY/9toDF9fjauHKZdZ1Ds
2QcHQ+XTywPGfzpduS4gLeoTX5cNDqY+qNYdoNle98ZXE5qlRatDNqAY86bMATDP
UJ6lFNfM+asDtVtFADcStg3s6TIsJXkqdvmRosnCUiHjqySK8M+unundQhFSTE7h
rY5G3Vsbv2icQdDletNzZyqGK2xrJNHpkAIEXl2l2Ljt9CCST+UECwMZZP8e9kBR
JNsTlI9iM08jwWVm5iPCbBE9L2Qtv1KSazJLSA7Q8LmEjmaLALphreytSqShhQy1
KjGtodbh6hlcWETgnBrnP5NhW7gntoPrcryzlcOxvxQtt7loxJWjymi+nbB6ebj0
2q2tB9MDftBPqh8/k0f4BuWSfmYEkbPJLEh2iObnVGKL8MmnRiJ+hV+9YOWXPkhC
+siC5Ag6u3X45pb1qJsVAHpd6KGjswsx2w6RabDCazTPMwVMkYu41UGLO6/2kuzN
WYpuQl3Z9koaKplJQxk68HDw2LFcgI14dB+Fp1UbQFzkFeyqgJCipMAD50a6CNW1
G1CeTnTz0evM+iqWowz0d/tPs0e1O06HjZpDp48md7ZEWR6t8fDzFD/QMyBXpDYh
0O7gmCT7+rn0huOYmSXO/V5UXjbml4tc67NWPuV/N4xwLpz3JFHFjuxlN3ffkaZL
EXkiUoN+hOY7K1CB1TC6RUHHvJ2s/5u0KUNZi6n4gWEPPZHdFhblrshp53G6a4vv
MxlrBlkWEeVXNvHHyJ551thRHsE6G7t/xTnvijRQogAhFEr0ZfzhA6DkdbNRNBFo
3CpC500m8i5RyiNJNafOqTu0uIGjlfV6lWLkxv3EBLtc6twqnDDIAEyRH00+JXik
sIp/ztJYuqpcWtJRmXAzqJRaYAO9CwSEUeMxLGbRmglYOzPbRpJdNj3tjuLorMFA
RaamCfi9oyDFmNPcojKu1BPBfyaZDig1bN5mphKzOjQdxg5mZ1Jw6zJsV6Ev8WgG
aE9lrUuChWorDTAv508yy9c6UJ+BBPspc7C+EUiKWeGRO5x1y30fzgO0c5eXCzLe
AVXXIlNkLoWEZJe7JdG0chkHgcpJ4anmnrfzPgJFS2p6NqFcNvTNwsGyCtQYZDGF
mukbNsoxAgINuAdEJ5mKBUue7g1owjGJihcO0PeLvHeLmnkK1O21/k09r9mKwCkZ
/9kh4+0lKYUIgVB8V+JuZF+oAFoKVhJdqnKJX0tqHGEl02SZ+uJyPGqyJLFimDJq
ZaK0UqaGwcv/HXfv6q9bllexosF7FqF2Ftv/5RJvYvGjg4N/+jq/tepoU+i5vNxW
vqo30X/q3CX32WW9JD3i0sztJsd/wmRXizA9Zyirc553k2EV9RM3tEg0KCS/r17n
HhPbq8TqR4XADJdU7TCf7/2Vnvwru3aSZjheFIwvklkm3ErKI4dkAp+MEAvyNbN+
vbxDjMxaB3l7t58qCG/9Fm/faPyiVGCX3oTKmvx5PakK95KS9Kl2cBeh38dp5mBT
AkasXrprzwaYX0Ba3hFhwk/Nmm4QsY47NcxN2AJZqbZx+ugOFfD3ZoVqHUp0DruL
u+o1ESO+pViEDGmN5g0s2xQhjCyBheiJ6pNITaB/3WfG0CyfjkVeDas57ja3At7O
58DrgI8YyySB/nSMdWtoxtL0Ou7hQNES8Nnq6Eq6rIy7twN0OGe+X5OwD9OXLiAC
vUsQ0EVFwLe7Pgvjrykid+MDQCgCf8WuR3cWE8EfLlT62czdBC8F7x8wm7JQTIIB
X73zebqCJNjXaxn+Znb7uDHKC3cyVapddy4VwTMMSHhETVYrzTU72UOd/apTqlxW
me2AZqTuBNcdB573dxjb1XlbTlWlcqsuwjI0TAjKoCK0lMYDPXPbco4AvtdksUUQ
TIsnF6GzHCDfA1t8xQwGIcPY7WN/b7E69OR6vQA/dMtrfeWM3NpnLEUcfz0MRADr
4QOpGEeEKxhzq5OatvpNc/0WvkNWvdILR9jz9DJaBg7WTItIAmJBe2qsUro253dl
Ka93fetPGaTxuSqMvumSDXk95ZKOrhtzuL30PY4jjyWhDK0xsR83Db6A/WyPEc8C
26dKDAm6tob0OP07mf5QxpQoaQ5dnxFCRIpKqoEb+6D5dI9R7pmcA1H9QkH9MiXL
Hdp46IYvSCXT2uV6XDC8wBsJgU7XQjK8rDoKk3nH83GWwdWeLaf4+756X1wD9xs3
+xpgN9H0BXrXyIOHtIuOGoj29o+6BgnH2l3gDI2AU0mcW13JBwxhCYAQGgPxcsrp
bCoGlebmLbB1ZgJ6P/Z7eZSMGoE6WsQi4ZJauXsf2Ozaq9OSFCce402jHWufMj75
EsERt776ULmbaXmtzV2TA4eFd8v4Ru1Zhz5LHZ05U7uuqVaXKfOqVxn1EEMba+GJ
zN6wVtIR7Wcqx/XzAw4bhbQ5c81Y0yV7VtCmfYLKoJIE2rtnLVfQsm+4fSFTTtZD
SBSObsbPZraNQFAswKRaf/vcDFqcpwBUqnCAc6PCjEvv/qldLy73yF8pz1Zh6z7s
uatzzwBFaE73eJaW1ZiY99//LTJ3Mc35X9X7nVDVy1py7XJlIB26zcpj89V/FAVJ
Y17w0V2h5u10DpJeOcfSsXmRzhIpNB8M9i27sIefZZe8tmc14/elCe7gfJ0xSuQc
RnkwkKGzuQQpn6WhBl+gClMzCfX2GkpAgXFKGLxf7aer4s8cCEAhxNAPMMyhn2tC
yj8lFeQ25DkPwUaT6t5z262L4CEt3DiQQUOIQpOR35Z4xg1QtacsDQzhRlxoGlX/
gzrPPel7wSKH5VkMUer63pckuLRLD1o/RmUFe91ztr69X+V2m6IVUH/d5YStA7Hb
k/bDnWv4Rf3PT+t+ukoBvzixmO8vj24KMmSbV76HsJlU1Uslb+baAAjqDohAwu+Z
rukssHFmFBmukHBMb5uOqqArLxQ2RyjM5s4/zpeanY+0Zt1StXJlzAg12lGqGUAK
vaVK9BF7BJPj3dJ+humrN7ZElXffrK0BGOv+45co4T+OhodwVB6Fk/21O1Lzzjyw
q+jsx6Zn4R9bwHY0L5F1CiPRXMA+7BADod207QxWZM6fKag7cz3/ZSdGBoo7SyDp
tDDWCicrlACr/fuPxqlIMpokln3jdcwRCT4H+7dAEi5mhT1yvGVHF2Fr63zwjfLT
r7Syg4M8X30ya4gKJ18XKQZkX4Y7sRPDwavLEv/Km6JFr3i5rm+Sp2D4KOzvMvs1
AIAC+lbO+uYbOb+TB0uYNCTKT3buSMvjZ3yve246AxQ+ZPmD99CSyquBQ1UKaMF9
/gwz9K6F9+fohIQcoTIA4+xFrKgYYK5wxziYHDzDkVPokWJ4BDNk1h4VgCVlYD14
LViqd5XAYiZshm1isM1Q7kgt8V4ErVYcbqPoqx+hjf+wpYFxBnbi4L3R+Q0cZTp0
+5laLzvyQNk7U3epdK2U/3S6kcj8v6fOiMHEJriAQ0Ibieop2oJbbJ4rMgOjh7dX
nd3ygr4fHUT7oJkAcc1zjSP9ohzIa+7BA5dKuexUXTApXC50HjcU1W3QT7BW9jGt
wxEgUJ0jlQj36H2/1SHpKBgtYjICISfPbSfmF7CzKUWmScZIoudojejPRlczpU9B
CvGtyeX4NfLw3n7KT0o7GFe6lmMLWF4o3BpYshvu+ZqxsDxbVfSPVlrPCqPfLi51
jG0ktasfQydxYasKYBgTTHciRY3grZv4aC/BhBskzLK7jRgI+SXD0FUFVaJewjcu
DP2m2G8IzInLj/mSM3+jQSGR/BxwvAnBRTsVEe8Dmhz8l9jpvx23HIr8ArjLYaiI
r4iWDVCXiixzv+6+p72DgF3mruCC8tn5oaxkRbNGPaDDfYn1pxM5xSfUrmzgvuS7
JPyQFj7WqliNWgMB89pF7hr4Hrh7IEh4HrVWergIF6TyHe/FmBtglRl+b4zXSA14
2Bq7OOxPa0zct1llDAeLczBM9lW9agNd87CFeLH6FAexf7EurBpCe/onYBd1puly
3Lw6CwcHgRQ1AcMulUWrSLvNzdmJHfJ5bDsVxBlmWzmXZoRag8ggBjsyOFOB8ZgJ
s1aycBsdCe3UxtRHOlUcg8orm84GllbG2jZJYyiURRJipv6Y62d8nYupEOYkK6cd
IssfQYGiLMAlxlUERVBy+Ss/MnA3bK0rrVhEsketmqtBpJQiV1IHgxzu7k+ro2W9
kyfSWgT5sbANf94wGqYzC7pLVrTPn/Ucctnlskp7XpihvyfSmVqm0jdFTmEADr4M
LgWdQyXbKpyUq353WX0F9MwHWBkalcFfrpKr3oGP2Uc7bNqzc7nemOG7tOhXqVTh
FNK+cYdD5YUKPqx/EjGRktn8zzDj8IrgpPA7FX979CWv8dfV/HYKiJY1jO0M3ecV
Jp6DTg3P2PU0BQlK7f8Y3hJO3HAVQQR3nkjsMNmHSfzseQBLorjzGY7bfal3cBoF
3x90qzw2QQE0l8g7FeKV1JsQGC9wCBceO3VlCBJz9nCZmQJWEghaj1wyGOandbXE
FnhOH54YBrmqIs8GpxQZDO15nqZxzBPR5GinMLMmldQ821++wDiOmdotgX6s1LWe
5AACn7mSOb1jDa4YFcsopMDfJIdtudjkMvWbOeBNCW5L5pY1Vpv36c8gbySyrfHb
nnYL9i5v5J4hbmNcNVtHBWjPShIZyGAWWLcR72jDouNoqlxtt+HW2YzoicWXTtwL
/KKIdYlDzbGupwkztwGKEGD7JVaQP2/GSly+CqJWpCW9ODnSe121ZWV1lTQprFTt
Ls/wgZ5HYIPYFaG1RXaKVsrL0Aj4VD+WzKONkFgZqyWGHmlCQxqjTxyFBDGdgeoy
MX+kv8Se84V8nbaY6Qzb/Gv8+HAnWWlYF8hRopjHjfrD891vS2m/gj1F+IoiC8Ha
8orMf+vn6YGwg90ZIFFxr2v7XaBhXi3ppqPgdy+xd0U+gZ6UkH3yprfH2MZN0+Aw
XA4f5yr6zHZaY2ZxG6+Q9YuenN4fUUo1ZXDhJ1WjSmckuVPOuKV0T84DXWk6kVeV
SVkCILlybjUOAo7EqiJdhpS+PeX8DeVuIVh3qGI4ebBZedLvq+dtVxfUmwO70OyR
IVZj5rrQm7AE58u0pWChKOtBh6JZTPE08hFnP0AehGGmsm0Fd0wZeOQINwdvclOS
B8hdjM9jjOnXDDF+Ep2+i/p5IS75lX+seJ44lXRILBM4rAeHag5ER0tIgkXnGKSS
K+REEap+EshOdMCvOv4qVzxXcOjcgpwSm5soA6DNfZSBL1m+V7Td4fpbN1AOEmso
zeEAJscN8Ovc+Krwm41JXgYfOFw85ow6FV2xeKYcpiMRzbx0PyFurzIJpdeZFiME
d3c/IW1NhpKjq/xdR7u5XTpC6FkdzN+JcgGbP4K4svmZp0iiylQ14mwO1jm7NpuD
TLjcAR2sjlt4ph0ljwt7ecHLcu9ejHQcjVOJ4mXCGtrLboH4MfxjEfgzuwROCF31
H3A3zGMYZ4HLXd+w9LeFUfHdlQcBmEg2o9Cbmq5CtPwNI4Nc6BbryLnizFmmB6Jl
+bXWc0BVDS9J8BP6M2XNYTCCmoFMF9Wn2yhFA0DO1y4sCdUeLeBZMEqEgHEDpGSX
UdV7h076oJnK5usX75l09IvOgj4TBhz7RXXoMbhRxP5uyBVM0deibgGuw+mbmiMN
OKiJJ1dTwvkeYVwZsuN8+Dj7qoye4srd9w7cLJceV+KKiOV3oXbawPmIzkFUhW/0
eIu2XlHXL87O6Mn9esR0iO41em/fjedzbA+0kNwaMkB9hIG4tdoZ7c6QtIIbWlJp
Ug+aYwZ/tCg9aYvsnjh9xg/pDqzdaEnAnZ6MsZSZdqHNapYx2bxRJepTE8ofH6oO
5DZujHmJLRmJKF86rIhMXJ1kE8SG8E9WkfInrkTLw5Tx0bLESqCTVoes2pB4VFuc
lFW7mQbRV34SaNChgM6UGDZIYuUys76bfiHovYZflyrCBARFTmjZBZpBlHDhG5M0
NRxgCfNO8tF9lfN6kyTIG5xAkzq9+BHxBwrTd6x3GdJq64beCAEGHpAlzj6s/s3V
rfCnMOxhDS7wpYo35sT9f+G2lyy4x5uBvksY5I1kSQY+Z+CusGs0RKxJ4oKv0dKb
f4Rcgi0OqOLjXm3VHt3kiRnBPlOLE+H/iSCuMR6lRTdZ2/sKzavN1svWkrsultjn
ZgOMH/QwjtDJLxTsi3zY/iS9PXaRn53pCuZTC35KPgeo9kZQ5PLN/rq4PVWirdNP
NddtPX83GS7yT9gZgTqLqocbTbOEvxuJMi14ydsE7O2YWjzp60LMMo1ycQn5c//u
tV0DBgF3S5AURgj9QA+kE56EVsglwqFKWeS0gAYrrzOP4+mjO+qz+1/s2Ulu0RLM
ZkhQa1vUVUmRbXaJlXqN3ewEV36w9wbGJjKsH1A4OlGtJCmHxgIh61cznpyDkNh7
sjBUPMxz2OXfD88GSj8M0kakM0S7NkIgrdcu8pr02/2mbHc0T4arNVIndPnsRUU7
b0B072NfI+eYEKhX08rMXeCt/Ju3/rEnsNApjkuHdblEWz67C3EpVWITJzvgOeg6
B1T+d5A2sKdy5XlOchJZ/YS8f6CnrLCLZ52PDhLcNp1DEwtZIODO/4z59A9mNZNA
0hBCgpygWJ8wwAx8gZbmde0KYbhbv78TXS30l1Xq/55n01RSJcPdKoFGXHQgTDNq
iSiAUnCRagDswz3YTg9E9AkaMvE4xl67josJimmXzkWok+tUlE48g1de7HqAfATZ
ibbdUF52ddNHvPqv6kLkgiHct4H2HaM2OM+zbw7GEcediux4orB2rrhLfHGKeSWO
a+tczAP7jGlbCvGyEizja2iD9BF8/VY9DWWnLqRHv+Hgrb3TO5tIakVGGngLrh2i
FoIffXK/A3cd0GMmj52gSdz5tvq7yenF3hakIxfAxKVrDrL7biOReepQLmh0qXqv
mGuxljwi/Y90bXj/c6d0u+Lm1Jpxrk5VY2lFfksKd+QyJnI8cziilPy0n/UkaM/K
uxzZjGq4ufqFB8A6f7Dp4pfCgqnip9m3KwVjBb2SL51vWn6blnsolbPvHKCSlFUz
kkyMfYPFMRHXEbRFGb7rVHLw5IqUMbtDMNW4w2Vrjhr9Ze/jcavM/I9zkj+MFhrk
eY8Sw4zxW1X7RBuAM8qa1yjBGfbjMZLGoaaB1RieIrzHryQHmLAaEq8D+V9cv9pe
VQv7QAa0Jcf3nAy3LNmsZQeiPDuEEMR76xw1b6s0mkAQmN2Lu59ndUvxPiiZLkps
N6j5wL8yySafVoxxeUV4p86Trceo1FY1CNVHNhrLczKEHfk7W9Jrqv06nPOyddJm
1T3DN3uigV3KveakovvAHU1c+YJiGs6/hR1etXCgDN/kjtbSGsYe5jzLbc8WCLmt
t2wUrV4fRpXt5jl6/13op8qLEqqwCWGQBK6MOU+30Kflo5brI4JqnPJu5xaR4PCi
tGM+yTxl8P9JYEzJbYOFFC1VvlCHUZmbENfjvwbPvlkah+uKxG+sA8xAwjnHJU46
o68I9XKeEVsTfXp2Z4XCfNWlUo4yfQkD97GahjHNEUjQPlYVfNbg9xFy6MoLvAXs
QVRPg4+l+S7aayD84UC9cegvmaQyaMGp45ClP5xr3OTAVjnJDYPQTbN9RX9vwChG
9vFTHKwHkApfu96ekdkyRbR2V2/bU8x9ZN9T+i2aS5gQNKAYZvFazXZeqaaoF26c
qzcskkhoU4gOOvCQ7RCItd2RbOiKegij2x9KrAG2oYKz4RzEP+tQsLozj0aJ5jCf
Nh0SBbW7Ib82LAed05d0J4Abj4A2TQLv9S57Q5fGSlfsvagWZMs+CSMOpCGIfNPJ
Vw7W8M8BnhQWHTyjbhSjL7qEdiK+LxqiVGdvcYd2iAUewkNXLfNHTkFw2epD4+/m
ddE4azFJGjy7tUUk8EM4+Gaxxr1FbQ+7s973Bi1ZniP8I4CAuDz/kb/KIApRzL4Q
iBE5IKyz9Q4OMcobNxB7TxiQo/8vf1kE6V9Z3Ak0HD7UAY5YCOyKFWAiX3OEAgvq
8lmvJUZ9SQJAoFonpFUFC8F2v+RmQm4gmb6cbmE8JqZqGT9ZEpnv2BAOoYEQgxLU
FSm3S4tRMPYXvVCpL2F6RIG9haMhf2lrolk5H/TnJ4dp4kRAxMlV1rYrgoRrp0OA
tYBQTmDa2dqsyYNmtVuteumrP0Ac9eKPUxdZOKZ4lcmJRwNT9c9uRVo7NaYswybv
Hx49rlZ+Er8WEEvpmEMt6Yk1+uKsNIxRhVLjqd6gCvcdXzKn7zGKu9At1Sde17KS
+2fHTz1CYSR07Fms8jrS8V8icg5nTs7bdaObOxOmGHAs8hRenHsuNZLCCvEWPd0Y
FSaIX97Dl8bS44a11E31D1WwFmRiyrTBKecRESqaomDmgV442eDIaQR3NEtkRwL1
F+t58fDyqDxR8z3dDO5Mh+iPpLidwGKabyj9k/hnRDFrfIHtNGml3FaAwtCMsKBj
K5FPEK3dT1E/bRZb5emXpBt4eDdR3eWwwh/f2VIbdM8XVg/1vHzJi4ayPMxBF9xN
rLb2UMT0sH1RW59KZaEn2pTnlguQKGG7N15n7GDfcOmVLPemS29/u9OVCTFDxLJp
+Oj6aDQefr/N+dsULTOPCstxhFf/YKK1UJytq2qys1E7IMXZnRvebvPyKYmE0+TI
EVaqH/hc55OSZpOUOblrXDCQqbH28QXY2Yf0qiCemnMu2LRy6adAVdYcQM9cEJ03
tlHqdijGQ6/xyQgdmhBKV4kLDKOStkAN2k/DpKQaYC54ZZr7o9QA4ocw94CK9A7a
fTQ2Q5mVvUBlZSi2+JpL0cHjw6cinZT9WFRXmexs7svjIr2pYKbEffQ+z2N4BKok
USnee8tJ1Y/DXRsFnxZzgdkFva9feZ2WJvL8/EEGq9nUd1uq/mK3dAApf7V7P02J
MQW6QLcfm2DC2mmhmeu96fitVq6Z7jeBRr0JSLzv/8S8eE33d5Q59uuaMFDIl8aM
w/VOfnzpeJVzFX4CcoZkhX1IhET1rqvqAomQZ+8bPy28xleR0WfT9CoC9vIG+VVQ
hJj0bTOCUkgbLw0QQc4O+pwQXvsMcy+OdbfQ3lMoVZFpuajLLty3Kv6+PfxiWqVq
bIU8STPsjktbbUjVNDVHDYRcPxSImdBMR/1X48foAA0783PE08zRZIHmg3+Rcr33
6Hl3BAvh9RwlWXGHKwNX120hkaU/cvj6iQLX6G4jRhq4bEhKMeIDUDfbqmOyaSBG
fqYqzW1Dxv0iYsr8pWmwD5wgLebGdnKTNFTWC4nOG28V2sDLoVbI73zK/DzEfIem
vy1HltE7Dq7znUof9faGozneT9uoTRFqTnvj+Y8wICaD6MU/orBUP9cPvZWRZsVx
O2ZjvrovLBWliHUDo486KNsW4FGzCFDRh7VLWDWuPI5AChaqGBdVAOJYuXnB7HKr
Yi9nPvqR2jlB6FkDX53QS1tozVvN0cJhZSUM0+GAT4/IAkDYEV7GHx1+heJQa/6g
pRL8VIVb89z8mR9oMWOVvKQlVGzUKSKE2UcF6TOlpiMI+rVSl3or4Z1qJdU6F1mt
cH/5x4VSqKu7pwFk7Po28XFRKzkQgetHYKE5fMFVAx+fLb0qzhBMv6AYs8fPtAiq
C/dB+1lE1AZuyQFav2Oj3ztpDKEFagjMxag2G1+UppJl8y+DWhhAIVwO5Djg6lNK
EENNRY3gunxCGnnRvKiq15XySVcqJm3YDP5qukNZRzBp3CgshAZectXh7vSSHKQT
Ui4Kls9fUlGCgWdIyMHAht2jyVPsVni9A6qOW2wUsNtAJeaiRPJqNW8UTJ2apEDo
4yisIKmm7q8WbGKEys9dF60nXj/fHTfXPgylQDUv65mPX053KE22wu+gshqijGti
wFENYwUQk5/AY+BtlTKoCz03h83s0DALsRDbzxKjbDCpBoM4iMZFjlNXs2lyFrap
1pb7dy/JJ3ROWY7+Vep6p4E3gf2makVlsCsSql+9K7xLTOrGZhwybvvpdAVuAGbo
wibX/44fmle0PjeMJDr5dsNCXUJU+8QNwk7DV7hUj6vkJ3AGwFZFcJ08thuyI4mG
/YErK3bLhibGtxH99ua2cBuqzTabX7o9CbIzKlDxD8yklW/lNBqcOi/7BG2kbNzA
YhspDaI8ktyn/Rkmwq/jbn5hJXlHYhZTUZIrWCaxMxvwA/GccxwfNgqrep/d+gIb
PTWM3N4qE59pMKgtnnqiVenW+nQi0yyA8NaW3Hacfz/LFGICpL8k7ypnrqg1zf+q
Nrq7id2t34iOUooP+klwaVDsnuw9IpICypELv3hmMg7MJBS7E/ekaZTSJKmKUdhR
m2Y1hBIBeR1kAo/lhjhzzdcL++1hwqdaTCA241xaMEoOaJcdlvnibEYhlaUvzv18
b43BesJADVswrFMKEDcXNO4bMl8wdAXeSharY4avAU2E+fTvZ+19lkKIaO+0cHGd
7wE1NQIfAIsJJMWF26g1MV1cponswiuaCv8zWO9hFUtTspK/erVCDvr3b+kKXD49
vA5+REdEtXvQxrthGln4DbprRE2l3gd5K/PO0jn1TrgXgzYXGNbiZCg2OC68iM3u
82n+lRmREQHkOA+kbLd91q1gdgU5+II58Ez55re4jTp1igj7MZC7jtuxd9AXeAz1
YQnD1XAva/EsyrcrRMIHq/o/SL2UyQcKiMxuLUYmtC2hlt9Q6I5y1RiQgiuC1j2L
SHeT0UDdxfRGILXX1Q+r8eMBdVyfW6zRs57v96lz1xiMx9SjYTz8oEKnZcam3OEf
ST4XQRjhWHwd9fejP7pfukPYNrkts80/57r/1fdyx9qVSM1ZJKcHuvOa36CPyh14
biDouLmO85hSpK6rdCJloC/8aVcNOMPeuhcZU2sXSBsbm/nnagUUMoGXqV6aEXGw
DhN11aYcgARYnMAT/iqfkLTlVvTj5GNp1rHek73FMIeDoejeD096RHNLSVYG/ksu
cbgw0PejwwogYRYDgirUaso3DvWxp9xHjbjF27UquFnldBDWYfC6m2DWSbnCGkR2
EPCn2BU4gZ/eXx7HSwVRMaC7TKbMrZcISofWkEd8aPggLiP+8QKJy8G/drhV2HHJ
iAVz/QEmWBNJiRmfp3+Die7WYAHhhxuMFNoIXcZeoOrKJFD3CI2FGIdlJKbHbWtN
GIoWL+3+lR1yZOw/eHzVD32/nGrjgrAHzpujDnGUn/HGNGsNBpXZ+ojU2v2bhaQr
1j48tLrf6m3Bx+IidHh5FfCknXE4hnTPq7E7BDMO5zv/09DRQAdpBbwt2beTy6ny
/sHv2Dh50rS4R4DWRJSeb8f1ars65Exk55/yx6VcRYeyG9IPPaeRnaTdPgiG9pZk
MbSJXWQLu7e94cunC7oD5xtvzYOXO4M14Tra6OZ7KlgSHMH4hTTQt1bIDmAjLPWe
gzb1qm6fqbtLJ+Ly1c17fVJ+TkGMW+BLnRCW+wuK0GPOTeNB8F6hkqI5T3c+nb0G
qII2BZzQXXthHzuR5MBFXRozhoGMRUXMwlJVTenAUqraQS+Yt6yDkbJjlUdYISBi
fEYb8ZvEnAR0Z9GWRfNqcHRnHAi1JNnNEFHgpGVrAQQ24dAncGp7D1XgGvqGOdTJ
IGuoOvrMvdJ0bl2JtvfJ23N6ZhMfy+EkiHm8hRhqC3pshrjCtAtQwLNt+yumgc7p
Y15iYAzkAboqLezrxLvsgp70Cb+yXYDZ4l+ibd2r76fMF38+VyZL56171CZWNwF/
ONoeyykMYGdXwFm2um6EFgq37HkgMsBqUpK40VeXtRwIjXS5kFZ4m2CfZ6QyMY3R
zAFf5/UJMNndbb4nPaUdOZlNmrrSC/jTLX2cM5YEXYdIrVwWMFybxR8XYbqE3//a
PguzC/iqd0lMjOsFQnbn1r5E0WK0B9//hJjQ7IEOQtvfHor7uoANYDEMYKnubEP5
cml/rIbC+5eeTht1aqVSB2qVMdDjlx+/SN8R0OQYjtKLqrl8nuXNWvizLOhx3kfB
PKfo++eQY+X6X8HUc0mmgodQkP3idZtdMznWM5ZsbQwX4ZybJBiPXSISEpV49Ki8
vWkc8cAlI9E2ahqpveYwfFgTfYt0/XlD9zeNY1YoyXif4QxQ+KEZkO5+AtBPHXTt
PLy1Sqc94Q+xT0MIPWICiRRoPZm4FzkqmHfDzZQPcqzwHSvpUCR2dkVK//sgq6lp
JgZorSBg8x1O2uFMbtYYT8B8pFla+e7uzNgaBj+FH6UsnJiwOjPoiBgl+ryhiqKi
gAzAR2XgmulRXyi6XgZnwa4SRWerzckXrtg3eiTEcIdNrAD5kEbmxFAyKejOxUdG
1kDS3t1jJUQEiYjlierI5KAXY9Wvk7VEl0gUC8NOHg7KhINTKlo/uQlBQ4Th8P9/
6M5+fDVMbU4OGnNGlUakVLHNmHST6ClMa8MeAWxGCTNu77SBGQwlu0Vm+7od847S
s0AJ6+FD/oA/a17WmbIlGlYLJKhBGWdO9sDmEwhOGohnDpt72U9+QrHqfGYfztVs
wjM5FnGMVpLzpkeaYp4wEezgyqV6JZdWBuHCR3WLgngOWL6g0YL8sxG3+Bf1yyH6
bEwM7tHr6jQZKtrMyzmxoX4KO5aAv2kEi0iu4gI4xQlK1robMTo7fTdyeBGNGJrp
rXqHOhvJvppvdRAczc5e72wNTS9piILy0hsAeZonUVfwdW6gerUVRZg73MpE/Ai6
RpxxHfj6/iqYjDqUtC2K7Y4JL33ZxW6gMlJjBTQnNhemvUfvhdlh1jDIPzXPOBGC
xWDwyBUTpAqAmbmeF+l2B1ytp07HgXmObqZB6w5R1bR5ei0+5fNwxnXSW+srmsbM
0dfvhVeEKWoCFwMS6G+OkiMVnIfkpH1zZsAGNw1mlzU1VYEaSqrtX5FamxKcM+jc
rLnhyCzo+H3opL6+STkVTFJ++NDqAiLJv1BAjNZMPe3IEk42VVARMkQV1ZGiMg3i
o5nNWsGMtEnAvvPOf45IMim4pl9QK0DBWyM5XDvbhcWlQ4E6aeZ/QTPzuXrs0TeC
mcrLBH47kDuPAhQwsRVAxZ3T/VaZww6DMu4J8pIJJ57pz0by/d8MZS7T1GxAlEtx
PFjX7d70oygEJq3QTos5fOxXRJr3a/mbljnLw/HAAsCkLoMykg3FkKafgY/KrWxy
oZPsNjswqsNw3VZBtEJHk/7qSqZTEHVraAomP406eXvXMy40EQHQGeJSEXa3XMQP
R1Tn5i4DtkuuwKtxzpLdspPV0JlfS5oX7NnQsfBu/xG8H9y+rU8MYyshBo1m8tbc
m0jrNPjSU1EzM+yHbhcGKtpOHUDR9TzyHV83ekEBOdaq6FOLNykvWZcjtH9+kqMo
3mzQnU7H37iKTkK9qAVmtI5hE0aHOnLUFgx8HYpqROPw5OLvnfxkRaFvPFI6e146
uN9EK5yE7WZ4FcblUUpHVd2DZRnnAn+zO5g0Tn9L1JDFz7yl12wN3DSezrV4YIIQ
F4YVeSqIN9pkfzTwImgjlsRVtUiZWMVtrXMtmzHNyrE8k94Oay+EtpBOAxJDKjED
R8YCjhZnGPThE7Y1bunIlx+iVz41A0ZS8SAGJN2x6CQdTcNhN9wKO3rrAMDpx711
TmdGnl27Q7rmev74nRI1geoSSg02iBCkFT/9GWVahRBeQr/bhfYZtMMDuM/iJS5B
v5A8MJV9FKwuf1PgpcwhUZg5DesBilQDh6L2wLPgJva87l58MFudtNDbdqdEi3H7
xbytpfRGO0wrAsa15XkIu4wbK0gytykYacRdmINdRaKSxNgGDnRHkr4f33irdRuN
0gUgMsc4pgCIRd1omsmL+DU7V+JUYWlE/4PHt355o2h8X4cgHfOOgsSxviAPUA8y
QcWUSPaIRuMl7916RT0+ILWOlOkH0v6KCshddBQL1tlXIdfqMIqSQ0h9hOV/8oGR
+All89f6q9wtezR1y5cqv4C05xKdP1yym+lD1LTExaTOnkv+fruoZ1RHcwvkyU87
qyUiT8S9DrUrBwoqbq7QojqG6P9KUoeBXq83hhhLQvEE6KUKmeggx3upUhkz7Ffg
Biqmug/Z1daY5HQD24DR2VzyxGKnfBBKdAkHid8+870OcsANJFgt8RXAWtGJ/2Ik
uE7IhCAyIwEg/vd8HnLhpaC7fgBNlwlbEhwGyDZeG8D6zFPIb9OR6mutnqep7h0r
G2kou10hkqzzREA07xhGm8ZSBlAHGFuHY0jrEah4e3zGASpftGRa9jpZTqsjyAH+
7aip31RPAjflDbmLGIAQtYg/4YeOHxl/lAFaSzUNarqoK7ZplNDIOTiXxDjR7blq
usSRHEQLrOVcz/1hwvgwH+/hB7+RjSvLRo2xEbSA3LOc0lJyhG0ZtZYPJuNpSvJ0
aNrZttg1RKfpQeHeH6WlLPQYOYpyLQawCNDIMmlrUmshv+IEzLrShoyMsLOvAm92
za/ZQ1HoQrve+dzpZ0evS7o1FMVgG9dt3GfTJfiEkJGurospNoi/MK3uGS1NMUA1
1O2yOhtgKTTxRHi2lse8hU1406URnEZVFdkmOJkW//0osQ63Clw1i018KyEmQaTv
+ML7F2p+JQivByElIoz/xTsxmx4y5AUVMl+1UwifMzaicaeiYD8m3UegzGGOC/jO
YfKpptEVhfofoZoF1rBgqBlTw5lSUdqLwqReqC9IPk1f6Ihnb/rcrWYIt7cWSs4N
XhBUOhWHqtgQ/OKZknASyHBED6cx1E/kZYt8yfmY59a9ubG/BjI1FBIhgp8ueO6n
fyqsNYCZtvmE90kkJKk3WnWyt/nurX6O3ghGWxPg4yLLx/4BwLyuMJmFqskBKuYa
ZIW0UhrB1XrDkDdw7/or+4jeBH++6SSLYyIWpZo/KIbUWGw3veEEwbj6h68AQlnF
VamEbJVph8vsyb9uJPLXtQ5uYBtz4M5+d0Vn6OOAXCUjewSx09MUJRCErtO/Daj3
jiREvmpwDWdDUe4ykW4wx2SVvbOkIimsFuX/ucaZZ995Yt0uIlyO4oBeXkxGEXN4
YhDBRu+yY+kj/6uTPMhylaqbENQqrSLzRNw2iBkqGTaghLZTaPPuz0tVNck/1b5v
k8uG9pdYZJvGWmmMGR5XvTbhz6wsBTF+E/v6k9CM3AlIMIBtzn8qSpHYpifNEIWZ
3fkBRaLoBr9osKR5RjlYnmuAfGOkI9+zMCj7BSmzX3zE5ei46LrRx/gaCXVeX1qi
xUmX+Fr/S7JuLYYFCwq6aFMkWkLRnhOxGTNspN31dqnU/gGNqU7o4ZiZywMHTgSY
SahiLLqhcw8Z0RXWx4YvQsZ5BFDlUX9f30trLpNyyTAmNWjXuvXL+bQWUSL7bBk9
TrXrzS5+iBhe/Use9ZS1Il0pviPPq9p3o/vDY9FbMXfsgGL2fbTzT4g4PHJ9egb/
SgdPMm//HaG5e/GAbtbQu6KLHfHKI8aqZTYYhzkVSs5Fjtmx97yPzAwlW5XLxk9b
LnXluTzAYM3vvU3x1JRQXqTLHF379x9KyIx6V+OeOs+f6jr5fMQnqVLN8bEo1gi0
S/E7WjttCUKtQ5W+sBrIJinv7yw1oxFxfbnRV3zB9CbuHu+KJbwd2FVrOFAwNk6a
bbr4Dfwk1venvtyGYD0mICkDJLSDHv3Xp47+ub6gFphplQHJ5IaewGpZMEUwNsGJ
LQD20kRmNA78xYlLLEoim4vF4TLeY7sG5Ky5zZO5sAibCdG3iG7NE0YPOuhR05w3
PtqUi8yx5PW08gRjjQkweVXYGY+DX9S9v1il+870QNF0yW4XcdljFbwj5KQ0yy0y
xf5drZdg+Lh2yyvWi1hSt7sFpoYy/Wf2Ic+0/rClZfnx/zPVXX2BRZo6tqnj08FD
loN0ds37Rfqj0mVoTYP01FO0lpzKxRtsnypeeJ0k60WX7MoqKl2hhLxnfIWbQjFn
SRuD5ItPhLPzpJKqFFDhsCeAVfNDliQc7TfTh5ZBCKZVaAN7kNljoPVf9iN0sHz1
c3e1hXtxINzWggsxr5Rcl1Ma1wj9WY5xcQgdHYy4IXytBFXUTcdcsp3gzEL08AQh
cJuybyFJtF/6jiCJ4XvebRVGC29tR2FrlHyC1/1wu3NB3vPmFR3cIkj2CK6K+DuG
DevsbXsklxiD3Eof4wvkW9Tpp+sC9eLR2YI5+Ph3ope70knLlgoCTrnkAgEQYJvH
5vbuFZKwaeQ0WFb1JVNVQJSGPhcEjuFUaBww0xQ2o2RJ1StQPhr0P7gujMb+GU+G
23rraTmj/v3ra+/UeiNBp+Ew6leXPRcJUiSozfdatE/bvRR9v5CGe77q90QPepPw
j7mZQV47JL3KeVG97FwZbymg5sS3DpAEXIwakfTa3YzazaU05xXwjZsZVKgixQSK
1LGmMpUpzEsLfEZVhRXgfsNK8U2GUoFUTrJH99Z9DxYgTdAkICo2XUPgAeWAy3K7
UGwSqh2gT2537ot4dphL86ORTT3Vz3RXw00I+uyuucYvCDO9mffh5Go6K8iVbkuu
EqQ85rvSEsxg/YyAwZGmPK33faE/VfXt9P1SQLST7m+sF7XAGj8yjKhNUqXGVnks
AxC6MxVEilyzd+F3MIM6p4fWux+XndoLDvwwrrz7DE/5FIj6icPWoOhNlZJSNPTf
S8Fz+yypv2+fzU3L1w3nCg03qAH403GXQIqekQ9y8v2cKTG9ul/9wsDCBzZWm3D2
SrBBYIRgn6VBO/GxrWuRxIDHwjahTuK+omjE9NgLqo6PziCAi6wr/QAKFCqbNfu0
NPfu5o2jlmeO1vTjMh2y2zrvEftGQn/XS/xW57ohVI5DsobwqSn+wkLkLTq60kn4
YnI2C9ML+bUHFyGgrEhifrCAesw+aydOnF781QuwMSEohA9sBWZol3Naj9n8honM
gMw8Gb9yK8x1WpIkdMaVz3Z/KuDMrceHXKQHawbk6faNrzTFeokGL6ILl3edOPLO
+VQnWbDW1qvTwFcg+W5WEP4P3kUtldFTgDHKABCPH5HG0Q5BpC62qlgvaGFwxctL
nIdKttgZjUYvEfkp9c4URI9GFLvznMdtjRwmzje1ZqlP1cK7fpn44A//N2qb4EaB
mmlZc8HkJKbR8tZAwvsuRlWStQlDoCmQ/+duyBtscDi9H/T5DZT+LWVwrZUwJKyb
Z+c7Vk2UrXlOaZ1oHeL3ezbv6NqQTO3cEGHoqh9z76G/EAtlz32aldB7rvqcnOhO
slwb0NboO+/sOm+7UYfWyu2gI2EVAV0C8b8cQsAkOTcv0kQRv4GeTyWs4dNwLWYd
dh/yMA59+EjMJdi+WS5lllJSoL5nCRmwPPB9INXSEK1Ho8/hEJK2rsTRrMRz9s9P
0L5aACzobWyMSXlhACp6xSf2Bwewe+f1t8j+I5uIlctZ0QtXd4zLX1GYkPCjL0DJ
Z23DfofvT58tNlJiWXGldtuFbrSrDOtoaJtUiTT+3u8sAx7pr22PJDeswYtivGj2
0ttcVkaU3Bztevn+euatWcOqBDz+1W4jEE8dm10/SAmQ86Kh8/vHuuwEJxwJm5M3
BhuY7RoEtVZq0mbxfMZY3gKrHq7jJOtd5tAZR9TA0r8z4mhouMx88xy3jpizqWyn
jFtQXs7qTjsiSAQI4h3A6Nqg2i+YqQTz5J/o2x7XmzDnbFBSujYBCBIile+wJNIn
0y5UrUDd7juiAkiOMO+m90EvBq30vas3U8GIejmjvrcik9JcowBmF8AU7PvBY+R9
ME3L2wJvrhHcMErRM21uWsR+SfypKU29ubotvnMoqkx79QADOS/Hp3tVx+vqtdYw
KzNwZgpFIV8MbSpDmwhgrccCNGhSQO07lhmfveeyr27zXF7rO1EnOriBo/w2601+
kiY6SovU77RrOREcNEXH0d5jCENjdSmfXNmOrvmWmd8OMv7SDXQJPZW0jPubSgYK
YMtUrPm8XiyFYawFQCUIDC/hn1724U4F9X7ZUb1po87Kk0jsRXLKAx8+qxxNbf7l
l+ZN5yFLOEzl7AWR+8uJANdGav0u6WUwyinppJ7cDj2P8XwYlzIPZuPajIo+Swf5
O86QybKH71Z1zykkk+Ea7IbR7yMcoHSnOn5lFCYYsriQSN6wTgx6X4o3Clz8hPgq
usUkevVtIuWQHwkBfNuilGTiH9SGg/c2/vjZilfI6JtOtGP1KWGTF+kZuj7SVoOz
f6+x315w2DkSUHzjjI342iYSFhFuNR1wbCGha6uwuBh4sjzIK2uLwA38gMAa9F2i
JvKxRFBJ7jTnlbZ1YBqEKijJFqcKU05UeAHFTek1ABFH5Dx2hy3e5xcbJYn2S2tB
5JNINjYoVneAOqj0QpHcSjoTZV7yObT94zeSnd79lwfZR/Vwl1AhI79h2IsfC3+Z
DXcv50rW5DqSMt+5pvdR0796soIicBBRoqd5ZNfx/V7QDdQ0q8+W98UgBZc9KTI2
q8UwDm4e4ztHrjZl3wNnMkZmA8K7Mo8RPwGW09vkH8xc1gn6BmhPTICllA9TM2aA
/PFbHBzfYrdztil2J3zTc8SqQZtOWGzA+36qhznGvCJpFwu9jyefmc+fX29Hsqym
QhMbfnajIVFHh1pMCU6ifrJa7wuPGWDPhZOF3FOcOYsTaWDG7e4MkW9rqHF41ZjH
ynyFRiMIJJngfpdEokTsx46nIfHx/9qAyRUGRRp+zlwR/orY9lsK7k+zq3k6j/xL
hc2lti3i+yoibQBRuNOMFkqDDIzsP3Dw20wUx/aUDoaUQPsy6W+F9MJvSHBVrDqb
gJBdV9CPtrvdwsz/u8FSnSlsynEBiYZuk6FN0y0RfJPC/awZ44yHJ/pS8JjKHFKB
T2CuNh/y8q8QnJfcb3otDvQEFMiEdUYG8JtGMCm5Jf61hs6CrOu4NnkElsXDtPRk
ewBL+QLk0PQi0KgwkDFnsuZ/V1J1KA1g22HKfTInsUpmDcoXiPRW5Ve41N0qfpGL
SJNH+X3IDpZnllsSdHNEkE7RgIDOyCFjS2b7mfWEidrdGZUPpOkkQoUSn8eP7vXg
B78TiPGlILAY86YJoxI0MVS37enzQczNR89xNGEZq92wSjvZZPaKoYeoGzOyx/zw
+L37bg9e7bKh2P29FYzEYprskOReifCxqkudIqeYdPRgc0mui4iWDR9q4Ft9FrAh
AgeMu7KQRq/cyPQhJ3feyqYziWU8xwhBI0L2wHeNcvH71M4kDpUmIEr5PRtK0//P
Z1H8P3LVQ2msRz7z35RpxT7hLnz7b9gHIv83oRP1ykXbYOcFCGgheJzF1+x85MKH
8pyhRU7Pqsa01wHiLk7xYlC8lP80GPTmpx6OFV1kfzVT18vV+sTQ063V9wW6/yYl
TuYZ9jzHAGe1XAzd0m+GdUlG9+lZN84sYAZBsebcLIHbTeRuHPQ49zw169Vt/uJG
xQOsvB9zEZWamxDKRGIif13ad3OYVpzKKJ8jNpNYOFExPVyFm/OGvQaQdTJo8zEc
ID34v7H9qj/lxcckwiUGkWUtIyV3ToAtmKE9a+IONAenvP+6hxdmq9WSnDd1kbW2
p4yucQVtZgyNfqJTP7Kf7gCwRnyxCAp8XIGmMNtjWwuEvI4Hdeoak/mkwgdZfHhO
r68pbpF9uc//x+nkXstssL4cBdRTwy9UH5NMxl+E/YKyEmrxhGijlvfXGaGWQ9X9
n5VQ/i81rHgeaxSeyHoJmfFQnoibD62hY3JCCwqbswosJbLXEB4Q/Skuda4Q16WA
SZdG8CNDNnfGhK6pAIzssbkeZlcg/I9NBmNa1oZq6jmLUPwh3882aMmcbWbymR7D
RII1OyjfHyPH9A79y5oyWR1qQfHx4d6FSptaRexTTXuxk6YuG7yfqnxCGYlDYpZQ
waEJpV+KzgyNMFsu1I+HCKHOTAEGJMwdnISwIA1OKnn6OOC6/tsGPiV2aByrpcGY
r7hByZQTSY3TqWEnytXorQ82StQeWHJY3q5bUfH95TMqjJXx2AMeQ8grRiHhko2x
r7AI/n9PQjB9JOzpXrNm3b5J2tThGn1Djt7MiVXQ+x3oX417w+EK5sbV5TT5+A/C
uqEtMmk+NPvcsJGyiPvoK/JmDX0VvgeL2haHzAEOFcTYk4J4BrKXQlML1tupKATk
ed6Xqs9V9WOtJCASWA0CtX47os/mbzGjczW0RDX9a2X2Aaa36UY6Kw5zpyenhjar
Ykc4/N+KESEqIiPLpcZgyUXIGSFVCGtID/lUel06O5868yox/1ZxLS9fYtBsQAxf
agwslFdGjly+RACyDfxMXq8hldxpQ+sKN/nIKTaLMb5/f39BB02AQm9Z3jN0BYxC
+B+rBe1da66vwiLxoIY6g/eKbAmyvURtLymd2+L10FVjQBok/PB5hNsKrkk4kpQA
U6Y+xRebf0i33SiLklAQiSWVp88OQx0NPnjx8bPMGy03QoL2gNJ6deuhJ4H55qrh
e5YaoYSqLwrTyTbyC45Jqsfw44Dg2Aeg6U5tyAJRxb3s8xL1+Hg/6xjslQKkLTia
GYYQAd/iKswv5YFIGpkKFpSYzdqESAFFvYMSk1XVsLaD0oZt2BUO4Wm9yKJuhtqn
60O5gXk6mcBrMYGkKayPRI7552m7FRjL73jY45F8jeLhmq0SVpH6V92fQexF8SPC
rcSl/FVg7OR8pwy+g7FuCFFQYEV70BPUnxJ8nUNPqw45MTiWayDkJr2CAmyaIeg8
o3CIbEJhQewvmjFYiDLh+SCWhdGa+DNWmwBRE6IQxYN3R+4hVs6JS06boMiyhiS+
fC328eyJctil+JwcxiXvo10CRYS9O4n5JUweK0Kd69A2pqXJfoMQXXcs+6JQz0Vt
GmwFHx3vxBhUo4Ke/CVWvotakPcqbZ7ECgGOaUbSM/aYC71x+8rFrviMSLcpxSdZ
2O7m/nsVsBpjGV9IhOVya6Dmvx78dpuzI/XqCilG9NE/IQjSwtELmeQZVqfYsHZj
KxMR5Zs/u7EGPyXWSwXVxGSbqXGPfp5Q6ZjRgG6PYZs5r2ytpoI805HYx1L9QLly
zxJNQmTj2cj1UrJez1RsthTfJUavY8GlON01rqpQTaJ49jioXqo5RBY8PU3Ucbq0
qA/376Z6j3McguX5aTpKGD07zxJsN5BA4D/f4ZPn1BEDsSGYUb5NrqmA3dHpU2e1
3TJFYdNpb6ayqKYJPT/75mLOuPkuD4t9uWUW2UU28lg1xxGi3Jh3zmtQ0D9JTFdx
72uasareFzKnn7CQzBd+Cu4NI3gGK4tkjLcHzugnDsc88OaSPwvyydTQvIjW6GJP
BIxcGI8cAsqB17Ob+ANJZ8JjyrHn+3/VbfyyuaqbuYXXyNZJ9Apcvz39XBNkLDJV
elLCmn4GDcLR+7h4swjwjVi0D9gzHvLolPJCglcMjh4SNUtNDExIqYj/Gt22aq//
05ZEWWOtjJ3jl5u/Z1MTIgMtUx5RqYpNX/gsOc2tHj0dvss/yxjd7cZp8k3YvM/B
BE7aph3At2jwSAYAWtI//6/nJD9wnSGqxcRRAccWbafMr+6cx8JtmHGoOWOeE8jd
9kEZ6xSrRJD3GD1hybLkx9MWCzkFXn/zA/863leaa0Wd0UeHd38FUe+NMqyEBb4H
qVLdehA0q4DA0x9Uoj6nm/4eDcMZhVgoCOgJFo0L2dfAMz/qjvLVnAcEdJVVvxyw
9qg5XkksVKLtiR8ALvBNU0KdndpNfKHGdfZQuRdvKu5h73KxfKSFTbOIroKhdVwd
JNvY9uvchfj5oww2ZsBDS/A1z2sxoIYWKovc5jEB1i3egpaAP+hux6axwQ7JPGnh
NckHW98Y5XexUrEoH2341ZQgZnJgKKtduq8cW3mF3NBXAq4ejST6VgZwVGv17wOx
B25ehfGkGtbq7mJBSZkdVa0R01yeEA14wRe3Ch0V17yr5eC/W+nS47HsuooAwPEH
IC2uHo7T5OZrSEwL8FMsYwGqdq6/LdKq6M6nbiBTRNP1mHgoFgt8IRbOyWnvMSbd
tZDAg8ikNbHg+VHDPBWC4e+RgtTSjutlfd4/cNd/vZk3/oYKmOcqoSjh6pggOciJ
ibuBFrgAnj6XoauP61WcAws6+um+OSHotVB6fAuGD6ZtyTzD9OsNHMcWkcuqGHdV
zyxj7KRSfU6UUalQj2bj+dF3PCZfRuLgeTDqT0LY8aaiR7QMPVf0dLQQEfdJCNFc
zI+VFBI4X6uj5L2oku3luPjjlN1HkCzJar1DoitdxD+/yKv8eGH9LD7c5jBDrIPC
KTT+dblqdoYFJA4JWni5u6e5mOnmxU4rWa6Y8WEMU7natRGCpvVBtPrkJVNHAs60
5E3QSn6poaebCjHTIEB25sJwV6vxS4DL+l8HShnD2nMfeHyRBRN0qZMbWykK0/Pj
gFvWK6O5ibhoUYwTepRvccBeNpSFcgv7yNMT4d9aWGN3Puddxj5zUXMoHm4CgNDY
UebM23veA0DKh3PGj7feFpTVkgEkzy9iJoiGUy4l7iRVxc6qZPebZ4viCs3YtEfY
6G/RLM0qNiQQrmk32rATeYC3ETHtU4D1O6D2po0l1Jri12dIjrF5c+8jtS91+ysS
xJDiSnIMT7zs+TswGv+1nhb2AJbjFJ9XuEIz+fqCaeyuBKcQyFLzqwTIZUDr7XuD
Y6WDKHT8tZXYLnvNPIXAQQRuwKp6XF6i9a6MOcdzdCFQ29GztvFk49nZHbthN75m
kbLbl24JInh/f/kbeZGorjDYEoLhVi5YD5jxvgHyUTzZvTYeWBXeSCDF3ro06sA+
E9JRLmzaeaeY0sIWFjbAjLLsGR7yGwC96vdjK4kCITfmFf0MvNikBFQ7bF+2dBLr
B0arw6XOI7kLDkxIYRW/JFuMEtdTS5HKIyLxv37M1ve6R6OOTYbuoMR37hEfipGc
FEgp3dVi23QDg6i/sjHZ3eDahYT3vsPBkdtMo2yWVn7rYrKbIv/4C/JJ0kcGvmp6
iQyudccns2BU0HTQTo/1vPSDvKb2v7ZAbJNqip7cd+Jl+Js8nUguCQXnWl/TMN7b
DpY/sUH5z6xA5jhL1b3e0hLL+9D6tYdbItKySuAFw70ktcTpmc19WOsBNOE6GnQc
mLMQAjBmg4SWqHue8xHYUbpD2FDYbAiis2ORqQfJkZI9o1QVCDhCWX2yklVODXm9
Nc23VwRkdchrvPyNm9sHPYdeGX6yl7ABqdj84G14oLoA1qFl7yVf3caqpHTkmrOk
ATC+uH3R0i553BTs+/yZ/iyR1R8Ij8mMnMI/YWHHveeeVlrLuyHE9oyFm/YdYR8K
NdeZRMyztiYKfGvf1ZLLM46CWM6+ajp/O6h7RiiKMcJ7GtQ4lXy1r24ufAG++XO7
Wfcgqmcl5Vb+VaAgwHzbZvULa3rk6oAS8fwlogRgvYhcPqFJXRlHhs1Uwo1Qmjvd
35E/Vnj+h9ipmOhWyusU8ttBUN9YsBHhvRjhVBbk0opkE0XyP4558uOEZdhuiC4I
kWMm8d6RRANzT2RNV2W3m8Isz1ib2nxAswnB7V/V58g/9ri3dhX4b9X91cG2qMLT
g8MjFv1TeZn+wXlNNX/M13PtGWM7SF29vjrDgbK8lnL23QNh1XK+cjhNQf9tATrB
hbVHzLgdeTEf0zFICsKVFQjE1EF+rnIp8zqIvp23WcuEjFlgu2X0dxeVDNtN577L
ZZFRULOg/O596o5yoOPxrdzQvbEIn+imcwwWiQzysJCHX2/HZgjzSGhifDruiYEF
qQkPBBmT30KpPAtOAyXqPs3hEWgkVB7Q7+jXps1hAeN8gqd6bG21aLB6wr1Budjz
6squZua2LgNTuxEWMaJc7NUZ60Xmoj3w2ztLx9yldlFGtRpsKyz18Lz3hlnLaSoX
e8V1cGrNFmYiRIsfxSwUAhHp3/VgzQVRq1Z3DBFaWAjGVahHbcmG7FqFczNpm+er
CpJ6LrTh+yM7Z4nmpxmVm3S0WWJDbZVPonqsfHD766XCmV8on9sWPKKpq8JSK3h1
S1Q4hVQHgTCp3IQuQXXEMAAaHU3Ief2kAB5gC5DqnPLi0jQbgNBalxmPnKoniCN2
cdWsJtB60WPx3i6IKNuMBhCkDYi9D4VtrnHDwit3AiTrvbiaKK5wS14H1QSt0csg
aDW4VlMfRZ4O4GSXI2gsQNVR0xXP+BZ2AAcYzHuWpocCy0148+aC7MhXx7v2YibU
k/efPj/+9l0NnUUAkAtX0+8wvoVvuJkbiswCaSYNF1sJvoC9O7F51bnha+NGFlj9
dboKQOZBhPLBvImBF9XmOUMS+yFvKw5KXe2DB80NQvnavqy6kGBJ0LbVZLPjBN6H
4E29o4nxDZWa4hyfoI2mgwFP3NieUz0QkzLy0AhsXK9mrRHNm7uCyyv35l/gbKna
uArHrsS8cfNV0ueFuCcDiNackDf/Ef/Uo1+caVZE3ZE/gjc7Rb0vFYkkkJqdOnNH
NS7MYHHbq4PGtHA63ESFzTEYknzowLUO/z8QgYOJhByjbXVfqK7o5KpAHTtQaCPZ
RgtXIxaCxhQTVmxz3gzWU16y7F7l3D8PogM7noUtPkU2zlaUUXDImOEQA/Rdu9fH
J3pQ+g1dTeDnRRYxfhIDbECZVlU6/lR9fbVhXlU4UPPwWNHAPq5gnC6VVw1iky7v
LmS0/z3fx0PRcL4fPcgo0UdKC+hGsd0swhdIqlwbQS7fGF3rYDT6J0P201Zrfx45
lZJFVUxDGU599OU8bydTDhqKGtLEUKg45AgSERvV/l2ew3kQi28exX2LOupmstVw
PuArPFjGAA8KZRyZb+pDgozJOnXrbPzu9IrGv1aHP9zC48F8vrEik2ldDGExjXk5
UlIw1K2890rQww0w6Mch0YmDczSIWDo37rlLfJXMKEFSXAJINbgD3WmW9Ul+ilDy
T4OWt71NJiCEJFKUI2C5Gc0hrKwdbXddRMwYOc0fsDV3kFANPkSBp8jRkONu5R1F
C2Fg9djl1gRnAIcKOpNJQPkKRn2ZAqAsSQ5GT7qGrYN3HwbyCCv8LJhqvpiqCS4I
D0JUN2uj/Z3U4GJNNJJj60EkG80NTSVj+dTmmK7/S2drvdrNUVrjWQcbCLYnrROG
7W5hWdDOdBsappa5R0940dbOrSHGuAgedQd6gK6E98BGGhTV/wG85fe2ir9Ccddy
K4KSF0w6dV14R1g/eB+WQSWSEbv7t62yKhPBrsH2k7ywxIgpxW0ey6A61UtxvgNW
rYltFgZokXJ9hr0+J2OndWGDvGPn/M4ieP3UoOucZ8A+ObUG6PwZRO6MkxyMBM5v
yW5figb4lmpb9RLKkeWct5L3moNsuTEd9F13mn7F5H+YD2Cz//wWCIrY3sJ0DeC3
r2dz6TaZYRCwGe1bLXNduG7z/2xlEtLa1WRVKYaYlYHFbVCOEsTne0fawmlZujv9
7/rStphtbyDYPx0h+qaji6oaidWlVjKky4hV351uDWFNmvJjqSSiHmVQX3eNRHFv
QhJkWvSVDDSBaQBYb8yULxqoKHZ9jWdjA6WzlXaamTH8cR7BpewzL4naB8nP75o+
gd0g+NUGIXmRV2NLX8/BQbujUQ4N9FhBm/ib5SAD3hYkHmJ2NuF3fs352BW/mze9
x325UPwhXniHq8nSg5iD+N182D/xsc+1HbvjsGV8NSfNJE9gKsD3FaWIj4VqQAJc
JjLWu7PBjANkdKhSYtoA2x3EW42gUqowYdQaIHWf7aLMGmcfIYq5t2eHJ2cp+tL7
kJ3bA3S3Y14tWongVtSEFxKU8LJoGb5NnlHZKCVZxK7an6W6IZx4ZPtVNxiF9Ywf
OOxbSe4kNCqJxNdTbTJ6RnyHgxrO7DibCcO0J4IDZ9BBuXGRkHRGfBDmfCFVQ0Z1
jIr2cfWc6HP9kdt1MMTKI3kzOTh6KUeo38dAGbaXtE7Hx95KEW2t95+dobV6UyNh
GrTCevMLjk2znk4SHez3+aiDK0dEL6HyGFUQOBSuhy60i1b6Dx2JURLM+MvwQMMB
pnlWv2XN60mTzIvjlnMNxE4uUscngyreill6dDyE9xuGHsG1oB+1ZXK1/JO0biP6
yLCOO6MC/lj2/3wdrp8gGnCZvOvSQGrvac2Fy4Ep67/yAYibP+GB92Srpag+mhu9
vk6FUNQSUOjPDwHBRZn0aOMnl1NwOiGA+cAAe+JKm+B6DZ4E6bAn31evpKA7gXEp
oKDYlALEboEh6f1HvTJXgQ3+7BRrCMLxJ2jjqiwPBWi4YoHqm1I0raYLs0i7qzDu
Af9U52irUP6B4VM2Ztx+PveZJQ2rVMtyjdTsRNL/TeWjdwqUCQI97wymnQU82esi
aMWJ8XDYWejd++VkrGGjnj8snX8NCHssCn079n6rRg27Ej1VgRtjynPM3xnSky2t
0u+415yq0SvjDnrHO348Q2I/beCabYxjh+3X63GEpI9VNsOYz7SZXI7F0Wbwb0Kx
IbdPeP4FF54PF6bQlZQNCT5b2ViHOWViIuafWP2JBKssFIAJrO7+IPaPOyx8KLK3
4p1T0+sNFi5syR9bfkLEWZtX6a5VXKta+r5OkvOYwlWJJZba+46SAv5VB3xF2Va1
RC/7nUb/nICpFyjVZnLcvL0xiOdmr9g4GFNS1tO+rVv2l5CeoyRh+R68EClN/qoI
9PSh9NXJRws4wO0/QfHiUAXWkuU5B2euACXe5Zgi8Vw06R/9UmOC1EsPT82Wun9h
0H6nCg2d1m07+j+aApwg9LWqbrBfAtKZn3beR2pbzTU72k7j5Tpe55tRRLQKQjMv
2d+YmJJh8K+BuAxPpAfgpvCGiRd55OjVX5/QwTHMXIXIS58NCBQ9Hc4WI58OaCzm
XixmkX/kcKajRJ2gXQm6une91gon1wTVYGpcCHp15I7BBtMrq8B2HQTNxZG7UqEQ
uRZTabcR7Q85tDtr0sWSXHpawx94FzCUEV/DNobGRN0JcYvY7Gj4RqCVRhYgW7z3
jJKy8HJ53MRbdwNptujmOfempBoXTO387Dzfl46CEPVrla4KuRdq5w+leT1/umuV
31QcGOCHCni07veL3TlDOu+Rqz1PHkUiowwJQ4A7hmbDMbFjT2GABacBoD4ZQ3Nb
3ffsUAv+/eQMLYRwhZdZhyGo/iwnRD2kJVK31i2og/XbWb7ebOOzCBP9jFlQ5zsH
iK2KL1675J5kShhDvK7thga0FxcHrAysKSyN99XJjUlBPzHfm98/oMu1SdeP3nSH
H6msV5xpomtLpEyQpwR6JH1DBLfZVHiDDEblAZ4kQm4otYZL/EXGwQIosFeFYF+b
9YHMC6QJ1O9Q5/YIlpJotmkjH/YNWgfujdaVV6eQ0FOCBmC7+TVJV5SgxkLSZPue
sqm9M3CN1qYxDrd5/aB08T274XjICenZqooZ5s6/dpOgM/rytNriv+u4os1amCNk
OH4YgRvNZp6LwjUiF/eJyJzFCUbTT+IZszWkjqFF6iXAEimtHE90rTble/zOdqCD
r+C/8PxwoOSiTdLo16RCnMDVPCLBGwOxZqkj5t26nJkvQLlQTIWYOIkKFvtdhsSv
16ztIAKWl7fF+OzwEVi0On8m+FT+3AdhDrr+vvLkcbtyyD/Fhrk+83YYn9OBYAZc
brVm3X/6X/cxINWPBXoNmJsWd/SKsrwBqEBvdys+tHTEgN01iA+lnf4ykLS+fX/w
WFwMgOOgMIXFSlN671x35aXdR28gmmQnhKSFvL3/vd9fTehbZD5ryBbfSV6bkwrs
HSVQ0Z2r+pd4KXqCY+OZ4/ib3i0F1TOzDgtqNIKAvU2itxJpImfST/AUoiEKGUSi
req8v6GXAs0sz55BIfq+fmAkRbEpHZCFwmkUk+/fc91dijb61aK39rFaLW1xGJhS
Cuf2xxxeXTw72LqkmLZfZiP1rPGqb7D9MDRdrlMBTQms5KgHrLtugJTLHLGWA6tP
/IpRFeGvJ5a2/+mtYLhB4L4flk8C8o3Aq4K6Nim3KkoIvuzo6zJJSBtVz4G+fIDx
4ROAjPYYUmjCR/JchIRT4cwnd759vOwqfAAJQW/TZC3pVZkLuF+Yqd81yYuKca64
mBiSPTJOGTisFKnIqpDxcX6BAO/Sga3cHfzWn8t9VzyL5xqLNsPbLnFyYQk08Pbm
O2RDJVaSUXFHDK1zTgNpMmlkGvzPSniwZNhQTXXKjp+dMXa3tSMzKUNe6XNUahKV
BkPzJ94gwbw0extgkrtUfBo65qRvbeYgvZcBB35ymFW3LC9cmvL2pQJXV/C2W0kh
B7CAGyujyYGTegS2ZXDN7FkIYvDOEGBdCsF6Cs9gmaIJfi1yIk82iOMzHZ5DRbyG
3yHICZHNuYOG6ky2klCylqW0fARluMFHdFb9mrPSryYhCXZLshjFB5oZq8tfdoNz
8AjTiejBW7unQ3XH8cfCaKw8xg/6Am0P+sFJLNlc7YaA9z0a4XBLb3HSpMot3p3j
nD1frj2M5SXBVyJd8lBDUWECr7rah4632d3lN4bOV1u4bsvE2E/4a7m+IjpE2gvy
5JnBa66A6wNcKdr+XkJYyt46SJEor1Y9ykhVTfKWqdN8GXJEdU/7JSwNIl3kOIrU
KJVpXmAVKr0oTMBXzYMgUg9UODwGHT5MTu1azg8uXTjH2/RVT/T/T93Z5anTMttD
sH0NPPoYGfiEy6aWLE3dBrx6GjWX77fuV5njOAdXxWtf3idajesXo/dqi4pISdv2
/VA4sgdFlCFhFYfdUwHh3zUhcMJYmhM1gabb9/Sxf6nelyLUe9lLBxSSl1eXK8wo
ZU5febzTzNNXtc017GyGqnf5w8Cc3Cd4fi0YeQyuu55jfi8cGfVA+i3lXuGmqRb1
qoX3iiW/xX0IDAAcuqUfDU61r2WdwPLd0cwYZuwK9fL5OC3bxJHfbDSnMYoeaaeI
ZVbyfXbGq3Nc6ueBFIiOT1YLHQHSjNHwc7rPp3F5FuTQm7ALAbFv10jopLrSknN7
oFGSL8XQRnGfXhd09IGA0M5yDU2mgs2cUAQzAxwFRid4ByEiviPtqn9wC6rdsyKJ
OJUxEp2uJnjqHWZ9p+SF2FgLjTQrdWViHW0l+h8CdzjIeOmbm1uXyEZi0kPfIKJ0
AI3QwHdEa91dJjRm41ZeUzkYbB8Nm1gQ6AFSSPLgplsGLJSb4MLcRLRsqHo07Kv/
k65is5QDyd0srPjdm8/C27oAsxPBnSru47edgUU4QjbgBjsjwSz6jZIbaOlLFfsE
cli5gvHW2AD8/iLsQYA42qDlNZ7T/6lSPFc/g1JeLSvyZ+b8oZ9qbcKotjiIPBCh
zry/m62K+K4oEpfzepTWKTUfMKwBHHl/N2DRU28XBnZmw38ahyVEgLsCU4/Rd3xS
Ys9qgRXMPNs4p/IBeuMolRYtxwYhGWsKXeGf1zpYL3BCd7azyaYG7QFGHdnRTyrV
jb8VLeGohxyM9SON22UB7ggFtIwa8N8oaXTmsAuXpyS1iFMK3HOIJhSiN8kSFPbz
s2+bNoqslmXNAEm90FvqLJn4diw2N9UNktHbCJWdohqlbHsgT2V2gUR803NCzymK
mpVhnO5ZfJ3stkk9g0YNQaJM2M3v4X2DmuWEFWlhSDEL72DgtBnh3K5XadKFCkgj
KPR+ug5KKN6FNRgoKaipVvnMFi1+PZE2bYYc05vuOuIq+etOSYNiAqcElec5bO+b
762D5lDGvPa7cX21vwLwNVAOgr8iU7l19cXhU0PCOtkcmz4MLpbz2aM9NtW0LiG2
HyUQIvecdszwRuczpa9TQ3sFEwA4j/mtpEHBdQB30bI59n02z0QtYLwKK96DWy/n
76of2gghXI2wCUMk95MNlXFX5qBMGVpUiPcIeni7Ne/qq9QtTDhZbChbqNtSQnKp
AA0dIgenjwy1Bk6GmaJtC9RohoGrzWQQYpyBbaKzGH+W8d63IwJIAi8VXIAXjHKr
zey8ZoPj8fTIEuwOm5GrasBJxr4kFXsgzvbPvIOJdjxaG+ZsQ/rVqYlAI+6jzGMP
N1pv2HgS03AOTD151p7UoubghbQjZQJzl2rag1jVPqNWlWbo3luj8buofEvwxFKB
860x2ZWG5BTYPjB5d4yobsETIe34AxyIMV9Da8mryfIQ1TmRWDO14PKDBYZsLxHC
J5pmfwmojpj8BSSSftSbmScKD3RnH/0nctbjfOcWkWCljeEhM1IGZ6VWm2GTcT3h
6SrGeEgZLlRGZEumIgGBLJL28CPBIt1Xw8ujIdLMOgUen+CPJmf55MFQPyGrFsbE
O8h64mGDX34OowiEnCh7k6ggC6kz6Bm5y2JhhWccvm71kaFYJx6Ygf3RsInsQ0aD
ZIfCbLOPPc1/jYG/Qv8VBJAT1Cky8A27J4VvckudGzQnKLAdoHPvNWORTMeYz902
d7kHNoZ65rH8ezrESxR5lj6XyGA4eJTH6Eav13CXrDq+kMZMvWR4v5U4vWZlJCQE
1HI8FpXkhRa6rgVWq1fotVZk/XVFoZHmFj65iiDwKrY9/CeLzVQ0C2gI46WHpIkg
mKdH4y9b/rwMhatPz8IEn7gtYWocIl0MW7/Wj2wEiXYs4SCSwkcAkB5GIgMr7ed6
2w/GDOsgfh94r8ilBgpIxl1eeiZRPrGc3spCOZB2E1s8kkNlm0Uy37XJKZISz9Sr
ooBvi5+JAuZLzCn3s0vie2WhPpJ7qfvbEsAAD3exKaDeekUEOllCxhiVKW2SgR84
rQvYCQCmPFwhLEMt6fYATZzasDqu3XbytVaqfj9al7rA31p2vE5zWaaZn62WIFIm
IZzm+tPXhvCjoKxvv/3YPodl1JzXwcNRflMhxfyFjq849g6yCFnBLlAbOFhFRVIo
Rle5AMs7Hyk/CTircdqn6l36y0ekR1i+cMMNF3R1OPJFiomwVBT+RqOrgG+CD6Mb
2JzM1XczjTqHOaAxmJ8J2IvxypbdFJqIdSRvs3ivV+iU39xnoeAeu+SRqV58FuIs
jnnsjnPnqqU2deGbyJqnoYhZNmD/T2tcKDG3GYI9PUXQos4txL8fai1BeoKB2hmD
cbdAVeMvyQDJmwHMUq7xNgZkGQDQMIku5h4wVL2nODiLNgeg7AWYiOxypILpqacE
VdxXYBethHPVHGgwbLV/hnXk1jq/bng+iy9XNxqpiqOGXJ+Q7uQ+Kdm2GpbZQGoR
+unRH1C/8Dgu9+F6j3HMDO6KCJ8w2pWKY6hsFsk3k8xHhhKYGfufRxu3s62Xuclg
1U9ESpSObAgCzb4vf/XwxZK175tzsy4bpaTY3nPbc+nRRTpSqaCstG0p/LIUDHC6
lePj2IiYe8GbJz1FbxNs0bY5fKxtxz5u+VKSdu02Ccgctvj+dRaHcMP/2fxDgkhc
QlrIBf7Rqyesyg0Bo/HjW5wVA88wuHvfCP5E2fum7cODVaM0KfbUhVu20vKwDWHC
rQcd5d0gi2hSTFHMymf1bi6nADN/dzzhHEkEt9plP4mWX3C8meJnhACXz+NrZaDl
sjlOWRwFGbI4zmoPQHProiDovKNyi/Iw8LbuaFTRgQxSX9CNQ2Mf8JZAA5MPyQwZ
6HZTaBoRn2L77/1H7gFeLHTKJ4KAg+RXfPp5G1uYN6CqkBR5bqCefunTJpgVJVCs
PGrg8jFGcHwgEQ67p3wk4FxGQPDB1Ya44I923aOJ/uoAHq1h2pKJkdMdFSw88Dnq
pPi+uHlSLQG4eGBRM7lzJS72Up/k5k0h/yuB3itK/QZhA1M199DdslmOpUEtOs1E
D3olClsC3+w4Mkc/E8ow9yjcC1mju7gOzZU8YTBfT0n3pvQLr+oB8tnUE8+B73zp
XxHtsQgS4k5N1fTYR/kaXn0jfZHmsye/oQR38/J4eL0MQBF+t/8h/gHV5LqSBz7n
ZRuKvggIurJu89MOZstT6v/iQCIqNNgGyWM+ZaN5ax9Y+rOEwDWmP/0XBaW6BYgf
QA9p+gvs7deFSHlf9s/XtXx5NN7L7YLU41AB7O0pkH/rCkE75ejmtTyAyZ487N4Z
MR+FU3oiqGTh0wPOtRmjOSNteQuZleYWFrrfN4XZmh2q5yZSYGKZJP8YAs1YIPle
c54D5lkMdvclzetP7ocMkpKVRicP+zHLE3ctY6ryA2gdwYDLVNujH1dMzeyy2wLI
RHKT5ScSqjvZEQW/H9nankWIhjaNcbOUR8p5d7poUuTultP8dBZYwiSexFrcLJhE
jUW1mHkUN7Z0FokpxFSB6yA5xUOF+jGCBJgOCbZicstqbBv2Sae89nXagTz+M2Ay
yrMPWMIF8gpDpEYMYtQgoQ05Sp8mZuTbo4eIOWcRy8hXZVQfX7zQfefljziIRrkk
TtBnBLeg2W7djE9dLYmPUHgPjjuTdt035uEClBQkuQhraPNaGg2xFA2b3snwLS+p
f24g4WMeEjA4gyO6fMNjc7CRh14VZ+LFIjOkE1lJEGVXJRkzdWjWUMag9wSiD8Og
yNo0SmYsdnjikduyZudHL7aofBnAlTEche6GQP/tzrt4cKEC3e4aSzOUUIocREGu
XCGRZYjaVYguxk68SUCTgDyd9EXvjDb4UQxGPd4KPdtoN5rV5zomT+tYzuEmgQRj
cDiqetSHiJ8cHIiju+NAn26jxYLEt11NaTWjJJOnGUQtmj34sfmFc0v6ASdO008H
e0jgQyKv/pJ9yx/NptOdAL/1CVXUwnz7awW1O37OJPaRh/7aCF6ilGOpJoC59aj/
LvXOtp0hx60ntyAvQkYiI+aE8cTbraPxtrcyTNjAIqWLmENoYRM0pE3hUc8Vb+rU
dGxPjX3bTFrOzp6oSJeFWj0XE2NYqMHyLCneGnwijGaZN7+OrK5puDqT4T1N6tZc
+hTjPJ3J5kEm9wBN0Vrk1EMMypc64X5+AoYvSUxYozaWG0D1cDKV99zDnfjQ3rcn
6RRRvG7KsnWSmnT3sj24yvHw8N7uSFxEwIwmihfZOZioJL52hH/BqLQ1i0asYa4C
nNJSv5jTx65sjV1TMaVBhqLixBZiLFOIZ6PrOvoRbM8LfhzP7mLcLfOaStR1M6Xd
L3imhrctGTAlMiaCm3vdC7oZlMurXp85ipEekr6P0Ap0id5cAgSd4sEaJ/2aOYX1
alsE26Yo0z+nvmO7pZA5Sk3hQa9CR/uTFeykNrxpn2g803hC5Eh8UXlH519s3O2f
u9pzFx2kcJPoYufIz+lAOucYaADWv/SJc1maGJ5C2SHjUZu6h8X8QzIRhzOGKmID
0E5tQZJYTyrl0YSLCn3nnxEjlbjcxq++fnMaB6VfEfshYf9qILPZwyThOOvzWSOa
m59lUxOLcyXs1ipRTO6wVzdbVjiULUyK6Tp0jUPVuyP4R+kKaZNDPcM0yOWYwkLV
G8fUcYDgvvWfFk9SlQTYOJxbZIwZ8WYaE6ZxKONvHz72h3J/LPaS3aB0tDEP7twt
8GquU4SgE+dY1WFU+6BjYrKqhIa2zfo07yxWkbUlu7XK/0LbeBWef2MMaOc2XfsL
toTAl2GGoNwFDpBTM/RkqKI0miom7NZBhymZgF8SRLPiRLNr0fPgf67WvZ4lgtQ4
l1q26DBpYb+c/8CuSPpBSshkwOyosd094dA00O1YrY1v2zDJsWUkn7t17+NU0ewH
zQWC6XKbnPxzGEVREsBx03n73kfhfdF8PAyRDTOlL8VOUv1jy4rh9HhIPG0W+KRe
c+TTt1D3eDTNAJwlgj4lq4tPmXt7wMxTpfWCP2mCltVZnnbcnxOtelFRWY5N9GHw
nbSG/BUMZ2rLtt8af+pZR16AgxQEGW7y+5usubZ/6GqSZu6nXS1RQVldHkZU/njQ
R26Bz7JNrICXXWPe3MpCHtTbNEjmZPN2K1Q+uOmO8HwNEBZkA4pLOqpW0KiCKcWl
8iBO58MoTOKcvzxi79ffcgRw7kqSZl0pZykdtPDcRlijo1PVpINUt+QmOStPdm+O
wANExSbdRUr6A5RfrOSasTJryIBapOKfQkwi+wRV5s8yb1KrAeMSb3u8dIAozfZd
QfyUcmKKZvQVElhkMcsQ26WYDdOYwBAHFpwmH1+ARW6cxLpNJoa0u/x4WZKlTCHF
U/Iqayv0NTpUiaVuw9mZwRy8XP16ofdl6Lu7szB0so0SHe5WS4U78qT51p4hv1iH
zV08FfEF8PpbS2yUFJrudZ9vDOIEFJyhbZPM7LyxBlsaydIdgqiDnvd8RDHDXPLK
JlYCkI70mZwUueh/dnbYV/biTDCDkTnp25Rp8lRXK7u3pQbpWy5rzoDskzYlqVEL
arrK6QUEQ4D8kk/ym9B0gYHmZ/jGv4qSClbR1NXdDGiftPAgaJLbZ87wlV9GgwPM
6hgPWKZ17wEBvYmiw6p/EuKemrsGbSm8aN61RQQCGTz43dUgEvoJfIjsHuLXKHXB
9NHLhtCFNTlgqT3sYybdIVRzkNUY6TEF1cEhRM4xnKTQ2sl+LgbxfMvuwY/HT9+n
+5kkYkIeKGBa1H0c+P8VF1nUTmVyCKofoI11EmqupM/ntwh9i28hj7P+SyhR7y4m
312Jgqt/7Go2COxsza27rZTaZ7lKNbY/tUaZ1Gw1nq09NEyyiRi0KByb60U4cYyO
QEnd0gzqWvsHCkqX1pLgcIur2FGt8sXWSODbgLVm+1RolK1/gQ0nUdCzx7LribTU
voFECoWxZyAIXgcD8ONE/PwG0gHHeiecNFFJcHCCGm/8SIZaZUCrkbdAQhAAOZ3g
lKRpieGTM4hnvukyBlr4PDDAJzSxj8DfO1gRcmTJ+fo4MpECmxqYfSQe6jxyzTnn
CI0H6UhbmlDNP7zD0jUG8TQcs0eotQsPsc8Gq2AovLwvlLgsB4ZpA7q4rEZUAC25
7cmpjAxCMLm0XN8ZS2ZxOPFG0odKW+5V0HHaD+dTAJTcvjRQ7PiPkvfyM9jwl76y
KcYZtXNM3xKNwyy/hprW3K3VLLC/HPjEh0CfZJtX6KDaQ6A6A+Fv10XVQgAEqoG4
jZb5kY5rkxvl1zg3UvE+Ei/cEo0I5XBjsRvgmWGzu6EtER9VlejUPDNqlUeDOBMi
aK/qnCXq52QlXxCzbbMbl2bdCdipDjik8jywBpkXOnKe4HGydAKvmbj0qQoB/CRy
18IBK+cT5biFw4eFNjZJgjgD33ILWu8gOKbYFYG9NsUCb8dcBI1I8gsHJZHuxcVo
HDX3FZAoSIyKaiKE18rcfyHGdua7dKXFp63uva4M/NhHSrLmv6j9YxJdc6SWvtLY
B7VAWS0b4CIbout0010s+oRnX5A1l7uVZJ1CSB47/YlVOzRSlJCs/63BzdVgsEPB
OFzV0TybLcTRgry8J2JG3s4CykFQbipU7CfpjiiAyVyPJH4tJqN/0tdOoFJkCzeI
gfASXQcPu1qxQ8TDEwWuQL3q/mCHDJWnmOuZ3pBi7j/3oUXDWwySw1S0RN6arcB1
HHlGoenhsxlPb1SAnFva63z0GzNm2VHHUij3dYQr6fYiVNDzmMPyZ3Lv90pqiQHf
sub6a+kb6JXCRgaZWDrtFcTLrjVjvArjOx82ev+V4PS8IglDUCGjMNpF2BXbDo9b
gSn309WicfvdUsGQpVVxAhQ3mPlV8Ep84oG2HjhrllyKc9PxGoaNCX7LTy9X3ylC
MgmSrn5zr61wwHPhUxy3qFE+jEeVxC/9OIHCp1QYf8PwYwQNavI1MiFMzsuQPgjb
h1argo5ls3ySOzZTYeUkSphPDELu7+nwRy4470WkEtjDDe1sxZyl6Dmi5CaaNHfS
oLmH3aF8r42zI0Lhd1KLpKpX725AMSTE8Tp99qNo1ATTwk+X70OV7NXI9DLUCAyD
Msl3e9YL3YG3/uucAazfpdvWK1WRu+qiuxLgr+bRoz5ZKOxdO82AvrUvYpIW4XOp
HUF9IDhfRwtokqbcZFoLzedj9AOZ8rBU53LmRkrGulin9LRXCv8sWxH/xkE4JuFp
I2Q9tfPwrnGq//E2O2tbvEl5qx/meScOJ+M5bUrmER/oLL3KSvK6+wWrJRd9kUG3
WVYSNDgjrxE9adkCHEIKNcMHW0+y0fURXQkWD+YyjoSU8Dfe7eOE71/Pg8KuAtw1
s7YLJyo6vC8EpRTjPoSJkbd5oKDRcicVqvezq4eTgGTcJ2vIVA7VxfqAQGbIgqSb
rGMjgkI5vRFQ1b4Y3KCd10eGBDV/VjF+XgWbp41iZQSzKd42+hzHnNqZ/O4OG5MG
FTJihq5gJcjbrOOYZK9u3wVZJp6zEGIlvpyl/rbs01/ogefSEODIBve6CWwkZn3x
YHEEIA6EXjXrIFXIehEBmTHkNr3/3bV82BJT/WwRsp0OX763Uf11LpoxdRW/03Ro
t3xaa6cWdGkWQCILXPT3sBhbTYnL3gtzz+1HumwFBTOBd5uH3nguyE6JGaSMsUiM
Eq0ZA0cXKySHms/FAszfKeoOnl4zaQOJJsCEKYrVqtvC8/qE4dw9S442EnVJbERX
6+/MhfB4kymloHW9bl73zgIgJx96tt4ejevbRF3ZLWEge2RPM7if6GXRFOBIbnSM
OpOWFxLrebPtZXSfIZ+oRIZbTIa2zGg45oIqW8F6nNXYs5kaH+16OC53glQ8lwBZ
AvFSZ/NbpRZMDPmc2ztgs6C2pSz6sEOTpwqKqOUeowk+RYIfYduS/POT/Q4dxvF6
iySfU6iVKl/jRS5WskvS7v2PobOxCMn7y5sJII1vDOjT5fq0iaKfrMMo+GRr/cSI
FzjsqudjHMj4S1mEhErb/ZaSmfjTH8gdY1pivFuPV2IM4UKvI4WVxHkyKm0k9wAU
X6EH0o5Uexnjyf0AN9GVaWlUSKNrJAMyMNYKp1eJSLNNT8ln6kEikeBCq9/FSgih
JAT8EfVGDB0uLZ6jYUwEzoptEMJZAvT/dquGv4lkrcBv8opd9zzQp2lhRq8LBuiE
g65FtAKJ/beHBRB30Pp2xeikMAX8D61f5eXnGkAuYSU5gZ7g32nIktD6DyAwXsV7
ZZUrdP72Mbv0w+TOPRaoMxiHsrMSfNF6wVtWh5dDAspM3gCG8u7NJSc+2dOU899h
GMCerS+j5lfNfeR9bcQUVeycjVVChlnYx/SySkpod899W9ftTnHs/DC8KZBwl7N9
S+7/uYmBfiZn2iVHxKHCn/w0CUMwI2HCjPQiG2EofK2BTC4otpiBIIP84xwLpZ6O
kTfdjbhXxbZ2FjQFwodLet23bbLfd30p7+gS8NtcG8k+RRTaLu6rPlwrzOO8AHai
heFx4MeNhxdS4kzO9L6TugYwzaHmRuZn7akB2VnTV/hGWg2zk9Qb1i4hIK6RIAww
GvdwW81U+CRFeegQDGKnU7LgX0LE+nMUlnZe9Cy+XFLPeRzI5ru5jXc1+3stv5qo
AWTEnrA+lMToKboserBSoZNtQTAwF0+osAOGUkyC1EBJLExehotM+CYFFJzs+5/O
PFQ+HXSErZK1n0y+yJ4g5xVu/RS2pEtQqmVo1L97ChAE7y+BmnlkOzytZ5IVFan3
i80b3RSmbxFOo/vzsxXUcKIVo2LBRGTFbKzlxDYoOdivRa4H27jwsAt+FenvkXqe
P5f5000ZU4BP+NFYKzzfBWcZXhnGgeo4tk19Da5W8MyXHABUPkz8PpE5Vm4uNLfn
PNrNAVqn63gj8p0mTw4Eif/4EJiSqKxDE+U2/nZQqqX+cMraF9ECO/IcRhm964a0
4WKBHVC8gmHh0UDI1KlRKbrkiiR7p9oq89xAqIcniSyKklAY25sfwh1kcJ4GG5Fq
VdGLMhDwOi4IZsfTJ5uAG/RUA8r5iJmmf1aSOBtEq/DX/2o0qGhm0TPc3Cd93YCB
OvwMTsuJO2txhiwulS8LW+/HkJQEiwWfhF9wRSkDVpPh8BpQGW+nTyn2SL2njwo2
0lUFVWVx7kcCq2Qt4ir2aM10IYgZdb6Qh5IuZXNfybxm4nPU5G6WDb7kqadB/hId
bklwPmJZI17VO4KzWe6c41F3ksbtH6Rxix6aTBOVD0iLMeLpBnkUTJkgceAe0im+
8fpZBqJFfEdAqDnSRjRM0LaVQxtYVASf218rtFAJJU14hAjlJVaD7ESKeA4JDS8Q
+ZsGPReedU+kFYArti0rcgQqEnP9RmHNh7oU+HC9fjk4r58AwwdpURieryoExWoI
Kgp2ak3rMzaob8l4RWt+FiyaxBjb2WMeuuLXB5ygM3srtbDdQUkIqwvqx9zZido6
PN3hbZkFB7OMUutI2ctPkjoH4r5LiyYX/Cm5CRfMAYwCcVV6MBAz3eQFNDdTqvRU
uIkqH6GwPT85QMAj7lVJ3CYtiq+xCo8ZL5LRf2VfBvev3H112qj1+0G4stp0LZsV
G65oR7AGI8V9GAYnI+Jg0cNsXuTOWoGQfcoWIoWmtmmFlC5TuyX2/K+xKt1OSFZX
YaAGj4mNXmPYpzlWoIeR3M76NvyRfbudF2qZx0cnmnh/urUwMhNiDjjUZmqrS3lk
S5U/uIUyQKZgz0i1NbZ62AIrP5ZTYaItRtzH2vmDz8ry0qZjL3h9pVjWjX1Kyb/e
AE0kogELT0Kvjo3CyhV3w8T3SEL+yj4Hln8B5ABxarbjYFYLXjj4oM0GsYPCC6u/
iD+uuOHE57w2idv0P9l/eLTSglAhBWJ46SQPdnP5UoSBvl+MD/Jod/6nwW1X7XOJ
KLLqZCJAdx+oIBwkfqptoZyZxOiV1CtsVzOaWi31qUy/RMYlVqOnEdxwggI+Pc4R
ckE9DR8TZc2biifI2Ar3uS31CqkpZi5pefoLrj544LzaqWGD9Fhc5VsdrzfUgxxW
/d4qn5Q+Jg5VLsZEGjMA6N6z542nVAgGqyFVM3UkV+URXyesVsixPIBGGpb+iHnB
PueDzDRfSVtvCONOiZG2ZksSA+z1zkoTsqjlOTdzOHw6XIfrK3eAJRxmaENP27W6
4S+LbbhyzBS7kUeHzmT6W9THbQ/gOyPtcW4zCrN2INATHntr5ewJuIISmhAy/kRX
x+9iE2RWTc7VUCkDkqhbm8mC1L2xG+97/+WeoIPLz9uRqPC+CYfJpIhk2pbx9kDq
fiG7UCotdaFiKoqHA1wIVNzk9jG8dcbn+1iY36b/COXdr1gwAC4KUcux62hvDKqS
XB1CP5GeknXyWQO4B3PAI2xl5LWiHNT+N7r9/0k8Mdu27D3jhwDKduChqj1U9Tnb
xm5dgJ9PK2rwHedbAJYod4WNihTdRbyIenVuGc5whNFV1yW/UuIDCbFiWIy+i5lg
zem3FJvu+T79e7p/CHJFKk3FSUCuHckOtX29zgyI1Lhjcb0AhX+Alg6csB51Epfn
sCfgjxKjLct5r4ufe5xc7l36UGwC31zg7kFESXg6u86nytP2QPfrbTz//lM1Joj8
wHzC/6IXwmsCxR78t4qlniLxnPU6C0daoOhbDDkwBPAgCy95BLUijk6ibSucm3ye
cJ5AcSwTHfNFJk6k35mO3xVTULd8Dk6KVYCJ/N+X8EilxMyYvlvhZcv8jjvZH58D
RKTadkcx2OBDulkcuLbJURgk84gisxDKEarJXly0ziDQ4WTeSRTIfUI7hCxHRV5+
Dt7gTk0aNegqjcpWsvX5nnpK3a63/TUP+DDXe/honwCNCpgy/KGRBgLthDl0/TV9
2mxiQVeRzvn6ZWWX1Czx7tFxjjtd02bhwmgmaFxeWLQHv7NqN/TbHInCCmuD8vPy
dLvHk09Pf7qGXFm5aPQYEfiOcgT1o1zzNTiu5jL+SEEwSHW3F30r1I86ImlLwgZm
MgEtb/LqUltsN5kfxfP2lG7WjjbdDt/ZqimAtu+4OTbXbHYpHKj0pV9QV4nJraPZ
2trK5OeHCwYRsCA9BA9o4ADzUK74H4Hu9ELj5O5csgGfJhIUmXETuBQcAuLX/70c
7/nWxWm/xN/ILTzszltBBl597cRlMGuNU8zWA0HBQB/hVqtdnCTUG7eIsF8tdS2t
C4h/lyZE1+/+ZhEvjYCr8IWe7gu4WwZA05/1ihEJOtHhyGrKR0N/L/k2y2uoNaFQ
YEbKWEEdgnIBFjthW40I32Q1phKhmtZuhCwjJaL+6UIVCUHUDuc67pltswByAma1
/yg7V8DPhxF2TMnOVf7y5zC0eilEjOPwjoRcpklq0eI4zo2Bfb+W7YnpyxFJO3yO
QW4CeWDdQN0ZZRPcdaWhNlaoIw1tizgirNYKutG4z4ArXYZvfyqpUKZFEFBIKCh/
8lI5uM3Hnjan2cec7mqUhlxX04BqYszW3oNnLKrdMGVno5Rmruy6Xc4L1ayQ0daJ
P8H8NDe+X7y8Rp65ALsqBg0y+wVV1GOICIqDvhCbAIQX8fJHyHFWncqno+YeeaKS
rJwi5zJPlhd9sEwc9vXP5i3X7n6gGyqMoPJv9ISckaVEK3KKGu8YnY3AtZZrdDMT
0XIDNvaGfgYJG3kklzH4gmzPYb7FpWUCm2hNqud0ypy6h+79cKeHnxolFxxIsZQO
lS4NKiDDhHajN2VZF50pUUchn4PMr2Pt9xhffZxg6WrX7UDWmFxMG4iU1VBKRGS9
wK7bq5EA/dTmdDh5Hp5PzIl7AcJSrE3U66YH+mR0lCbdLUYekkBmAZ1kv4prwLLL
FqbdQcVtLnPYUUsSH+DHhJxdEQAsRFNbg5pNRadjQ3UT7cp554Cfb529eZRtXtRw
o6DCOmO2GmRvCo6VRl4Tv87Oh6sPqs9Lc1f5XwaIcNR64JUBsCvnZUDi6fqt19JU
qKbgXns5ruOWLd1OeDjJBltgiAgWk8syGe01idO8AFUj2m9U1jlhnRkHvWX6ujum
sU0EcvemzyyiMiduIy5gTQTdkU+y0qDt8YwnWbpvElD34QrNO+E9kCJt7bIG3x50
E38UUk/tflfCIvJqC4BdEEObJAHjP/QZulfwjiKaEzmwemWOXH6YQmnFaaCDa2sq
1ymp1kM/teIMU92oO0m3UiJBae7r1CU9CDx4PkES5C+6boA/3k+zcN6VK+najetK
B0xUVyym2hEslLIEZaRrNFKkbY4ss99T2QbYQpr+FqwcT2iwRDrY+ZO2M7B1ohju
1UvN+XIDwFwFrWbodXa+8wp/ayqyQD3OUL8EsgdP9HyAb1GLVqBK2CK5LV/PJWzj
oJLWwy8cNavxcyu60dbisoaazX+wmZotjreYh9bwu4B73ibhywNyxieBDpj/P7vT
x2tYqJHzSUIOjiiLORhotfsv3kpqJXN2/hsF7vAdAzfxnpp6MxNgtUNAwxlDOzo+
xjTYgB0CMoLKIfkPoQbOWsc84DP2FkhKCtXxa90jRhB2tbgWvq80D1/JTRMpwfgY
ECVd8dSHrYqmUMdgb29OITmkGHC/9YoN0HrsAbDnuV7+0H3sCSK1WobOT+jOsRfC
QK0rypSBJRaYX1ZEHkuwMqzsYcNm6KRJC2NdtCIwOvDb6Yg3vb2pfoQG32cjpJCQ
dztebeQlYytmf5nsg+8TY8wNbkY336XKX0ugFEqT/ZGWtVuhnE56kY5uvsVLKV2e
P7EexYr0nQAxAjbZQlUjxgOOfG64FFArx5lJQaau/X0ysDrQuQ6uJ0vIWiCrxmJH
UT6dPcUTTFqm2c9AQLV1d8+t/cOOMSM0XcG4o7sNLyDVC76M9m0qNt3ailMsMmpL
43hjoAc3fxLWd219M6XnO/kbq9o4niaCAV4ugLtaazsXTGReJ4vbzpNJZiXcPAtq
TWhhBOVhRZQovM6TnVh9LVndbpbUEqGjXRyxbMYVjVDVf9UAn9+HkwdYrxXtnsJh
mxegbmA90+p2gMqtM7/3Qny2LfkAvwoJkb9l27yGvXwxUxOVTjKvL+59/cj+nLoX
CN38cCz/BiMZNA/NxTYd+JW4eulDm0pMbwTkNnl/+wU2vKQjrs8tR1nTs7Er4382
oTLizMOQtNIenvIQ0ztFe/p0nWjw8Biu37oEF0uw75uMfESSuIpdxv5AXoJ30C6m
TQzRAi2dlNIw74AsaYdwkL5pjuQZDz9FoR9yoykbA6Z6v/X4UJUaouT+QjJOZ2CC
R/S9i3uA2QrI1XEgoiUIc4NOWscJ12d/8p65HeQt8cSYeozURJQaCWqbmy10ed59
so342vt9yPplG+kQ57lEb7HLEYKNIK1T8oUk+HlgZpAXYhGt3xh+qZqm4+qMgbC1
bVUGnfV56FeFulYzAeCv4eIj4IgubSsJjKnOV/azszBxyb7G2Yy7v2d6ajEw5iMx
0N32wbPrOBbYAkfxn0Bp7Dm74NQZzZgPiiZDH9RXMWLVpQc5A9GOw81bsx/GGafP
6zRS6x+UD7dxOmqS1cCDAUZBugkPeuCF1vwTM2hiAXCnMos5dkuQgEmwlS/J0rSr
VVoRK5qTvA/S0us/QP8bx+0k0RXlWUMkZ6avxjD1mDs1y3SFCmDUG08oEzwtdifU
lDdodH7kqGicPd3y6VVn0EWhwrnc0Ws5lcxVJWUTyku3N0uLKGYhhyqD+jwm/RYM
LglkDnwf7OY/Hvqqolr9lBvF4KcI6Fmlq3IiZ3iZaZDBQl47vgeSxB2WeWtCtSUC
1Tno2YM6id8r6DdSu6CqE4I/sgCwfx6vrcw1ka9T+9uLMozZRb9ETTZr1FIG5qcn
hriaX4rAQGjCbFCgD226tGn3JVWOmhlCiJpFBvcXDtLsOm+l/6yyM2QUVstBXxv+
hA41waBSc0b9frpCBRhqb0/o4Mwk0Xho/NS2fRMBViTTGNHPbgZqv8r8YskfIa+R
9P3tNzHpcjMFRfYKrgujwJDIaJdtmq20hwFxxPYrIoeibqcbnQGF0AFPUT+eSVkL
J/GmgVY5BvT894yTqv/N8p/2ekSCQ/yqwTBWVLk0fMFingKB7kaKm99bg4V6aHR9
7A9WGyMEJGbCgBxMNIVb9nYHqWSA3J5bDvCZT/MgRAo+3itFjAIHb6DTB0u8LEDX
GY6nqEIC+zm469rL1HdSTJcOiK0VZcrXBnli5lXESMypWBilvnuoQxQqR1/dGa3y
xCVeqJFSgX8YpVD9OztEoC0hPNoE8sisTeCyUm8hSFbINT+wYYj7Elw0mlF7ALr4
aWwOWhzVGJOzuwJWGGGY/L88El3kZ3rCKVVyWjUGdOTkUEfzh2L90lJjgGuGIStq
bfLQsrrM1FGmRqVcY3TAIVNzXjnwSCjr/7d+qTsxs4PxyPVmWtJxcr9a/YMgbIoa
SpfmbXDEBcCOevgPWqWPi0GjinsppgWtQdv8fnEsvfRxFEsZNgfsSUk4EC5Kx64u
Y6jSHYpz5E1Wz6QBujmrV/JCRpGzyKKkY/nf67w1j308eUQHP0iKpUM57hyniz8e
i9ptWzl+pvTjnf+YknL7xIlTGkidfizUQOrjab4nSYP5blcyGTrJGL4gA12TxHzW
B1ghMQjlCABYLSTkAHomRqWcoqT04IsgdqsMDg5a7hIJYnW5w3ra2CckZmk1xDkr
KrUNKCeKa2fJHJfQklfCCmNVSygL1S/Q7RekEBeJie2jx8jTVy+zJo5Shp0RvGFu
tf16UNld4gqNrTNiEc/yv/JVYqZr2PjaWSqQv8cI2ydUqdpq4wap31e1r2CR2Uww
ioiZpIy+8Ll97WDiShEiTr2KGOPJGB7kg65VKgGYSHD3/2mf2pXR7N4iTtE5GEFe
ppDvUWvY6InVPfvk7GjJqVNFPaCCT6LSLHUY7gGto7unXn5QJ6BzPmuyhvvMmlMl
6xVegLTfHuxNzyA42LixlPlMWyl/25Jt0N2KmDfeiC7tkrR7QMu9MlWnApHKF+Xk
ud4c8lX6t4X4CNHWeUC1rV/VabARnCNQlczEDnxueNh4Yg+8X38f8YbBEtD+2YYO
KwPJWdfIVTW2590jXThO88jsCjOsuhiRMONEn2TZHb56jwQY7XJTNABgbE98xQL+
4ZGxY1rSWdL4dS9i6A78gZ+ePiAlPi9vX4Lg6YPLK7V1I+mVP/ngckGp8gw4y17b
Td5xhzBySO+10J/Ck5HsLi1KpjQCxgk34s1HDNnqSvflF6P5lQq5eS0DaRHw0eZ0
hoRN5axUfPy95O4COX695MPkJUWMn5kMAIhq9dMwpAbeTGdJLR182dM+4E5M6mS/
PePEuoXlXP/wO2EvEH213wIULWKbj0gQA3kuGi/eqmiL651XCfohHTxPJid4OTGM
eLYQfB5c1YxOc1s3PDvHFr0urjS0U7kYHHBoZNT0M4fCdW8Hd6MvT/wlAbYWzX/P
xBWv6509qlnZL7TzZgGp2K7zh9HOTkk0WMtw07/cUa+FyxtnGRgMO5SRjrkwwZ8G
BhoQWe/hSvQ5gjnDRYj406L/zXoYyWGen7KUU3ALa/nxv9//PKPMlrNNPd4s4asD
FGPVaadwE6MwpvzP39MpRbEapccpUDipKKrMXs3wjImQG3DWagxACoJ+2WGVsegW
Nkimvuiqqcl4VGqpix5ssweF7SLR9fc3lKkitcZkCEVe1H6RXsKqsKOngIf04IxY
flXcTRmRMS/StqPCUZpihXAUtndqmHnkLaFNlm8Jt9mzrtE3CnVDBVwefcbWCEd3
JihAMKY5hL6UbDmqi3dZnl2zLJsGOxkV8hnMw/UWzzW00V7SuAhpqpj+x+ujJEZT
GbZERF17gr9UYfQMWKD25tTm6UYsBZs5K/mnTspPvyxIVAar8TKrjD7XwTkO4+ME
IDx2QeBAGupLoIDasxRmokmqrgjUb5W/HbquyByIDxEE+J2F2iq+Pmxo9k+XwqeO
u5P30WVHYrB8VYvNYSmZpWfhZwn4hEngk2z9PFKCdS/H5ec1ZdGcrCYdYf7Zse5h
si5FnFBDNR99EMt54DD2YsokR3kMgl1rcwfiF8URcSwrUhMfKzDDAktRYP1+diXK
XZ1bId0b7XLQgB/BapD/J62B0Jl04wlObcn84Btvu0kvxLp1l01N03eB8z27HWWm
crlzhBenm/7E0oS3udeITo38GTMfodPOAmI9DMtZojGt2vRYoe7l+Z1gTVga0pFV
1QfmNmChD+SykAkHR8RBfu+ho/7LhV+E8Y3qUBs48tj1IeEWQ6VwELvr/OhrExf1
XTXqDGXWQOGwwboNtR0jreoblpDVwdM7GtFY+KSU8DJ6gxDNSWaoO+a+CChJK/zV
mSn1wat8ayTU4pKpF027Nh+3m/reJm9/svY7oGh3v4Qc4O22qPaUa1MBvbUn8DaY
kXNFSojfrEyMbPOjTjqWV5XKjxDnMVo8Jo1ZnDybAFhGnDoHAxkETGu8prgYG3ri
F9/ur6CTgf4ObT46K4+elP73YzsmE6aZBoz+zgDMYoPP20uWfDK2gvrVmNB8yb0e
HBMXhENr1/Lic2HSV7IrklsvLkeB+wCGpllpT9pzVDq84dTMY+GWXMDeZRIBklpU
obfsFB8N9Jcm9iO1PtNlanXh91AT0ZYknIk73dcV+Obc76YRkAydBWorX85P862K
I9/oX4OmOL6vi87+3jnxbMKl5KYrra5iKac7APlP9m3YiW/e4D2OaUoyYSh59Jzz
k7IxXNWwRIfhxhyclmMyJptVrSif4gvY2GV/JoDRke9Zp/m42kE+v5biWAIrM2LZ
3YLPAtZiz4Mn9KGwT2sp+njWY5bSPUL163aLTyOYiTzsSLr5qCF79E6hr6UjCMQB
rhWAn7UqIYCqRxWrnP5JEQexFAtsbBojCI9Qd1s51x1p1FKH25z4rOLCdwBt/Kih
NMmqBdp752ylOQQ0RfH7hGCDZsU3sQXHhkAVD6G7R6l/FhDxBclLgBncKQtXLlxH
Pm83SsIwgyQPM1tezExrwT+Yfox3dC+USeTX54uTDu5ff8W0wysK9xvdEPOTEV0w
8YPBXRN1bxCMvvlmMydKhsKMa172e2aJpg/ONS1FuV76bkFV0HZrp6YkuMLPTdS7
Sr8SHrj//odiAw/eYJ4jnRZGCTZZz/IV2oZMQ2lhsMcMoaFODFn02ffim9Qvpq4C
BJGeOVrp6smYNFA8LMf6VqMF5W4rixpl0EWxsJCkGw5ggWdwBkcvx+FGdcPw8EZM
TWKerXr1aMDiozzRqxH+KCI1455n8CQfx/qTwsFccEzPxJw4S7SF+Eg/1vCpeCF8
boU/gvSBbOVkU7Mv6UAqS44QoX32FaySYTAhLxp6f/beDOSX6wf/mqWhT4F2PGxs
pCHrJPc3pbaai+GF49x0EU4u22d8TaN6RWdF4fNzXqI1u6+To/CV2dfcUxFudB4y
VVRAAo6sCMf2UvyRebwXtVoSkRklSpEmo2HgJSj477HUNM6cKuDUwhKAx2fFxvLt
3YgGgq4mgLF62aarkzR1u/U+J0lFRxspZc3j0WuvrrTb2J37JPwdYG8nq5kKL7k8
cw3dDb2zg68xXhk42hP5J9Ld9ccToh8lUj919IbsDS43Zb/rAKl0xX5MGJ/Cmj/c
VpfvOX/UpSj/KJZjnRoS1aDn3eV8aPW7gA8uPZk+FBkj49hVw+nE1+kolV+t9bkK
nGwTRhcnnpEoo1gqKyTg7sjhnDia6ONsVWaBGdD7kiNjSp+/NDkjn4mqJ24UCN13
HFZ/kxj0Z0H67QkEfRMWU9O2U/C13xchEx4hbhVplzWU/BMtrCDYmJFKREuikODV
Ncd5VI0Z1JPf537ki2ymyL+PuGUHJymsJ5mpAJytbXxcSsJzNfRSazgmaDgQ/eSJ
MPZlCX1ycgQBjDWceXCx/aleSL37xHUXl1sh1bhMedBXeHPzrbEfOmEQkZ8aktpu
T3oiCjLRShPWo3WnhjthCun6yO3kSJj41w5kz8wDdmJMzVM1TGJNFyYMIDYX8Bti
N9qv1BrA0SLXhTV+3+B22pMATFuBADwSPptJi6Ox8bPCVuCgcY81FEcWiS5Pd0tW
xCR0Mf0YFVm0UklZ9EuqrvHkE2wI3yHEh4ptbWNUO65D6CDHJE1CMSdId/YxRirE
eaC4ocHoFgegmCE9ORiATy9R7qQ+cD82h5PTPJGoj8NvKURzyh3qOCP06Lfq9P8y
S6jyJn2Afp3jxZz02FGXc7nEiYZ9IIrcWrbETZzN4cLEOB1aPBRkpC4xf1NQZkKr
wq5nWVqoS/21/Cx53XwGx0n+lblCYTzr/qNsyyVHUsJHum5cYBiu8xy9l2t/bZvp
Uqgje7rpuXaWYR/c1aTSTZiVf9xSVGbiO8akU1RZBgUmLWZlT9qZ9QHU2wpUnICs
Vheq093gdBmTI/uWZ2OAgjz0zZvWWnHJFQIYXJjFLk4DmVDEMNS+VOQ0bv/T/0gV
lOprlyS/AxyC5JC5005EIo2Dfiz/FODWD7JBM8t3nnunngjqMfHTj7B1n68JVJ++
UxIMuyeXnR76B63L6h02x1tNy8ZuWGUgYjcIqOxIiqidzR7bweyZtvJmQPST0a2e
kxATvCVHnKVp/LnhbjZAo4OOij7+rr7GrIBXoleg3DMoGRtXzqTSnT0MAZppsk7A
nrilQv5DWC5Kg0L8uNN1bvihCEHpW8JNaGdXGLgGFJOGiTF0NRAc/qK8BvxyLYUz
eq0zLj/6Zt1/dqPWznnXviiqdjKSuWIxPn2EFJAUO15b0YXfXM4CkBLwlqrgaXMz
EOnxkplFRgi3Rwv/yE70niYwg7vMbtYeWIeIiCpHcLyTxeUJatLAabrk3uun0Xi+
uZIy/mqHyHA8AsyPvoaO5+DQwrI1R3PTbrq6gj2PE+NpCcxczaQ+5J+1318X2Zcs
YeobCNtvNxJNxtMX9d3oiAWGPFY2Tupo/LOF52r8+eU/oaUqYFgmCq2D4AY2ph3B
XGxqZt7XFYeOWiKdMuz/yzXOt1nKzkjDI+R0kqMSx1sSlw9ZXRcQxmCSnGt3j5yQ
L0i2OrTNvOj5oXK7TtH2jQjdNehsdvRDirsldCq5zZ9fwrDOkaozqRV8m1jUMnO6
sat1Ab0uAPvDDit3gvJLqVTbzJZwPanXDC2MX/Lh+wm9Czd82bHy+/8+DBcbqP1h
xaTfBgMpif7FY7dn6ISVdvmeSKhT+JBP3atWLZjI3oNqDVxTQpCTmolT0sHh+vBd
CAZyNO8g+lOzr0VWtxPC1hF5LYar2h70wdH6HsBc+YYEfFGo+PQmUy+8fZfVqk4N
QcxST03D3IJk/HyhwpGKjfGlWKO+bQywj5dkDtHqtBPhYvW6ZDn+4b+y7Gmzekik
r86/JTB8ZPpo2UCuZpRZuPTbu7jTihBzNI25VYW3KrI8yaQSWXBsi/Y/nsikW+Qq
p/2g+UgTLFN3pDtPc8tuu2okja0uEgF7Lz5P3aJ5IGbHd5u1PGdSVVw+F54SawAS
biwZJpzOmDrqtD32SGS7UBIScE55lMrvY43DEaBgtbf4c2Al+7iXLdw/H2hCDfuO
Y4MqYfQFLAq2EvMpNLiwDWVtyHbTjhF2aEqF1WnUf+LKDMbk19Y+Vq0/5MZUxd4w
NGM7POUJwJycIQJplRFYwzn2wkVz65Nb8aNLa6ktfu7tgFMsw01vC1u45gA+GXar
FwJikBBo1RYmv2NGdfGQAOdt7BgyYieb+gcUDBSXVwiS9PO1e+sEciYsRMUW+mKz
PUkmuQ5aLb0wRIVjm0GH/kN/bEgF1cKD3CoIj1Gpke47UMiv2MZFHXaJO/uvF+Xl
1Hje7EfGXpvaPq2dIUWTW7hXLCL7dxp416OGOngAVNkloMmqmHxBWlZ8zGDj+V+F
JlkYM6KMF07gTR62ZN9uDSNoL/LU3ovfxZDRN895m/8Mp7H6GY3XyiaGins9ZNjx
BFGHv8EEFxh6nopW9AG72DVa/TKTHfk+4AD1SuJFQ0zBHy5dgVIi46Elj8XyxlXn
pLNy4iEiqVwiHDBiaYtpiNK9PIvIDyjo95vmWrgqxPv8jiKa3JMKZyS2oaCE2nag
4FOZ4vPOXof1D+rDwo9L6qlQdAnI+wg3rTC47JGIDPd1+pNj40OsxoN8n9QRuTxa
ZV4AjbarqPN0WkzIx2KeIe5PjoicOG6AFDR3os32TKgF3S16Qqxa3Ozq1T0e0M6n
ODfayoT68eE6mtlvhpIw29zbZG2CBxbUeF7/UXlmZdZWx3V3CnozbT6HAlCY1z8E
CrajfFcSTKGG+cGCo5F3mHa7F2P0ZmrWzilNjb0I1Ss8hPFYBTDeEAXqZ5lLG6dt
/FQ6bkpb4TPZQMR8+1v3rc58Cti3jIbI+fznWwT+pQVYzO47u9nE9FQTTIJEbdAU
8XX9wB5Hku66RW0fMMJ2h77511IV7Dq82v5Cyq/o/IamryZmJiv7j1fcKxGLNp1+
9a9CNXBzgi8eQcXMGqQT5Y5BX6mDu4Ridj5YPimRq/tQ4vO0x1mA+j4YmkkOa1Jh
VdcLB1HxEp8RQ7stV6X12Fb5I+TwZE+e9rsxXMXKGQTw2jTWxJ1Zh8RfIwkLQKK6
6fMUT7TbSyGtupwRqbuIJ5CQ0mXxj5xjteFEPk1oVtdHd72O/Eas0R/A7UuUJ/W0
BrYu+i3Q6Ql3TJdh+Mmcpd7ryagWO1vnQRQ7ltYN0Dw141SGmfBLO+Me35lTOvwl
zqbe+5sggpRwmjNS8uu2mNE8p0yK/qRMO41fpaWsIcvETfnxOUhj3EaLOE33SHkw
9hA1ULyrHe8h7ZNfyNvZHAqfDwmUjhNHtZKXlOgDnxqW61nCqQEpW4B881QWskhf
q4ZKaXocrslbmhDxKlogHKlrGwYdkalAUyULFcA1vrsi/YaTGz91p7wlgdEzrGL4
fSVdzKULYwIiI/7IhbxDlipDgc+Vpy3SFwDVhmvToEGKw3all89/hRRw17tm4/GQ
D2HIKFDK+zjTaKK3eCgDa6YiRGu6VS3g60PoZ/xbj5ADnfBT1isp2SMOwgIQITBT
wr/UrJhPYpfUIGyKv/UKHrd0BMVXZiGQRRSWnQVjuwYEmLIp+zTpvxAnJw6G4Jtn
uKSSChA1OJuNH2gEhvxkcLoFOfmdwOtjCUJsAx5pR4aN28F7xpe2AgrFTJ6zLDtl
jTphJgxioqTuijbjy6XuEqcLaSKC+C1UIZUjzhTP5IkGBv3JPdBAa3Vp0KWHqYQc
x3KMK+id4bVuBDETce63iBVcbxyoUOL9UARH8Oxj0DKSSykz2J0rod5jeqm4lyk7
CfMACwVfNRRde1gi6gLR51CL91P+S5T63b8smAxjQbDXWZChHeSjkcaB7YQfC4l1
gG7zdvMhrQEXt6kMGM7jaXuFRJodHN3FHMjKCUV7/AOY7lV3Of5tOc3UvmXGWSb/
YzPI+jEGrzRfbWPJHHtHTj0AnvgkbuQk7G60Sj1XoNDA/vikVyzLwHPeojgmmMGB
mth5HO7oQefQTJJwzFLFOCcDwSFC1uZJLal11YLPcsw1icpzzrZve8egqo9GNhEG
5KAydBvC7n1rCfJlXnY8Sk7zxpHhG2Gw9STuDUppy/32eMqnEtYUqtKb0Gy+oIS/
/uKbvmCODeYDdddWi4WO1jADCZxf8DtRj8hXg3S06RCPePOSvqMoHi7/crCVvvxY
Knpvbp5ZaQe/R/RHD7Tk2LIc4XUVFAqt6HGGBpvgg9uRIqJGGivb2TeDbRJ42T5F
4A+33kzJBSuVgwrpeJJTrS65nAlt/fVMkCiwrokD8qL8BcvV++p8pKeOKUpIa7XZ
0Ytovwm8d+PcCGrL9TypOkJF6y959xrrJC1L9xClx8vQk4uBbjhc8Z3j73z6SgxF
BZoq7shZyN8EVulfcxmLm/9MxdWAZw/XBIsojNWJz6kGAEJRzNRq1+A41MHZSFvl
T/O3EtlKclPep6b6DIYFVB2ElCdhs7lyiw6PDiF60R2c9kOF7URb2AxnPMElrvPd
yk75NAocRSn95V5HN5XOX5X4zG2myr4nLzFUayIqxmfQbnuUnMAL4zUoHHIjGrJY
zfUbyWIF2/UcgP1Q8mBiK+tdaft1Tq4Dxw3Gm/EjB/ZXJyN+O7ya/KQFMo1deZx/
Vrqd09FPJV8E0LZvzRhSEV/qjzvLlyJ+c0f5sM4gX5I4hSH/xE8Iacs55LGKDoi4
Yi48QzSbNAb7juUeYved7gx4bdway+JFzV2WxFq+XprH7nSR0TpWke1Y8I4uoYmb
MR3ndQjpLfDuHZVrb7nKNVJNjbi52Gbrl3BO3NkzN1z0rT+ER1SKOr5ROE/UAUlC
+XbRsFCENf8Fex/0Fnk7w3+JOibBby18JUkWrjZK9w15R78+ckYBYwmukAGXAu30
6SQbzHLm4HA4qs/0PYqP8hbM/7UxzljLqe0M7a1hdJZ0m/wGqrFZzLvNabJ5ncvr
O4eN91Y76h4u3lRJ4+SKvfZeQQ6SS38hGeDv+XaRrtvH0T2T8O0FSjgUCawSw458
JKCHlGquN+yUmZ3hF/2+mmeLT+89jiPjhdFo3VbxBnQU1ws1oDUSszMyUHLqlGh/
Ci4pvPisT8uRP2GZbbsnl4D1+SdwJJpBvqRJp65Fq1yoTUKSs+FS5zEluz5wlnH6
zGazBD99L7RWiT164nEAnKJwdmImeqA29TRB6/reWQqrAVWhAgK3TCZNwzzsk3Ce
0prZJR+C3QxQXyt3pOXmyF6zwWQLze33pq9Yejcpyhrz0WHwZU0M5CdG/V9QvDo0
YG/dghxnvFoROtp9zRlffSNvJvP86jbfWES3as+VR4ulQhleeM046abE9qWG6j3G
jmQzH+jYUhUmzHri77ojbXeqCA6WjdGJey4lpsofqdZjgTMOGBQVH/GQtLxSc8Pn
pNKFfP3/wM2PLLNG9vNiPqtwsyCPDjK/S8mDsGcdllVlf/X26kD3NEfxa+MkCmDM
ujMWSGLKIkUm/iGUA/IJM/9wKaa68TleB5ZrtfKapIOWOI9bBpPgv2Ol46C+Fe1P
Sl/sGPAlBLvwiBnSWNHABXd8zG+e+AxqPm/pme+iOMC+vj98XUGCD0+s8HJt0/6B
8D/S6uphBnxXnUyyVJMOMLxx6zOf4I5+EGQ0jmMKEZw/fYUs9AlF1locuLTbY3xE
qtJx0NE6h+uYvdZ/eDT+swc2PPcLdPyChEZXRSLzG6QWzIMfLZ+uxwO9R7uJx/Aw
7xFZW6APlCY2opPi8IWFe2R6REd4T7jT8vAJwCJHRI/J/IFX56IIBWQNbEHS1viX
JpwPilci3eBqaX+goVHjNuosmgUaZIYuzICrh2plqydbWVDRYZ7ELVvUHtRJKk/r
dRQFXylzMjl0qwFkrSONIJdhKumYrPYcgCj0L1Vtbkv7RBfV6AvP+HIhse4Z/k6s
xreWRSZeR92pLZXTy53CpLhcKbrP0fNCWKZf805UIIOutCWMyNtLzObZHonfkmNA
9VVi6XzfDzaoWPypQFQScxyk4cZxp+EceJAhp6iLcg/Wc67YgxRGNDAG97lWDpuP
9ceDOF5wjHwr/crQN/VWdKM3F0PGBVfiRdJ2owjqrTNQLts/fi3okgHTyaZ3LKtr
G6wRTlV/flr/0Ew8okUDuZBwutGDvAZoSWaxM4DW6xtD6tlC1vyPUGUBbHmtcHLu
`protect END_PROTECTED
