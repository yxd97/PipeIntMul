`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tceJLX9P2u4fBY+c5y3oO1GKbYBd1wIZHmSwz+s4bh1QthaJqYKSrqHQl/wUU9s3
JC9SpXFs4N6dEHE3OXmotn6zQmGK5WzaLq52mxA69WkgQ6ASirZ/UnsikQ5nvKQP
us7y8YvkaHVnFby7ZJ1ikJ3b7Yf3LEDbzST20PPaAA7V6Uiupo00cIMMOMG+nN7Y
226cKOHw3iYkuee1Pwgw5Q6WBroMOhFhzNE9leb+g2KxGMvmQ4ynUUlMUvbT9efg
xd9+6siOCt0uJmILv/cg4jRfZBcGt0prJkXXVqqURMg6yHOT+mK1eJDOlo0VUxJs
jgJ+DiFBw9RAT6q5EgfazArDBwVXQMbQRFk6H49SwpmisS0pgXnWg9NLLdc2yyZI
bFkBd2d0UIoq6O0ZIFJBkLaFAjg+/MUrPaBOUdmrOeMFUKlNLQVnmpq6y99gximT
jUt0y4UBUVTX9sEyvr3Z749jvNaKa7DCDnIyeMNDAeg56hTwsbsAZo5riBAhdrYi
aufNrDzZpq5IO3c+6iRtm8EIub5VyQAPEeyVWtrLMdINlMeLdLK/Qp6SsBZeB0tW
AVZKN0zu63T9QKrCu8fWQIeSatnh4ZibSJkFOxwkrTuil87sR1z1N83oHG/Xc9Ux
MDYru53ER7MJQ21ANfWzHZPyKIGKj8wrpOacuekoFQl+ekwDFtI8jtTnLYOb7nMy
3ADhZY187lraIIOVrcsMYZY/SHGRRiIowh9f5UZNUAyg2Fa39NxkiuEqGZf+mTl/
hHrC0T/DQewUYgWZYBBV7FnzDxDitwlH5Jg4Ewcip5gRuhcFGNlrNTzmdyZyECfR
oA1XyAt+9DKmrEJfAcVQXg==
`protect END_PROTECTED
