`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+lQU1q1/4fmjqoYkdJxJNgb8u5pedWjI1LYkP1l4FKQkw8AFZ+oovGx9bRQjNmyt
OE451l964FU6RgnkZKtCioG8RMY25VYu7+0cynBGUzjeWmclkFVYc3NISbA4hCK9
BrqmekpOpzZ0BtsPcGhRDThEPd17AYKD6Z6cLWVhJuZ/tfOa37wjYzTjYm7pkJzn
KdnNgAJao1fMQvrgxP6r8jfeI3vhzqauYF0tLlkr6VCBN7HPEF67SGb8wPzwe3hK
hPB33ClHjig90ct9cZVzkYyD8fkWSrj7pQgRiLCtMtEEdbzXfEhJ8bkADOjZcCAn
axVZXmZH7YxA75AnXkGix7cVbYNKbiMVK0aQYcwDtcmYDpzbFVipVJsQV+xalQMc
irZW7hGkNv9tFt9ApcEMYGd3PyScIPjenGsMNvZ8aMvv9QsLz9tn49JsIIDODGTA
FI2lru8p5WWvoTEaKOEI0zxhASuhDMD4cmeyXSBt5c5TuFfzsR6b3PQIH0nSps5y
qUGSzscDVvsTF2ixuHQsu0k/iHlJAUT2AvzARLtbTzSfRss3k97s4fu3t65DdzSB
2cmIFuYVDGKLrnJRTAhOhWX6UPE9ydnELobHmih4KbE0e9qlLv8NoC0rIek8Epzi
fDHaL1KcMW/mlFUWp9zj53FUJ3LI+JcGQSkqZ+WEqc0Yp87P7wF3BTucjQg9STXZ
agmLr8nI5YO0uq86zemUhmJH7165/OCwlFrio2jhsEE8xjAGBicMeuvxXJx1efdo
uyweTvBaT1wNSS2ifVEz7Mrsqrp7U1N4/gaaJVhH/g090MgU2hrHh/RTo3L+33YH
P2nFmTXfw++MOYUU2+nqXZS7nO/WkE9+BAH6B3UDGLSsywdazFdWXycw5fcGeNhO
9iuiaaHlidzrph15xfKM5jJeyuWwCfUU5U3lsruinoBwqoZugwNt+la4gKAGD+jo
yUeDPMMqtSwe5ATNd5ejSHzh75yabtb3PAgzIEvefJ7okBSMplan87Vy4z8bsQkE
kVv2dvNu/CHWLht3pFLA2gA/ZyL0s+dfrISa4+i5Gy37g8bWzK0AmjLx6MiWTkBy
jCnWgUfd7kT2Fh0VXAsIc6bRiQ7NARO88T6COhXPKjEWmhvtbHazXPrJDdC1xYBq
WEQdxzgcuFpzHWyWi86HtfESzKknRWjVE/DaXFPBF1o/xCZ1ClfDAc/FDqzDPZEx
`protect END_PROTECTED
