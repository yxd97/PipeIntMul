`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ABtoL/NeN/WsAdABVbHDchNYAE/mI02ku38eNANHsLYZBgM7cDdlOvnqbX6vJ5B
WynEhEJqxZJaLVKV1Fj8teycDEP+d1o4klZeXj+t0S82CNPxz6CH5fk/+LB/rmIT
8eA0L1JbqugiT4K8+LE35tC3MaRB7d/hP8xyflpn++km+o2eak2dktejOpFyeqsH
uosc7Hp2Sl1i6yFQxyREShhT8ezQDYM0S2iGNyf6cLoHtwyom2mJNTh9EggJyIj4
FbiCIaO/I5BMDE5VdKs3o/oNMoDsud6SO3NTX2D7EaO/KguDFqdXaAcW3lyUPSfl
/DaYlxlRQok5dFmUFauea2+2l98rKNa/OoVoSJbJ8esagOhMyYJYitNWvCaghoL4
BgTPuhyDKoykZ3/QDd8RQKUmuJOm+doqcK5thf5vpYTWEAL/yPeVUHyILM7VO0J+
jVRNgjug/R2zBq7/8GabwDNntg/4T8OFJj75Fzemgb1Ua2gNbNpFEWj1yXd/CzEE
Cx13n/Ryc4dmo+12ypt9FDlqolZ7rgHYR9EXnz78Y+IPMlv+RuYuQ/srFUt9P5n1
h54W6uTKFjlTOd882JLgdE6Aqj2MtJUYrG40R3wHAgRQOwD6rbUYFKCPART/ahHZ
JG/+rsM0lWCmzThz85aipEV9g4KZLFaynESCW8aOpL2gyd5Z8Bk54cc8qJ7JTBUJ
8UcP3Vt91pT7yMETjHLkJSS7z7yixEqi58J8ciOGjA4md8suDiYdmNSxp0Ef56bP
GXlHewYPXLH9W+pknrCVlfk3O1M7SjEBoS3Uq7+F2B7qIgrX3oFWB7bkiPYiPhHm
pXQm1kRE+ZMbrghBkIsMArcn6LqgTv3ujWPhCSp1D0ZrcdleYnWzfpdmi+Wsqol5
wJloE40hXxX4Ia0roxIMWM2zAHxRw72oHAMygb0C8sZsseZUtVb13jk04cqnLaMI
zZWDijoDJ11rKSGy0t3yzUkClpt8aBMZwlWnrNvky17izSph8MGtSTbVGvaJUL8f
Pn5+9iGhpeZiPLZl/Mf3tkIbbLYOkjXdu9z6Dg5lW6MOFeSRdbS7z6PhHecxJD85
MDxaGuLbfscmsNxWqTOwRRXo0Wtnyf35vSLzANcKzhfV19LLFw1/95CwMIWR1CzG
4m0rBnD58BNUsZYKJwPq/bJQ7j41vl6XormXBfkDVmReLXPdP8adiuI4GPs/dJB6
Hf9J7nSd+G0ioQg06g6h5pMflIyk13B7rOVSCAlCfJpO4SPHUDEe2AyeKQVc4l10
7Y959unAIG6YESdRg6BDmtmG8FEJ/uND9xmxD9PMG/3vYlWR6gIErabQSjryO/ag
XUYNeyvvihck0UgCF390PkhRWYGg6RdbUDua97cF2/uLbNKrOz76f+TINklEv61l
OFzoPeT2oplPXZ1UAh15Id5doiBiNaG0qY3GI+XGmMA8KcB49lMRq7hwff5cMGpj
+2QPQx2EefKhDPVpwHWgyAYcTgEXZZ/I95p1PnVbFjrxCGlR2b2PJmp2g8wsQPPV
4dhpVxklQJBF0SFJ68BsL+iBSwIFfKD+4k9SeWVtot5RVbVZdBrXCOx4VD1QYdKK
wkTMxRsFjEq2+cCURzTmj+rHLxJEqEncK2AcSX7aYxEI+/V7PDpKIZ+RFkq6B+kW
cvcpKeQgkPe0koCT5eZcSih+MPRFclDBhEt7dOyw5f8A6P5x6ETgZLtd8ZrstLdw
KnTDC1lxD0ZEn9UuTtNPibLDN8RKc/NuZUEqkLnPngypoTJP15MV+5EAGHlKOc9t
zsbyoedoxrIeXQwrVd51Hqi7oN7J6NYyUTprXCpjvut2hkepg0fO1Rv0R42Wvgg/
kZTwhCyz3bo9nVEwBKDkRZb72Xs+L2QJ6HBUgL+iwpuEtUUQR5mFF/ZiRgMznc0y
i2Mf9CPi2PNF7L8ZGEkdJwzjbdyFAUbruJMdWaR3X0grv2TZ1N5lxKQVWEm3L4UM
8gLjCfjJLTK8We6NDiBEP/wVc5BzuVPPuEjlqHJSm9qFMXl+dBIFNqySvcQCgbcQ
7TzDqoIPbIPFbr7mHRx0kCm5LT7oBTQSrJ/nJj6585rB52hBOvxRAmgw1p+GCmvw
v7ZjJZ4xNM3pOZcn18Fd3L/Hg0NMtLKdKT+AaWhffNkLhqa5YPCC2eYtBRnIlzlf
XtWY9F5DgospQae/Ye6ven2R2taJ2CSTrIPbELfCyW5kAmYsyTXTaoZ9yOAN5fge
3okS3zTsh5NdfSf9ccIUCpZgAWiv97iW+8oNOMec4vexi+oAFtNbKEEIezlIousM
P6TWuxKJwdDldnx9msqjGLXz62iXIqe7+43/cbZer1rOFQ30fNxO+SBrRKUdnPUf
ZKTpRt9bipSSDcm3hGXPUH0AlGTVEQ+pZUxOYlpiKzF/SW/mTDDtmMOHbVdjOoM3
r94Ok05WzHd97mEL3aiRiHyu+RNXLBi6dKm+tTAWeqU+afMU/opfPdUzSji2o1/u
DFG2sGoU7mTBumLmJhr/G4/fkAD0SX2gTsKDkxeD9clZglcX9AORKOXG3MeP73Cw
HXLIF6ixe7Uy5LPOGvGLADI/O2pFcunmCknJ40ReKqqA2p8ZFbSKYoiKhA+3dt/+
RQJsheHmiIHG4DTCqb2a6Je6lYySmYoXFiECj2niz5w1HrvMSZol5wNM0d1bl5ED
U3qEfbdLIhBxw+47qEZnPcGz1Rr5UVWIKTYtlG6nTRXL+vTqGzPxQiro2pea7C5f
NCQIlo0VrMMJvZv4XyyAMEVwzpW7Bnq1BnlRQSW3Lcyx5XvQg9VL/VwO45ahOWPd
mzB61j5CwXcucLrv6WMxc2yjc5EOGFJ1HAV4BoCpC5+Ky3c87Upn/Qnt6L8OWyaN
2ljKI0oXs+1VFfYXmNqnFY9TKKlqaCuWrdcZg1OXMbEiE2tPVjWXoseeqaXwJ2+k
jG2lA1wNkov2dMu8q1A4RvT3ywitzvKfLkB2C0h1hfYAYlTZRbU91dsnUIS6t2Hw
g6LYH351/3eFj3dYW6N2arRXZ3RtCAhdDgUtyQejrqBXZbsymL+xQyp1rNoDGqdU
Gnv3UNZoojIIEU3EGmxRbilHs47jsOkEmtmdr8HjYNDQZZJ8+txWw7YMsW9l6+4Z
fT+1AlmzH6PLJapwuR8I7RlI57Qo3+AbMr36rnQ3cqdKOa6zsSS/X57BI1kvqhUt
4FMyfBfJMNROL6680Ja7M3axtoK9/Q5lioiCqpQ7AdaB6DjMH8yUnOewUzwxd1OD
TGpdVy5Tr6hgTtXeNwv4l2VQ5WCAmkAJyFYnPvjIpVLtURCxWWv4XMMMFSWhDGOx
Ptq0UyGIIRBsNgHMPOpQrJkQAfsIwNiSZq3br4hiXTRnm8RLjst7lghwK5VO2VF+
7bxvXbv6fk+ats7llfp1bhCa5BUIORg4WnJ8GvDzA+tJntlVF+biXA6bekeYlW/E
PfSUlfOivBmKsMiApO212i6fimHFLT0xdzAqUoLicjiR61WO3KRAjtS+JNw8zI3h
Imp59KMspv9mcoFy2PEY9DW5Hgvd6OeHg5xeuursKcQk231eXqdYR9ZZs/AccZPB
yWs2InSoK1AmTQu+mAPFhuPeSt6I/qsYNIRG8gJZMoahx8e53sxiToV92FRtPvho
wHDpi1VKdAIfxz68cyS0tR7/UUM6RVrzNn3895DEpc+2ncsYtar1SqJkFKHUgLCs
3JW2SP0SqxxcSitdq/fop8ENUHJZV/khsm0w0xxW+LLXYgJQxpEyhgV/hg5VcOOf
Hw3/LOnDAk9nmzdo9GW9WVYOVZNMzFCYKYAwmVLcmsr4/lv9NdBJjtvn7mhGP2yU
fS0xmiaFDUnOvREpY0dEf2vuIF15l+rD641rEoUtRZbXDBUUhM7N8uTZD0/uGEGk
gTW/7OJ7Moe/ztvJIxUlgGc2J20+XtjQf7EDdeJDEDW6+QOFqQONr2tSV3DLx25v
sXRi7eWGvTXNdqJjiR/RXted+LhLgQ287tbq+lqGcS+j7I+zr1qEfKMXqm81pEBM
7WPONK4bu+d8PXfurneqA0dk3IWwbEInv9k22Mre7wF9yl8nCE6soRkbN0UO6k4H
sbmyBb0+MBUmz8mhMAAcdfALEOBGeZAiVWRWnRW80083iDgwEeSz+nxXHZxLw6x5
vm0NrHWSPLekb87YBO9XLxp0ZrzZBUXCg5wDHPrrQ2tyz2xtFLsRC0vSF/r48Cws
2xlmNvAv4yu57CwV7ZpuYLTikydrgq+mzcvilNu3LiyXAYAn1j23DYxhB514qXbP
V/rmc2Pc7om8VRO5jQaojFfazX6Ee5Ro0MlwGjf8j+iScwcUtLxv9WOOp4TVOrQo
3Oeeotsry9A3RCAx1gMo7hiD3qpiomox0b3LMU4noEO4TT1WDIT8kMVJO9ZFLVNW
xDe6C91MmesaMbtcF7jU3odSBb5+Iq9dYt/IphX09IhSnIGxif91a6yXZn/iA0gJ
436FHXXxUBXOn8P2j631XUjcy/Rv3TLfUoN36t2ApVT5yslzH/wo0W+1ijwkDTa2
SlNxyIAA4c8l8hEYSbq+3N0qwckztffm+iPnpUUEQzPvMGpFTZS4Pp4eB5leR43X
socqjgEtmqQY5paGeluBtOPb0QrJ3mmA7yIo3Wv3tOCHNOuqYeuLE5tMNfGlyEUa
DQ86eXeOxnLXV4VFxyqKkQfWZCRKtnuY3Mg81ciXMyJ0L+CS/uTuxZnMbam1sWsJ
wQjRJnYduUkPU+xBG11xQBu3kfz/rbP93bTPt1pAAT7ZCD6Z6iNDOHqFIpmF0peS
uTwUD9Gm2b9GJ5c3U6z7sATwt3yE+QeUR/AmVZ/9SV9p9c37pZZTjljKkWXfPQso
kzk2hsCXzlpS3VUdnrIRLjfBwsoU9Nxuyys4jyLW3t9KdANidyIy/U+aGjcPwmu5
UzmrC7VGzOHJ04+7obeYpGwyWzt3Y/chjdymhPxAY3hWBYMIpIJDgzhZg4b8PAW0
jWQig8jod7dCQxB4DNawf7HLUDRfS5OvkM60RCvc16AiBCpKZarfEAR72/02wKGG
xMLthhHDxNGfyErCBE02pT6vbvTftV1YXhwSZ2L233l7ZAMq3GLScLIeI52r+aIu
MlmvcO59+uZaE/pksAO4IcMIAlWAngV6X0RJjoff3yj5zuLDVl60STAkLqFlbxgx
YZAg7zkTrX6U3+Byzqvnf7/nMfexr4yEF3RnjuzsIy5MEB71EejR8PQx3wOU7LwF
nO/4OZjoh+bbCXLLNflRUDa5iQYkwHJEU7n09DvxYb1rUwMcyZfAogSo3OMOaY7C
rFNGmH/0NXMyvNWY6vSZLPCQaJJg09leiRShcSaunCs9PVg6vpJRfaNIpvB3C/w2
gol3KvYE8Svp0b7sBD6NmjjVBU3g8MrVXmuasVr8Sg1P8NFVDchuDptwza8On+Qd
cZDb4Ijw4BPQ4AFuNyCCIF34uxmCHA1lSYXgwQIOqdVgp7DahOfZ2mN9zTz+z6xv
HkFwvD5/oxu3/YABBwYYNEZx8jrARmPAAw2eU24CGCrVHxozpWa9IMFOclc6rqzC
d/qZ/h3wr1mOePQNPJbQWR3rqOUxwazVFQH+y6nOlzJ6H+ed9uGmviBvhoZWVjCj
bNqNrA+1XyGVTxZBYizaFXdpDRciLXgN229PaS39GLa/KgsMlVPeWCfTrsI64rPz
UjnvW0JYy3Fo3li5IIGhb3RnLT/HA80X2focWqemC8U=
`protect END_PROTECTED
