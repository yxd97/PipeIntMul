`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tucdc/TH/cvm3maZvwUM/3je+7Kl5pD4hA9nHoEA3fimi1+v18AK92A73gx7br4O
D3AzDhYcl3wy5ZQbYVxOYlRUoNqLiBpI7q1WWiAJqzjsTS8oiwNKYTmjrGqGFdbI
drNU5k1HpLvylVmwDsY05yebZiJY4jR/DUr3jiDA/i55dZfH4ILDSUqT0UC7MckP
5dlC+bW4n1LrQaqJAB9d86DH+c4czLnSXQpgFKPFZ15EgwOquBs15/p6GU+frjnS
9kFa/0/UowipgilZ0AMw8ZtnaeXg5NFHiQVZPbIX32IwG0z21qge15xeV+8cdyUk
pF051mPUkhw9DdUFZm6HuiU+RKMzGPZVzoXS0rkAQ0wPKmTMJWcLSkjn7KEhKMox
p5D/QjeAQzSOLsihRCWOWwgbb50jjBMeJv4pz8nQAvl8mjNfID2uiWZNSQY7Wt3U
X6UeWjsVwWvjEyCPDZBqaMujDXgVqaUjMEvPoWxkEokvMRll7GJ45h4llCfCbYUI
fP+KpWg+nbsuCFzWbCX6ejBJpnmCXwokwwYfS1Ef6XDnw+qEN7ujXW2qayTycQoK
/t6t3cwBU08pHCtt4gBecyNkToNimADrEpZK8ljR1/xXjRNX5BxbShTS3T+YIIEs
MCR9Cf05IN4r3v1LY/FLzrY1PVjkoLb+8S5fHGqJuzkvxTSBzgUVpLpzhWkSccQ3
Qo6HAXzgA8tH0GAd7oQvWWXY+E3eLR4IIUOuhxzUcLY+F+HHsTx9lXGOgFAB1BCp
DYiMhVZsd6B5sXFYf5LPPRgIUK/3YlFqNUb1y93GumQBoDVZ2Oe5HM1h4YGpT5hi
4GQOqOXOciSXXgsByWQLiqljkKvbQeY1/vq7tOMqurgB4qc+J0XpoZog3QOEM6D0
Pv7yst4fRJs+CmoLw9HWEHFBT2puaBn92VbC24bx8rVXmBjGD7JF2xiFc4f4/ScO
bD6kjm9EqnnY8ABrPifVe31gTeNe+55AmZdy73UBt6LgdDnW3s5kj+wJKoMB6qFG
lgdA4etx7bJsDskHfF8bohf37I7Nrf1OjdoUvwLTUm5B8MD89E5iPAvaYTQukJuA
aJP9OfNUJ2tOaKBH580uzQUy02HMfbWMxIHbFltyMW+RENZr81HbqsOKn5zjVuw9
a4rx/FzmO+JNkemmzjuOHmVSoEn2sFg/L3XoSFLQu8ykbud4wInsvP3URQlMGc/n
xaLFA0Qu8TA9jTh37RMQ1opA+0euvFFUNofJlSsrvI3gsy+6+Q8nrtC4PpH1wdV+
ZPPUPf/HD5T7lihB85Yg9YRoHWMPoHF9IZFyuh0/f2fQXrKsZxXCIV+foHeCx+he
9esvp6YuIiT1EJhdPGH4wW+juWK4J7ae13a/SsJLYmC31Q12cMD8/Ji84UE3jm4W
eOaQY+cg50RN5CEr+Ja4h+AFd4n658oHtyhttwmrc0oO92BCFLcjPK+/Mw3UBVPB
6uZ2Zk4fvrwWJ2uQXcBSaXufD46IWo2n8vmY8t9kEsUERc+Tcu23/wA5x1AnWAmY
v1LJBqRQJ1+bFGcbQEOcDm85O9FB8cDvVxS+vv/XChdTqdGFe2PM7mmRjsUEeH3L
31V0RaCG+TsF3yY4ZUNgwtUuTXw15/8UjOIP3BmGU0PgSnSO/6SIUc2AoU8M/F9J
5lftzYK+wdb3UbIfhNhEpo058bdAbaZLmdvQu/YNicDV8VYUrRjiMr1JRQ/NN+VN
1HOpKiI0KhCsoyttllHuS9LR+jKjBOGCLgUezsuvm26VaatuJLmXjuUpnEUi02VA
zDKBVyFpUHuqEDzCaI2ow1g7va3KfRx0zRsEOEsJ5FeaBeYpw3pg+hNcVSOlY1y9
jKgPEGFGaEpzLcqpRUi6ii/gI7fN/yPD8Bu6PPyUuLZOKPfcGjcPW0jabtcTsydU
U74brfjGHqjN0b9H4ZJrDblR8MZxrROoKVYKjsd5qj0kSAwwAgLtG2uDmwlmIT5O
fYirElzlftwVNgv3nkXJEFtHv8RJkGR5jzlRMd5IJJN1D1GRkWCYwL4VeE4dk9cK
eDL1k/5BxyBrkETprjNuLtE5bPkYqUnTq2tJ/Od2HhNU2+XEZwAS8I+rXlr38Wxs
8b0pPOZz678Loh7+URFjEpmJpgIwqdzJFFZ2baelhYkVPAGA7H1RaIURhFIEmbwc
QMSXuFpgTgpf21wXZHAIleDMDeMTcspRPw/3SiR2Z0C7GS7psX82UnTupfDcdu5m
iKpY3Wwb/BE8UvgPtUoA/C8YzpAzqghooQ3P6g2Zrhh9nL+MrQi443DvJSo2/QhF
oAE/3nW0DSp48IuV4i7Acj1txQCFTztw6rhr7qkJilRoh5SXpNhf1UK0ub8e3rHv
Ecb7yyIhsyRGuohl99y3a6QaR/wxvmm1gaGmtYU1RQBMM0o5u5MtzZwl4Xr2kVMT
FLuA3AQCOFgqn298uYnd6m6RtFXXcwoRhcP1WAg190WV9i0Ifsj9WN2+osJyBTCM
rZDX56NzqmyzrzOrntg2F6QsIXzAa+2J7GikxpXK9n5d2T3VrilzJ1GvChOUSGvy
34pJzl412m08ZMRr+spRnPKKmCGUwzvCAV3ns5sfqWQgQrYab720Nz8taPykqd1R
XqeTNy4fhyGz2C+9aN5j7NZr4KsQ4hy0QI6LoMjd1B3vCsJM5e1rOEK+tHk8cbd4
0pJltGmfssuUeLlanC9sozs92rbvf4Q4YBK1RQLQecZHNUG9Dgq7ffugTI/k7qF9
esLK9yzukzlRTp5TU0/P+EREWUQkbKOgIZ4HJSXcq+IrAv/3CQ5ylt3Hy/+qCQID
UwfCsrSrmYoKKgnjPaJ33skqryCy/5hRqtMXaql46whtbRi+6COpA+JHwNHLN+Mp
ZpA254xcE4jbw7dY/2R+eN7pig6k2bUAJtnGfP2APn8K+iI6g1YEJs292pPdstK8
W0Zj01pHelvK5z3K8HMACeMdVqDw+z34Bms7XF1kIo4mngDPdDy93+n0JU5gg3D4
nPQQLPVGZoNBczGr+I7/cota268X6F3J94yFYEmGJCLY2tUvT55z2tWeTKE0IpBm
Czh791bfdzjhJwU9CdbFt0QJK3eDaJwlINFTYSjKOGphxNJHUfG4dv7abcjT5+Uo
c6ri2mxZLCUVyGpvOSd4q970d3aOC1NRwzBGk1mNZ5IgwNxt1lGkdDwBS2/sOnV/
xsjeKTuOrPtnRg7FWGULZczkOuqIuyH+E0pOsL3/N81gd/6p4iFOfEPio4NA1Oyz
0Y3UCG4Nuny5heRJRg17CpHLneE8PoBwrDnucpShIk/IoSqO1os77pSi8DUk4byA
tTYhE8fkRI7zBPaUGEIrETRYCNucojWCiBEIN58zOH3dzzIHUOIeQR/EUggPEroZ
IEgZmC2QRcQ6+ZLpDj8cLb1o9UQpepuDzzGiXn4t7uH/GBm1UMj7cHTaCfKoTJsB
csEsuHnMIWh+WvIPFU8PzNKp9+wr2piXjGQO9LlUUYl5k78i2N43aZVuMrYWa0Bh
ZlRxKCl15gqdImHTwc3COvIyW8brBJ2HId+IP4bg6drbzTs8A7Q3VVdEZ6FpsrQa
loqcHYSixZ9S9rfTIq1owHp+rUhofCzACvz4bQPHU64gCsTd92JogP5lihD8X+6p
NddWQ4oH3cnxDcM+cRYxwR1B3PUdLWUaqzJPAWFggL5+38oj5w3ZGiHEURBoGZqu
jgXAp0WcuoxoqbK73bcSz3RXlNdXxUTHjnRGo56MdP8ElyCkzgv0O7dKCqjRf/kh
Wq0G4077eKkL7QPbDUJJDjrgy65uJsMIQZpFPSTowqQvkAuEjfutBVmCVcmkLSpN
EhodTA5kJbBuCAejBtnSrDZosCa4rZ5bEJzukNIdnQXS4mKmPbdg5egGREjHK29o
7zcK4UUMZjVlScF/XRsZsw==
`protect END_PROTECTED
