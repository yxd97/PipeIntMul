`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
muI1hmUti1d699IE5w2cY5STaHHaoq7I8cvHv5ZAE09K/2w6DUf//QjgWvc8EYF2
tX/nkO/vP1eJm4apPKlzTAuVmiESDTzffFW+8JI1pe5jxn/MBJa2Ant7Wrm0e5fH
iYoMhmudATjXiXIVas4Jf5zB8jU1Gj+jERnMXds5qWWHjGhReYbFmyTO36lKCSGZ
H4+5XvWgpcPv7y6q+9Iz5KY1Mq1zy3PJ4NdLvScKqPVjfd2VWKPSulT5dtcSWvAM
sk6EwTCAwKnvc188xJmwkeFbJery20MSjFfBSSCYGu2VXjybMY8KagC9uiMPgaMI
8xm1x2ssXET5NyLmAGvBaf6YFs2uxN4PoCrfmLh+6nuTk3qcshouKj0mUpSr9uZs
9Ehgo0pKMRDojkx897iwU4OYwILItlrWJP/8QSyJw6jfIXYdwX8cDwrYtGOxtbO2
M3n732PKm3/UqCfB4cq/SSs9Qe1NS6nHDI4ufoiswHNhKSRYYqxeUrYg9nu855dL
NDWPS7jRkuMyCMJl3mE6k9f/Sf+CswxbizFyZMhkgkjv+cKOSxMXAebC4DDDZ2hU
`protect END_PROTECTED
