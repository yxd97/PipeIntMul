`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7o1gtp+gk/VqYqfBPv77Ui0v1IlCm5tjjahJOvaFm6//kYeBYD/slqVNAxeHNEZ
rSwH+zUrKNAqOwMLS1RI/q2BQqMa+c6SkT5QZjDYpp1WqsLLtgISFbS0AYsSQh+K
bLt398OGlXWt95DJ+aVxcNnQ1pO88xM1HzlZ1YtDUOAZYwy9/V10BySyNr4s5hZd
8CVDWz57wG1C/PzKeBS2nQ==
`protect END_PROTECTED
