`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p5fZPCSiC9QrEfL+lZOncGW8NwJexivj38MBOhMhA9aEiTFW/pWrmaEu7VRNZeJ4
i4kq876dm8a8nvz4hNXw7C8ibJb2hVnUHOWtvOkMCbLymOdFkNGtSAC2XHJFarMx
8skX7IrmOIqE2p5MTeGeOLPlBUSfVZHdJP2YSH9mfMLgYNg81JT9aCFE6dncETl0
8cMJvsZIcw+jriTkccxOKIlCCBRbb20VQGYHj+SJSKd7wqTOQPQSwFsJCO+Lq0Gt
GvqDIuZJNb1MzXz3rBRtnQUQ3iOBLsVjWmaFp/YKnAtKMr9sA4MefCQR+nSsM83x
6uREh2DSmvxqHrXeO0buvToCtOO3xqp4ODx+lt3lhbJy6dTJG4bigR0l0Eaat6ZV
Skh9sY0WcYVeSYJ8MxFGvC5qnsuuW9/2jJWitVHUM7WcIVXshb7M4mImboWmMuNa
TsJUPdShmO2ejSKzwbLlKHLEL5Q5Tr4NyDL9h0WgE/TPVor3vA/xs6//hvjQ/lIR
+rHNyzgiQEwkxOuCrEeoBCcQtqhNSDYrn2FK/2uC7yIj+9IoakpwH3Mjk6Cjeqwu
douww/XvjxnKWwcgTIMizOGELdYZiRDt28Q9Raa1LIUJCkrOyJVR/m6f9674IPZx
ApAj4Zkrr/UPK3Dyhaw8CCboRzUtYOuUBYiA3MGlCYIEPvlpLeYX9e86DCcnmPia
+F7HFHdcVzVo4UypemrPd/QMroxlJE40y+YouWeTHOY339fBCvA4Z1TegIY4lSMq
u3Q2lV9JtVXyJhrdY5boAwk3qMm4AIUYdZPft0PRa4kJAPWNZBiiOrpu3kUhdU8s
vj3ZVh2Qp+dIRA6EJSF0lyL21WDx6hepq0f8dxYCYcTFCASeXVyXdoCEnJfsFwCM
C9KCHh26+8Rf+OhkEMSpvlzjtPrjajXzlInGuAvizl+0zeDOyR6LpxgJfeJuhA4P
5E/hkIpQCq/Bv3yFf21SoUqlD4gWVeoRBqkNp4YkRhcKj9S05b/FDrC3YEgOrzUr
OVbmV5pEPLc6xbSj2eA3Jzsytbi9KTqFE5gCr+aG9T+ZuPOK4emMdAev3/Fh18qO
FItUS1xKGzOlapMolAk4wBpsSufvrLgKyxnjx/djN1zNxnK4Bsl3xyBhJ3gR3bFu
QfNovhdQvORRhhbBAltq74vW9dYEoKU1/7qVE6RhM2NcBDtxqDmRve9TzRFxUm+/
0LQqI0FqnVnvk3Vd5wwr4Lf015MhiEjk3eYJpwiol6WVY7NaeGJDkYAexj4ZM6Xc
6E7kle/MpEXreTsFx5A2xPGZ+0EFGv1hgOGj857h6UvofYsrpqmuNfDU9cj5FxhM
nlLQi6jBXAyWISxUvN054CEGc575a5DYZPBzVo2y83jMJkVc6mkj4qj5CQi7JvoS
7+sXUA6NIFOYW18awosNRI27OHi1KI2Qee3MPOVFtU2WOI0/1jUAPkthB7DSVR/L
dbS73RIPqZ7BExEuAPDtm6AnwgpBYohyH9OMu3OI2DFxrNfqsVAn1Fcwm+E0uNJx
6mC8FuSADvfXUlsAeuoygazTYKSDmmSXEYq1r0ZzYoAEn8PMI377zRXW9jyYBGmX
FSIw+i6PCKb9aBtc6Lr/APOsPaKm6jCp4fmz0crvZbUS1N5r+VCW9DeDCYQPiaNH
L/XKnZLTA7M8fxEzRTBNYDc2nUY5JW3YZrg+mRm6tPJCyirwZfXRLUZ+zInfgccJ
1KTVWFT63vnTa+tTakeJN5gCjporcbemMAmuOa4/MzowZCb7Lfln9KxREillDf6a
BTEwyfmMWnOH38h6yx7JoVgSrtRj+j1seqU8z4D21xfpl1tOCsdhC8BmZZPJ5ya9
MjLO95lPtJ2mw14ygh3DLXEx3rlDk9lgtJniIyFzNwvCPUokLBCGimrZjWNTxVU1
QWxwfhQ9eHrySnY853M6laNNMWbZB7VsBQFrAL4xQmbj8fLaSrUTrxZM/ZmmmMhz
0TSz2OAEN/pwUFo81au+uPtpHudxdH1yVi9/lH8lEvbUzQPnHzcBZK6GnnOIWqa8
gJdup//8YgeGZ8/TNgtwpGNnwlEVQIB4W31sAz+YkbJUfigxemRHjCRNYLyOmcDM
36HbvAmQ4tEbcCAcpLZn0psaRnNx5JqEz43REd46TT/0OA4XoPvw08yW9ZpQbTrK
zqXbR1LMYQmpqb20romOcVqP/bbuPNvTCu0/be+JeCLQadvGOvcAZecc5r22z8VL
+tc6u2lCNDJqYATkyeib+cU0j0b/3yihxVayE25U4cHsYMV/FYBgF6usOrqUhkYz
evkpsZiuxhq0u7szRCWPMKt/rU2muvVX1pII/mSEEFdrH0TRF8DnvFr0YEakqsLa
WAunD1SEqklJvjmF8Q3/8gEOW9KivDaQ1wVg5ZlAdFwLYTLdk/2vSZLyJdv/R3c9
ZoxyW/xrh1AtWMkph+4OlsKVyfQeppiff2D0HmvxYRv7YBmMp+n8Th7G6CW6EFFF
lazFassR21grMInvbg26fuggrZEEqIzRphdxmd0b/NM5rJLp46JfezRUy3nF7kkY
dK3/NxfepExDHVXtwwIu/SaTW6JdlgnmI/5xIeiRTndgdaCjeQ+lrBvbN7X1L5LN
siABoXTTCDSJ3Z1UJxSd0BQs9D+aGeMP5V9JJh3ttvyU0KgyIfaGzvSetuOeDqv9
zG89O06dHCO/80auHIrZPm5NsAySmwhzBx//VCie2wcWECq9GKJ7ErP/SJENWDwS
L3rL3jA3XumX2VBCrFyY6Vs9fBVrFqpLpVFi0J0iSXmx6kW1WGtmacZXeoG4j3D4
pFwUxboKpITwn6kCE1MJXamqB56/Lu3zZ8/tCPdyNd0rbL/Y+1B7O1hhWPXZNTpH
sQ1LOMpwJdb3rMxzhb8kHuQZl1i0P1kYqP7+v5GFsKLOPBa3l3RCgE0qfGYcoyw7
ZyyBAiusTbugOkCoGUobLRcxaBT5174LEm7tFtZ/5Cv9rqfgH7OJZDt3At0iyPIE
81bpdKCODHHnHeCTOBSyBuNxRfnl5oHAaeZN0UGELaFth7VDr8xMIy8zPFh5HnKv
nON6WX570CPL7ynYkG5VaaXmU6yc7tLGsO6u9Ec5hs+mH9q1bnohi078QqMj62ho
3XNZKVPkUa0DWSSh6GN7G7+eHoD/iH+SoDQQTRKdoybc1jfB0PTDYSnePTbHMD+E
IlP2K56biiZbOVrtrxlDYdiOztYjk7vsFqpAvWyJPGt0rkjTjQKa2ETFwkEWv/UF
LwZ6W1eZBB0/j0BCoyrIgTua95ej4KGXjGEQNJLyBXvdk1s7OIHH+ryDaqWkZgvM
Wbn+c1tXiHeTrWxBqKoRu7PR8Xy/UWTGyQccFoZelhFMSa2puC4aFNsd98cZFvHG
6Ir1k4GC5qh7MlVnZGhuJA6D9oSPgufyIw0YbLAm03agxxMESCGnKYLlBpYP5Tr1
ER+mEOHLdC5LIybuYw3J4QQamPjEaXFV59UFF/ZJfhcN/qq5rbL6CgH9rryIzVpH
Tyj6ARVcwOFFML9lFIbyNVfgHi9hP/nrZX+cyT2pKWgvZfese9/mu7ldYtv7j+NV
8MEoIlvDpeqY5Bxp/O4I64oouaJ+mZobvaK/dvnE/HsFOee4KFkSHfD9fM33csEb
7od808syv58tHMzMdZGUTd/8u81kTJynfIqnHIFxUWAI1QXZwVT1Uvp8lyXNJUD1
6q7s3dsg+pIqstf4EKVYaeef01UXIHZuMiqsN/7He7tvwyxO1yxNHU6DHtA1HboM
RwbYU078kyZo6B3ypP2j0vn7gvotJ7jSweJXvVbVK+0nZxLi3piuJeN5TfCRv0sd
4YnevVymh0oQZBMnwWYWNeygRaMoo9/K6wGWDixCzcPoSN2416NHZXbjbk0rvt6X
NmLj5djpzLIwdPpKgwGGRywOM/sqrTXMiWnoIjgfVpULxNYYc7E3GOyHKSXl+5ab
lLtTE7eyvDI/aFzsTSUaRKR9WlkLOsCB21ChrfsXp8R1X1+orrNq8viGLK3hFG+V
fZ+RQ48SgMq0VHCG8tLdRUgrzOX+kvbVFta+oik1ykAQR9LX3SfMLMdBKEpSlBFr
IqdfbK7nuSKDB/oxtplMJR1CJPQv29eUF89cM/LiXQ7FFCZocLr/QOhtgQN51CDu
C6C6wPylaH0Mh65ifgVuIrWwA2uZnXZliUS8rZWEWOHq5MgFZVM4M8SLc2om9Qkf
Ln8C0BNok9pLmshXB3T0phE0rb4rZoMUrJE5fO9bL8AovWMsn/wVVbUi+Acv5Tn+
EAbdK79P3Dfq6hlNnSGIgpQG3ccBu4uDdQm3MrEsic+9lYDcl2h9PMzUxAIzcAar
RqCvOy0Of45CjeYvnXkd+Bh7WUvrjZ65wMCHW/BTC7/E1UakyExWbBQQO8SpQZtY
TWZsLYkiQ86boIlNpf20EtIZCnkVPRnZXYarVHRodu6NXBGcIE+gZ/2cmZci39mk
jI7wxu43QofC40xwxKMuQEA5MWN7k3iE2PnwGXVg5asniFK1gGZuqerxSaH5jbaJ
fvnSHcgjKSNEjVB8Xb0Fy3fHAgWDRIPbqpTopFXJDqReTvXIODl5SMEBonO0bRom
Jr7W+kswVeRwyZIVzWxIZQFu5DCbcFO4egzy1SF68PXrS5E8AcXmspuyYdjRcf4d
an9KTdo+CLg6Ff97k4fyCipXLSwRN+ZncplinrsgfCPoIxZOIM6lXqL8+s2k+vFV
/RT/RzVhWP7ahX1E/tjRnY52cFajbHkVO6wWkoLUNIituG30Y7FHs4CS8QXmfosy
QA46Tkw2esEBI0CO8wrq2Xc6NQlT+tYXatMIYI1nDGGaxHq7mcRFq0EyNV0jmQRA
8cBuc2fQxczoPXX0HENXr7HP83eDH7AEXuQOeawHaJpY8gb4Y/+Pws0W1JhSTfQ2
Fs195OP6aie01hSICfcF84AT5xFtm1wrqz18cqGJk0+jiE5fcqqYQnNbkUiB4mjN
0KuC+JtI2YumrSdHCwn7AGOYI3YEOebruFseRG5K7VKax16zjzbXQbjYacr6ONzW
1RuiqCL7CH/uorlg3HeIkC2iSuTGkVabiIVKa/QdKchKEpUDtX65vKXEJIZ6LRH9
8b2r6ZNS5baVZ+TrD4LxRlEiR33EBQkaWNYaCKXSnqup79FzeL6mvmZ7Z9aAq+F6
XfERvp5k5Tu7eBm83J3buF1eGlNfnjcR4tljBWPu5bSSH2Dusuvo22EfACfUdyhF
fhQDAEMCbnLQYybjMwLj+a9YS4KDeQ/Ge4KmZwMdghRgmE1e3aCHIQj8mDZhl0P0
TX/8tyTCiytNV7XQNetL1T9lVXTvSlWWTSRiZfkiRA2HArVWMQsG59mM5PsmDOab
CgKD+Lie6lhwS8XxN0sh2BWSYXq8hgamZWMNIh3EvfcSOEzdnh+82x2XwwY5PU9x
xMYyYszVtj98tjJoGEL1lnvi+ndkX2IoF3cy34iv3wA/lC4eCLDyO2tToBCvAVqc
URdopfz3bnu9Nsie8vteHnTAO9qBwEy+7SCOwoDwWN99cz/soJIgIJRf/b88LAmG
OJjkOzG66ndW2dp329NLziDpFPTBGCiJ/nCpeRwQhUcDuaJ6nzXXsgqSnO185QZ1
gryHdpGecdKxj7XRQa0kIgcQbmc3vTBFrkMdcsAz8/vjeQDuBMfohyzqEXdwGPKa
VXi1t0oG6PUIRLOtsoP48QLhsPm3X074A9Iys4InPtxEAXngpn4NJMDQDBON5AvS
u+l6BL42DSmi8yLlJAQSMKWo40c24FZ/mD3msoVvZ5n3ldX3Sa55CM10SZQly/nP
ANq91H0QFRXXzq9bredBLnV8QX1w44xEZs1IcnuV/f/32f7/uUoi0LeS90UQXYFJ
XcnNvhmT1aseoDa4Q099iZq4D+ujhl4Pz30DtWTrhPPQWOdS5mPPB353gEW8bOW8
vT5fnMozrcn31ntfwflR0rYGMlckeLTOQ4G8+rwH1ZW1f+ZyllpbwFQbdhhbxaq1
CBpXjPq8D5tVFmFoe5/RnyejzQr0vzxlgkYtKKUaOHXiQ5eVNb/oemMqOmwYyOmz
bFmQWXM5rRQPvzXE1keIRsiNGu5WF7vq+9SgWlluiY8dw8xgc1Rj0VeLwvWtIeQ2
a44JfnavhZXq5Tec+OSLqQ/Zq2/e6oXmIDBnoeNM7Y08aPWN9PLqTpRq1uyNejAj
pR1uzBz/cBuviqN94itmzehGZpSLNTpsOuiIODBCf8fVE0YbOe5PY+a99ZdlBOmY
/NC2oFxDGlwhj/gsjvFXkYcdzye75NErQIE85LMQ7aZf9ShqTS30oh3aPJS7phQt
vVlVVA6TUwykG8mVxvguRwIGoKfokojdUDAocP/uhp7WJqOGhXo2KmAMiQpK2N1F
MHRwVpesWim2lChMzI5/bBAxpvUvAWPcREiq3ddgnITAVKhsnSoBcorv0MopKtWq
LAQsxxgtw7e8jCrw/La9Cy95PoqLnjdGmCv5csfCqfOY6n4bKoAjGRuGZem8WiyE
pMpKms0Zmun/RaxTnQ39GDVAL0Fnewsxsr/q4fTXEhpB1IZeCmS/TpPjeb9ixZaP
WyWpyJUSWVCXk7pIY1CgFsXfhaNKkblZsqJHiQQYpj9Ha7Sr/AyGCAALDrf+1olL
m6CpOffsmoo3BmXFU5WOFrcPVg0yOgC/z7zg4SKAEUTA1T2ogf5jlG8De62qugwF
RqPTJEPmctDm6y/HhGavOA8tuSgr2MOHGQ00VbvnCRAD+Hs99yes/tiNvF1JXi/c
FXz+uXokVIP/ZOyuOQ3AxCK4T1mCwpleZLL2QSgGMMI/nBBqRdQmPiOMzlUAxIIv
S2FEF0iC96hR9mJ2wbHSyNfrUkQNp4sNdGcv+WIk4qDp0TOuLvV6956Bzz4Nr189
yEMQ7kEKjaQDEX+d55qhtyrwOGh4A3aqtHBGlFS0p3MoeOU25IAGfzO1dOw4Lu8F
Fd4Ak3obR3sb3xd5c71UIaQZDj28eY1Z4RryZd47mTEt0kQsMtjdKV1mhVrUlHwb
dOgB9jxSZHKTpZyz6adtJfRn3xKFsSPya0M//6Bj563Xu8zSGVIRBk9MGTRuRksv
CT+awey8nbJhVDGF5g1rbf4zL1BM7A0Ur/hgF6WBf0EurXRZ1hxC50K0Z/S1RCTU
SwgskuaVMLHOZr0KR7kMO9tZIV5kP9QGjAI5BhZtvmHOD9Yym21FsbAsO55TvQXG
hxzLIIBhuOMJ3Vceg4AxBRxtUU7wWHSECHIcoHXLwWjLmsxpsMAl92Og5A4V+twm
xmt501/KYTUX/mwneJFtBB2ULN2ra6szSVVNiKUYR2BuGlSogkxnqfxpFmGpQRlQ
MuzrTFjq242p3jwKuwUZ/s7NV+Bhsmtb/CR+9didp0HuyF+kyYXjJt0OA1cKzcNi
Ipg3TLBNNUo3JjiaVV/rrfxEmHwla95whWDaMx5ZoJ7Ep5n2o4jLX3nh0Tz69A1V
XQPGAH/3c/RQ2w20xkutjUGmyUPmouwf1QQa7XpZ2drOaEyuEqj5ERSzYtstTGtu
YrzzYVhaQD5Ndh9QRv8tQfA0eBV9Ek3tSHyKnCD68X4Jim5LNQTDm6QMVoAVm4OC
jrT3RAL3cmO6wIWa5Tl5Ge7S2X9CCrx1JTQQ+istEacBuYw0Jq37+DQeduBL0/fH
fT7NY6BQRxZlxRJRd0eEPIaxgEvUpGo7vNtyxmIJdVjnCjGfkhTL0HUGO5otzbH6
4R3YP6X3HZZeFgzFpQ0q4MV77baQmCY+SpljjIVqSFJFCcsKoourasQlp4h0FOBN
lQcEAU+vAfIgfXYaQYPdXpVC1N9INeOfz0HHoRMtYTxLNP06UigIkq9FkulE3UXU
BCguXPriZGrfxl018lLvbiH/dJxoTqRQmsnwArWPIjaHB/F8wmnl9fvNOVVEMJHg
Ug46wzmnamEYebiCSCtgzs56k82uwX7pwKLA+qnN8lRUNIvF86SqseuJfKpCHpAz
vahvYzZ4ipzsLpmqMTtoXb4ghjhZs/mDp6+RzXlvnLfJWVRGdmnvOPpyQcaoKEYw
NFrDshWJ19pap8e9lQ5M3giz2vXSLTKwRkuw0nDPsHOOcBfrZ0bbNugkEYep3/fE
F2+ro7U7guA85EtzSmdNUD5/uxpEEs8GD0yuikNefV0kqj7akZj5lem7eU4FUS+T
x0ETMXq1lgeha9qilv+i1XltqtXOYXFFdGqOh2w5+JTVJ4AeRupIP1g9jN0pXw5S
7V9gO81d1vKixwFdaxpLjA2cid8LHOmu8pe/AzvRPvcjGJxBTudRG7bMYiCC5NF6
1b2Y1IAfu4OSOgTa1Bpzu+k8LK7B6UG5m2b9HcRW+LsZCUvp0mCHvOoWrNkJ7YDe
R0SMckkkqN1iF1pgY1fPSGdOPD3yPgHMoPGTHrbbpVwtFsznVBXZ5yNAaYxD5SxE
zCDK3pfqcOb0zurjIesZK6G2ldjDXCPOBiWZ2SF5vcOifBRj5PzEpNJmNemkk+oF
dZqYmxsYRDCucNFy870A/K0fCEEySOLNLYa+CGwRcURPVqh+aGHCoYy1xo6gASvy
8tptZvgAjSCGmUZ0RLlDGi9WjJWJifPRMcpTeB7DyqmDfFNFtzzPZRyZ3PK58VhK
kdmZMMI5Ayo33j45082NzB6CQ0O1RHJtevoOxyG5tjbyMdP8r3NHezflooDdqaZ9
sccDyzdEz/j5b96wGJKD14eBYSfaVqX/zS9Md4VNaBZSRx1jg2Hi4LKCH4TJKPo6
BYWTPJsGhn4eIzANSilW2BK68yhpyw0snudnhHpNDFK8forPkp1U+bSqL/PHloDO
IdnHkzhaZlhT3Xt20xt0mjM/K1EzvY1R2oASQVwPkpGdFBK97fCCV4eUIvH86VdK
5iuhKIiRurOOTYRRD/PmPIeV9ArmUA/ud4QLX0knl0MtrEImO9Tkkce1ZqJBfvXa
2uX9mKqaxKv4m05qfnvrtDagojgSO1phexiycZuphDKQefy6FKBlwM0ArFgjJaEa
zy8WohQSsbTM+0eBsTdk+sbIkTmKyfnrwDylNFwL39l5jG5AKcCUyRuUDPDIRWI+
G9XNvq3qOjPgJodaWXuGf6T6GxJGD8NdNJG3dI0AYMoU/l2clskAwcpWiiayPW3G
WNnT14fEVxtRtjlJIGiQrDtXw22uhWVy8MLa9tkueihfMbOexiGAjPbglALcdPR+
10JFVncO9k8hjI3oE4EcZfwCAFJ+N4XTcd65zmpaG0JoQPCxQtTfc6qmjXGRtiMh
pYdQdUzk2VhBUe++17bQ4wRTE4DXd7Azj+LlCuW5rvKoO0s3TDZGlnGDiSOW/XEo
Wunkh+O5fi7KZFC2C4itRCEyFsyAEz5A3gn4e19C1FPw+nF7hb++ibdOCJROQazp
rcPkNABTTVAWBQCZu37gE8dRAhkaAEe5pJlq61yjVE/vZJnQxtNTE8l02ayM5Um1
VRbmyUzZzHNG71ywFIeFzTVe3iNFFBEYU5va5cL/QtcPjoHI1zRdCxTLxL0JghqO
UW6DWWC+Ivomsp2/ZUaJMCo3w8sP93XqUOKKjQ9wg08nf9h9zhn9i+M0QHghOGas
OZOWFw2fBVHsjuusIYa5pBd7PYTyz+CIBip/KZfWtC2kb3ZbMF7cPL6A+3fzWhRE
uVLcATCsH89i+jI5XB3UTZaECKXQGQ3sSCTP/pnXPrOcrRkRvgIPock42q82EP2y
WgeYY4hgOqRa1WWT/k0U+2fr9DD22H4VjR9WfCUeLRl4FG9Supfm4eVRUeLfpwoH
4gvAjaKDoz8zMfSIDkIyeyzZgvqdQqlJI6BKUnGc5K+nookWI3pm3CrTYDrSmn4h
M2zI43opVz5+pJmcG+JcSvZznV0U4KJvgl3LlcQoGpp0XDWMWxqsjjdzvEgV5zNz
9nh+bb/TDkijaja6Q83QzKx4YR8EPXj9uOlPowfnYlkz9fHnRXcOpvdEayy2rLCL
ZGKAFc3Z31G/FoU3hUCQZmIpAN6h17Cnp/iCPimP6KO9X8P4sDES9O1ncnmP2bQu
3plab5v3s8a9cs0IcuHDG0MKU2S2K0r9NK9m+wyKsBJojLaJHAE5ES3+Se/V9cqz
z09hvcmx6Sh3o2mFkTjQRrKkJQqv66K5LzpGh06ro0qSmLN11O1CJPsdoxt2XCKy
SYP4777yxMpH9yIP0qKDiZ1fG1Eh4MS2bEfQDHIxKCgPhcig6ufeaznaZ+AF7+7M
FJUatl3F6OTllImGxt8hqrsmcyGsvBPNWEcidbShlL0E39VnLK1z4Gqwc0EsQ2Lu
drqsfC4ZHs7qJfSsuQAVeEJ0d60y7kY5dwA8yoy77P0yzt8CTjBFG1jxmzgL4HNI
T/dkL+PBUR+4HiXgW/GaWe4k05ZM6lbyY3TxQ5WN4BwupRmNAmODWghuRVtlPqT3
+yNk3YoqoKWkasBTYZy0z1DqcIjeALoeID8FCpiMzQR2jNgWFENPks4PcB9P1Vk7
nOezjeZotd9OhsPhb2oQEaiKL6236DCFKM5HNhdrrRw9tRhFQxMmtxDI+Y62HooB
Vyqf/QM1ORRl2b82GMhnG+zmP+E/rwb5okhT6BZ9AjQJi0ph9oEfHMSvxtgfI7Mj
3Qir4OPI6L8O4Dq5cYMohn6aZrZghQg3EcUcFpUVzFDTqcQ2WXkp8+tJeHox+BkL
ZeeRlnhibLTzJjinXEeJq3SeiZboGIDWzwli7v6i3e7G8SsuW+ExCEF/xF3kMd7d
oDQvMB++Oq5ZcJT3dA7twYfI5oK7a4FM5nnlxoefehB1q242sgQe3ftpE8hu9EhM
cL0bFae7W+1CnjYjn11MoVDq2nFgDvI9UA9QBakGd7gsXOHF7XDn75QeRzDDG+4x
eQXtGpGseQYm075xFqEu2O5Jm64IQgcWnAzSf/C+C10ZzYHB9b6iATQc3N/ZMyMO
m62X4CWHsS0EyxHxOKmBPP3m7Jeamrz35ayShJoZuniMW5sHWqwR1BvPg6cQp+FU
attCBdmAZZR0BAn1wU69DkfKPspeZ6M3JEH4j/jXpQQlQbzPFOMP+4Vcmih3sLfW
2P4ul6a1h+Soez6Rbn1JKphglWP3SINfucnm/DRvJIa4i/kVCDZME865cklDBUzg
91QNu+Dx5kNPWI7ARreX+fpgPj+X8GKlecZOnVyBPMEI+1tc741mm5zIj5O3Ib8p
4Dr/Q3kgL9V7op7QrMLEZRQ3DfnJd9Eiitrp+XPX+hApVj6PMIN74YNY3qQLnbRo
rvN3lqyKSkjmBGLHMj9TFgCBqQ2rvhV7NgDbYeTHqoOPE4fgRodhCmlu06/6uCgn
wjbfiz08fIN/DCzMnBsiyyet0EOYtpzWXND5DD5t8FzIm6oPZpxH7aKFngonVLZg
bUxqz7Wdjg9Mik/FbFbe5EC9rS1pMTta/rZbvHe93a4XFbX1XbCk3ZYRV6TCiKo+
uBBxVzQw4YSAmEADqVKmZh9qBTCPrtccE22uDFdI+rYOeqH7l6sgEgIvmSohOHyd
1+jFzMdhFY6CyWRU2wf/6lpfNEtOI/XszcWjF8ZhqXwPxBwWS9I/8dLqXwm3DCah
CRgwAdnM1IYohd1LNN9D+V35KCZpWZ5bnPUhaiwZw09OJSmR/Q2txKs43MAbJN4A
QGErzhl6LLN61PD6Y3TUeW1EN0TvZ2eZG/oxll8WxxKffxI5+WowxWQJVJfgXUO1
kHm2bRkQq2lsa9G+CoDKJgpubjK4BGi1LPSe1iVESpTaGLLSgi5kzzjSRVZSTB7m
iAElDHo4u4N8SsPsFvdG4uP4ENxBWVWkZyQHW26QkCUwKEl21iqUpTlWeOIDKiJ0
n9iNbS1+fLdePSYoslm6sbn0R13qbX68BhSKVJDR6lf+3D1h2dkcow93/ooo2yaA
SvJKC0vLJXGQpx2+ogwtpHV4Hq+kG9rLONcWAgVltGiEPsJkWJ1Y2ZdPXi21N5a5
cSOWosRXjlnCatvobZfiwIGWbx6lpRS5XKSp2hRtvOQrg2DdbcnTSAl4ciRSOmPj
EK4hc1fR6i/b9wjvcgXxJXRVgc2EXylrfMRF5q/rkHh5qEuSWYY5ZhsCyEA1YFr5
Bm3h5VUrgNyQXthQ3+nHzieVxayhn+J02T/wU6ADkSq3yn86ZgVR96LgsSrvuF7c
S7nxFNo8TsYyb/vvd5iq/jZsypU3+piaXXlDKGsiPwIOFe2D1RqJagNZLTxoh8mM
I0fT8mnRyr5wTSU2s/5p0X2XxsrLOLj6eIN02BDBV6LOkI0sAhc12u5gL2Jds6ox
SvIoYDpdfXo8gAqf+4aRi3V0DMUqJMimbFYZA2V7RS0BhJD6zm8PLSK3JE++abLb
uzlcSRn5Rpmk+pAO0uSsUcoIVBnK73z/t4Bxs6YA/4JfhVx8Ka7YVjro0ioS6mPo
qD2v5ZUxnMvjpAurXTQN2RQOOdcDDeWcOd0kn34dVXzxwli8lF8sLaeb3mmLtKdT
u3NhhH2/OBAWYgdWsl7YHjfbKxELhEq7MvVymEf0ciU2FBt6Ku/tVmmb7xUeMheh
dXxoOer33BklWgxEUkJN/HN/K6lO5K2wkoDnZ+Ln4ytsVC7kL3ghcDNG0+WOtYOw
I7cIYgBLyYGEJnxxp3fB0shK89OoVJN7OFIRKn9ZsTMS+5MzOP2KontMb+lrOiIH
JT32M0JMsZRafEgn+0bW+wER6l50mJqN2hL/AOuK1CCZF1co5uUHM9jUF4lEQm+x
qjCd9+EoOliGnkglXOo4o/o/RFqOcxOgBCxyToqzLb9XeuCeczZmkDeyh20oahDY
usz00eIhsH+HT6GGmNs3fMnvZg3C3exDNu7eR61Dwprt49Qo5Wa6LQ6HpFB6/DdO
it2rkwVPW3m8GfKfaVjlkIaXHnuX3J7lGv1v9UPD0hvaouYTBar2mfbA/tN+hEJP
sQ6f2E9310FeHujVsnG48uMIAs7FHFRBoazEG/G+wFFGi2tQaWuIu9wE49t/gr9v
VCS/8ApNtRIVMleLDQA+6Ux4JF2xeUsfTpi2QGYdiohhNzhOj1wU+cCc9PBU/Xfn
Dl80Oi2azp8v9indCzisw+WNYHbQFM9c444gM0pp8Hown5C1KykIS6ySsznXImJ6
AXhyBkqz3Hev3CG74K7QYGfqTAoSeXv1/jNPfRkRJSrmcyfF6cX7n876hgUeBYHq
iA9hFDfdeQ2zo/mPvTMZPm+vrMVWoDtoAbJsMEAuc9iAs7ypTRopC8/Mdd5HQIru
i6ay/NgKk1uQmLgAWDiWY4p6XO96g39yhz2CwoM7LrySgHzIVeC9w67dtfJvDr/k
q0NyQ16GXsotNZ1jbpXp+GOStworeyHpORMtr+et4nazESzUJofXHp3sjY5SNWcg
gJ/ehECuvI0jmKfaD/JiYLERCUJl6cYG5PnC81Pfo0JmGa0FZaA0hM+av2feB3kp
Dleq7apo7tH3mlbHI/ayMOTNWGIXatmgjAvpCCzc81UxNr8YQQHxHYsZpGjKfMou
asGIhtr6kPR26/BQFtKVpUBnJcpUZwb3bNiEa5Dv/gzOzjIiYKMmaHw9ut9AvUge
E0KqWxlK7i6sFc9ZCmWEJ8mTTpvaxB3mj4pNIep2E6RzEUjrGbAeK5bCNsppJqfi
90tQWunSNOEwcCDTkxFAVHJ6Ml1aVVduJWeLzNDeWpzUYe0SjW3b7KPpR3bm9TEI
i148YHevq70UD8QTaFgzZIGJXt+gW7MVFzFKGaSz8BMF3jaM7Ckdgk2Iu++ajZ+5
k27PseI53bkc0cz6N3vBVvGLrwQjFDdOjNO9yg++9W7anvmY0KDUD8TKdamLcq72
cvruLEcTA0tovut+B4rekfhAbXklGfmQoatYRz+rqB+6svh6kZataRGGh0Iprby/
bWUQYJq4X5d6NT5BZJf1WJPolBegxf6QqX9iXOK9YvXtQd5re8lMXnz0d+a4ofOk
KnwWbqt7rXzmlIvGHcaJzVH32aAarjFHxRY1hWwPzzlDpOe4kHkkK57YjByE6NkD
Cu2Ed00OrXo7F50iIGeRff8KgGiJ5HFgSmA1gcbfqcEmd+u1GOUzGGPjqDx4g7R9
tqEvh9OULL3X/OvhXvtn/Pb/gdNTv592T3UnMU7Li8brcnokgg26nIvsTtEIsAcc
wNai59j2mfPE7DeZ6Eq2R6yXjc2tx5bHiKuC2ca1yZg44K+O3EoyMzGDj3GkCT7E
X81nlhR/mgTb8FxLN2NSUlsvlbZlQ42rhYaDARZAOTRqYycacksFVTjnG+JP5hff
xryKx0eysvNdmRTKw2Zin8/bH2JRYataxq6J50ChEf1EGkeSRiJfVnVwwG02wuNw
+fl4RMKUGXbKhFpKUoE0PhKREgy9GwbYAntadaQAgi2JBxgo/m/DBKop5Ef3vP1X
inG9VQHerd0cnlHhocPN5IJcEkV0RdZkXsdbQO8ZnFrd0oc9riXJufzom5946lEF
g+5EpbVTPCvW54SCKZH/mO9lecj4E2JhjeJMVWCZ9oBwwwmwVlerezIa4dE+VY0j
vV5+7PB3NwaR7ZsP0ci/u5ZLtuHLzkYpkwgh5FnAMdL5kszuaMnjOU8jdTPfNhKI
mA41vTHVFeNLn/LWxKHE3TNUdMayx2oUpbxU0xr7FFf1h+/ufwBVPmA0spqLnDDl
8dOZIDQ8PBVI6olmTyuGTtjPDvNmCJj30bpcJnISSyPT6h6ZGwdTPFj6mr2G1osk
39R/+fnfLexpLUpjGu2vf7I01qDmqukqPSG5LOSjhKmtZfNYYr7ZeJdm9wg1v734
A9j/cExnV1wvySo6ekT/KdjBj2Gh+ozIFG6hGLBtUwVdHAW2opDySIEMXNCP1mTg
V4oVTLSUQHjbGGey5ap3XBVPJlA39zTrtEhLTUBc5xPsjTA3jzo9ScpGV/8utY7X
aCso+2kxksqwml4pCa6MtGPSBiI6Jq1zQxDc+KNL00gKi0P3LMQsKLEKxjMJNR6t
2kVOlTX8u7u7kigCYoUQCDcx8b369/EnfQnr8kNmMOFcp/DQQ+CVNUbb2R7IGXNR
dN0OGSh9z0HE3kncXtn1g+qTmeKiGWwEry0IyeAykl8OL5npdLLCzsgdQSpkBwBb
HzKL8DoqAm+pKjL/l8Q913NvJcXbxCaYD9T6fJ3D44CUwy3WqqIYkU3gYA2FTFwE
S9uyp1w39yH6b+LlUY+/PORT9akwPTBkerVB4hXkiXpW/U6tGsJ2fRn9x74Sj8Q8
yloeBvkT2wE21MPf+tCstoF12/5PpVJcTLtQsuV2OlHI+zMSBwkyrTe8yfGZgH91
eBJikrribPNdr4JhCyIOIldTOPjXO1TctrTvqOwvQwoUnyMA+/M7TCHzsU7aE36w
YEO+Lr22Si4SYpI9TlIg9VUeZazYlWpUKyFICMSHKRCQYfv3yzMLfaaYeYyYvgpY
jHy19+vyebcUPj2VmD7R+zEVVlRrfJtrCr+NhS1Ifp6H6+vWCnvbWMtCx1qMAjLy
6LAZdDdBIwedx1fi2iLxLPpBJka6SH8hgQl4XrJgbXZheUZlC/TJ0Vw8xFuJqmfS
wbM4aNFix+7FPhRNe3rpwxsO9mUPHO3Mhhh9pr0IZvODp/SZAtDbw6M+YPoBx8rf
UP9a8/ZdbGFudrtB6wS9btXgJ3t7erezoYz3im6dJBpdUyIkkTvDO49pRdULyfB6
SfTPbf4oCRa6pLfG2I4WV7NFcxFH2WveaD6wzhi92yMYF9FWc4MSM8sODBcMMzyt
bDipUIDHW4e06kUnR1jx97FU5qFbaXG6KMcHDWC3p/BFVPy3PSviAT+HIQ8v6eLC
gn9ApDn2kHqUkqHoiHr+nKN6SaahD9sD8hRS/uh03fLUwQHAQ6xeNae1fFHkgZm2
oQPnXuF9bU/esCiEy3mKFsyPgTkdGLzgc7eG56CaDStTq8WcSTQtAaSL4xPV6oNJ
rzBQJJ3dFFZ9rZIl9mYmVC8EaxcN3eS9gCiHJam7rGIf95Jc9p4Etd/BBrCx19MW
xQL/LONnM/wnHaDYOihqmjpgoqh7fa7JWuAC8pS0IAeDawQ7HvcI5MeoXmf2JQKW
/5iO36Dr3uCHfAtrubtL75W2rZiAOszOmFQDBMOiFNCWYs6vQyIlgploeXjyHOkU
98xUu6ubHzuJs+F0wZ4aNrDoNAAX+XfqPhWjJEQ/I9wYqNsg943LrYriGg/HDGGR
KG8CYqGRQbR1E3d+BFl6Jfj9duaDVOnYPTpDkLA+bxhnmYjsyZ8Dn4jCPw7qi0W7
pxUn89K2Wpj10do7PC5zapp7D4RD3Xl/sOExCs8OIY2UkE7EdXOqRpOmEgJ6J/8k
jR73lQF2s0wlh2XLr6ngL9P9nx0mufkV9LzJ8s5IHkjskbCIkM49+BO9L03I+Lfb
D4ILbUx4Ozu1jjg3hSas8aOvvy62DNCkoqI9hAD0SM1pqJbHReEwXfqedAZ8xuF9
lqr8GRQYIyMnU3/idEHdVntMx5ffzhxZVvE5y6uTv4Hb4Hgr+vGv/kFvVqGBrj3d
8tr+w5XvW/rDN09lu+0JkLm7/OaPKaINKru3OF9WFYe/+aBAWeGMjcXBXXghWJR1
hLOZqI84Dlfjy2txI50RvdpyWMtKJmWYSZu0K7oFcqlixwFWHiCxN3SmbN8vUQdc
37ZSbNv1AXRAb0rWdrgOBUgIInSvYORk3DzaRuKXnot9gDeNkQJlJQtgnPlC+Wyt
quqDPsppuhgPFMJoDIGedS0iS5jwCP+N6XTSLalD0Tl5dVoBMNZrkzaNjlW4XO14
pNxAy87JCPGQUSPdJS1tp/xhfgZ09Tt0auaZXUpZWCg9qI3wFbFDsvM8v7wYT8WN
Qs9/C0AHeo+ATIRVO4LZvrgLHnmMiriibem19G9t1xVPfKq+q39HV0r84h0BOZWZ
Yi5P1b/zPb2vvKdDHp3Qxjj7Z7EdvzaHP5Kl1EQYh78UTXuxEcBIHdKrPoXF948N
q2pQTSGw29b92rBiuUyt9a3cma8er1DS0bB5FPOo0imOhXcgNK3f2PK75F9ykOVH
uCNTY1Ex/UFlh03VMOFRzPmycApQ++F4IM6kwvSN3GdLQKkFGkGerhQEOwtmZW0b
83H+9f1M1zT0coZTr9nxrzdAkSdJCalk5dFv1WbKhImisI5L+J+ENOxkcCMII8th
CtWHeL2BeDdSUeh0P3I6NwCNhZUcdRxkLS0jn+cj2RrHa0sKyARyoH0q8UF7eAR9
erpeZA24QEhCRy9m5EWoQ1TItHzxYj5FT9X396AJlXeNyyoNNjrQcSdbxr9n2Qto
DfM3sP0x2CRtRJc+FkxAH8qrNRVbm0sbybsYaNH8S/wpH2V1dRlOUnL3d1PyYumX
xDti7nOAgY5PIxKeHvjN0tliItv8nCIfS0Rm9i8ZADYZd/UGie7jWd/5+7nImXOj
OoVYew/cIilavXeBzvydVSZGYnKnk/gY7SsZPdIWIVKADS7qxns+qCs9pjFyGLnO
x+Pe/9tEnzLMQXzRYlyDuvI0NY6B9Z2/73rtbMhZ5QA15OKswbBvHWcAMdMkrS+N
jhv5NBmL/PajCSx7U6DLqEn4wx8CyT81MGqLY7NYl6MsdqCVHn0PYrZ02lvuilYl
GJAK80FcIhav5BqCtzE05oxI8VOGVoENKZOtSiDiptuzHvfQFn5aFdIlou9IVlb7
k9TEq7FTVTYcxvP4Bf5chfoQTcTDWiUgb/OxVk1hyhYPWHJ4Z8R8KaHxoICTEWJq
4MtLnle+WwiJ1jHxX+RVBWWs0IYmw4UGypSP3XyMN/gMyZ2H+ZklAQD2Ya8djz22
tKOltE9yXVGLGA2j6Wl9ys40+3scYYQnoU5fqdvkIkOm+YvcAbjKwU+3buW2k1rV
IMiRKIvtjH6WPiwveSW08QrgN6hFEsLSCWcBYGerpL+AXNYtm7ONbNtutEodacjT
HlWO7d1MXAbc6nY6WoG/kI39pV/xujL9WnDbNivkyHI+bvqkwdmeEtX5MdbHbaUA
0lEqewPXN3FVRpFFmtEWgBE3wwZ5+Gg8BGruixEPUviZwuLAwTXPpMLrLVm8d1U4
ZSa8ltdHSQJdgUazWT/p50FXVngehyxIuTpEv+bqrba/m+r9MvdYHyLtry9L7tLP
IwRJooxHVptMuYG/Va24YJv/gnWZByt+TlMhzqeiNhNU5aMZtR+BZXVxmrneRFij
s+lEoGsKVs3j/W1nczrdWO9hYN60hwndEo0LCDcIH1MId8ivHKaTCO2IMq2tFa9r
aZe0RxT/efSscj8v/i5soZs8Jlp4zxBFO535IU77+XILaodbsj7zrjV8dUXsypTJ
jjfb7Nhw32FqfalylLeLMZUWDRvBh68DnJZxmODuxEHsro/Vi2SyU01lb+ZHGa31
4E+vO4gYZACWsdHZR1SSjDbdOCwkrLlJJWISB2Gt+pETSx8vHHR6luhxL7/64R6w
Z8yScbQDcPRviH2q60xXtEq13RxECgwUzwZNz18IF1tCGL8nfORZy7vSWvu5yLNQ
CVnzzaq55fATIzf4MSUE97ok5HQ/Nqe6EVWLK/aBwA2UN7fD5mxpd4o7RhWVY1aj
bxoInXe2ldI0CtqTRWn9OayQ3CHf+7x2vn0M4N6gA4HnIHGUEc7f8tpXZD2mMVYK
Pp+8Zo32ZoGDTmTT0kBpImxOvkQKU5Vxxy4PZHGO7ebfVy/BS4ZT+l2LfRCOeDrU
CPu70jFkH1Q1hjiQfyTQR/Vu8ETbeWk4zbgOr8VIAo+7gam3mTdi1nJSPIzv5YCW
GoZz8BI1NNSnR82n0FynYSoZY/g2YaxRSDViuJkpCwZKn+bVOTNVslL5RSxvYTNa
qLyiXzilSbpXV3d1sXlqTQCAVoxngSi2Ae41xtB4EtEU6ZT8plhFeAPUsHl5lRBC
H13+lfDrCUZXHSKJw98gkIAGRner9mo74jkLEIfAOGlQtB3h4ohvYTZWQ6UuvEKY
5JXMzECZoBU2BMZT24lK9wD0quEU+DlFRSeu0dfpMqOufNDPWYNDhkzaeWSzEZku
yn6G+HgWxq+1eWhhwm2Canhs78vxr0ILjvTp3uuZ827Xk/oGVo5res8aR8ZhXlRt
EFEN846HmyZ3rhRuTd9ogkkLSimDWcPFAaYbzXo9AIE0lRCVRw/pkPPW2XUDFPUO
+ZuMwqz97lXWE1OMl34xDL0C4mIG0hqJfQXfIzdKrZAxkEwMeF/D6PsCEJMixq4P
fAuEiZUEw8nq130BgyjBZ+Hu4Ha2kWU84sdZODbDp519uLdU8B9XNRrCcFkBy/q0
KYvTzjZa/RXGXKY5fW2VK0j0zRUUde4Rneri6oM1ee/QV/dNfONF0t9faOzMQ5QN
oA4/b1KVNTGym0oCBTB8csp+lOUMab5LuJjchDmGrB9kA6t1lD4zRMY0X1+U76Do
RRgJlclRaD/+bOyTZ4cEJRR1IhnF8dvY/XFSqBFFuehHs9S7fEuWsz7S044RrJX4
IPVCcmw89XrYQIIGK+8BdGftgVfJnxkZYyGAvvJPTdEKbTxiOmOxCjmpkyUQOKXN
3LPFRZt1n+bxpffL9R7PD6aFsh6+tlR5w6Eszfjs+TRuUvDA7KjrCZGzui55qSXG
vhspHGoqtFSddeV20t3Zf8kBkqU6ZXtsD+iWT7E9DUEP+gLDKtejqXBFQeH8iW9a
sfwQd6Hm75vTrDITOyGsos+7BRsPhT5t1DI8iuc37vk7aO5eEMZu2+7zGPLS71iw
Gpc1844FdYdvLgPtFh/714pB5gdDqaU/Pq9Zq36INrXq5JurU/b2AvdEJv2AVcDg
DrOF6LJEsgjAQpQZmb4ODsnan6P1DqN9PM+d0K7wVRdMkpijBTMu/zavXkR8/laM
TD8YkNz+uaV7WHRohbbVxa8muV0ZRo7YUpfG6FFOey8TboAj6/EnJiDIeDUx82VU
9cciOHBxVmFWqDMOeQIP2youACmZ7EDvH4ijF4ZHoF491DZzH6fx4PsppCPE0xbR
O7HAbcT3DXcEe9rZhro6r1gz6m9zZHDD31pxSoBuvF9P9fgMWtyKoFtIrNX1suZS
phuY03CWwLRvthdZzCqWf3eOlJ6BsV/vARzWF0D7KKwh5gd3OhVEQ3jpwSlYvjHd
dstQe8Ezd8EPIcNTwOpl7WZiCeFuXGlvy+w9xQksvLkMIc116rYaeDe/ObFIUBc3
nNWIGEa3JseN72JhWU2Cgf5DP5V95HEjyYyVB9nqWsxFS4pwthcHdc2SgU2K8DPs
QoA6xcuPMFZgaGP6iE4Ke7VVT6EyiukHquXVMsLOD+HVOPRaoiz8hz7wmuV2vOMW
W2TY9BgjpElBdAXcmBUoDr0Mn3AFxUkMq9cNOafMrPSQ9w+S3fe8k4xK/wodoq3a
3wlQcAafP2MgA2P6uxgMrhPIXcve+KzR+OgxLHT/fcVHjhd+TA6QuMF3E9oH2HiV
YaiBV3h/l10tjDu4z+DMaUb/LJ5TH6+6sJRerdcooOK7c+X4Zqi4D6oI5QVWyWDU
FkI2PJVbgp8tBR4aTKTrAuIM5yXcGUxZj2zWnpkgrbqn5sR4HIZcqOaCn20HPIXr
JuVjJlNuvqQ13mwnBbDGkEJVLRSGHQl3vKJi3xkQknG8AgAXLh5pjGMdoSg4KODE
tI4cQ431xTL2HyyOssERRzCvMB5hyzkMZJ+vKMhzh2cX/f8Fjhx2+VYk5KRnKeY1
245e75UmiL+CR1+Jq4ZSRTE5jaY1ukqSv19SP9GzbqBdC8vb9BPhCn11dofTZaxn
Q9/tz1xW3BiYP/W8Uf3Qr6Vfc3pMmu3KJ+8GuDIn9UDfU0Jrd9eml/xyh2AHgdeU
HgSTqOhk9MXqTotfA+B6aL0zd7UtldT/ezktzrQAbNDfABdxW5WPTKZjG2ELZx/h
LXXLiE0IqkP7Nf+gzqpgGcE1Y7Fp3FC2ViMIg1ttHHi/+v5BhWrcRnmE44VNHHsh
B/PGoznzNlvePodSHEZ/6shZRk5OdVsdHUN7NA2h8CKNL0VQbE3z1AcFLq+jRa7d
PR6EGhfqH/g+FyRr0DfsV3c7pT/gTWSmDZ3gmhGDhiKy8QuF1q9Gw2ZAqgjQ2X/6
0Ddh+98XgZmu8hLhrnftXbW/2VL7ZrgT/5Q6aDxCRfufDDuDoy+cJZ0cgBL9WtP5
q+XzrUVPxOB+ztAN1hKf1ggCCAlq2hm87IGAiJ1XsTCZsLZTbGPmiTIIzHF8fC7W
8C6NMdxoi4+zmhpVQ85+XePcLmdf5PCmWwkjWuGiear7jf9fPznURdFq5BsVjJKT
vlcRs+EfCBcuwVK6xf9vsr/16la3mru+/CSkiUhWj/SiZKoDN61xclIu+/WbdKkk
dy0sRi45FsDdHun/M5LJ65C+NDozGfqo8JIccWOnsBVr00il6VLBFxq2e0jCygPf
jkMCP8A/RZRViD8ZFqprCDi+eneN81yRBrbK5PmQouMvmeb5F42UYvd5HcoXZU2z
+mQNhbgdu7a95bT2/xTimzVx0Lr5CPuTIcF+rNxMAUd0KEC94xbJXVYgwgbxZurw
xurzeQy8IMLp9Xqbd9EMrn+cYtBY0qM0V98jZ1wo067WBsfQafmSRpN99EfzfFb6
72oeiJd74+R46+imOFl4Qb/xi6VYpGjmMqHZAwxXULOVNEsOuzqpo8qW+ZDT2Tp/
q6EB2hRx7nzpzLBdYsJ8CMEqwWfLBRyy3fvXSVQvw2ZI2spBbr6jJ10fiFN0QQMH
JI5NDGdC2O5UMXZLVUSKsuyTdTnCNt5o5xd7uuOpMqrXqP3ns4HHzDpg56fSyoTB
+yNRk6NVjo/o00WMGXi7aLYKdp/OWBJ7bNT3+36ITMmhwkhEi4bKrZPnJndp7eE0
y8GSkVvBGfwJp4eVdrGMW4OkjmFjn7SsfPgAAavHK90uVx7oq6Wk03+AobD8Lbiu
fYi0Pn7034b7i7OtWtm8N/c/C7OkGW6lMt+LDGVxjpXCAxRpT/JoIP4uFoDubeBb
ZbLyZRcfYHqt4k2HHNoB9ZCg6xcb3WPkHvWm5rOHrKo9Ia4hBJgHwU47oSH96V6h
Y1oaNWGUX5e7P6+drHqNvok0s1T8Y6vK4PFVticD7hRMiCpo/y7m7esJTppkaNqF
fa1LAaTkhymD/bEB8o8QpjTrA/gNhf9bMG/gYR5d9Y9RRqGyPeqYcEShqmVDypcG
sXGCcb6mztAQbDTFGx7WwISuusKq5lzewezrZJDNW9ThrHfXlOxJV8NGkMr2YUCZ
BMVscUiFg5D4rUYzcIHMkRbS+estjiPYSnjETo2ny6dir2vsCxcn3Gts/eGU7/HT
+FAlIcyjVS8/jRMi7n/p9kAn4I1+1HoB3x7MhBfmsGQczOfTGU1uo1rO/vyMQnEA
8quG65M44WijGDmJMVrcCZH4/XXa6B9Uic9SZmjwMGQCdmq+ZpK7cUZP3HMIdRP3
DwsRIJU4f2IsFyzbGbBq/6klqvdZ1tzn/J8k7KEWgWPr6tIefg7nMS3vzS7gQb6l
kMQsLTke5WilrBzMm7HB2HmPzWVmakpVfzIUlp45l43hcXQZ/OM+YRvoE0CLjwFV
HZ5v+OCwdhqb/QRinycmt0iKfuQ3O1Q2MH0dL0FiUV/WNLoO6qd61N5gq7Gg1ZaZ
x5gAbClCIyaZMnEh2sIGQocSnNwdy2s7SQNXn/zG47mR/DFb1LnIeg19K6M5pMc2
wVb8UytAjIx4qs2GlhCMmz5UIR/FS0mC2pOMK3SE+J7AImOs1LA9IwJbuZ4iXfdZ
HYs7y/vG+ubZsgxW81uVW/6mqYlV9BhPh0uDZ7C0o7seYP6tHmG5igK5K1f0ph56
SvDK+ckDZqCMoAwneTrziF57SwN881N2Usbj+UZPXCV9iu958DQ3invsXob6M9Nd
s2eukGfyqjIyx5AHbUiPvBjrfxoLVLDpErQOAlqaIbSInJftrT2dC9YccLlKMUhx
PQ+gt5YbkTKtG1rBi7xGBN8GzDVXU05ZnOPCNcMu5rnqvtWxc8wkiFTT9JyMREnv
t8JkEVruxbDYWSNvZEZdC30EwR1nwHJqX2jLMRg4HAqKUnMaw4VaQKZFRJn26Nf/
1bjABc6Wq6gc6tTiClDJ1X40IaGqH67WY/ya/1sCwc/wBCdFKwQtsi24AsxvaUNY
obcNLM7d/Wfo/bttsOrdxqXMa1u1LkCM7tWB/rbzVMohUmcdHBzWJYOIIQSHaLfx
VXIYograkAwG0QDEjyH5ZJk5JrxnZ6itfggChcJnTPxHLBjXoEbS8MGOWMCZGq3p
Rc5/KsfIw2HPnY3SsROQkk+EuIC4v+MIr+us+NpjgYd3CGSAZfT9dT6SGFni9MFp
TTSb1JXZN71LRU44uv/6O3KcxEapY/442Hvh5/5gXn/qbOAByZ0FUwT2OEctHDrA
3OSC4g21kZhJiL1M3vwwtQxmaRnxnWwk/YfpipG/oB9ky5EC6UCrFUTHoiJ1O+Ih
Kk64ebAoPI+NDj2Slc2Mh+BAmShOroN6OFzTnkK2hjSJk0R6OqDtxZ9mc0TykQG1
30TRgDELiH1czKc+uFVeNzJ6+cXYwg3O14PPbySt2ut+uNB42HmqXYA7RtAj0xoX
/5yUeJ/SikmTYpB5GkQhmIPK5dVwEZAa8+UGysrVW8UuIYZuHr7DrQxz4Gd10v2h
6YGoIatSkOWLXxGfzT8nwNTo01KtIKt7XLrq4Ya2Uj9Sgwv7zV8Qcfbxd/d775hJ
OkHhbrJ/WnctUVrjP8jTeQ5qfrarM2LC6+ft+uGgVEd3RId5B9KWj//7Go9+9mcp
5fTd9bNToP2SCNUuDvZeOga6jkeJddbAZSA2pSzYN6Yj3lDLdScVYpfXvhhV/ad+
HNThBYAXEtYF8Z5tKRZEozcmjCMT9svjrcTUke4WSJMdQN0leCABQI2YZZJsYIgA
oSxPJBokdXkVurzymWrOtUImZPHouF8Up/dq6WsXBApYqUbnQY5cKgydaDfqt8ti
7VFKIyOoSrT8glp2f/NhJG0buC4qZITrcBtoRwhABuL67rcbtRM8EsX7jBV9akKI
fyxB74Gdpjg3bdBtM5K530ZvI6P0fRVvIhj6ai1nD7HNyBvaMzaGzyRP6//tN3aI
rTLXb2YnT9xvtGe+1ztoc0aOqb8Rd8KiwvoguVSBECguSX5JxFQYxN7TUVYiVIUU
YpZjXKNBEa9p03dRNfp7Rms+c997uevn+Tn2bM8/wAYUXZcBqJPZRS3lXcXZPb5n
WpNMbrKdK3xl5ur9WChuHwgJhWOtDffXiovtDV9SH3g5F4mvxnYzxEFs6k8Gc/yD
zgXF0r0ZiU4xiNYkKEguiFA9pMp23w0ABvak4dJarFnE6VMSKu6F2Q8bPNfVSXAZ
fFTL1oUZpsc1H959PLEwuDprv8lyeCAFaYMRaUaHZzTGFxXjhbsItE5PpEVpgAGL
V212GtzOXDzw6+o/o3Yaw6yuybDIvOmvjHUIfiSCGc6IQACGUMngCTK5e7DN0woP
V88RCeNwUDThHWLYLiwVKfTZRu4P9UFpHiAuniG5t6mzi3kXSfXHTB7piIzP6mlv
bwOFJzeVzpmhwyBRT5GZIPwiSoqifoN12SiXk0/sBEAqsTZMYIBSaXvKJ5G7Wpvb
HriKcfCEELUiQA1SENWUd/YukBUE5dqxgbepGptwcDEqfme4YaboJ8yiR+0kCK3g
mKFYzasVHsufFbdQMoJCxE+ksQVsBM0DE7H16SDD3JeVc2K9qvl9PB1A0udc0u/R
lxXuzFKkZ3eRlGzcVrym4guLPUd5GXjFPnyx7UR9WejvpLeL/41bblpXQyOqMNjt
5L4gfaHM5mpEK/JZmVGEJbRM3bp888n9V8DugKAA8K9Su9NYx0/Hxg/1kNlYK+Qi
+q2Yj+BSqbx8zNqXYezTL7uSFow+0VSYpMMopMKklN1LcBQ8rdpj2ouQeZFTx2Os
gmypnfXFYAI5HTNmVCkXbEYPpSrosRhpFdq0/25dOSGQr7QFHSsz9gv20jmufE3t
CGWkuypq5qEp1xOC618AH05UoYR09yHugQIF++WGm1gxtnyF/1DcUnlpYvkcACFn
UBItwf1M8ffEi8bHsPr337EzOZuwtaJrydLsgSL5DH84Qcc0ZAmWJ5v/Nqe5uXS7
056IVyVFibHbec5gPYbhT+fnLE86KeCOyyZnS+rox7ut0pNCAXltGyNaLRQa2jym
Ezz8YWmIvZyWvIjbFrFZZVLUlKZ1RohRw/cVPbRvpTo4cft7a5VapTi+y5U+vAZ1
vEM00IxhoJxXCvI/jykipanl2kJuax8LF0xwtjUv4bA3tlYp+3Bz2DOkpYH4/zk+
kMhKpmbfbip/2UMj7oRBmKQOUUrMDbpcIjBrCTbZvW0keDJtw5GZ3GMO/bnVLH8G
QGMGq5hUhmJmi+VEm2YuCXUBMuguF9d9/izzGox7hoRWZjbccaP0s62b2inWe/KG
GK5yVkzRUkIfTxTcSW3X2Scb/f9LM9cYI88vwJujU6IpUiCgatH79suP3ApuRw7p
OCfgNuuZq5XDC9uTbnPH9cbLxbXKd0H1Q7tc9DrR0hwrhJWtw2z86bt+fsGgwrur
PMzlZlYv5O++4HCBUDeQvrvx8xhyY3sFjnu4PalxZ4yu088J2BuzSdhfSp3qjRT6
oJ1NTXGIntImsqOJ9Z7ylsW/Zr/b4hLLgMog5VxP7SI+ImYQU1OyDDsHWTmtr7EY
Jk25i1CM7fLtu4SCz7VpCP5gXFedLmfIBu24SRacGT1x9qfz81Xb3jBGNdXPAPhg
56PVmRRxWEA21ffalVe2bAqTO9vCLV8wshT8CtZvQZfMQi1a6sRlfk9HIpeDqUBE
c7DjrUOzDzQN07HbSJ3beoyavpPyS10AsDjASuiB9kcmq6hEWlD91U94ba0sDuOt
UghHNSZpWxA5ebQ2AlLO4IkZLUFFTVC04WEPwLuUsihE3Pvs6PwNiX91gedajcP/
MaRpooPpSt/yb/9dbAM9LKPUSloyhdPNoqR52VSqff1IULzwjVZ5beoRaDnPl8g4
qhN4MxCAYOwlJffn6t2YX2O4hlL5CmgHRqDs7yDV67sFFNfwYdy7ZFMXPwPSG4Lc
R4pSZBuNWTjxDhkHjO0qWPnQnD2hmPSUvWzQ3aKFAEMZFnjrwBAxPCqM74aWofWX
LG9r9Ml8yUnk6z6hohHQa2rggzYCmQcS6zOMo17q9UshBnZvG0ITSlGq6cZNf5vd
LmVZEiepcufkPTfZ/7XxYASy1/B7+phe9STmLSAIprcXP/YUsv5Sbn6XnSyEWJal
b2xsUX+pOMXNlxl7Gcvu8CWtCDJ4PaEh0FKZfi25ODx345BfTFoBlpleTCuf5t9M
H9Bo6EQsucInL4OwC/FgYK3VTEF9nHFFxyr87WlyhZJ1+HpFXvnDqV41/IAp7e5x
h2vr53DQ0QnmY18p5wdAcX7OY8QFGNXHWpqr3eTJF/LS2WRzsB+fsmvJSi8g3dw4
HOTP1tZj/Ol5W4Nu/v+b6MDpmVwEE1ymAPawWdNbXDOYaFy/jiIHkEp3Dr6YlSNB
SPCjcoZ37NN1Sj/Yua4aooj090MaqyXGgWbWbtNB7BioGBn9btDaeNsCRdT75WK9
SFw5bVIduAuRwDvX5siNiporKNLTIIwcb9J//bmH/sPxvPMcYnKc3hmvcwwPgIWo
QXJ5j3pwqnnnNmSptUkJo2VdZpKVKdVYwABWgqgHVs/FHzMXssNsqPYVQ7apSs2r
pV52PtB4PfZeY3ifx1+3F8Aq0dGb7KFkrCeOiOUGUS+B+Zt3qwiaRwZSTEkrPAHQ
bFkcKxkesztUQDvVkHRmM6irIiAe99FawulOlrAxtz7IMQ6Fe/uEtbuUQwG8kZWJ
6lSTswuc9gL6rA15OAh6whC4jNPRLkKg/VuHm18iWeyu5frGBS4hY+eEzYakBD0O
Lu1Hm/ocWufm68GGJVFZJGhcy8kWd0VZj9a6W3lkTW3h/++9VWIrrIZKgLX5m1Lp
acZ+yLbnEawI6Cb+tx7B4UX824Py3TyQVPm0nxtrD6d6UoZQ6Djqg4nsU5YqtZeq
HEuhmy1vFAx5RjBDDQaa8Jymp0kRsZ2+orVnLZ71K4WBGuDhJty3ZH6PIsl7nVw1
FPoC2dBYZHlE3CKgMWBmVv7IyJEDp6ZgF4tP3keUcHUBr14965yL8yKizo7N/T27
zAKnLOSCXWH3trNg++SR27y4ryJbfA7cv7yicyS8RXctU3nK/4Zv6xvGGxlVVpuf
+nQg+9e6GrwKyBVoz2fiEVCkqac6qYhgoYv5cg9DHvXnw8/rvnCJBqf3OIx8BFJe
3D/jhJk9jeKa4I+IrLo507NKZHvVFx8WwyUEvmA898/UxgYn4wgENO4iOl5AMqIr
SNr0d66che5JqzqPeADfT3O9i9yrrmmF16NWGM2wHLUaK5WnmpaNOjD4+Z0ZEtxl
rglUErzYCdV3AR6lcp7xfMSL5t4OYiXoa9B5s++mcjpYn/0l3EIjEO/IOmYwLOfy
EKArkh+gAekbUEungq26aSgm197jvBJKkU84WzLl9BvrVRdq0hSyjzbvmfJDgEYI
Epg2XUKYairZP7zQfaSUy5D07Jb0Hsy00H52wfhxONckB2qgfFTG1loznF3R/D4O
utaIc61X0ZKnA+jZXh/6HQHE26d3/OBYASjpyDLL8Fa2vq7LEEiqkPyovK6WOsuA
45kQGsoJR6/b8I6adKvWo3KFgiFPfe31ppz19aikyINNet9iPJctk64p254lnut9
vX35pxkFHrV0ymroDh5lARX5Tw9FC/tQj36++2f2bkMSC8SUApePLATD0RCtzDQ6
m6ueLhOXvbYIHp/GFLOMbygPw4ekt1Qg7/tLnXqArHmgMFS+gOxxdeBOrFlTsUTm
bvV5rhGT/0HqNe0zx84s4X13P70BLONzH6RtGjxLyCq6UXwiPUR8mtFgZ7V66c/w
HJtmhtWQd/RSBHTsQHdTXvZbSdJMoQSb+eSXGUx3SJTD+/fdoNPcd1Q9tPSibkvs
Cy2eeOdKNuCYDOQ/XWPhg8eDQVHQEhnVN4bmCDGLAfdRx4Mp3OY4HziFnazX5K0F
5JFnzCavtx1FW/xHhlaaYVClu22iHGKKXesSLEYKMEHPgS8CfFSU81bjO9dMnJcK
+lInthjUWMwipXNQhVDqRT1eg5S/0fzrnPD7HYHPZkVS7CGdowoUsUbXMvRz/m5i
DaPaACYTi6C8xiZg+Y1HfVEwcrrxRHxx6Qoz4YqK/FIjZgt8lbDVudxs1l4G078I
/6lrXJ1E8RQfVgENMYMc5344jAgFmhSfLnu0uVFlot4Vbq2zJ6X/SF/ss4pDtrWn
Js1etVj1i5h49fSDeO9ZfW5qtwdh7sDpsBhGsIbO/Wo=
`protect END_PROTECTED
