`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mUqbD9xGj64KSl6B5bgpzVYQIEoEJD19kdVm7uL4cKQWRg1T5We3KEJImP8B7+LM
xgq3iSxFyiFAYElMxLeP1G+kfWfORxF+9SyP0mhn+L+vx8qv7BYwqktsACbG1l3N
KyXN/lcv3pmbBDRTZsv7joPSFkArO9neLJPEWAiArk2aKyztGOplqvE3W95VYaup
msS/LV2pPCuM8B549i/vVCgyHjW7K8WrdxvXgPY09TciaULCgf0gAGJd1d5nxo+6
/2bpAwVuKKuWOpDfC8feb4GOeK7z4bxo4RJZ2qsYO425OdZYZk4QkL6oRXLFjkM0
GMsnPQGGcqJdGfhtJ13NZPopaf/5T6WOhmBuq1G1bMWSQ5B03LYkQ9QA67T83rja
0EOeuvt114AV82Mf13/COHYnKHSE6VbHjMWZ6uaRhFo=
`protect END_PROTECTED
