`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQmcJoxptr77vDxrPm5oxj5ptCrM9RFvfbZ6VEtVF1TFlNXFv6YpzDDn+/vxOrRq
fH8wTuFQ1tW+tecym+fpTUPrxopLgCzmSEozMk2668B0Bt+3Pwzr94bn9oSJzlgE
Q1UmB0ZNwWCKIW4WdMovV0B10ZWFWwSeUoZRkYunstpi/UL7C6dxoOz8HfTPV0uJ
cy3hoBzOhP4WSKK0C0e/6fGejhVsUy/RedoPnf1OGsD9xVbQO1bmuW1C9Hf60QYy
D0Sl+RuEfOO3rGbDFYyRvMHPF4h+0AH/tPc9U20fJCvVdW4eUFJCDeJ1qANbW94r
Sl6PkdhMYtI7B8AS/ncteNPPFnU16mQGTe0WlRNIJr2zLFQAYTycupTVYH0+GoJJ
ZCGDknU0dCUpJWq0AQ25ZQudA9jp4tnJxS0SD0SuSzRVHnnjueMQAgDhtqDcZH/H
GGO++DSQTN3zF3xHvFasyJFlyRmsFemAHlMdeNRG0UAbiWsakueX+qq5+iqfYfrz
wVzKPMSahL5v/TjzzyInSmbapF3JlgNRn4TgGdbCjY7WZsRhGjv4sgKfi3i7zKvs
c1TcT/Wa9Vt3h5IhE0PYwQclM6+FRKGSZS0n1js8XtyR32I8ElAqtpr7GHf6+k34
pXK3C33CbKZImxgo2aubvyYawq9kI2MHG60xtc24X7s=
`protect END_PROTECTED
