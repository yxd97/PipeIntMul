`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTt1PTRISWL+A5lo9bIlWGAvW7RNZm4FkFcgh3khBVeSYl4u2naW0bqZzcReJdfe
gpdCzCj5Kj/j3VGZd+7EaihEApR/orvXlOb084ak1vbuX9loACWA66ySwYMVU6ae
rspvXRkshNe7t5a8+sEGIvwWrFW3GGkjkD4nHK5+dwKsy+Fr8wzQbt1XYb6AmEBD
nfZkBoEQij9Boy91/vP/NaFa6acdAhwdbeZIygFtwPzghfiVSlNA7r2EwfokmcV8
iVm7M9W5bvhfrYeFp/sdiqjEaOLftCoSeAq11vgIJ3JNmbpl5Ifnv9kF4wJq+5pO
5kx5JG7MC45ZOCgmeIJdacyWDFbLCd2sPLpiMeWczEzBtVrLMN0U4KMjKwT5O+Yi
`protect END_PROTECTED
