`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n8qkBkH+TmYJmnhiUDoC9inOY+fZRzmwb9nWsE8ajNyLFFQJfUtlydM6o6sWhxzg
VX6yv+cVY4zQCKSGgzWgiIGL0NPJc7lGciVKhVK3EqSBawXxntq/az9BLJDR3V4Y
zVWqZ/h7pDSHcqtlh4LssXqFxLim43buWlXEOsyk1ElQks1IWrppPnUno7zrjDU1
OoY202FCvQVQfwGLgG96lHOKx9Zmb7ijRUnnONSjF59uZJKvfdGNRBw7pcP42/7g
yTcRo8DXj3AJasTtimLSJOAS+J0ck+5xUsgQ+UFeZkoFdUFTzMHQL9VRH9u+myuj
zNVO1TnbGLxLvxMmukRyi/aWnpeCDlJD80Jwy0GFUzfhSWY47oytL/xe0Pz6pa+u
14VpVVkbMQkBAYJncL7ZEuNaYK9WMcHZ5+Hej/nq7/ybY7WrpLuujBTClfpONYGJ
clncH3okErp16cGsL1QpuqdmEhMJMfKqod8vuPYB76OE/IfCTIF125vXnn5xrxWI
1AuatXmxUqFlXjKF+8L8Mke702GJxdzwXOueFR+0UIkXly7Amkb4zzROpXZSUAO6
qwqN/+cInSe8Po4iiqMTkVFMztz92Upe2JRsNIic32qs+OwOy8OrtN279sjnfEJG
a7fBTyeXNsZvbOwuNmbRA3KBH2/yBAd2EC/xC7xNHPwoIUVjT3Au5TDG7V05TfaP
`protect END_PROTECTED
