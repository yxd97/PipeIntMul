`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hlHZ/0dipseYFTAnsTVjt8CQ9nVcWK4VSpKioZwoUYqvqUDXl7jbBZGalDoEQQi
xRBcfLxJYXBUcK1SE59Prgy4zW+5gi6NVam1areYqR83UCMXotEy+W5P2ZgVGQm1
Hip5Hz7iawiR/KIOMrD2R49f2xHA548wqbAuKzOzW5Paxjzvhd+J1xZK4XgGA4PR
WxlWsSChK+8WuYahzqG4Lw5Kit5VxbK3ZqG5uS1Yz6SEmKbYBTS7GXUhGSkzI4Vj
fls5U4rTUQ1obBH5zqfcjg==
`protect END_PROTECTED
