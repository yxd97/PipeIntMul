`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6NMQVcZfzcX9k3Yo1AnRhKKqR1jXjhmYrZycfZGSjso2jQ+wxjE47GQgyJS7DIox
eQQ0wAB4sPjT2HykbJhmNjflu03nPLDkS6F40tg4gybOuobfaPDBw8Amd287qwg7
+OvMeXknoTMRCucPAioF2GJMVyhDxWroGWxmYG3bxuTEXBpVxIxJiUcY+olz8mbD
aweNk1uT1AEsrN5lwJz1QquGt5Ikj9sBwbxk29x3xYyZ8bhJiMBDrQRlKUwig+aN
p1J8gTD4rsdK5NnRbmlEZYCg7r2XZcm3Tp+MMLVn6DA=
`protect END_PROTECTED
