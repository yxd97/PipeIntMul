`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LQQwt78u7Yp/T2vsSsDqKDWh9hOXCrNyPmZkfothFrJ04xwjwoK6CLo8bkYE8xJe
40e9hoFmaCxMwJjKsSZCsu2GOquk1caaiAwCZEMRvrL8/B9j1WyqSh6xdbZ8Okx9
QOdvpES7tBM/TDxU7R3Yj5o8JI+RW2UhIeT3/ekVPvqIaHyo8a4cWKokwX8NrHIt
uNTDrF5+vK2PgEI3m+tUYbhRezrRNJm7kw6Ql+NWhPhlSN9pWvbPifSYZNnNdCtp
IXoORDlSgbqepaZTmwFAWQ==
`protect END_PROTECTED
