`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fzJK9oTThaqrWuTcCNqpajsi44pKhWy41UtcQFUjAB3fl6MN47Lh2JJnQ2n4HnBR
BsScxKp+5M6AQb+BwjCq9hVu0TA4d0I1MWauPaFepEPO/uzr6Ym74Rtw5RhiDD0P
WvwknPw7cVk+iMl3yGuib2bpyfpxK+uh9dIz9P17nHI8IffapFALWvYYMTlQvtaz
6WvS81krMYEKi/3kLsAlnor1M2bw7DN9RhvahyEuVhcBsb2WhZ1u0waY+ZLrVMpf
USTyc2kvISHuHRwefXf/+vVGftxQhzmn3zJXVKqJOxgqpNx3rQzRrxiM6Q8CPn0P
k9Q7WmYorHrtNnfpZvnjxwTReKDnel/NiBbheNiGLafv8yWMBjtqZsofEeGUb3RP
Yiw759OOhoO12/K1WT9bNyuZ4ywwI2cwDUfZTGa/45XktFSC3e8XNLCDtf7G3qFz
a3vt5/qdjwwOj+kLHIgFwfXXG36wbxzIzFlunPJC8KeygL8IIkn3ljDY2qXi8nkO
n+CeK72Cavo9F9XiL+l+7A==
`protect END_PROTECTED
