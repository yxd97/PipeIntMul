`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
274w7ya1wuMI7cbXEdxg1obsWdJw5RWFUUc6061I6cNQC0fnK1nFUkvYdaabgOqd
vorhT650GhWjye0iZ2x/LnuVy2gETOILZ6VhIkdzsdOWyBEX/usKH9oQYpwWZNTm
0SMm8Ur7eEFsnw+UdD8nMRBgz9VZVDaTlJHoD901YZP2H2U3oL1Kcpj6KVAnw3Og
cmzQadl/LHVbce5o8Dx6gPOiBkqBXvcA/FU5RlvEI8JEws2CZuQ/MDl3x19YkQT4
A4Ep+Kw0q6JFgnEUwAtGz6N/9p0HZLS5FaiDjoI3CnN19I5UOSOhHtBWB7NP6IDU
3H3edTrsOxipOmsS2Z56xZDAF0zB+WCdl9Hyyo7GUoO4ERfQpH4Et9cT+XM95lHR
CP4n1wD3GDIpGo/DQkOc0ZRNSyXFE1DkUh0UGCBNTsbjf5eoBaEfWdg4+Jq/wKUp
ai1nDJGtRHUfOoVVLswhIMWisSO58cEpkBypjLX/vTQokxQdhdelKAIhUArWGU66
r18bohDLnJ4T7+1QENsXinedoVfR74MmfeIU5om/Ec5MmWGjpIgUu4Nw/MRtI38s
KzsNKMkJfprGSbEahLkLqPbvlYcWqQhZ5x1auVNICqM=
`protect END_PROTECTED
