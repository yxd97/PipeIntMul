`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yds+rMpve/WJYTcWAMdp82Gvn2XH4CtvXFDNSbVn+pry2Yf09UxqAb12ttDZ1/wP
clVEzWJDkKO/OyNz74ydEoQIN4t/BuzddoNXPE1pilK3dF5r5o4ajXTlJu/JUXQL
mFVMEJ+BM/0ydujtNF/7QBju7MsZCj/mmzE+kXJUs0CbyJxkavTGwRvG6rDuBFj4
EL+YkAi5ond+iR/K9mHC9ArLBAAazwoJV0Gj0dGWRfT5RGLLlzA+ZRtjfGGE12xq
fB01CPBbuYHHZ1gqhxrBnMRcnKjiWmO3beQyg2LCzgB/zovrrDhpBYUFx0uJIgvm
1XkZxOHDRko+FxUL39b4eQbvUBs5a9VB/RQNTCQyy10+LCm4uHK4D1GhyBsrZJBu
+aPsNvgQUYA/aQLyinRObA==
`protect END_PROTECTED
