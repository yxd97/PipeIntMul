`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spSzz3yVU2JV9owVSpchOoC8XKkG7yaALDt7p2RuenEVqfIEjjeuCOK8CtOsQ/Nf
gwcfLsv6l3kWz75rDHtaiDqbwNTQx3a42nrpyffUE1UqvFLP8NH4Lx/VjGqaDjME
qzes8X0n6o1GayBsKLmoYzlnaBQV888ceXkrCyli0/ra/kvSXWVzOHuIs9daFxCv
xSX93jbZGFs61TMHgVjgThBVu1rBeOJBpjz6KuEMrgQqSXHlP9lC9ltI6VzHiOjN
1pEOQrtRAb0i2bV6Of+lvQ/pLYfWFBFDVaXJtUaeumem1y4IMp78jT/uyYUcNXXA
jj6Rj+uKVVxyLudGHvCoZ6CNAlD/cmQOK/xn/fjl3HWLEBaQNVthg6uPDq1Szjj6
IEqjEohtarDE16areQutScdaL4eQR+sLFjirBEuzSdvLIdaPK376SEPZEumD+xBp
vvuLYnYTTV0d5MX5TEDnQxQ/UhkdX/FCupCDM5yZ2P63jhgqMV5LyIaW3gUMThKt
8hdplB+0F5IfSkt59fHxUeiV3m7wvMegLAoyMIMx3KPYeSLgG9YpW2kZl5d/goGn
mXpRLXTuU/09Ru+EVivwLHUtsyRLq/KLIghIBThIUHXtTY6sbcfMovfTKqd2DnJ5
RL9bK/rXIa0BKbWsgLCOCWSVoTi5s93swRmmIJ8jCMi52C8mrxMp/3JBD2FT8zKq
/29PY/pBus2jKVJAlqwd7Q==
`protect END_PROTECTED
