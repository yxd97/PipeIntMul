`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWIMQbQOx0QEcG5yY3oIm+kaYKlswTUoZlbYRo8OWODjkCZTPFEoleJMPvK80h5D
HBx2eE56V+JCACuIYaCZQfRMQ4hzAMqYc+4lpWhzD6NztK3wAB+FNlEaZz3c0emU
VXv2Pcfp9ZMYuRpkKMeyMQfYM5n6IaByO0O5QTMqxBBNV7An7xhJcEiren0EzzZ4
b7TFbc6aK8Vuvr7BkjElfbb2rpe+J4FNvjfa+vOZ7jiS7G+6ehuZBRzWQwTaUOhS
R64XC+IOElh4HEP8I8Hyau+dyaEbsC200dxNWZNQaIpocHaNHulvNGbvTObBIB53
a7SNXuDhKxe88yYgd8Q5IB29VysJ6v9vXRMyrFh/lQ3Rv/4ERtynNC/MgqNONFUf
KxFKQGvrQyXy6k9Slg8t1a99Yl1wHJ2Tw6PkE2JAdtXfcpd7pQw3c7Zahxd4VnYv
VOBQVNk09zoW0OVCJmaJzFRiz3vrD5tmDtIAyJY911+CgbW4TBJKgzoAI6AVgsDL
EAk/WtxWDkKVudIP13fz8K7hyvIqmd2h2T6Ntp3gMZecWpaJ6ZmTgw8ULnEbMid6
ltc5R9CqxMHWBE0s6ShVbAvO2F7qYclyOC/gvIQYn0Tftrt3oJ/Y0H1YpAyIKCmu
Jpts6XxhAdsE+2evqHh2U18v0qBviQFNUvjENeSSX0zhaze9fnGxJJOFgbxfx+U9
C7Jr1PJAu80MmOW9AN+wyH4zvbOdsXIWLWQO1BMnCM6ayAWZTZEbSRmgTcV75G2L
rP7ESAHosYMRFYWRPu83QIfNWmuNbiGjvqcACC/OHBOmutA7xW8oV2RzDEVgaFWU
AP6YY5YQkailTP9CNUCYLumTLPYr6x7pkfXfNAKAAZ3M55fSf3kc9Rob+1G15epJ
cobFhNuauosreW9sTKeNjS0iPz9G8nuQZugIzQ9oYILF6GuO/KNsZX4cIhGA2Mac
gJX29HophOCsEkznqoR6wTKSWajZMhyryBS5SBFWmr8/KvZQjQ/rPQM+owVvC7gJ
qNuDb/Xw3ufI5nr/IsJk00G6vNgvMvIcgDYQJ7jXeuk=
`protect END_PROTECTED
