`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y7zvw4A+QWGQoPTzTW/oiUrcUswqNlQfKmAGgn3ZRbIi5qRUyG7AnvJigt8KbOPH
YfplMcpWvHcRRCAT3qJD8U9f6QsW2gUoysQvLd20mRoXBpHBn61swwiqGDkCevBx
oSBchMU8vz5hxE4N3H9t6Wn2lLezckYYL3H3Gx+FW6BlttGcs/t/dam30njcp7Jf
p1TlN/GqrPSpz/FninTJmDWyfe1Ini+oJdXQRRsW44aLab4p3bFUmYF7tPIhMJxj
poZNQWsWz3Lbo9ekZX/NFszj5KRKRS5XSwNkc/H3oOS+psiD58h6o1MlODkx/soI
LXp2v8YhYdJ0P48VUncCeeAHiO/x2OZZyONVGTGJ+J6KENNLA9WApD29mGIHkxOD
KUeTXJ10qe5RTWYqMTQ4FgurpD0hYJtVuDw3cnG2r3A=
`protect END_PROTECTED
