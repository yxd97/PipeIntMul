`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lglb+1BunJHMisxq/yTABz1dMiiljYhGg/j/zOsBCXy34fvxwpS1sDW2oO/2u3D9
TlOAY2m/KfhHXr8t8ntF5g9IRyvvjs9tyUYF9ir0UG2bKH1qTs8Tk/pf9YVHehig
wu8eEZ34S7ygmQ0wpepMC0SuYaVYY86+DjVDaVGYwGZQ/ILL/0HL3EEKZUx5cvgR
9IW3CoxBGWWsLowvU5HkN1m7T0gAx7WPkUy6D3L/Ub6PfJiFrEQsqMGW1aM/CUHt
2ffAwszrAWUEf9ScjefOT4i0XSoPbB2miTC9Vmn3s8wRZQOJgIerZXtqTTA9yuMn
AxW4+B4XhghB/EiFX3oU4aGNn+LydyBLe+giyrfK9fW/Thm8xeFIN3ZRWYe3I+4U
lOuIWnOTZJbXaT49Qsu0OdloNd5UHNia6IaWkOxLnKCoheKmME2icPGiO9hHTHhV
gLKFJsCQjH5tdtvr4d9QYOjmWWmEEvoHj2i7ZV//qH/kbkWIhl2X2txKXmNzZBBS
`protect END_PROTECTED
