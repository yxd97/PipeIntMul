`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aax8sg5ANCI0dE9xXab3nbnombRVofj2WC78RQrX+JUhZM0c4Z89oDa9n8bU5ZkQ
oD+2d5uMHcohgxFYOOuDts6QE2GSxTGAttewcw3NUEto/jny3JH9GvRo1uuTeJBR
FhL8L2yNMXNF1qY4VuLWEAVN4naoBImysM9yGe9EJpE+RJIyHDQv4qzgVrVkMq3+
U4uejGW5Rd0EEmHmCcdwKvcqBDeUDCgVYmKrOkpz18WOe2BgdvgZQrsK8eP65kK4
9KEbkui0Kn2q2sJOTP1f3Xw2OR2No2E6/855rB3c1O1Hr5cZyisFOCczpEPooYdk
pgXDytueij8F5Fc3MSoM40yQdoI0jWcd9NoDwSIR6CQa8c4eJdX4V1Ys+rjnsIIg
l/XOfmWJmn/OzUEP/umpKLFy7zzCUHyfSq/yUMytq/pxWsrWc3Huw2OlStxira5+
z8bJJcYifEGqiGuZKi5g59oajSgxjaY0k5LShyHJNyresfdIGZf87i4fegLu8+1u
`protect END_PROTECTED
