`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VsWzxm4gxu6lWytc9Jy+gT6rw9QLgUwN6O9tq4yeljwy7pT8slZXe1uiQuGwWVyq
DofVxKLJWlzlNtVoPHxyocoJ9+OLuACEhXGJjYHBpITM2kxpEiMzcrrLHQ1Nt2Hc
bgUc2/Z1zhd2JiCLKPHl33oHxCDayliX0n4HIkdTKT48+jigNHpLr2PyyZXAHspt
nf5AMfXK62MsiNquBjKwOuEXeUoPQKXWAxPIVmeYlh3sqGcahyNKv1ET6aAaXHQ5
oY2A50GvuWX6LBEfEM3OqciTHfPbTyZaRfnKRfmKQlPhw0zJER9oJn0z9CStn0JO
n9EuM9DdTrL2PS2Zcg6eTnamMy23McyD2xE5BIWuGucIJLXpjEU1VGx1A/WHlY2S
JWbj3O2pb6tG94o0fps4W9DOfBM3K4Fg7+wE/Y7vCKEIKAj186qDHiJvl9XrJpxb
`protect END_PROTECTED
