`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yRKOALMj5mB8RW5mi+oz3rthyh3rcxGbnk3nibjhuPndP/jWesEFWHXH/jvp5gmQ
MjtOMf0Agm6DvwVT+IVA+Tqcld5+PHvcd1N5jC+3GTCbrkfoOX3si5/4AgHNCOh8
sqC4aXsNXi5hJuxsUC4Jcc0GYwXPWlBBgG1RHDDjuUXaZdDZYs1PwbF7GHC/KwbS
JIT7IE+vFklifNF7zs4rK0LytCjfIf3rgeq3FiS4ibiv9R4gjtiLN7iHIgAFOl/d
PO2HUyHvpSU5LuolflJ7LZSFI2JyIkPb03YErETs2B7xh25a4Zz0wqygd+ovzDoY
f8NLMZsTmFS1eFztJ/aTNLqfaRpx+5ORKZQYEesdJNg3fg6ZJps9NH7CwYUWclf0
hCuwhBHClvNmMLL0eXaYmKVzdCYlXWdUOLBFgLyOQFCg6n1KNoDE9pVVVtt1bxYk
xAFanAGegaBfud8qcuIMvHHrgabRdov0dhu+/H4VOcxLwN27AEpY/6tc6oI34yZN
z4etu11KGi21bJu9wFO0BQM1DMOgpIl4PokrDTTskIY=
`protect END_PROTECTED
