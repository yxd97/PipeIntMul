`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Yv31Fwjq76cbEoWCAaDjBHJZUNY0Lh0reSM5eCgTZ6a8BtpkesW6xj3uBOdRz6K
IKO0qRVgmzjhfD5zYs0/wpwRqM6oICEYQhVvuyHZIOF7LFX89FWHTtI3hac9KdaN
wjVblt7EfgJmz2FnKl8z0yX5J2s9P/Iy/3f4DdyzULV1nQto5Qo+9Q7SrxkB2YC/
IyVmDD4o1Sodd/8XMwVU9EErRzQG/HTKmptslT8g6G90Xtn1OO8CB+bDt6Hu6ujx
gPLPvLbPEqvBK25L6iuRhQXZORCsViSzZFh8HmJiK4jMTHUeIMrAsD2ScBiDEa9K
01+VBSJ3g6MiBxAuNHer7KbS2mzRz4r8gPFz8lSInAlVOxU+yEI2neCeex9yf/LI
EnjD1QqNOG+j1w+t1zhYGsVmVvxWUUQRnnPwXYzeioIMkAy1/zUJY5Dku+2+6vVa
`protect END_PROTECTED
