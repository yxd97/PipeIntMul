`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Udb6yoFqyRhH8sB06UGUQBSPmqUdgR6GrCUgrCsh2W/DfI72Yjcmq1bJIp6dAthg
zf6iJqDdNjvM1mhRVQyQA3IGl4I9CKhSJRvCF6QjJNuIl7f8GTo2KnJs4R281Fnb
Ywli1mH3hIkNZmZIwDWI//H99KK7um/qsZZUYfX8Jz5aKu/pdKVCTX9MzXZOoF5H
YQyOUpBMmXhrp7DnkXTRExsCIWfRJZY/AT/SS9+P2TKcQY7573HujrYoivZrAocT
08fpzLWQRPYSzKOk3/uZEg==
`protect END_PROTECTED
