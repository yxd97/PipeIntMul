`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ofmmzvDNZJzq9Q7Ly9Td0r4LyIoT7ltjGNo9AmJqQtUr1R1AmKawwUoxmzSPifHn
gXk5CMdK0uERUnE50zJ4800Fh9oak8e5tCQj/J/CV+AKSvwP3n5objAHyJgeXcJe
s55MFjnPPrkBXiKP31rVVc+tDuhQKw7gR4f+zwYf/LUelXqffi5IeTIMl9lnBKWo
nUhrODNpjsrNOoX8zyYfV2y2c27VeWfaKE+4SjRBNeGSdcY1JpG1k/ZOh0xjsjEt
cR33PRBTQKD/4gAYav+cwHHcunBaJcrbguO1qDBQQsKo+jPq2nZgBnUuswUdmB9t
XS4M9GHvhNu6N1loNTCKPjwFmNw8TI6w6cKMVDYx+4fHsMR+k8D+DNb0tNHUefKL
d1iX9AFxZqfsevVVp6u69yk++hzr84N2zR7Az/4Yrz1SZxMLE941Y0fEPZEhwpyx
nSsHgaS1uo6IwIwP5WOzeALSJlatf8YZTZ4q4zMhAdNwIhhr14YGlYSgFA1e4O8i
lPu4pak47pUdz1t6BybTZF/pGdrXPfv1E7QWuinYvZkikdzgKW1N9AgrZ0TGZSoj
tU8QwE1XNqQk90ANKOPKPsxPzt2QFxoP7WDhKI4Z6dbT7Y6JgHNTLvsb7FOjPpUE
VYAypWoLURLCnvVdgn89xiThETaOG1pvsLNQzt2cp6EilpVg86b378r9BIEn/Yes
IZODrLpGj8SdiW7mguxA7XbgmlIaru/4BuxlbYbbOlgDfWZTaBgnFAOT0y+eQ70l
3YjBmBmbZE8N16L8TOf3TA==
`protect END_PROTECTED
