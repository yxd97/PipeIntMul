`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ac9xTiKq09Uhn7o0Dhx3vI7/9Q65bZ9vV8itpU15DqQSScH3x20TGqjP749S3kBa
d5IIoBKKaOgEiacsqf4fqH6GE8ZVdKASFzF0nieigdIbwSrIH5sHnLLuHSzkEf0y
Lkc4p6drRhmBozs+mcjLTPytFk1Vrfxv62jZsxXwZbFqUTMkWTVO0SFWn59mDIxl
sXEjaxr4U3EqBkUQdLoGT8xxAxvbQtr+TUjvaolNOo9e50NcyPPvzrL3KVq6+rFc
pBTG9cp1KiFLuORaVeTXGJGRC7syEPj5B2iSGOR3nn/CkaPjmuuQPfMYhjWMEv2L
CeA0uTCOCVghGLDsdT0pK0b6qge8NkdEtEUEPIzATjQQpbHmd4di+/HkOTfJ/xlh
OVMrx+jIUaR5iJ3Wzh8iPqkLvc6A93QJCx+J5skBv9KovZNFK4+R7gydiVZ4Bm8P
ccS72nE1vYdGEeIjDmwVklHZrNBr7mL8GgbHWWObxj4JNGlaP0j1QtXnRY8Icenu
m2uqIS3oHj9jOhMLbsiisCp7nmc9TQviEekLqq6CP+/4EW5Gxb84UvFTdyGPpUEl
EQSecEff1YRvxxhetOWuLeIAxiMUIRY18tVRh/8nmiCKMkD/q6KT2uZfd03mQkFM
N/VbBEaDrz/On96lDncOwA==
`protect END_PROTECTED
