`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRn9jYTGAJ00FR2/5JnYq8HJ/09uW7YTe1YqFd4TO2oSxLB3ZSVcYiQFgR4G77Qq
ixASCA7NBL+J8ZFBvvqm4QS5uS+f+wbUifkKkJ02Zr0ll5wN3K743mOmJqMlyGZ3
/OgeVQcEiSUUT3KaUbXaGUfRvuN2V++kYq/Rzcd5CwK9G/FbGbG0DOstlD2tXYb/
G2odQC7jCKJPPPIpPmaiOxAprC2fw/2pDmLVTVvZyirnUMpnRYhavwXmXDoKnaBQ
4AyOx/0hr+Lg15W+MDqVy/OYwHkhDMB2oRktzz6+BG6T4SpIcrF9t56WsTyaNViR
DyHPDpF/aEEpQvHs52nKh2QqrniEJqhCBfKdbihtfnbPWUIj8h9E4vRZo8jbn26t
OOveJEdYLFVOWuPngbifwD0vIZxnjL1Mbow00k858tjjERPLIuqZlmvMIELKrB03
5kIUALeAcveUihiXJOBE/T85ifk63/HGjMZd0fM2OvP71qT3fkWJggDkvpUPDqbH
whk8K3IG/enkbhp1vh4RYkDssDDun5NjzFbyQ1cuY3sD4UDH3fBaU+7WS/9fZwD5
iJHz103CNSZ9aiaU2FHjw+LwEV7Jg9rWnMhhR6KmuDJjtYeaNcp7BH4uTbgig1a+
NgxMO7Cr7OAB08vlZATsrrhdMx1Bx3WSeOXcXRlMOxtpnockrIbXUNeFy6MhPZUF
CF2+JRe3ZfBydAwr1BtsfOa1PbG+jmNPLshPphAgZo4Zkc3DibEcV+KdJYLcCcBW
9xiWPnyr5EXX5416Uo7nUfiGyBlWgcS30OzAT5Oa9iyy0bHG4wf3re6LHuXz2eAQ
OmiDodwvjV2TIkA4GP6qdID2oExd6GXHKDhjxbWEhDo+8SOIPAKx1Lp32C7fF2uW
EAc2rRiR1jNXPlbam4Fn97ezVGj0djZEdSRfeAGdMOAvjvCOmyNisJ+mDXHBXZuG
VfBk4lfKsNCQjByg2uEIRXYgpgloi8nUMKnXusvE3+F8BxodbjbUYz/mvoxAPMsW
NwIeGkRH9bn0MePo/K40hThCW0OKBU1aDjg2rTguF1huvStkWcJly+xIvhXoc1+7
pgIUFJD9mVAq5JlT7Tt5CMFYc3ESkrRD8AI/WlZ1fle0F7QarjF24fIzhEMKr2qk
wgIAVf8NfzcBF1KTgCo3FV12B4C4Yrh5EBIs5D812YJDUvg+2MNevr3DYp7quJ5O
Yq455cHU489AJvRp2E9RBxqs/DQNjqoy26l7T33JgM07rfde1U4sPM9Z+GxdY4T0
RqvOjOqko42oI8HaCXwwUBd1r9bAlppiwxcMq2Utc2SbuIREgf6oZ6ZMi4a9m16e
lwD48NVBw7GF3E271wTCIdax8Xf1tQji3zWtqj4vdJrEZcrAcvTJPeI59I5nfKbY
tXWRllurmtzrfHB1Uw7wgOEwVsUCw2eI7Z/EX8ZRXYBqtMap9xuHUJhvrLJM0ccv
dNK9m1n8oTk52OruNFOM6tAUld5wNzNuB3E0otz+6i9huAqxAILbbABjE3UyDskc
Tk0YCihpVCcmN53nyW7gdkMw8nRqb2c8CrI6BCou39dRytp1iz4bpVx+22UezGN5
VsuzsPEJyrX/cnsdqLotZCP2PRElKCoF+xu+4uBWW+Z3OJ8VoBeKk0r97krVJeF+
B/FwINCSsGcfHn2QmzsjtA/RKxHNNXB7X+8qKbmsMhVvQwvwgLpZosrgJQUKEfpb
vRQ5DqILVogbXTM7PDAlIpbBdtjVEgn8EmhtJaJrkh3os/94SNrZE+BiK+WlF4lG
s6/YD1BtWgsXDlif/mKkje3DJmRZcotllUNoW/MDV9gpYR5KWNG37OpgmhmYExae
aT6nRxqll53pI5cI29Xisca2JiU+X8354kAyIokoVnbyhgwnIoCBSNXfY4xH+sgQ
`protect END_PROTECTED
