`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oxrrnar5umX4TknRxCJLupGyCkULDpcfSqgCoe51IUvt0UJDb5GFQyPrhUb5osso
uVjFx8VHAi3bt3V0CAgNOsQqmwZloMq8LBMfeMAfeN1iDEe7NISqhU2yWlxBUG8V
3Le0FtskncEhqaFZYCHrEnhmguLfxndNYPP5lfSy7WXPNLPCQEKk6xezOcp+ss8V
EoJ1G3aoD88W+gYIXsSZDSxauHYA5O/fcbvBKNPR7TZky+G76O3qrvr3l09NvFzb
mHQLo2kZnAlDxng6HhdyrFlypW8di9NZbycHt2dctLv7wWk4TpLDj+0xINsvg3lM
pQIPjkg6vu2gQpTbQ2n+hPsm0iPA25m+lVcEjopSIag=
`protect END_PROTECTED
