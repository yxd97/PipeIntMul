`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jDu8vDxBaIydHaet5+pkP3ucbDfPHLUzJXPOvEkxeBxx+957kcV4xUJinzI6RHzc
vxV82UTs4mnR2p7dNZzSeGhNX1k5W8tvcTsiM3gtCE7nD2riosIYK4Z9G2HxDc0Y
b9RwMd2ROc2yPFF+dgsVHM19gzf2NMSCyPpP5ctfT1GXCyq7bMpxTIBxk4BdaE+6
u+tnNMaYxvWaRNbhtI/e6N37hzPyB8pmlI+ViYRdmuDa/wgWHhqG0lXXSccYI75j
0+hlau3OgAFQTBVcwn1JQ02LGBdsvhD3cgl5isXKiGvvUnfxhnOcTJL1sSdrET0G
mwCe/S5q7ej1mkNjz3DNC6fdQKN8BJTZPmj7eSzKrzdGiEDQbIeCz4rOt6HyYICO
XZridOJkGzcOo+oT96mg+w==
`protect END_PROTECTED
