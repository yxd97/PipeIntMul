`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7k3adQFKRMYGlLAllWqh3Ae0SMOSmndCbXq7HWRMnjWYv2t0OrgjIHDI93Ley+g2
s2IDdFxElfFAxsFWmzzdJQOogq2+mG0PSVoKvFH0+HiJ18fvBk41irrT2IFQGZqs
44w41zlFM+oXCEXmF3Wj/+uDzBUigXwxarCEddWHXZMmVyinYDVk28sPc9jnAw71
HYzdJIcWvj7r1DhiWsrtYZxGxu431Kp8Q/SKNQd7iEs4cVj2I/67ILgYgwS5weQI
5F/gbi4aQUG74H/vtOb7K4sSR8jOYZnahb8fTDyF3+8KwLXEdY405GETlkh18EGe
jq/f+tzz+4cQ4UyZ39lS0xT9+gVmBewTPPo5xqmPBY8AXDHCjOgApYkEpmFUVo0f
8GLcdA7BJhlCFoM5bNegWUphQctfdSfXbT3d5jhmKpk=
`protect END_PROTECTED
