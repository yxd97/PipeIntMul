`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+JcuC/cCNAwNv1TS7f39Uh60gabjpJ0NwWkWMOU3W8bzhhLqIVJKBnXFIzq9Njw
RAAdfBVX3frpMmC2cwjqW5EDQST0dP88/yUfTUe2ju+/iCaw+H4d6UOhOEaGoI07
t67Fw7GEJ1Kt1mLTsg36StdzKzZ/BBF/l33vJ7tYd28xUsEmFU4w/h94tsbZYvkI
DUSI5mkm0qxogcv4RNLMs+AlD7vttwZ3lNWArzmr5NXsjcYvLvWf6HnCS/fkb+R+
8chNTKTFROBksE6uSJEO9J52kSqu1Q/tcZz9HZyBNAY1RkiZU1weue3j7Q01wmUI
hZ4cywwN72IcSBQOzsw6boXFpOsA29ldC38bh2Fixv7h4D2L69EgyP3C+HS2t+FN
FvNNJ1GPnpSET9TEwecpB/Ao/FvZ+HNvcBG2Pkg3cTyogfUA7gFJ0y23/GVHtT9W
zmit7P+VwJSIoIsHEWNR6MR20B2yhffbJdrvbwLvOO8iTZH7690vtAZ/uusZWEjO
StbHVmGPjBwHZ1mrxH8pOHvxN72yqYhGQxTVa8z+3DneIo4+RDrV425KNIiP2JNE
ylWncW0DLKcL2jVhM9ED3gz9KV+Ux9Ifkcb994I0FexltFvOLscKbpANblpo0ClL
mswDB3JjBlL5eCydoMnzjRZGR+S/LuAYyEIil+Jgc10OYB2lD9rUmMb+LYbJEJhK
VVbIuQYH7R/eAF/D/yIdcIHBWb57jMigYC2sIo0mloFmD9iCUuH8PwTvVkq5N/HQ
zLvk2CxcsYzMz2jV9DTtXvMrLYK9LBE2YDnh5primTUnFm5F7vVkfWHD5FQP5Oll
CHdJDEwI8u4hLRikwzhW9z5ffGOb1xE2kq+yWqiEj7lFJTyKCaKAqgeVeOz7emLr
9JSBGIbSe22umYa09CHjXxptYxPHFilVUssFhDq6jxVq9Gb+sQuA1a2WqaUDPCoa
wftdsep6bK3xb8HVUSE7s2cZBbiaPpuhq4WpBe7ZWn4/ZrJuwRGcHpwM4D7M6Pn6
KvxLE0N8kHz3+KeZVn7t9rrXrXHvJ0Agv6zNe8TZFwYDm/+8uKSzsMKWuFv1MAp7
gTSCT1VzWAa0Dp/xiwRMHnDwr0z//d5qhLxQwkymV98mbQBnEVUlfNuiod5ol72O
wrBg10IekyWJOFgfU81NAvGtngbceQOp8huaGQp1mFBHVZmhzlLN/DJpnTPy3Hyj
R7fOrnJbwENrJ0ouwseYMTnU/yVoUprfRa1ZSDTmsrG8UMDs6WPFjb91dieNfLUk
lVGs1acw9IPSFYrLtpS/hFeCciTIWS0zbIy92bUu7P1E25fD7C7ok+0IpsC73VOg
/u3gX0YtlK/6z3iaWOikx2uZLE1SFmmZHuFCMianllA+yCP40U9EkUgi5v0tllWV
uCMX6SGezAKOKXyOPHQJkCBnO6UyWvw9R907Cy34H7DhFJhxtYb/x/ALfKJTAPxP
cSwB89gSfociH+RXWqzld+G1YIfdxVWHGUjh1F9p/SksUEoABd/7eATRFvyXgZVd
1ozugfS7uQO6AYJkinzTxp/tzhC6BX0OTeHES4cMYFSe3WIH7AnWI1myt4BAzjur
8bG+pOsKjFe946ITZbBk/TiRPcKX/OIrbtIpsxm+z4YxYpWHZh95M02/cLM/Vsq9
Q+SoEysPiI6IvjOurGLGVntDGV1G5Fz8oA68zmRQeXbv4YoLoR3zO6mFFcntRdC4
1lN+1JoUHU2B8htWOzPS68hGJSMtMwOjZG2qxcwBDvyFznOj3qR/xdP8oxk0c7ln
pehKsxYU6drXndEurxbnoHg+MDm9sj0xihHDSBpMjXZARajHu8DCmLjxBuLnCaeD
OxzS75yFWM4jJ+abtLDhsROtG6C8UNygv/ZBKbaUofPh6DYA1SKh57k/ylgtBaYz
YnjV1RmtavFCdVBB/OJSHe7wyj+xUdtcAFfLU3igFUBtdUg9No3jc+djlUJb/IzJ
13OXnuuVTz1CGpZlPvd52aTloA78eQpiZKoT7+GNKycfOlW9h6ptzpATf7xAfkwH
E9Ga8fs3RMh3oc6eG4K1iUEh7AZO2ArMt7SGeMvedfZh5/5JDeiEAX6xS6F0+wE/
SYs1oV4ExNYvh0YCqSVTzzVX5IM/C0fOBwifDktTCBd/zBVsM1T5ZurXr5B3EU8Z
tNdtiVeyp33EtReOjuzWT0lhM5kLagHXapvosz5ajDCZLidokGUM15+KZkp4Ttsq
JGX5iK41B6KCxtcwi42w7nT2Df8YgfKIUCpPjEvFJZEmqE8PaEXnGaIJQEl8Xxlq
RW+Q1rDPKX8knmsmKap6I7zga7RSWjdHUSsUZ/SMGkv7Tn0E3wS5YBYhuJdAF8Jr
VcI0qg0AsYE8vDicG8MTdCHmXzNlA9iLJLazqdqZORjcFYEtlanq0lO5n+zlZ+3g
`protect END_PROTECTED
