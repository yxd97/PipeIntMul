`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9TILlzqTb7Idx0mz1K3MDwba+iPmFMKeTUA3TXYQCOeW9bNbrL9ELNerA5O79Fcj
ozK6uvHjYujzSk8Rgjuv/PiIfDqWdG5qi7L5HZSBW2Qrbg1chezKaB+UiFCZrAa0
kjWCsTRpsAzrWb2r5tiSWZM+KjOlmgmL+kDrgS6ifyWNHJZ470A9qBf278OF0epW
36RNbuOqShbw7TWLsh0jpIIfzVlzqUN8sl+UU+K0PDF57HmVYnHITF7lT69Riqbv
DLhxjsDuHMFKSEhNqr6KjR4R5F3tjRfARfp/dr2VsJYMNcTZWLSDQZkymW/cwILS
7XPbSIsKRyZvSweKxmHLA2TpBCXUVPvbiJ3fiZYtCBb96b9hZfe1HFQZ7IM13Raf
dtqZRd5/J0pllth9ZNHRv4y+CNxWxUfHJXRnponPbrYfJMp6Xbp78SIY5lIjPydK
fvdlIJ3RLCV/tzgvOC7NxgoMteQ4ylfRRvwjTyEUzmJYP1ImsXA1DlvWFU398vYV
g79+//h2kndr7Ze3K97P62C+Ry/CGU5K+Pknqw+xXZnuwpP3//QPEubYXAxG+OLZ
CmVJVjDB5jRHwWXlyVCgnoDp3ctOeiHV3XEn1kaCH6Voh7czzw6zMd+2uBOpRm+x
4tfSGibPqn5LW3DPrKY9tbOp1icYPp5qKaTzws5dE5LbI69g7Xvfh2xc6ic9z0Hz
deG4HzEYaykDI8tKiD2FMWij1Wz7BlvA7Fvv4Wdy2TR4EA+n8cDFUnsrMJeLGQXx
HkPQelHjcRiT688hynjWBBakte4+9/ujWU6nX7Psuwa6GVz9K8dGm5KQ39DErzO9
HqI8oKc3ee5vpRArr3d0ynVQiTlh1MJHZABi3DS57cxz9DPTfQBdD+08qdvtzY7R
0QHMTn03JIS+HoqasrYSyB3imr/DS9eSs1bDaWdnp+M=
`protect END_PROTECTED
