`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bXXlAMzkbnDLRg+WCzgH3fHRohk/a+iRrJ3AYLBafY9IzZB9rTNAQuIM2vhNrc+V
6IHWJ9E1HYg8ryTfDl61zejIz7k2WVTddOu3QKb0tLHI07U9FwtgKEd9/+o14U3s
HgwO+kDUtNmUnAjGI1kT52muEhMKj5f3qJIF0s7+wqmXpr5DWC1QTS1PPWpYzYDr
YJVOdnJOt9xx5p5uIqa9bkQE0flpcbfluDqyddfjbBwWCZRLCn4+qgrv3xRZHEyu
UyAYlxQmZ+rrsrgyW0y56U0Zot4H+xqOpHsPIGE69yX6bU6VGCNfkxXp7i1Hd2qM
+VvH2E9b0WCujR+eN9/R194qmeyK0q8ilym/pRG6oFuDFVZcZuBc9vS5yIBDGZvC
VYmFdLXeNbBc6nu5IoS4HVAFI27rKrbBLHFX6eg9tk7x2SMsfBDJ2MgJlELq7Q8o
1B+VG+DIpzm5lgEhByqE0Whim1hlrWQ+Z7YsKUiMDnoA4adHrl4WGRLbxhAIMa/Q
cd6Elek/O/0vnA4oA1gz5/pUhfrl1LTnXusUnj/g1v9nKoOQpZmoPXGbViWywh/P
Ro7xLJQ8ctOVSpU5zajoB2xa/3VdxiJBmL8HhwmzsDcMSAV03GMkdClUfncKlWWp
FICJjdKEt6DSxlYlNxE7gKFNvtv9H5Ni9XQlsXfg5biR/7V9LAiGFc/6ImLpyQKb
qdOWURJLnG/2WyAn8d/YzbRJC82wC3+YIcDBVP04fAldctmpJzAkJcSOy1pTMrx+
MFj2iT/S4LrmvTrf5gnqUVDNshn7XGmkqwrxOqMNlwiY5ve0dsl+iqHrjXFaLmJt
zl12suSYS7urc+IPp8mU8gL63uTqTb+Tpk6gG5H3U+05twyiUs5NvGoeG76cZE5k
w4G/NRMUVCnh2maWfxWPjCWf21arV9LVprpBYWWBHSt8dK63h3jdbINQgPQh+oF2
6zxYqk/JtOtERHKFDjXqlCOSeRc1WHVTwlbYaJdB5Rd90MLiNGoXwo/CPvoNS6bv
GlqXzNdn3CKLliQwAuYdaKOSueHqbRFodUSBt8vjbr0pSXToHivjWlY9gxAMApfU
Ituy1NBqy69o6PPmiTHkAz6HpvoX5Us0mTMWgbAHbjJVHh2ghROtk3fGdbMgDlBz
pTCx/8s+PIFiHipjlVNgwZHURQZmLybm9Q2pTd6a1e5xX3pXR3x+t0nWk74us6s3
NURqAgOAiJqodxAPGjVAtTcDVd/LnfmBYIHCWBY/KqpVg5xpnptwWhxweIwrWhSL
DbjT7Lzs/4ypokOPpMUWsgubiINfNCtk31NRQ8bBuBbe45tTw4eYNak67qaO2tmL
3XPjnW0AmVX2aqAbM6inPmOCiFPtt9Q0K8yZ8b/BkYK9333iCrIAO5zxVRtsVK1/
GvkzKmYzq4GGIMKGnawjNI8+Xo0/N4gA66vkhGeLid0Y4eThj17NdmoQ59smFjD+
26fKAm30jcKejzPpbVACdJ4UmF8M3SalBIRWdaV5xp7bLq3el+XOY7dZuzqXC6Q3
qIlPbhvcL+yqpx2dquRwWz1IpUkGETmNPClnZ4Rk204yLpJldpzbxRpAV09uuGUr
64ap54CcH+eRtZoxrSEFsjHIYTme0Z5WXN0HiIVcmHe5x1Mwnn29Hx8eCaBUpr4W
HH1Go9kOIyx3W4RyTTi4lj6MXU4n8hLwRQUc7bJ3zN1Xou5rtvcLE2euNyQ/JggH
5kkxredEUdJSBR+8/cEyCPDoIzw6sJqp7V9Jvn2h4HEvKWG5e+0+LEGmwqNJnLNS
s7BcsJrO2OJ2MPZlytejVufUwAR7C7kKjroqFToAFFtsjl95dA/doVP2KO68WqXH
xovG75O/XG/mO2KGjj2yI9gzATnVymPnOt0123GnGpTvKMkGZX0TX/EtIhdyvb95
G0BKLivy55JbxXgJrtYh7r79jH1Zz+tr3u+1vrCm3fxKSZSK+9CwqUf7PGm1yD8/
YnOppjnCkJm8DfARtEhSjqY6NBadRTeJcB6DkNUKKyY5vmNLMBgHCzmmyQDNPYvJ
M+g+FvSnb923BvSPi/EJtzvPvXlEgqs4ul4lBZRPCv4hDcAldPflPoiJaAY1U4LW
pwEyFkJgNuP7ssM9Wj+xIeW2qdFTrnrrJ1wKJ+VoA8zecfitj+tk6zTlM1/H/AYu
TrMtfHWjj7strIk5+YcC2/rn5ujdm5o0y7ovld4Y2MrFkb/0ObGqm3fO2Dp4Rqiu
ce0arhpFGz02+/MYpl6BkTxgr7pLBk8jUOjy+RzdKImDHxf3Bx7jxOvuKsuWt57d
Zh1Ibpbu7a9PWQt57uTgvqz3CsIrAU7JnMSgUcz1xt9f9sWhxp7A9shU5CLDd92d
S10NgN0N3xrqheqaOneSMeKrBhigTY42L+O/8RFNHfS4uu4CYwncMW0YcgYnBIQv
lYRzdKBuVo2sMsljtBsePtNPlJeDlVkPxwx2mOfkkEuJQtZ411yjN5qPuCfqF4Hl
iHOh++jiwTcRTVaa/RM2XGFgkoKGflxrjPcNtbE1qvjUpUheG2sBtBb/d9QhIxlT
6KkAzeGyn8EOvk/etCCKL4rK2/rc9my3cicm2Q+KW7SecSZ5IPggCgFKZyEPWx95
tXDeH+vDBY65ZwTDynQ+2CfgSDFwo1IbxU/ogLwrgSYC23aBJyBhsGStFWK7arJK
b6VxFunu7cfLC3aKKV01u3dBxlBZGwG1jaTzwTS1HukHJiTexy/c4FNiB+zEC3Mh
LyPgdyWn5nVXYpi56kl+wLXZo4x9DOg1kjftYMHZ47ptU6vaDCjwjrrx7MYh5FJQ
UXfbTxriqCiIPvi91O5hdz4xwlqViMLrJIVIDKlYE9VKYKswuoMNS4xe+8jWN9q/
Dm66xVEayPilQRIkFWaebLXOF8lRaG5tR4k2D1qT7/6PuRxF9cd7MjLrUU1Ykwiy
Cc8B2iZkkADh1lr4z7S4AMZcgj04jn9C3EtHuFJbvKczWyhmkBpV6rNiie3oxRsJ
2dh/S5KhRP0J6MIBdamJ7qSzEF+em4Cn/q98t0gcVwwkwx1zkxqh+CwIXtnGQE+X
I0HFManppN0XynMKWYp0VK2Qmdws2YVP+BhsL6UVE8LueBg3n1gEsVcF7nvie21m
aRrN74ht4T1BjuJNDHrj/d1iQqVbqPjP2R8Gr04u6JkmjUh99ObGE9KKjhtObN7L
7JtV2kRIUl4LNqDpRk0rtCMnv1eBqyb0TSI/WRlHQbeIiDaV0Mz8kVqMUYYCoiph
F/rhBkIRMJpcWQ5IykyE1KKLBz8AqDStrB73X9U/jua9i7ROzdY6dq88OuDy+Aoc
03doPSbtR0Dbz+7vA2xttPK8Ik54hVCJnkHWMtLfj80kXWRJKmgHuZw6hdtTinH+
9VsmfymzUce/UoZx/5rv7+He1oKl3Ks47ahctOw3XT/ZnBZMJKy9Rqc4oRb5TACi
qewpNd/SLskKyumL17w3JJPFZwTOfzNBm4HO3i8EXs+rNgNeH08V4A1DzWcZiqvG
5684FFijMxe6yn2bUefNlND/uhOst4o2xAUwfBO73MHZqLRBowcTErPqpPjTflPz
AjkUFvribeKs9QvL/IXW2h40ZJIiSSQLqal84P51VIfs9PPwiCF5BN2aqcaituxB
/KztphjcMIxA9xwJ2vTAenjPlaF/9qBp0SZJSiUaOK32xbVYSn60xqbjo6vPPJBb
oztiH44CVW2RMIbzQE8GTuw9uOLWKABLSJ7qmP5r4k9FeBPW+1qTS4gG7VFKCFt/
4nbnd+Lm9ddRCnmAN/ArxZ6cXMwZT2lUvNKCgABR7jnoz90BjgJU2ccwtmO/GD/O
2tTi5QTjDPXr0v9X+f0ygKBEPsokLGK2P4OYtpRz5JjkJI2GWmzAVhCpr6vgFu6L
aB5UVRV6FlWmUaPOYmbKT8NVnmd9KH3PqWLlw48+JQBIeDXASN1Zfv2/ZDoqwYuI
MYmOFuhHEjUPzZAMf/ehiEm5e/kqn2ls0Fo8Jy2aDmo/gzkn/dooXB/tMf8DirBZ
DEkCIy68IngKaBPi6TsWaPt+cNJdhdn7fmJ0uGYRTVZUf3i49oB1IepdNu67WSRJ
6vPpTRGpPtBXqJgfzE95J315pln4SKp4rH3TkhXyvcXdo0ZHOCdhWh+0xMWoodbH
sanywQKYCFPDSJ98wFtg/afy6LCuCCubUxBmuLoQYCe3K3Tso/l9+5etTQmFImqp
RhQ5dBHuVNQASFMCSDSK867TMix1A2njeglbLA9HlI81ocZK+yktvO5ieZRrpK8f
xG+TkxzeJHXtAE6NAfryciln9cR+XuBkaNWiXhduEjnL1m53EXfYZ0OlC+bHVuM9
NKpuMPKgPYjdSzjzNFg/wKL5kUrVsZ4w9X90oVfzeBuaY0gvWCOblh/EoyzwySuH
37Fp4455ciH2q3GsVx+w+90JbWOlYhgB+3zLB3aVsGa7AhlmRD95ia5RWJpwVEFF
t81RtwBhxdD9+kO7x/M0KNdw9/8Gp4NNplg3+jO4VcemHgjOKWDTMSj3QD9Yx1cQ
qOkluRg1xvfVlQrx6AZVC77bVhN2+5XUt9yhFWEWTueIxnoFzOp4I5pr2WAdog4Y
H+UcY5dUPIiSo1HH20xFMbhOCTXjFR2gVnXw7BTBedjeolBfTyadfwun38hu9kmC
FB/oc9e3mKeV4zvlutF3bUJ7a6dtY8nSVMi2cfh67+z/BpJnrOVH9b5V8gdRDf1A
h0rFir4NB/QlvfTOJNzsKs3nTSRDVjJSGPmMQ7buxxplUr5cGJNenYXpk/d+yyjr
TujnmhF0ELrMEgvwmlujEykyuhR4WKzx5TfK3roT2gKYkCFDczHGX9rFMce+NyS7
MkuYr7vq0fMOTan0SKZzfT60hNLyMbMP9aoXW2LTXwRjVF+4zjjmjY0LE112GWoE
xK2aSfiqAVAIZY/1wcOcskTJ+AdOS8/wHLnf99VMuoWWEzPf+2XHBk/NWbmiIvuI
dPwvbphRNnSDtW/nZCu5CdzZ8Uq48oKaGg4tRtd9OJIj/cns1A/WFRpF+oEk/+V2
+W/oSM7GDfYjV7e2FTmD0T7sfn5TnGrsGhVyTGMHT0QSEy2qwAnPkkedZwQl0YGg
vC3nYmPKCcr0a6JlcPJyYrliBAlij/hgt7BZFj+Nten1pM/9va0L0TXcUdoEHwtW
M723cPvp+8wXmVC2on+C0Gz9JkGDOAUzRE8U3DRV1N6CKaKkbbyXDyx1VbQndI8a
1eh8rrD2Zzmj5WJO4vvJpXOeJtYBXm24ftnGBWlWvkzjuJSr8G4MRH6v1UhwWyzh
3fwnjY4WA6658HbxozPoF0u0m7aB4N8NZgIlK1MeBMMWEtSScWwObRamweW93hoN
sFuN7H4fFc6QgimopO4yr9zwMsnwrsvgRQKRJWQIKHDF6IcJYFcFxmptIQCP3Ihn
p6++mHtBnGUJCjPmDJDF/kWGZfEYM10pJatgc88+WFmhsVjdNNuw6qLpdA0wF3tO
JfEHl/TO3VIULl+3w59UMvN2vDc4ThnhCyxPQ4pjJatx8GmCUgzFCDsfHOJywEXQ
N4p104zeAcpJsWz4X474Ypb1WdXtXv77bERMbA09uJiYGQBmGpqZZCbEL8ju/xmv
Mn6zi5mIbo/Epsb3jboOFG66aOX7DDtDx34EjRrTcDiScRYjlJRWb3H/U2Jc/vnv
GgEhJcnqJjUwpI/hBEXUDm6UyFFqyy1XNlwN6QOdnrkx6XV0sWv+Ygjp4I62cT7q
pq7dFCtOzVieGhHod8eDWBd7nhx1zIqTY/toWI/JVNaK59ZX2mgK0vPhmtad1GJx
DvNNRPIoguTw/Lb0IWgCNS0Dg6nT8sx07Dgxi9i05cUl9uwrUz5KU7/KKHaAPzJM
vaRzRnznwqUTBe1Q3EN2ipVl9sX77hXY5OY0MfCpM5HNmcCF9O5+wi+1FzwhKz9U
WMCzDwSOv2l1P31MC2AW6vC4sd5cLTWFpFrye0dNqjv8vl4aBswsuiA/RA3OilNx
EUURtt+u7oCxEz6oGr7iL08qflbTjq1Gg8NtGgA3q0AoQJeucf8IXMQimmmTheLe
NYgkeN+rhoGZUjVANEuxIBqPuxQf0VI0gKcw+aFFvmXmnVvZeJI4O77GwS/ffYy6
6iUwCGCDc/C8tq/X13hSLA3/0lbmRzbjVCLyocAQ9zV3wbQCvWajnfYRy5ScrVJl
Y6VmhwV6KW3LRHRe60mNbC3KJ9vWmk6YiCPFN7sxCWl6700viVPRqIqfBMDPdMBj
uML8E/ufHc8rLDKMmMub5GGumM0XRtP7OUivQ+mULrXEfTiLLH2grUd/qrw8cEms
+KXKoUsHBUQ166laV0wQMbybb5oREz6fLHM1l9viq0i9tnIvkn/iR+2aFdg1HAqZ
YpUuk+hoByjpEzwQf7JV21aKFWNhBulG5DjWvZFMhDxN/isbhVLDiKGAh+EIxqQ1
+H0LJeOP/sOBlRcxsX87F6zP/DE1gQQVt11jethjdP+rMFAZnBr5b9v7APTjWGpY
N/+wqTvxZGqv33FMj1XU2lkyDRTLM8Rm4DX1HBfAOAURQhDQ2wAq3uumWAChD87o
zwrv7zJ/jClFTuo/0578xQdDbPDYbbwSfqKz3mlpDRM8peOr72+kMEPibTujLjro
Ao6NFpywlsk7Av+8kwTDtnCxyXRqCOM9oj87KkgTeRis2hlTfa0OiaG1nU3/l1mo
7JePEwvJJo4W2Q189HT/C/4PTt2r/fCItZJOVQ9rtgnFUdjVNnhOuZGqN1zGM4z4
sICeuhVE9aoKKErxWCfdLFlb1bPzhbwm78OBW4HzTnEWmzPZ3MQPiMmOqKUvAQ+f
e2ElxbF/XuCcliKBELGJl0SO6J6G4ncqhls/2xAcsTjorD5v7/L7EERnp6Wzz+ij
L/DsRorXDj2GrcGQnoYLjZJ68NFT5o3hE4dsxIHpRxNcm3XiAQLQ2zbch+ukPcWg
8YFdYmTviHBn185WGgk14EfitJA9+UGTlXJNC0982dkAk7b2JvvnxT472EU8mA5Q
b6/apPUclBWG+Rs+/JQZlp1J2teQjyFxxtTWiXgs6WUoQ2GPqOrzyyyf2OnL6/Xf
TlWmgnSNMGu3thOxyhRfmz+ooPmgcNxGRM+04YU5DzALUHwkyKdaZtXnlvxFoKEx
qZZ2fPgF4Yzx5w0tYJ7Arxt5dT1/gVU2qLICot0ULeb+bBykiuOgkvuI6V4sRJl6
NXTfEhu08SKlDDsUvyOdgwP0HErCyo3Dc4lZc/e2/Cib+kcFkIO88ZukU2fkVUWJ
/ccpGHWTeMwqaPIKrOXOTY3bmNh0Olr1pyF0uYuLKo+Vghce7cWlxJL7IBr0yn9g
iVD+z6Y0vZ0Tv+C/jIt3qfmRqVw6Olae32+dh817Iz2W85YTVHMBU2sDQ8D7l11W
X+5gYU1ezSrBq+Ge4eTT0KlHh9+hOkKcSvGNSkVE6lRCRBD3cR3SKGm1wuOjNjvh
IPipmfT2WNHGX4H0oEs2ZRiRTC5OhutjECYSRJs3KtHeqB8H68oyVRJyMj6/qMDq
cyHVYEUm6D1ZK8A8DfvlkFqh/9e2MOAq8ihC0nTGB3Rd6E3bH13HeJmaX7V7NOH0
wy9wrPUQKX7az751phIZ3AcdcMIrR+FfQZvE7C4HE5FQG5GYB9xGH1kmAP4BFlGO
wwwFRJyIxd6m5CC1wBSObbvzjT0XRFtkl7bVgsR4IrNyuh52BxU+RaD/xepp5ElI
hN6prl6yduux8KpgaD5GH2PnrM6++Rv6KY3CuSseAXvYTKNKJcKPZixTFNwbhRrA
JAKoiiJjECPPouSDmIvpnzGHj27MN+T35BTHjAYPh9eJ0m7EGNI2SlWARjigiOYP
XAPogHu2cPPTXXMJKXtafB5752M9wdyvZcNM4JaRif3KJHEaXc3IEb4kLvTJSlO1
p2JijKltuvd19CZV0yjHO/t58U79C+G9Nn5IAEpJzfKpxeokvbNnF+2ciwX248D4
3sKOZQTyxXDb4TmlHsg5lIjSe5ZjrSmXyTaObXc4nC3RUNMLaUuQbRDINRgOXb1N
As1jlUBiu4ynQJt1nHq2Gblsos/xvGHHN4F3YgMrkrExyh4HsKRJVjr0RCJue4Ph
+usz/cpD7fNm+Y5jE2fEMNQEb8v28l0/77JKA1worWUzAWJ3f2B5jEc2uSRZ7Ehf
Xi82+7YFlpY9RdBshFjT5/naHp5m5bMilLx9e5SgHBmBcixE3T/Af30X5da/1AH7
b8lvEAISreqsGKm4Lwe7M36kSIsnMDXYEvVXVikEQ4IrtSrFzH6ZRRDvvIrQdUrR
OAxGfJs87HgpWtZDNg9vhzkdIpzq91o3KrlY61deWWhWjtCdOso/w1R+ecgua1hh
BMgIr7emb0vn8wZi8aGe1Uh28aDi93ihLfXhMDzJb3WJFS2qdIbGGkA8rNK83LDX
aCrFtwfpiUQiqtUsFamDIDuk7H+2p4MIAnT9rpK0FNVZVTi7jkrB0xxAYzL1MdrE
IUxaAsSnHYosESrG5MqRHMfxW01JHnFpqWRY//p4C5R2LvoT2EDLHJPxY4T585Vv
CgQXAz0n4Qd/1Q11zexVB1pyJKPaiEiG9BOA2gfnKEAtm8p+YdNbOcuG+cATy1JH
c8DhAP5fI1lIQmJgJvmyYpiHxwkQLcAUTZ1aJwq4jaKtgs6vGSgsiwbFw8r2vRWT
ctvJAStO/YMshx7d4PVG1uinR3a+sjDGzJpCI8/L+ssSCo4bWvyH0hYTVybZ9Aeh
tKKLkdMZCIWqYDxmEDe20NTp2HgWq4CUpKLFiBbE1hA9kvg50NhlmOpIMDDKQlxn
5l+YbtIwZxMyc2gwlxXnCHoZ1pkY0cRyUK1KLt3Y005ohDh1rDxOE2h3jKfOGKzd
4RsAxxlK9z0NJVY+rQupVr8pstM0dAJUsheiQErNxl2obDgVn/Qj3CK73+SFF/KS
qGA5l8sh7thsUm3jfAbklEOD94Nmc+bZLfnGHgvId6rST0eJMBT4eoIiDcdNpQKV
Sg6D9mSzp/Grzab758eSL7ph1QaoTrrmnIDuZtDRk5lXrdgvly2qpmq7dZnRJFjn
Bsj8M3IGCBSJqyHQQK6kCM9OgVqDFwnGJfXfwQDEpjk0ITXsp5X1jYpintW1EBwF
p2o/HSf+UzjPLamhljMM3GHZHZ8OQO4COXg/x2xlfjEudHTN1TuGl7mlcw4UvGY3
qjAZwGVNqkLOFUrO2PQUH0N2Ng6XXzRdaMHSugsnlwG/pSsoX8QuyjrTbdGcGnSi
+92VryaYZNN7MShsXcS4mrfGiDmX0fMLOFkHsVAVqT4rcFim5oe0+LieqA7mAdEv
5VDQ3N7e9GNbjwU3TM+Kq4RfM9pCASwE8UIu8bElepkD7GCwNQ97jnG5gw/VtH4H
E9aKi622rqvKjT5xqZDLqF96l05wWKmKpX0C2BqF64q1SwKYaAhFNjt0FYqdUzs/
o8KSd5Jc+8Y30jVKbgg4swARiQnBjuUEwO7NjqkhZjMWVl3BFeFbiQxv3ZODYJAL
eWzPtnesMkwhqdL8sK1iQTY0rdzsoDc8pwTK2hIIEnd9l6n3gcmjpR3lUr+u+/pK
oiFpMKeos/lQ9TRaGA3/k0KK16NOjl+bFCJrL7UL3LebYN6V2WY4zGGM7G4CCKe2
pGyis1+yCua+yq+lRra903n/KEPaPdquSDxaLVQFJD9VIgrUqnOTUBnUn/sb88GK
RjiwbiZqTHzUGuzie5KkXRWlICeHA2jml7uy16t2RpG4c249odDfR6hfwSM10vv8
DAYjXH7QfJV9Kk8JgETorVkxOMCl4D+nOjLorUhf7GqRHe2xCLibBkCxBjVY5i+U
YvNoV0DUq35JiLWRs12NjKv08zbkvyJQcrd3ZLjkLfzf7UvFZ6M9hzwcZGdyJF9k
iFBfNMcevI5uuqgcKydqfmfz/Wwia/FpmJmIZa/6rTtKCJz4fQeMBOI9d2Aqu0Cb
lnOgvhOm4D5vyL6otMwnKcR1sij/PQEtMFsaQm8kTFTIivYS0ZclaSXmeqHwaV8B
ATb/OgGPT0twD85nUlKRJRm2ZGCyr1lZbMSovlgKqni0aZhSTWrsvFAyjWQ90g/w
5K10AE6lIuZthkcwCqYZRKP9WoeSN+F3hgUb0Tp+A/YCPr8q/Ox4pIwWfoY45yQZ
UlPYOjyghxBDIBBhfnDf0f3Bsm8NXo7r6aB1s4paiJ+U4lZ3PHbLGOHZ1RHhvt4q
1LpU7khSxI5ZsmXyj2r70jc6I8spaEosPo4G+GqYdpypC5pAbS/agl+rCL95gzU0
j6Mlc7vPnIEZB7prSEgJg4oH5afa9EhlMuEjzF0ofXdou/yvy1CJsXGdJWeAqpun
JCfqtECa1uLm8NAuF0e4ninbhRP3c6hkJmDN22xQD7/iLfqTQo2foE/UhhCsSxGB
16MJxsKd8xPF7fQVxDa00XQuXZ3cn1mVyQYIHIZC5dAo4CHC9/iBcC5k8oZf/FYa
B2UsODHjflsYIPKI2REm2cCk5mcoq48jpOIDPoLHe2th4OOMcye0HUf/dA6pjGO3
9C0gfhwneDydrizjkOvHwjMT37mffuyttiOKZLH9d+u4N8wmAsNtk1yknQfjTwBu
SQhy1/fFB04C5/oEEw6LtfUErZfbjjuJRstCo3Ip01i2eONbEkL7Hd0fBMLDZhJy
CYxwHYt/LH9UM93t/ILs1EgR3WlKg8bVby9HuIQxwxEIj8IeB/jpXclwvAgBEkMv
dJoaDOlFjOVo4IgIQem7P1iENL1L0Cluvv7b95CYvQH/uYGDgo1oUrPs6/7GOeSD
M2dEq37JZS6sldqTCOOdk3vWmlE2Xgo5ejVl/oMdGgW4UHFTx4FXfZPisPZOsPHX
YejEcqXCvzrsJciZN3Qz8EdqH3ZvC1p3ncJsORq34fzOmT3AMX8b+I5eLU+iXZkN
gvO6YzIVytaqAZlf4HKF3QIG6oYjCbF9engm7g3YACGkD43kFUKUnIgrCdpS9Qoj
vvuCzIJcw3Xjfr/iqojidcU3TRJkaotIO7ULNT5twsfJUkfzNgHWJSVDmwknRU/9
xIF5uDsD/5gdTRIRKtMuilWYKZYFNxzyApzrsuz7BCbCY9HXpNjdIW+ighqsg2Ti
MZb9oFJd8aTJeeA8Izs6Mky82jE6cdP4AR3dbgIBLCT9OTYCjM7xPjjoTYig81wY
H4jBtQMtEf4nGwx14VCnu5KqFHYQNFmGXaI7TImhVJmJCTIDBi+tdyaCO6LvbIkZ
cwowO3KaC+awAMy7ozgPtudp2d/HvoxF/wnuyFmKKZfnizXFiF7BHfnt+cFWd7Ph
M9NVeCLRZvKlQWPn84KsFeSevnLWFr7ZZQ3pqHM4tQfvu0mFdRLKLBsNH0O0X4bM
wmSlxt9hPW56V2h+1YyZuH3sYJzDHHVXN2IS5yk+G2Ep2Ya2OEz9diZpxO8/Jhbk
aoghT8MKTZS8u/TCTKKzBaqKyegha4ScFiHlVW6ZZCDaYzW2a+Jxl+F0vN7QhnjL
iGYNWsiwTgsbnjtaQMZcz+O2fqD7GgKbdtY/i485PgVJo0a4o/Ks1s3ebAxsIJYn
jkQ5GQUiIr9etutmN95yHL6QjYNkv199eW/R/Q/zgoxKwZ+AMbXnrSswllOdgl58
RGVguA4Vjd6xUB/R2fmRBhaIKJvQNBm7zxsrXFq4YCMvInmUZc+dbiEN8XhSg/Gb
sg5ipyIg1qwdFvU6fe/HNu/AotMZ1XFG0y1jpm4PxbgxoLnG9j/OaKRYWtV5acDU
l0Klz7YRp9gUZI8FbztX09qL0jxVTXfYj/uP6i807sN7WMQGOagvU87XIjHXV+t1
9h4NiIPL94xhBxoGz/+/IsUqYe7y/NV58gSQumbfWH7FSQsBtZAIiZJn0PCITwXa
BZZoljiUqzZOqzf27ufd3W41YX4PpS0+1BfEfn6lQsl65/xa4QLHwfRAddVj2QNp
q7esmzu5+TrxErGD/0RthguR0WodCK+GlWKUbzEJzS//bdfKKRKENrtzP3GyTANz
YxzwF7U+giLcrTDY4W5re6tk+wCymmyIotxbVyx+CbXPgGJauPHLExrmcJggchhq
bYkvAXvVMmZLu6k90+/g0vQoQvDKBuo8EFhEGrEPA47+E6czXjr+KD7A4O4CzifC
TkS7DJZXD4SIFcQj3p43OyS6YMHwevvMjYLIuVPHB+ku5GKa7EWM5M2pQWjhnCWU
EFWqYoC8MUGXqRoFJvpM8SghOKyT2XX7/74T4+dMdFBZ/dLqTTM4wl9QlXGJO8vR
Saqw1XmzzheG7CpPwNCJoPt6VFPGAPoHcVsP5eZkLUXTre5j0EyFOsh+tK22zD1F
Tb48/eMqePX7Brps80hVUF3eZ8NHY8+0w220eIijMFMb1/YtArVsoAlhOHim9D//
efuLREC9J04GOtRJUPEWJ7Bko5OEQ8qvLUiKp3SiMve7uzPrY+rHwHDlTWzcUIwP
Mme60zx+eDRivEoMN+kpGCt3yrdICytHyaiThCODkglDTmR2PQxseIQpwkFdtcr+
8SZQ6e/EYjofmsDRi2OHTfTfkcV/A45ARgMi+AcX/O0Z9Uq+pS5D6k+cauYEaObR
T/MozcaPp8iaVSfJ9oiK2t6ecqf/3c76A0/RNr0+sc8otvrWLTCzBLwx+gcllkui
M0w629emC1WTWP6llXPUnToHAbgAUvUZIsnF/te8//PpnjY39N4iaHTPH/yPo/RJ
WDjXOq3aGCH8+MekoI82Mnm1ZDCc8QnX0F57Zg/xuAPNqTX9///E0nuhmAETzcNU
vw+vN9qqHJrMPVBl/p+oBVZ1jYvXiSa8FcVr7Y8wrAKOGTg04GDyWr2sgxuUZaQ1
gAzxlQSMcGtR9vWvH6/dEhWLBQrVkEdL7hbTuEO7zhFkd+ai6FG8vyiw+Qil4vVO
S1Q3o4/VQgxp0G7+SWpfvMQGQjdUSfroPInxYqvaG+4rDImIZqx9LcHnBKELQM0m
TuH3KTqFR1qixuJgxFMvsvF3N2uWMjkJKYZzf+sEKZb6ISdjNSWUxznnQ/YiiU78
oLQICOpg6i1TPA1YIbJALLkMkBSWnKtiOTOWVpNSIUr498GujC4Q6uf4r+s1mVJE
fVdy9uY+kekKIQJvbt9cIgyj1umGHy+i7tvNnrgu7s5v1HAinPt2yYE1Cax12v9x
rfqtm6ID7qJI4yy+Sp1fBzqFvp+NNWb4ZWHCoii7CUPH6Dus6hVTDW87P/sWQdzf
EVZyoLEe26adAMTsvjk9fRsWwX54biNa2JVvUtE8jFVD/9Z8qOhuIIOc2VA/jLwX
mfnp9zj17bF5ibH/P0AnqbmDj6/9we8Z1AUPnR1oOyXbH+iA7Gd5S+rXy7ANREl0
zXhgH5oEflcNPJfX4qQPBAksoIV+BZzZ27ODc3hylYubUgwhVarFAD6dbw8hvTpj
jdaIt9g+OGjrtOAXvgRaAMdKMnTIZBnyn+ZV3XiKJ+K/XSmaQcpWaCwx66kzctf3
12gmvMH3kNC4ViYiGf6myN8O8hBlSHFC62aSU+1kAK8iKd4rFEYzsBPi5NioDQGO
OykSLw1Mgug8eyMNzWLZMXjttwWH1mc09zWMg1ECjjGXwIi62v4v60RVOtozgFc3
XHp9rqXW+v3SDFkdrq9zQ89zVfDY8v2pTGw4lAQIPNv4GCx0GA+D5Mtsaf1U0CSO
/dZg7VemU9xnRl0LrfzQUwlxGjO5dbFwiOnPuCYnmS5qzlg2hKFdD+9GQsrjKucL
v7Nc90qbmWPc31rkjVfebRzEwSvfPMJps6du3vJnKPe2mwjtEGL6QlTdLyktEByz
REVSr5sDxDs4yc5HVkTzALk5jarjmKqqZsqc6TMvGkDv44KJz5dwwZTkyFC9i1Ao
6GSoa1WqkEJRC6KtIsbFve6J2sAz4MZ89KYr4UDUXEt54EvxjiLks3Ee/1LunwSp
8qSBoBqsoEDocsaRhM+LBfZYXmtcYXV3Oa6ffowLA9Mu+SZ3vdjZ9y6y6PzIrhyH
vxT1Cg2bYJum7XWsaB68fNs/p4RpmG/lFVR7oOeSGnI0RC+zeXNk+xAthqagM+kj
KjZ2sDp7caGRb9tu2OewbyYGB36LeYBtLpNCtdCuV7+NbEahpu6ihLlEu97J8F+c
9W6iisaVE9YyUb4o6emaPfhnOigKj4UOxALM+NI46Y5FJ8XP0yHEAImiPIUjLHc0
wbMZVFb1alXvJHPC+lnGtBXoovxHcj5+/zbzTcpoXIRC3BXp+mq+dWbDWK6QWnVX
XFULonv0+QiT6OeeAcOFyXBiHKysUN+jRX+69pO0fssvs+RSOoajBBQQR5Ie+sQu
LrYlEA5+ZseFh/nl4AewijTCCGXpVPB4YPLqP0488yNQ3nGdcNLiprhnPMeZWZds
ymkoZk4jsPXuXyvUr7dNEZRYgoTC/Z/GIOjdowoGcN63px4taHEnZJ+TatCGd2QE
OXk/0ugXLM4UAfZO1TRrwVev6k+A990XymdFTmz+yCOKE2mkzVcIj4pz8B2oK48j
axohhGtVggWNkRkTR0miT/EDwJnrCLVeKeoTQepwkt8pK0e/WLl4MQrtwYp6dnCA
xcZRAM+aFBVW65XCVhwFn39+mS5mmd5PUot4z9s1ZejKPAZnysX9DZHT4ZTgEBeg
TM31U3Phnb1t9KT7EYa+++ZlzlI887FvPpFleN3c6a9zcvNpfMXHlksDuoCdrDai
mHiIwpP2EzReeD9m7BsKJRQXDFfkfhLZWGD0K+3Q23uTYzxWivSralG2+BTeLtq8
9Os+p3nUkaXwLp4D60qkTnsvVSrP9SPMi9Zxc1W+bLNt77aoxDwtKQZ+tw7pl/+O
YtL+YkhSK5jul7m0f8iwipTiyFxtNcv3QPUhvTV6EH6/kKmkwFDIWkxYaD46ch4G
lTc8ToNU3IW7rmSXfFl2C+eFXxS3l+DDazehXcGgr2mGyi1ww948BUSBRAT3rsZc
RKyPokwI6KsrgznG7dSNlBv1lPFaq+VkA3fOkuY80qy6OCrgTF+EiGed0TDfjuHL
BrxmGMAE7KIUw7vglD6PUbst8acSiK7LzuKNIe1GmuX18ka15WuPBWSrHKIF5bmY
5pbLJkN6TH3e4iNJsHBHXoSdljlkhrMetMwLP7WwQvtqF1dwkYCXQWz54Zw0PnDw
eRAp25a0fn+mfDOxN82fWQVzembhGppk3fda8Fh/3PV5PHCBhh5Ezj/kft5VulpW
+JZC4+SHFbIdmqBpU4R1CpqkqEu6n9b0Yn8ohJkt44XydIDu6yiDVTTL1toteH2N
OEyEG6dergg7ybsvDITNuOlupGvHXqek0jsdJ/06fe9PyaipJ81lGUDWH1cyW3eo
d1FniOijU755R9Kr5vKr8lwwp5y7lMgOeIcxRWBtoTHxydb33peTPnNP3ZaR23K0
L/rqLXmJEH9G9ZAp1XDhS9m8qmZnVISyeXyacojF8IKwvg2fhMzUCFcpUIQ2Bq5/
ZRkqbrky4cuRYgnClXiQqP5NHtg9h7S6WTDxrXf9RelfHG000gH/AFfgwgHmBTV4
gmQ1En9920tYqeXJQuCj274ERtFMsJgPurbp6/9K09JO1z3pJxnlvG1gA51xt42a
xbkHtdnr3bMur1OWREY0+szunRjd8liZDnPrY1gkm5omcm+d90NzMi0896wyWUs+
rv03lMv64kdrgH2O8umDpRC9lavnD9mny3Eg0IDp+VofaCUdCsG3yV8Fd+H2OOVK
xy/kSgE/lA4UjqC0ueIwp4vHzarhvWA5M1K9WJrCs4C95UVOS7pVIMenzPGrhDLn
GhuYwFPGjbDoRelqsSnhAceMs7iVp7w8vCGDsxZEpg/u8prdit4UGmxerJx5XSSY
Fca3bwNFqkfNhK922mAdLhiAh+Bi1YxZZ7BxePZrfH95vKgWR074GUWqZZaTM9+4
Ukk9ZMCiQDFmMZ0oOupKnTnXmO+77gJB0dWRMfKx3FNEqFa5jHP2KF7J254DxhZ+
NOI0/ILaDc3afxAksXv7VdMJ00gJL5yq9kk6AbpUs5yiJn27jbwz2wX5p13da/RX
yxxRSq6X96G/2hUb2o5dVRiINGfi41aou9eoC6uBKlcdzvoNBF7TWt32TxfbAHO6
sx3MtJGeyh472j5XPxm/CnJ2zKGXJDGulXyOBDU5gXihNPP9D/MQ6lr2GjFYDz2R
SQQ6CWVH6Phx58FyO3GA4rq2sLSVzCm8AiyqCKE8zym374azNExdp84e/fcS8tKq
7b0E63DOFYVXABJYxP3cq5i6tDQ9gPCe2aBiDJoZLxR7wiE2KyEKVQ42sWr0Do7v
fpDVhl4vNRWyT1mfslQLzj1tXupfHCaI7LIrZLaPONFU0+rmc5b2R0Mz8/HeznGA
cORNi5bI0pmyFQEt1IM71KFweeXjcglsYRs4v+UxrEXwtbIE7cY5gftZXTeBj/B7
Ys3u7+VWPIIdzTCVVRZw85VJqNQIeNs6u9wg9pcWLowH2i05bXDDR2jyrS7AxXa9
ULy6fkofw0r5zKCgDQWRN40dODKU8IxqX1wqPDh9fp3ZwkISisAH35YimWQy/s/v
dfJSNfS/3ec9oCpOThdsxvRz+wkvJS32WI5P5+WFoX+u+Mul8H8lXkdKSwv8wW05
0gWRlMl4RjjVP0fEoHcd4qT7EEOVOXqe3I0CPcCeiqsN0vBgCtPK3RJNyXOv6YeA
RZomLHV84PAJILiCsFtwwpIdplpI12WSilNrwrdNr9q2cyJ/rlFloOoJFZtBGKX5
Ky/TrunhAxyNPurhWnkbDux0fWf7ftftQeoTVRuWen7Jeo4FKvRS+lndU2UeE4cG
3BbyijtFEocDm+dfBsaUFwKfwqur4pXobQLu5KBf6Zi5iXSyvb7BGDwFP3twzQnR
aXob8R6fKne80h016iYfxYso2r3IZTbcfQLyUE+9nEVAnVTED3k8eKcqSzca7xR2
wDoaTyUvdtLSYiEH5om+OBkA3oVxp5tnetNqc7m9NTqplWjP6VDCTG9tRWx+TI/b
j1/Ykgdlm6wPvY/yhBCRLmhB/dT9Xdv5gJsHsQbOZMRQ86/LBvNfP+voJY8D2zJ9
9DUb96oGt7M3EAlsqGk+RqLro73shzH2Osfh0julffxfE4UK2LcH1ihP07+e86Ul
qCVXIyfMFjgsLmShJy84QYJy2T0xjL/49NNb3xF2nYMfpR+CxXW2pXQXcFffpH6L
XoLF/ay/JUISPKqJEjXUVUU1rIkHAm2dpv4Zgr8dVwViCoeO+QyjtNZFhOSoNiut
UGxZQEPJjNEXbl8kAkX2qsJElLxtpDQHFikeoIuyBXaA2LFbZoU30ZTYkRrKyKHb
4RxDbsMkgQaEp+k0goAxmqI3dj50P9GUrRrNwx+XVAt1u6DuoD3E+c9K8js/MoV/
UrgMKjaCnEXRdURnvpFWH6iMrYmuNA+8mF+RCVS+2guzDvCgKGmPCKS9TliNGgsH
nyPIRzxEdajF+MXDKQGbjoRPasi9YzdExwxxQ8J4iq3y77GxAqtkorqafsySXpgb
SQjfLrZBqNL5pXFSTuWgkQc5eTcdqTylF+LUJfx3EcFIBJol+y3uLRZk53aqTeO1
+tUe0Yc7igmS43oHukSXTQAzej2f9+jP0Zr6aoK+UC3fSRrJ7sJcoymuUwD9fVX0
Yc6rhuuy7PrD/ubF5d7rQ2ThKtpeFWrZxorFD3Kx0lRgO/tpCz5voTiTaKc43vdS
Ff1/zrwREyqKwts4G8FFGgHa55DiCjHh25M3Jk6XRiZ9FqtItvgYeu3EvoMfyCND
wSpp/Wv/Q4UiCHdeKeICWVobjvHLilt0PhBZIim/TpI53iddXPprbWgaoQisN00p
AbKtEp3BjeggP5sww1WaxBb6U9RpuIvNjaQFRsXlkQuv8FJRe4Nhc39+WLz2+WJt
bZcEDoj0SRICKEed/Z6kzMGKH1X44UBVJds7QXhlwxtWE017oIv+Tk6RVj4BUR6Z
v+73gx5BeIBG5fUQk8l2QcyepQeTv3Ad5DKmd4Ka/2/noFfOg6joI27at426DNDK
QI/4w2QrulRWgucT4/2ZI6Ebntpa6xRiR2pCq4vcovhBFCCD0iOe1mikaKsQv7fQ
eK9rNPzcIDsTkf4VEp4xHe3BKbLiyEeO2gqWHd2tw4AsIth0+z+g7DIuSED0pvoT
iJkzItbCL8+0YITHceUrbYcdif80vu9VYCRCOShKiU503ZIMZ5Xdzenm70eH5lLZ
IkCn0lJg7Gnad6xF6pP5UsIzUsiZ6BSX7BeccAe0kMvAXUGCcdbWSgHXhxO/lIG2
c+XO29spdtOal0hpbOeJioXMcU1acAiTnUkVEipW4ux33/CA1anXxUw3gtk6kOgG
/6pEIgmZIAHhmax9Y3oy2MGH3529VpGxIsC8KFxVdiCXmyzY72YYDy9zSMSrYQU/
FsNdhUZvMrraKtj1LywGSQzcoyr5hXeF0UgGfsLC7KDvEVoac7ed/dW+9HS6po3q
ECTA8IVyhAzoXI9cBX39+UD6Tfa4bbpLyOFgzaU1QbBjH4YWnobeHR+OO9lFVX00
9nzbIk5EwEH4N+1RjSrkor1Vq3SUGvzIKuArt1cMQzxgxLzRGmSHeqUZSv/gjgV/
1EdCzTmu0/BChbBPBnjpAblt0cas2jH6pbEpH1EokjUYfFrZz8MvENykhb1bPetn
lL3q/CUQJEswprbFXEknmMTV9OXgK7ukk8KHegG2p1EkPhCvcC5+BJF8c0DGgN9T
aJFy0zB25BwxM+5oBRX2l/Hnq2UmT77o5QhiLlMmCfBT1+C+WFgiPqb8kqcPiELD
cKl+WA66J62qeBmYIX77tpWGISqAWuAxej8jXPnC2MLYO9SHGCkd8dfgjD7mcZjx
rVAWvtOS+Ba8WJnZugWAOppb1J39Zi8gMXPAPKSSArEMGdNhR+Vuxfbp75QPhx5+
KPJiqp8rNKqfajM8spGaLw7UzTqMAMuGYgsMl04gLHl8JXFFqtMhA8xfLsf4DCAk
O7MvtpO3XPvvIv0oD1HlmPTJMBPCXICpapH0X8FfygGqEXDDXXYGnzbiprM1wx0/
twii2sFZgr6gzDgDDxYp1HJyTSVqGgLKB32zcNVDbIDHbQbWscqkbWLPzBgRfNXL
0vjOzLbU/FQXQYugsDqUqeNKi/0JbkzgaUyADPe0mxPMIFSLzbq01QHIhPZaUKkZ
KmjorT8J4lsq/wJbf1UkeqOLM9PKL8rcQnL+6u7ey2NgrPOoFzI+9+4MOJRxuiBX
HMxdvXl1KJo8NH9/5c7Rv0ikn0qeYgNPmRyaNCtOIBg4/qBbd8PWG7TlM1+kVN7X
0oHD30rDiC0F3j7bw+0yKqB9xy6dV3XD17bM3awr+9TYy0AgYvZYj4INACNJWJMM
uhzjf9XF1pDunHxkv22ZxuJFky5ThTLLaJ6FF4EWQSkrQAHJ1fsMUg8mqHF5Dgeh
fQYHCR9ftOkASUeqnO6y1r/UtXTUc6mhWCIcqg/brz1WHNFTX+82+p1LWlhFWlcy
zpXJoEJwQmqvJrYkRZT3k2/nl8ZEPsHtBDwNI2BUXgHRWNQ33etbZGRycKVQeR0M
FVEdn2X52F43NYy+KlL41o2WSoA4vvxpjQ7EAQvKJFD1QosJH+tRak4ACP9j9KfH
qjUU8OyzaMBOk1XtOYZuT91YDZEzu1MVRbiO5TOhqN6o/xk4c0P3i1PDtQY5M78F
XcXPIIRjmZt9wEsl3IIIuO7N+Sgp7fCQXT43ggF0jGHAdXdX/t961YJWYJREYLlj
/l8wMGprCh2Z7vOuLX4LkTScw2/YvvVPtQ8SVQxLINzoy2j2s/Lt3PdKHiJ19TMA
Axllfo9JAglf8k0bFNdNKXeOuvSB77l6DZrlqTk/JcZwaCjFqx13Vc5P1U4PQ3Uw
Y697RJpUNAYfGDsYLWiExN+cW4BEQSS1HQcANJwzrMmZ9JFfrBcPU6+YCfFqjT/7
2vi/SSZT/KgHKrBzlDVV6rZ50S17FZDs56NSqpjNZbk6AuYEU0upQkiuj8Al7dUT
0SDR3r14/l7js3JuMUKCTZYxhBxG5vHXXzURRroFFUDl31I9CpUB/mPIgzooRLIY
idz3EbZHq6OKY798F2r7LSZwS1deZ1LH8LxDfN3xpv/j1cRAviW6T/eAIpkJANtZ
DOPJHDN7yKpyX1TYCLEYrTIUn/lvmGOhkpAyyohfawh437k6K5nvJvYsLd0hBGPv
BuBMk+e9B10sUjaPzJDttZZrFKDDhf7WXw3bLaABAhLWgvt9p+d84i1rgcBFXW9z
zOo6jf59MPkdppAatY4bmi+qZVstcX8FTSFjypybkH/csPSenqbgD51B4c6JYaw7
SdFMd3FaeEW8sVDK4UOX8F0eyu6z2y+EXqgaUQt/kD/XQVW768EV2a5g6+400s1w
ol8mm9IHfg3a8Ic/z70U42gOvcrgqF64sFS70nVk1T23xgKgpKV0dYztsC5MHD43
8IS/Nidh7fATg4en99TT7I1pTqrJDyJtkEIxo9Ia5JrFdbthHN/qZ6dGC+8wz5kJ
m8d/vApbWqVAHdnMpfjPI2PDpEXKSUfiTZa6KEglhua+RGBTVPMBOpVQCsKmeCOp
g6TfcdnnQKqfrOADARMPiQg560viz4LQtpncw6XBBaL8KCKo+vnlg9wsEHqcKU/I
rNBc/bHBGij6qdYDVmdA7WOMegll449tDucwcJy5MHa3pUx4G+VHJAm+V4eIBbT5
RqwwxoGUYXZJfCbOfIsYX8KiFXIACms2qkm3dOgCPQw/qBOV0KytEZZgpmfZ/Tsk
+QPQcAThC117P/txoJvYN33J54hRnOanygrqWJkW9EGiGscrxp/OjGvvxlYwzJi6
i4uD8xMbpaF9cLZ5OuJvP4izaTEi5NQF8vY8ZTMQF1K4kP4Vxsrr00PL6PRqOvHi
i2EJzGpDVq3Qp3OQRFt2ED+3kdva2I6u8MAhc3sUsWhu/6uJ8SHjM0FO8NP6/d+h
sgcm92KbfuZoCjj+p94AHjEtfJe3WH4D+qBJe9EEATPVsPtwz1zpTem3/by3y3d8
46V7MBxkZFzWQhAktn9CWVUlFITkvoJ8+iphgu1nc/XKFJGfFJnFMJ5gO66GK7Fc
lZvdX7muMpWf9T0U52g6hURMeQ5dRJxry9CWkNZN7fn0f2MhAoeU6BqISt0HePS8
wi9gZsmvlBIvOyV4aPXwoA3SMcpetBjeRH+9NGRucFCTBnvbw7DzK0b3BHa7fpdd
AgPWbJ4PbAEXrq7A8+ZrKEJ1JyolZ0v1Vsf80dn1KGLcQO6XjJFIAOZQ+zCeR64K
i0IRjqUN+j+OgxvgbrQZ2IwdVhdAypsqm34lllBMbehjknZvP6y7KQTO3lAbIHWa
e09XIA/1Z1+laosTyo/E5xIkiWtkJtNJQNlOYp7I8SSw6RSMO/wyMrvyaxUW/X9D
QlmZEuGEdmE4kc/hI2XtE2fHIfN0wALbdjEtQYYeZkR0T8tOCk6vEcFkeTqTORlD
wokQ1w8+lukCVFqrbwixrtJy0aPhJX1acwY4OpklbuNTnq1rg+PHvEBWMMtMYeyg
xejd7T1YSWQZiN2hsySFbRjKveY5w/JhoFKEMv40pv2zv3Zr3WmuqQqXr+Qw05rA
+5jcLmeA3DeVdcXJ1a0j02owq7iSV4jPTyVgzbANoaWXzO6NopgYgTP3OH3G64An
LVHdvsbY0izDnuYahRyYEpE9JZ2Rv6aHTPdowt8vQ9/OBPTGDBwAS/w7YTbWmSgf
sliBYcHdfkrJdva1aK9bqE/uw/SC1RssR6h9D1pJ7KRntJFB+yskSedzYf9PUDzb
oHnopFPNTISkhk/A7Hm57NJiVssfiL5dXuHE0VNrbrulK8mhNTCXR+XsWgvhNyEK
NvuuHO7qNLNYsKSoHY+P+SlOcVLXEtUjw0X1y4s1FQHmQj0vO0SWRWrG4IfcO7YU
NuEsez//EAPXp3Yj8d3D135fWOeitqyvjXqg+xi4wIF8AF8srA3wJPSmTbI3snGr
AcoltSb+6HuZU/rRaVYaqqYlwYI67NrBqjJus/9yRerSP6r9uZkBZh29fCayxW4w
jrjBJ4Pf3Ofvs55SUwdGEgj8zuzpCFVUEUcwklwPmRTDgnxQyPk6lcgmLeWRHxd6
KZn+rIT0c9kqM5Mtn2YF4CN1GzqAnqtLk9JOrh8uNmwX1qlPXs02WLqeflQn4eg7
LmIMs91OBXTbpNfDBDYusBFTn8OrufvjKM5lem/d/aWyxchWRsapPijk54QwC9ik
5CTpAz3cTUtpoTEkmGVZxFaYBMvZP6DErYap5pDDioB8lIM2y409See19y5nZXiv
dp13mgdTPfr0R21hA00jl7SIBFWjezeYQXnmPOPg2FrnIqluDmVjkwd181jmazKw
fyKCEZ553iGaWZYTpQYpgHCLcxE0tJgawGn+FcQKB7YVgMDW3SGzxr5Npi8gJY0w
fNrDXnss16tBdS4ls+2lwdPGGjytFfTKnMynqG94Iwd5rc0ZFDljKrXR0mcmsren
cK6USDP1Qvpt+VxoVxruDz5VNGin0auGtE8lm1hEAqRDnh4HgyS7UggijVZLgx+O
QIPsaC6dt4wDm2DAdLg8vkZc2o9njn8pl3op/nQera3mHfqGYY41dvDHrJRAbHf+
Vcmkoh5XRpTjOeAErPz8fKD6YJWVC+jab7WBfCCd5cD3J5b/jk2DA115hKXQEqvE
J1X+Fp5UCTm0q5IKzzmQo6Oh0GON816IHhfRq2tymKFY0SWIPhbf8NTJII2Nb0XR
14Gd3JsHEvjR7YGNR/24e0JDlGTzrnTw8sOfjODzm6IsReb33nqrqdYi1ZG1TKNH
ZR98vnPwd4lI0rTjcQJ4Ze04ak6juKq2RGsDj1mI3mF+nvrDWYBnKgeffhHNAGO6
ZL5z73twh2PO29zj95DbubDUtEGoQuG74k5LmnhsrEgUUnEzlrqqhwtr2xNJH+dm
1s2HQtQfC9IGAnNN0oFH9Veqt9QSva6QdIyhYwZ5aTlMWBo/86U802TLnM9U7sTS
tbquIWk73v0hDAYYpDvteo3y+69iExO0Fqgbnkhl0hrCO2t64GdQs/1RB5ml4MIg
mn9DjKfbh3nuDAxzQrIOrkwj5HI+ofQWh1UcrnpQv29215dxhSko67IDe74FdMzZ
XPRzI03yEPKwmF17W7qxxo37n+K+VxZmXD6u7TTDWNBlxRssamAKkQB3kPowVb4+
Qa/jLQfejIvhVtqJ16L6w1zLjBTRltzoMko9mMVDBe2O7EekHeWI3yfCryDCz6ac
wQN3ymt+PYEDdAuzDKrJNijTE5lM+x5Ud9+ESK7+4b1y8ya43zeIDEYaFosuXq6j
r9kD3guJdw1ZHIkjktvrzAGkDdVtG3T74Q9iiv4kjoukrfVtmTIVQSwWIG3XvU2K
pCNRNtCgCzLDx+APqgemqSsRZ1k/sYI+ODx0mh+BPyV5QkEiy0gCbNJQhvp7eEcw
cEieEkujiyzkGM1ZuF1tnIEB5xQUApLIeCAevHp5Z+g4XvozT4X2A0EXBcL8tYKb
J6O/QbbcaE7zSGBiP0KsgkPLeMnkYfDQHhRJjTaLN/ZL66h1m3jUaGXxgt5fwHo6
GOdQDtCwE7lQ7e51HpfnhFgWegXMtijCENyzXD/jw/gqVo1wMvYE/vdhwmJEvAk3
cjdAb09xZpfENU2JOLYYN3bpEN5PLTP47Rl32QH/2LSnslfcSCxZZ4L2v0Wieq7L
nlkV2hSk4cUtZ+KzZyUbHmUham0lpDB9vhYaNAWWPXpQUV94hwEb8Dgy4WqmxpQ9
Anr5S4I29TbxFNNxd7gnMqKm2nA3NDAcdcsHvCRJhua9FT8nY/majFjYyv37Tf91
e6AGxm9SIoBoGgPxJ7g0vmpVw0rJ1vOkkarUj+BRhY4SYAZhB75zbeoxDRwKyBVF
1I96xYGy/BaandcfvMqhUIF0kh0yTTGQFOJAYMMaYr0AYumZliudSNSIjOE6Aaoz
9q8XZ0gWFslfwRiTbKWEkqRAj2zy8XsSEzn8csGLFkiXWIJAG3cn8iGD/yTTTrld
2Zuljbjn8+TJOiYOrNOeTDZNcRhOm/P5K07WsktxpNrwikWyffozJllWtbUHfmJS
gg/0op1nJxBzauTizT26ruH6ekLbAZsDodeHbLFAqbBeuUK/jEP9aWYNo1n2gHic
omz5jZWpqpt0lw+XvxoAFYQFjPFKP4ueYNGk3qLE7A4j7bZ9wNdkDmemgVxj5mOw
iN7w2nPHE1cPqVHcbV+YOnew1i3ThlgooXmltPLfGcvOKAqfsX31izd3Xxur3r8g
Epb4X48uRLnOwjn6NcKOKRuSf7Id43/QRxlx225pUgv+kzYD3Htn26lyOzbGMZJn
VO7pKrZU4iutIe/n8kiymXqtwf0VT26GiCX/FdgwAW8Miyz3tXTz3AK7yGeX29Q8
3G1t2PzEKw7+2EcxzEgjUtuV3w+9pxWZ4X+MIJZQFD/UerCFNx66344TktnctpW1
giaqLFE4FY4hBc3l0ukfUu7lEtlx0ns8Z5aU5YYavYxWzima/Del2Oby4jGXhG23
Bp0xC6QVw05Beg/m38Nn4ndTEWXCNcLqJA6b9auKJMA2bdZGwEZhkEICvO+OK5Fs
oveaXgdB18kjup6fB2UnJ/m+IB6c7QswGkEjylGLSDYnZKscPixZOV2rpys3Ab8R
oy8ySobQAnuXRKo3NeuBcEhmt/H+03ulmb5Zneb6BYL+nFpeCrnYFLxKw0WDBDMz
g+nmqBnBecHEGhZQr1kdQgNlNbpmNNpNkZ3HdrXqKhPyDCOsfhoHbzOHq6w9fKLT
91ESwCF/bVmLRRk46spLg9LRW+VRQBhQ/X9A2ADvqvTr9OaxVvUo4gpnjBZ30i1C
DV5f3kAbOOtAoPqzeOT+8J+P2cnGNdcOXJXyckQQExsS9CA5qwxFG4jMh1gB+2bU
/60mqs3PFa7GlbM3yy+9L215IaahgpO6/wLEfvPMOPft7QWnYbRxsExCJLf1d43e
vHf9ihkgYnPKu9qYIAUidXL5LU86fJLGA768cVIquDUgDjChuI89TqlTN32a2a+l
3XXpRzDcjObIkx21XWIHmh57uup6yNWetW9gvAn6k4io6zavW0qwHTzQoIyd6V/v
B7c+blpmRdQLzHZ2LsPro6f2VVgSi+6VT2rjipiZ+mjGZWv6yxSXS78hhJgL4H1I
YVeOmoU0WL0eVxe7sLEpy6uPqjQ7/J1H0dB6OPQ8OERcqLgrHDxy7ZQF8i4Zk6Ay
QIYCvn9AmYsYmTSPzddwHzP2f/zj/2cY2wp1OafxQWodvcTvgoPly/YgDzuKskIp
8k6B7Zi1BtdVns/xjFa2AF3P1k05TZTwkvvJpL9WSrfoIjU5rgLi54df6vhAEGb+
h/r5mouoH2YOZtq/se+J5/3IfY2ZnTCI0xD8aKzyPWLZVUNvaZotYAqrm0y5IfpZ
EPv9AXiLpsaLhet/Jdf4LcC9uhlOjRrFhsMXGHO21d5zn6uISouCOy1WnwCgyP6J
NVGkWJmHygW9O28qdWBzCg0ozSfmHg8zXrwI2G0vdNwfY+W2IGc0If0RE+eunu0H
qyqoT78WHn6TOKbUIhvLWADkZc96wY1Nu719MHWSBra5xhLK8wYc7COf5pYMLzGO
F1oFH442rXJTqCIic0BccUWG33HKZ5bIk+C4VKIW3H/873uACD1ADOFRxCkhAvw0
4N3AU+2jk4RtQDzmwC9e8Oj7tNmMXwupilf+ZwKzRzp050/nmUPot+1F6fNwqJ+M
tmmZX6H4k8cIXJv621xhRq8fE9pC+MvnuVjUj/xul3TfZmJFXrCwrxM504OhprlN
BUyy6mWOm26YCkGe33PeiiWIsZpSNTo8HGgJBdasVEyQLl8ooVhe31/k+KLPRBGM
WMqKzpLwUclT46Apg+m/mCI4tD1fU9g/wUCl9PdJCH0Q3C/u93swoW07+vFFqNCp
Ja0ONmEP292jbneAnL4acydZe3nIuuHrnugjAO5f7t2VihaFr1mRKGKf6fepq16h
Sy57RMo/mLCeTETO93pJzevjqEEo0jSJelLmQd83UxMIzhtMd1qTfi2aweB0DXOy
D6P/gT+oN2y2bA92KWhf4W3ihAJhEad0UcZsXnifIe/55RKsZ0rE3GIiaBiWR6yR
CTccs1ogfBwFX5gZbiTUmMeNQf3ztY+3AVSLxl5XccFvb/z6jlgfPpgFxbhZ2mev
QquZuHdWQeSHMxyMBy+wFl+aPJbwGtbha7Etn+63Z8YV2hEgBD/DnlpCt/bFEHPQ
cBTs75ZBROCEO8NE3jDE4bRs9epX6w26iT7ZUL6y3U5xL725znwXpRNhow21ZnCq
FEJG78O11P8v/UHVnvqpRY11fk+/zmRlkhqY76TvwPIg4oAPYAb/S7sjnGWlctu6
BBXUP3YnnTgwuT8GqGSVqZ1HhM7Y8HcdSzgDaKh7rQfiVRPNiDNfVYVKYLRIAWG2
lUbufKsmdfmJOaMZPj9FeI1bXXyJyONPdPGkStz8zCMAWI1VP1gZrMEj5dG9C4gt
hXBt7X/AtaZmrRnV+rgBiduJBtP7EWUt1T6kBbg1RLHjrloDj6J1Z6a2vDMSAD39
Mg8AaHGQxHpCwU4Bw6QVMZmDl7BW9Ag7ApjT93bXdKk5rGgfSJd2/CSIasn4KWxs
YgLhlglWvMJKwg7gpfHlaABvDnKpOvpvTsrZk5uXLCIXbW0DcaWc0jn3EPxQ6BUl
6YGdpI6f3U6IDP5DkSPVW9E9mnK8VfPiPUO4oIqEDQpwYj6/OeSEpFTprh7fPtRS
pn6U6jxMjU/lNlYFN7yh7oAukcS0yA8hSmZf41UFSCn0aNA8GZkVQiOqe4J5pF8Y
H3XctGlVz3rmGLRwOeo3pyz2PxEXgRpC1LgobZH3MEUle/wChfOzWqO3NGaDFYJO
Nj4AzddMlIuNyCxZl2pm+LfBzSI8VCfdmWECR549y990wkaTaXJvq5uYF2rMA/n2
kmRF244it2Mj1RhSIrm/OZIKgGkBD7EbeM0H7it82kLFAl7J3NFRb52etzY/o7pG
NcLUw4Wz+m+Ax1MNf4bN0/9aQAf+IlIf9yoabcyYLmgWA/lq73fFC8dzh28fbPJW
UXHcZQkLmOYuQ/a5r+wfRrJoL2sK3KJEdEnXE3GKypS2upx7XS4NhkubjrzfGjO5
d13bRTX7L5Cownvbb9VpctD0utyW5Y6JddJNEOgbIE+nijpy9fuGaaAAMS8WKJdR
TQsCiB50SkpimsmvF8ORH7jD0dCzyPHFjKrbQdbGuYnmAlkAZbFJOa0CUNVTRCtE
E999l010oIX6N/OTjtcqrBgOlJyCQmZ6bfRlARjcfaswYu9FDwgQCAR8v+rMVDkZ
uqAkJyiAoYeWXEV9kBKtSzY8VNZSFOQKt2HCvhceicOarkjZsZx+ArvM7rAaETEr
azDjGF0PQ/c9sm+XSSudEvHSxCUG7fNvuch/CnfiSeCXnuFP79NJAf8iOtzl9AnU
iuxDC3XzxSgv4tbx1eBireiArZC9OMeOOcaxPBb0a0EtM8xMM+s6Nk9o+NoToBBN
kEZweqMkLBkWDye1bmt0gp4LnDGAn8BXjej2L9mx7vaXFCBp8bo2hPrmOhLRPQn3
5ATJRcJkW0GMNGxuQlfdDlF8xZWoUv6ModyxhhvuzusnVVrxIDKuJ13vEkjySlbU
4AacCHLY8IxDlpv0t4NNHqJxEdQ7xrbw6M12p3AAEWyeFErvKEwY1sJTWYHduDC/
smZA8wnuMfUvw5I+6N18nhNMKhdwSlH0QtfW3YjQtkTxdA4e3oDPUq8Gc534tCwu
tP5ZSlPJYRXs0f7URd5F2h/BB3KyaALz4NcnwWVlWphJm2wUMYjOqpfg0OODV4gX
VaKglBbOfo5xnwXMs33ae3lxCLNg+B4yYV4WznZEogYzpUNmuMYNkfEj7rB0l0g2
tZOXJmyJjTKgD51RLO2Jmeh/dSaiWlY7I9RcWz4TdU8ixk7L0cuL4pjpCp+hoSN5
/v7M+vgd80rXjAQvs4UEGnuNSDUb79rIr5ZfRKe2ZYNem5ckGVPYlLG/K3aKN3dO
96WW/lS4rr1Ic9KtQkUiFj9bsHiCWduJO8jqwEkxPt3/ZZ7lsUp+MDZq2gdrX7Jr
3PSlNaQNo4L6wp0FYtHP6zFfb5QoQLi/BGOFZw4ZN3gmJQEMOc5zx1TDsYTzgv9F
ba7R2+g/25bP2t2Be93SR3nAiEJbScAW/KcFJL8HDu9nWBW72wWwP2Nph1oZ/R/Y
nvk/elkYa5eqKTGAfJvkpkbwbChwaq00KXj11U5keNBPXkZgHQDXaQks/XahBxpe
Po9SFcpCBNaWfEEx1QIjPv/tJxeanPXBB5hY1c3SS5of1xwLzgVWJ5YtU5CGkZLv
bAkDPbjVtXV2FUCR7aUkTMTWl0kLQcNICFUWZptFjE8bOh1rTp1qeAy6CaJpPGGw
v64LlkrvP0EBcA0QB9yZv2twd/vYX7h68cWKeUOyRka6tf0KURTcCFGv76eOylkW
oTAiihlZ+dsOxHWGlpPjwwqT/63IAkO7ksizQhTOUJSDyoKJZ0xQCI4EEbDLFo+O
30h0FaAJSlfKEofODoX/I16sDoKy8doZq93Tasz8UylsJHiEYCO9fRBvWsuXqhnb
qtQHUu1hZr4TSyi7Bf5GaB0hXS/YPi8M8QG1QDAmyu7X05sKmAUaSnMmsc7fD+u8
VKUAr9UdoYz8LVf5Kb/XZM7mWq109oC8kvJdjMcIdDHlUXds5OZMnonNWjR/l1qn
gxc6P/XrZPQ9lGbfgdngyt2JCt216rhj/zF7TnEW28Ev9NYsCH9qGwrP/aZXkXBT
kmzRf9H+8COL/KGzGUlCVN6HSLS+b8MqUh1iOnTS75SuD+XLDXtn28BUv33XdfY7
tollGbdIdHS3acv6BzdOE1GCCftEUUaqx4c1rajO2Bii6Rz7oVsqJuQwlK7epZMF
by2ezNpRjMbPw7bu3SrPmlAvCt/KAXv7C5un4EYYpToOJGG8xKe/ylxndO2umM8B
vhxgaPE6ujh472ld0omVS/wr/OoRUT7IgJCKFR7g1jEBrwdGtoVG+q4HUsW+xu1n
ENn3LXbos23WNvaAe9dkEIPMUZvcCcEjvCfOlj/1bG62jjPWLa6ULk7qF9IUgI5M
EzYTYFfK9RhRUq+2bqFlBtEprTC/W4eRFpBy5WdDbyB7908+708kVSqAlTlmhz5S
1CYqcPT+OzJqV21vNaUFJ4g2n9qyOnfKyPXn2GepxnQDjvCGLwAjfQHFUuciv9aH
U0uU/tahzl9V3W0Tkd08AJsPWF8WtMKBZEN/5Qs2lPdOwIcmRZyMnc2qA7aOxwQH
PMQeunH4K3JohBzKu0dKnMdB1bq0UcMw9+MV/vGlWVzBEQPzhfpMIC3wVtYgfIQt
6lH1akqnnnBtKkkSLILB6B3fCsD9Ux+ENX0nXNkXR2dgJzyftvo6XJsRJP7Id7Wa
ugqsRrgKGP3L6ttzVnBuf5qUihRZM6W8LK9z2wesmdDZFN7o7b5Tz6dAehnigX0W
pe3iFusTc9cZ4qiBeTH6NeG/wNq2jHfIIl3XdT+I9zebmLecNuC1RuOcX0ZIk/DZ
BHxBkLCf6+INul/b/yHy92edF7qBtglfIh45M8raF0qKc4JZpTyr7IGEIayYX+Kx
RTrefH7rKS0kiUc3eTnqBeY3c8b42dVN7bytkgs+u2lID6rzP8IOnMJbDdf8+SRQ
R8lB3G/rphmGxiSn8cYcEDhi63lMowPOhI2LZiQKJCgv3DAavEOQJGY1avanCbGA
pekRBhtBwLkLEc7tPn7msACtMEfVbgve/amX7e+dAD4D6/3crqce/dSdJoPRv+fa
K+8nExVsm9/ELBgqUgh3bPJjGDHiEHigPFRakS351hFn5TINUlpDUkATekLbhYGj
F1Skxf0lR39L5DjUBLMEAfg4LHUarPiCb0YdbxDuvr4FDgkY9KTaeflJs//pjgpF
BSDFXUo/T6Z9HzU+XEef7cWMx6ITMvZ8eQ0KGRrRjiV/ooDbvZlQ2IlmlikiHT+k
AUdC/hMqfYtyE0SK0QvhJ0ifNzJjK5j/mUkgC8Luf7du0AonNRf9A1arm5dDx3T9
Zte7GuZZpGAlhicBqQ+7cfgRKlAEyaHdwJvN7OZtF1/rrc9Tqp80hIY9MWEeKlG8
1lfeLlKFg1c98s7VJr4kGDcZDjWGRiklvG/xbL1XRJEdsHLskYewFJP0cGPhZQkX
ESY/Z9iSop3I6e8HEXvBmw4OYehNsRg+9Vu4OJrJFW7Spb0f2BAEe+jOe1qaLdsY
9i6ef+X1KEC/MjyZkX3Y/mrsBfWVyFS5xWeTb0jjLI51YqXTkVMGvLp6Rlyc4ajR
1t3MfWK54rf0vAvQLZ/7AxnQ4v/F+kb5Us8mxYEeg8K76CUPmnDeqv9uT+lCNWwU
PcnQzS/IvBOIuTML2BLraYNsyzK/gPQHv3N254jf2W/FIgDO6HD7QIGNqFZLNJOx
GiIiV4TP9cfKDl8Mm4Hlm0i1NvQpyUM3e427l772VVxjBn4zTDaYS/+dTLc3/0zs
T2bPxj6m3q9k4iK7aQdi19ljXbJdXdTcZeHBwnsYG25f5E80zZ8eDzPHAmj4dFAq
3QLOb8X744W/vrHuKmT2+t8K9BXpWxmUi1eTPnv1RWYPL4bdlioQ3lQHsihOQXgS
QOGLXshe0K3WRGETRdDpW0Aq8c8ZJu53ZOMBSRhFmC5qSb1LhxWdlsCCheKtrjFK
sA8ZlvltLRVikBHSRzIyzuQeDH+8pR44Os+gt41xB3gjfjP+gvGA6ee/fH0ZQoQR
a3Ztbd9Js8yDmyuKRUxBJcDBoK/XRoRULp501sppND1Aa+Jw1709rEurClw+YIuB
et5EbEPKIRTdeVU1XexZiAHTOJRLuHD0DEWUa44lCq15zpGaomNdeflYxfYnXldp
n5JAKLTBhNAAKS8uwzbI2CDUV/pk5mJZA/keVpFq0VM0ZnPa2cvkeEdLZUAtPHiF
189pnHJ+c4k0lcMexRYX/mOSAULaMb2BqpzIEnuNMC5tbr0/Xof84Znm8x+fFENf
vNQSZBab2EbzhzS00KFtugkgg70kUPtxi+aFlGW4hA2+i+zUm+rVKHt4lfqAVmpo
8TCJrh6znmzcPOnqh8anFRqsC7b60pab26A7EESMVTo4Ed+FRBtHtVyfNzCNXP3Q
YQO5wZX/nWbA1coO5HEAXNI40TW6WXQ0AZjJWgsAeL7CVXL2BXCPdXo7UkglpaYE
5O3OeQVeSP//BXuIpHkxteiIzoV0AcLwnbPEtplyE0iU58mAQEVD3bpyTPV0bQm0
W/Gvr3sTeAw52Qa4i4/EWzrs66c9ncimJyClfwxY3D91CXzp7lvi7aqgJXJTHphk
qvibPaAOr2F24bTaybCzDSLp6QenUbjJWH+qFlFyIgJuSVPb0xyEOf9LAkAv9plR
mci2MFraqIP+UvO3mh0pFkGo4ExZecwVkOLFDyeFNHLWsZHD4BsvM6oqH4v+7CHE
sYk2tGWNQDTqEfP5o3Zpqw7rxIR4hRivqILQhgLi99W0FEkmI5gHcyhTxe+wv/qJ
H4BwEbDjDVu8usU9gjzE5RYOENbB5CC6xURR/cYY4sv64FZ7OSYm1lm2rdL0nOnm
ptzKg7ll4ct+GlZCti/kaIAjExaUZsDpzGcs6e16/Z5FEFp52iO7zpZ3/lBl87GA
fuJyOHBSbkw5gSnxH+YUMgkn0NdP3umGcogwRWYuE4hMBrqNWHcB3CktrEZKi8Ek
hwptLXmvE6iRht1EToPwoxJrAJh/ZmzeGjTyvoILIzXqR/M0M8KKBkWuFbkiZUUe
6QzpRjvdNBZONDh7TIGXc7m85DUuQg/X9l6LbVBnQPI+2VeyNJUg5gaDEbn8b5Lf
0zAHshp3TBpQSeg3nGZoVe7BHTWsAo43D66X0leGNFNc22mvBqJpLfjaU50nszzk
wJhgTDRCR7NUvDkps9RQvlywIDTALa4jhGOOG/qJAr07qzG3oRHYX6E7QPWt3OSv
5M1gRIdhyhiijluILNfQDkpcE3X1KSfKkL4V0URFmqBtowGsevL3wVJOF6uH2HZk
cpl6oYLXxU0M3LepuV+PqPluG+IMPwnrq/eBbGaTbsbKWsm8Pf8E7ZxKEfeAw3ss
DlohzAojZFbSHL2NZhTkEjzdHE3niusmbsg3IGkEOlgw6xxUjJP9NRqiqCvfR/4S
oVpaOEglMiF45V90OxNjr5/MAFc5IqNZcjSQpEsPZEcHQH0oEx1QtrA4pTCKVbeD
0VSQoXk/9+8Iw8Ua5k4s0j9kE0A+jrI3tGCDfKcBAE4UHaqVnNcfibj7XefWZpz7
6CK4p+0Kw9a0hkMFngBjlCPTTmmlYKRCyixlrGOQjfqMqzPEl0uWFZ+2NpPfVj/C
yRRZIUHSa67dvWPOvq4SGKJogUAHcEn32zenm58JvoFBC8qUrdGthRbt6LRKifVb
Pk5QTsG4BpmMXcLLt4fXNxTc/WSRlO6H9rD20agPRUQoIA/E/8R4cDKFiJzilPxX
tWmj79pC7GDLPWSSM466AQ6JaphcuGKkxmd7AIb+FfT174Roi111FZWMe7T68jcL
7kGZgiKOqyCQFI24GKAYncDOr1Y1LA6rTOViLTbz6MPK5VJOUIIgKlAK8wPIU53S
rkTssCdHAZoIj+znngFWow2mIIj4aP+aRgiI8sKIRFdyUZfofK+5X7raSkkYs3fD
7yJzRZoAeUrhUGedKfk1jtjGn3xnYXmO83M5vHvAku8bQ5JDJG/xKhr6ZNR0DqmX
ub/ZwBBXemzpGMNbkZuZIozFI6BzklJ6E5JkSfD6vNVYa+YFDuCqEzVik2wd//qd
zO8qxDOLl73BbfPMjRquTpoDKIwFuFU0e7oCg+cApqhXg/Zn6uBUZf6U8jM25kKw
n1KI642bZu84ReUxe3leUf1rlt4OzO+80DLCaE+C3KA/1timOdEyvpX71rpL1e8L
4umQjlY1P6oB+nGM1LgWV0aQL96ibqm5R392IkP+QvVZ4SgWVsUM1QUSez+KMc+r
NSQ1BDVWBPYsVFz8fsJhEloKTYaH1DggNDpbYPGPGhEWyboBmNW+7DMSAawYPRUP
iJKrfY4pznfVmjKSHaY+s+9d68eDJCwQgPop7m1t05WlSjbMoUEIeQb2M8c6V/jl
jzh8Ii7XIiuC6VppCb1OnmghNsnTbyPxCyNxGVqr9ZXG+iUHFpFm3ZgoNk5Ip0iV
e17RLjhHL1bdg697oA8f1aTivlNbR0jDSt3GaP63LgXejsToqkO9ki35d3ru2iVC
mvTBjLccvSW/X0J8gIFOpPHt6N6xb6Qo8bNuGrZHUO6zq0CDMkG2R9ADWui3JxwR
pH5K9RBXLDqf771bxcLc4swhF4Sy73/ysqZbdpP2ogI0JkEIjvDEP2Xd0sAF7BbU
p5/Z0ek8qUpVDQ5rI4di2e+hBbrjBVLA+jQv/+poAqAVwoI2drUlHPPT8CCkM0sg
RX097IPEf031xEpqsW4vHOmH3UW8NAcTCPImltlgvZm55jV+funOph9o/W6WxiUT
LW9JfNv69YnE7up4Mi7KpFVupYWPrloI17WktCn7FdJ92egQHHyV2KWla1LMu7QK
qLqegP4HQLq8WjgL6c6HZTXB7npWIcN67b52UCp4Dv/cZuG60AdLgyowhcf6Akwk
geGU+7WO5GncpcrAv1EgRp62g/eDkSIo9nf+g1PpFDDg7pGkTInQshTR3dxz6VEP
C7svmr6b+16Hsd/TvYrbx7VkpAobvPw6zGlsbfHmDBAlsoN3PEQSk91bKTvPlerX
lbE9gX3SVl2QNk3tFbkgrNvRoLH5Z/zIZhxc3ES44Joctb+sctjKvg4/Zaxpl0hT
zyJ9MsKKcU5MpgK0hiRPdnDaugI9oWRMSQQ0nWsrAj0y0ZVz7Jf7dZaII4QWuYHo
NDuab7peNwHSBWOarIPo3wLS7xG24e3Z9dneTDKbqeTTP/AhcIhuSYbEG/I6fSw4
9nKk0mL78mIbgYbeXnzcwhhowRKa3fh0ZeqMl38mrtLQeq2wmiT0PUmWYfuB3jND
oGZQ5tU8tJD4JtuS9FgP7GDElza7BpVIWMOLnWmagKokFIXHku9XeQWspLL2bIFC
58qmYFtdYHl+kS0Q3GWMcBnArJ7OrDoNXeDeLppYZJe19JCX1uU4TEM+1thjZYk6
CaPJxVqa0379cUy50yfna5i/LVOOi1Lq/d5nn7psdPvkw3AFTFVPDtYSGYVEbNG/
7WPTUiSOxiqd46+QD8PZjJEehfTtr3r+BFAC1thKQQmxPdrAJn124DJ433URpsG0
oazU6Z2M30RNaBtPodh3g5d6EZduaFYQZWzBiTByHAxml65LXQsA8LIxpjmkblnb
ouajKdcbaSFqxq7gH5NvNvx390Pu1PgRJWLi0oNp2uZ3P1iEAf+l2qXBkFe1Rb4C
nv1KximmCpVWaKDLcPhnCdK40LOtQ1x8PdkJKMe/3iKj4sqUSMZv8JNEzAJODIA4
C+UxCC33KTObs2NsUA74mjhFnWj8eaJHUjXOQAsUmr6rXcQyv1FZLmGbxF0EbtRM
7RJizZQq4MUpu1ZpncvJ0c6KlkPB8aU8unw+4VmS6JiGGm5RxUIssPCVjZks994g
KpI2aURb8TFehiJXZbQ98O4cNbfPtvfGFbp9ZwRqex3lC2Z90qhxVTUQRLP2bQ1f
b+2KSY5LhKt1wyMarfFe5PG85XaCYMkH8XrGNlKbOnxpMthSu3qEkY3pvkOt7+i9
wooJa22SFDV6JhzWkBU20x9uPTD/xNWrlKkr1dz8B7+NamV1foZkm+k74HwkIIhW
q2vxLTqsK/mTtO/tYQmk5nm45vkRl6uG7ICDgcay4sLaeIGAksJZvi3rWJHcxPBg
iDLEHF5eYG8/hhvpQKbaWiyI93o28L+kHNbXW7ESnp8Ik8CT3ovoc+L5kKZouLYG
Np7PVknCz5nZGD/Ulewmavlplky2sNObspi6NIatphJ8a+mhRB/tzWiIL4egLAGf
HU+3t78+K95Jt25RXjRVPDgPvH/HvHzrBoxj6lR4mS6g5Z94lMvyPfIBrRPO+Ejq
9LwqHp/MthNIUlwtLWEKO0xcMT8wMSGqsuMp2XRJKB0drXJIc3Xx/w61MP+u9w0Q
Ye6cJB2f8m2fwXxBl/c/f+1ZsNUjknTFba13vi+lmi1iFoQ0hS7nRRWvn8B7yRQg
N8oK4U6J6ILRhLcRzikKD/z0HNi0hK+4S7kKvCh+0lWkYoHVs1QqJcF8/mIscml3
7EgY57OZKFWg50ASERfCgzh2g/2ceCLlG0m6olr7LAhO+jpb8azId9fmYC53Ktqh
8R4jGH5O8nDXUlSBCI4RBpkEX2rvFiSSu9e3LLyF8Ng+vnBiu90lSelqFjxWa3ap
jvbKpmMZkRdqeftEKSVhBc6SZyNZmIuiSShbzbompKm1VD34wrtM3aYXZhA1tvCb
ebOVi7qA0mzBBvbKI+F5r3zN1Ifr8idy1XHRvEVtnsENtVqjSF3KCB56AUvjvUxJ
4DlYZBATsMXpwkyggD1Kc7VoCAEweoTikRyBFRXjihOBqiVJ3FUhNvIui5lAvaFW
72MkTCgx97jlsKVJMXHmLdIey/zps+yOIjVK72tsHQPmshJa43wOJINpC5O/Mmoi
Ihiv/PiT8wym03q4O0qEmc29yrMr/+TABsbIyRIPZ6ueobtqnapcTwiijSs/Wpqw
JncwYhC/+ynMvQRNnffloF5Wgb1aZHPzlxCfriego8Cq6I4ii270hFLYBltJJ71S
8rtfDGHOhj+WEcZr7Id572VJxII/E5/AL9AIzNowRHnaOhEqE4Q81Au87AaokQPK
3/m1Uoj/i0zXymW2/ecwhC5NyqUMPUZL9027/RGZVkFZSM2d5ljn6Ejav0QdNYSB
fWJVRUCeprlhKzdrgp1TreAU1sEPCuQnubMGEtTIIwVlP+6COfQiuZEFPI0nYvOi
n4rl0dDsYTdT/htXs1Y4tWNGaqzDuS1S44TolHvjMS44twiE6m8oWv4A02HvfQnM
ST/HReWHIFyxKu+3Rlx0e9I9ibiWDfkWZoefCemFsYbbIi8co1QU4ANzFcaxiPA6
JAoTfr4eFeNJzTNO6kuWmzyrmp57uEBbFfa/PDHBqqsV6H1zYJn9uOMG6d6yftwx
+LU/BTWSa7TACzmUpAydiGuP10c8yJlrK+vBhBNFvR9wz55R3CTrZ99fq8XatC4b
dFIoN0kmOt7ph+DLX3bu85lPvPt0TOXApNi4X7jL3EzQp3ypjd5SethV3GXQ+g4a
1vXX7IcHg4x3naSDjw+ncnaoQagLCNyPDyn+KYonrTChJCgcqJ3mf2bi4tHKgCVi
oGwM0GqlZJ5/syWQnOkbaEIEVZ2VAWHJM5A13FxeaDFZRiaGP3bKtUYSaNIH/zie
S6/oV5eEF/iiG4XAFFQFaqQVwQF1vdHnSi//ckfLUF+IXF30W+ZAyUB7AH4xK809
S3kS1uC4xYBizoFcO2jJfZUL9cUMEvxD05IhGq+GfqiU5BoB62M4YCvVxMTgKMx3
STnbNS1jmzYQT61wIiFe2MRY6+nR92qSQuC3glBlkoG1dqXxOWuNIzO0G4y8Mu81
lfZ/NxsMfIgk/djn7UC+mUBjyVKU1JU5OERuLxhbWVoFPnRIIBbGqlu2SFcbQgnC
UFljgiGR9aFXIzE6T3ZrnHuJrY4dJZMlG5KfwTZIoSNAVWytr4i9oKDTBQt4/R3y
SlCSx/xhtCWlxmJY7OuliDwk6mC3zk/tQ856vZS+xvCXscGAnJdQlIlo0AWS5Suo
a0rt1ZGk51cqGt+q3RFEVHT9+4oZQOVi5wf1iKB0mxVxxZ4sHVSqAI13u0NySTK7
NBPSnv/tN8pAPn+Z1uSrfretO8avxvJTzY8FfWzIEhscYG4Cx7ffbuR6051SgVnE
K/V7dZIABrdu2dzmdqgQHSC5vp/D/fOJsloz13He5QBGlQC2PkyfgZP5sZVmT/bK
kLPaWJVzGCOIlyKZmrz/tFIWw2SX0H8ntfO0YvD92S8juX90pK21CsSn01NFSHR4
C5g0xVaXJJekGqKdNNsZ64M5NdLGBDnua5t0d1/pUVZuF3XeiUp9mkT6eHwQX1qE
bLNMoGT6sCBcW6drJP5IHqvxXrb2GYTnl+h8SyscwXENtcV9bDl7XRYuwcdkGrbs
eAq8kAgjUZDQE2sCYElpBscFiUEX8vjl54XlOstOBk7HmoqB7TWhZ3JikWvlvYpR
z6T1rgrlSRHkvMZbdTScaMLW4eQqgmngULmMxS6stAkJwhI/hMSWYe6D+ZInp9hS
wHq+aOGh5iv5qH9WAYkT54B/u8lnIPM199F32I5IvTgU2q0UQBxOhZxGd8nFdneC
ptFOT2nIoA/hzsN65GSkAgnNNPq2AX/zTDypbfeuiraCeAdk51lv6BfYaGSpmEcN
BE2GtyDLH6g7RcWoV3WN+XcP27IbIgOLdHfGoUXD0Qjii2R8KRdRrfKmbHY6y8wb
LNMgGhEtWel3+8kADtdeZfz/z3XM4XB136H74mSMzGRMNLkS4C0GbZreYefpgjg8
SaJi8jN/mnT8drMzzsJIUWjyDWmjKK5IyhvGerM/DHbwSNo/XuG94nuDFJ500RZ+
r5udDXyf9J0uz9oJh49ywyoDghDQCbv15huwI3iuhlyLM01Q6+eFINo354E5Aaay
DNh5thda1lWBJXcC2Qhs6IH1GxMzGpYQTBtdQQOF3OFmuWqaoweRpZuTbKWo/A0Z
GWW38ylR+3qY1c9jW/LdLJ2krLnQPH7wX0f9a+USpaTpPxHMH9ZsEwbZJi9wJPBR
BbHtj5ssoSatNU1A2GrIQxz0NWOL49+h5b77oQ6FcXe74+kIZ39YJt9mAacmm/p2
8tVPsI1F1xoHrYImq9o8QfK1xqxeG7PF1wsOuAxDDUBVm7LdItthCpIVjj8UdC2V
HXTWOw2oeARCOSxMFu05KAuIiItQgoEEvyFWEK71cijLp6LWaQRzSj+vkrFg6YOt
3fWiR+NF2JH3YYmLPiiX9gjQHlzMHGpZA7ah0XMxBDkJNHCvaQXDJJoJLX47gzv+
MiHoZdPTQ8ZQ4MA243O6J3GZWQ37sLggRQMANKDJkgb8ndCTem+uSHhKN+3xTyhZ
S2DFtDnV6EW2kmMGGnWPsh5QU8a+IBKrh3+TeFsvGJc7qrri1RJDXW129Rj2cCAG
trS3wSYaO6JrHCxQ0LdGlZZ6XVU2m6dTXb7tlcSTAENtBlpuMBVrIQRJ69qkmcyc
F7hMnFFIYgURa8+v04fhIo0WxwGvbPAoNZjsbSsz6oRV0WlutykW4IPU4qP/OlNP
iOKTkivCrImgAYZWSOGLrxtBhK3LIWu5JtLsGPOMc/n0+J/7fQ+zrhvMPLxWrTcq
8bArGrINWfVE2DpAmogMYj12KUYqJHLS2BC7wbwfDcsK/NyaRGks7Dxn+1k9y2G7
GI2t/4QYF35zGazUlfceEPXoJ9DlsZJyAVnC2/khL2cvqm7/11DHn2qmiKZwwhiP
aSUd5Fw6AGewsT/l/chWglfuRu132TNvHZndLZyx0kQpmf4h25iMF1kBlT8dYj1s
w7/ESn8wnvgNNoQtfKv5wLhRPa8tRi4a7by5Hhfuarqam6xH4alKsl/OL7ECcymL
EW6kIWCOpsUdURB5xb4VuDEDfE8kTmTmzUdifgRs9u+xMW92icwR6s1KMWiR95Wu
Y+7IVjQrx3Wr5lUyRu7+/hFmkbdptIAmjNZJ/IzsXgh+4Q1XqadxY+U31dY9ZoBC
J0ujVJrqCQjXgr5wwbKpylD8DdiYhYGnPM2Kj+2RAbXjuYTQmx2gciCE9WXFdWJo
vbBtFJheJu0o9DkxnkW7LBd8rdT/2Zfhuwb1YifPOmQ63b0D13ZruhnwNp0tQV1R
BfN6qpbNF4NjoiOZNVQjRoec2N3W9sBD0TEgqAPqqGpBkT8CbqLXHMvW1Ss/FrW0
1TdjnVE9xhukVqRNM2W2nNP8cZdI2rGtqiQHq3glmFWFHxFHmMkRWox7POLd5VYM
20NeLp8Vqr5qHXWM2HqVGYemA3qmtDd+YHt+nL7nyD8/QXduiSNGFWEzdjs/1445
rFN0ux+SXpCYFUdPDXjbKFZrETfBVL1Tm/qyyiVYhfLAlsL8pfNU/RjyPKS8+vX/
PMkPQxs080xgNsT7dTnQ+EV2dJZSzYxZxE7iSis5TZ726Uv8dA4gPyV92+80n9Vw
zpAxB3vs3JjkFAju2ozeOExe05p0gNPUJ8/XQizMreofZYjxZs4aowfE3H1kjqWU
GVCXAEhncaNLwTy59T2DTloUeRXQebu2jRFSnfQX7NVmpJQvaxMdaU2W/22jxWn9
19EtQG0Cn7wt6UkqOi7b1QhIQY+ExT8wXlPkiD3nkhw7gZbM6+jr7ltoLwRM7dAw
ZNGEiy3mG5lqRvlKjUVvq8GaVNs86bs7Z2RhBjjGpZOKjUVqAtSF+bjZpCL21q0t
qBvmlEO2esuI7jj5EhHTddqpo2IrsxpH/1BEoHy7qfOfZk7BocBVlBd4Qp23s8ea
pSkW28s11UMotXRqawMrdfPP+lN5EpFTAY1rt9CvViWja1Bat5GZFJmqv5vQtG9w
N4gdMnRpixk6vUWl8J0LNr0ZfFukNWSuDhdLGk8wrJT++WyfTOvlPRxu8+HJ1yA5
vGwLGn4Vhx65RDg7CjOckAfCptoUntSGcRqy7cECrrYi05Mh4iuHKIr6OtUjgTNg
C4pFfp5dC6RKpHYNV4FtrRFIv6nrsk8IR04CmWa4pUmfUBrUIX6jHHON0VIvhxUf
f/ebNjqLR7zjMgGtF7yD3mZAdAgSCmQe5HkFdgIxLANTHOzn7zcVBy0a5j4giIvO
LBSZQ1nk6xFHpfxM5ztKpOcFxbKeoeZUJJccFJSRzdJ2yW66mma6Cy1GroNKmg+q
zMUf3AOrk/X3LMkVbIBoZp8VayxE0vN/A1H7trEtyeRrDgwGktStfGWd1RiduiIu
0t8TDkzn1C3I0oNfDE05Ss2C9poHofXOp6XGKJP6Vi12ne14HkcLC4UeGSCrxQS4
HtLT6wPQGYbY35Z+af+HF8xR7pRa1j4pr9yQ0ILPMhgfLP6bpQfITJvGKr8YbLzw
xUpqXk2KJBnYiBWk/t3luZZpKUnh+nLyeYkcBljELnYtLxTKQf18SdZsMtWxgB9c
XVnWTLjXJM8CtQqDcxKTytB6tWCkJj85Fps6lHkRzhaHLLKJ59GeBwBZbyN8pciA
ClG3x4PWdOShi8A+gUSoOs8bCp9+zFhFOD6z0JvNVib3eglzYJIwtoTYpBKlD7RS
ODatWqj6QQPK7CuddRaKCHeC2f9tKf61CTWLk7LQj8PkfuQ1k+JjpFA1FxJi2rk3
qNu9n0ybRZmc3IznNlq2YMaE72VuGtXll3iaIsMEXd1kzeAZf/F1RNm85vth41af
78p3wgddEtqgWXRhMAxrQuLrzTPYe7ile8ADuusuE2OJPi4i6p+E0GJ171dtaieF
qtvVuUGjNuDKOfwPS2L5vyWGMETswC9dyrkv3VAgKitSHm/aABzch6K4poWT1SiF
Sx6mH+c4IACqh4Vvg3rYRO30Phmi4T2xTsEbzlafh4QM7Wg38ENSmPXYUKvtJ0Bz
7PlLomWb8ZtTm9Fwq+EmYYq8Q3dbTa9wAlIN982cEbUuvSq3kPMjIwbjcZ/PihcR
n6eV4OXplLCEavT0EwOcD1KmzvD/2dR0j78FD6USHjhWPsgUoAnLWu4Lf1A8CMk7
KHi0Eh9T4udrdVUuoG7k0cZmxVqWtc2PeJ5h4KW213/tQmNXS5INTFTWEr4/xIUz
WpeJhQEyZUc2Hgnhx1NScxMQ4utFHYB98NnSiYpEr85qDKf90i8dXeWZ7Byvpz5s
kN7AJQldHIrs342KOHZN44R3BKhl9ewKfKxLZR0+RpXMamvQPmtdKGV4flrTEL+C
WuRFYAFRhIkV8aaXXRqI3b8ls/aoBBcFu7Vg6okOvFaC9ULyCooy6NQrs9szwZPv
b6MES8CZ1OVd4o6ta2gXgjuYDVrE6FSx4vLzUKnByowQrwAFTzbC38DI3GG3+YOR
x/cTBMq5Zm5OvnFSIrNQck5Ivz1KOCLoGBxpm+8pyXh1iG/ED1knBX1lwOsrrZJl
Il7gPvrvv+4591SQNbYfcqDfDyZgmO0uTc7TaoGbTJEBJvI9Z6aZKotaqWwswCLI
al25u/FWHo+aAsZWSFeVeEED5sHoxVwozp5B9hRge9YYfoGzflqFdZTHi5gGD4sj
KiIiSf6Mh08VjC1LwpdVpLNTMaoNEip37MowjIViwVVm2IEeptdUOpvYrRuXsa/k
RP4rQFRFKsCZNXgSMWO4lWL/4B/bHHoxLX0/ztJbpBJ14d+pNs3AL3hpW/einGhA
X/GnE9bqJpBQaAkL0RN3MHkbLahH0bWCALEZ7jBEBrE/MIYWzjuca61Y6Bnp6XrD
JaTWxFcAT4st0J9GgLQUpmDu0gsySK+iFMJTXlwp4NjZu++lzxuM4a/qz2LF7vrp
eZwDXiNPycrQ22eNJ06Yu5l+jYF8/SLFRlBWLXFlEGryLXPu7sY0T64qpCp4NxkY
hIcV1YwvcJmeLQH+HfBYpjvXH0qZ10a+/vy1PFy1V41QXDkWejscxUKA6yvL5CEl
L19Y/4LQtaRkvrJg4C1zc/tgnFc3SlyFAW5sTcVSafl6lSudF4VQwNRd1PJe9KId
SlJQm7BKA1Sf4iCzloMM71LfVupEKFUvGFX8Kx+4T8+wG3pxOIGHv+D7EyFkas1a
1Tcw0a6oTk0gnQPR/wfnY9rFGN29uQjsqAKNeqBivJnpKrhf0MKK6SN3yPoUI9iG
3Q3L9K/DTrMK7CBWSNodECpc5GOqDDp5wOXGZ8cqdiva5n3S/PDFYA+2GvYjnBal
IvzpJ/04ZdXE/Rsw7QOfyWQofVAZVCF9whMJj+XfmoPGk0/a43Qnd6dxqp5qqEav
J/Z+Q5VnsNIgDFJ4+BkO1nk881x+z4298eys1McAUsNxlhy4J7qZZQGoookZQtvI
wZ+dr+COJ4kn4hyTQyA1txNYMVAs3xcNh6aPfjgFGw46bzpi8AYzwODM5Imumi8M
OyDGCIdskB/erjM/bNXpFUj+cE6g5CGrNOBM1A68aLhPMsW/v+8RER5pQ7nLQMdH
ALpdJotqhMApv6jDm6YhINPIe6dkOoxCp32Xj4vnP6NeODLiPRGEI1pPqVWmAbvS
8KeWg/7ZPAW2fJgkd32CASanc9+bubhEwBHeYQzCUgM23gnxsbZX3ssyDfI7NcO8
1wpXLA4+dgwcsEotCJLBbjbDokEHEkxabKXLHLiNa2cccwCWpqWjcx8cFmDs+End
Wy/vSL+Bh6bxEC5bEEBEcpj2n5DpL0me4jPapTpIGjK/TjFyEbmB3FTetJz1wIsd
HARwPUg1Lo/lnANlq94GhlLGjh//hhJQ6/lxGCB7RVuqDrPksIsgMrHEylS7t/cV
HYiT0zH40HgYZ61ZnlsSbkhjWuKYMzR7lGW4hNnOysLnRlyZ6794RPNrfaNGZfK4
yEp5yZ4AE1/b9OWRYedvyfRllmkmerJkSr43tRNwS/ypgrOdFpveUc41Rg85MyN4
M5DYQKGBKd6yV7GkFZ5C0n3wAy7sqOD120kPb86ZbVndtK9h8xJhNa3vWJAK93kO
PXjhKySZ5Rf2LKus2mKOyozrmEgx2oe0fhvzrKDIeXgqhZIG2FVDGYuELPTUlH/T
5TuAJsqnFiNQd3JqCELX+1PNFTT2kz1mocL5KelSIDfpYOaHa7e5Mi6M7ggg5aIc
CHBE25bbUioPv6wP37O3UiHKuKgd9k7h58wV3iPa3Ryc8pHp/IJF0Pi5/b8GMiSO
pM4gYHyd8RraYtn63GlcJKoUed0k69ohta2c29E3PNZySLO3FRc+JPcfSRscDnON
JpwojIBNsHfKQ3RZQxlWSzdmJaYG48pGXNbCWf/2TR4u6iiIbxULpBphsKmE99FF
8RTRYXWjr5giVPjotrqjZ11GcWRyI4hzl99fULMY6YfNOGgvfbCN1DRSXL/Sfi+A
22kOy/7pQbA8YOtWC0N3Sgb7//gLwD7Y4pxfYtiDMAnCEI+xgcyvYS/S0vQoL3NF
p5YJk9+d7WlRElgRuH2vQysqzecD393KtNwel9rCiCd9ldBdyu/YOieU360iSa4Y
PCg+NdM79nzcCfs85GHerIEZLVbMkk024IOdeavJ9jKrw8paiJlybXGO7CaCZsaM
ZYECo8oeZ6D/YdeAIg/zAfe0ixYGoDuT18Tackh9+Mt+CGpIdm0WIRHPixxYcSAt
4uvATRRdOoedHjaj7Wjzj09DfHPBm5wjFNCyX11+R6jDOqJbMefUZM1dz9vKVsQ+
tiftmMwQnD4Lsa2ngzd/rhYubCfJeb2yuPTXCP5iUNcibpR9z9aD/Y9nDnL6OAdM
76x/crMIn1vCotxzhjMm5yZzkGQagOCsDbDk22oUVITwLCY1IPEFu8vqNKxzrpZ+
YuIvDvuZAkFMAbQ8NHbv7XotAoVb+2IdgSBEiHPqyWqWO2+GBTELuGRtT7/u/Dep
+IB7gp758BBAHTRv8yRWuKpBeN1ivqdZ3PyRxkpUkEGwieH4NlN2mR9uMIf4fc3f
gNCcINCwLmm99Y3V7Hvjlvm1mO5xRC8r5X7gP6ltzjN3rywcODZlM26GEovzScbY
T1lc6TSkZMyoBiJUO3YUflEO22PuBrMatS8HK8eM/Qduxdns51gxYraohViBvoTG
pXtRpIvqxybpYi8+9zcu4kW05xUjo83cZ2zJdjocnroyAJG0Lsck6B9O9yUeIhoy
oNRwAKbDOARxl/Z0fUdGC6eQTueyaAxdJymI9E++tPMydNARLhlVxwytHd9eJeKq
tHybPvzdeO2i5jBc/+UPYYJumTAIBUyUTZEPHw2XmJbIMuwditqEfYmEkdswZHKR
e92c1TpzUKL5mTrJTqCpGi4QuthUtOGueMcYKUso+xjMBeuDTuWAnVmA1kpg+5tw
slb8L/GkmDX3WCziVfb6dWySakLdyrKcYN/Lm9lXG427oS7qFLqsp6jnH5MuIt2L
myQkbAE99wunZEGD0RHHsjQONxfu76c7aGuzj7wF5vBkLWbYKMZgoJKGz8+kycXp
phFJ2SHCBcpvdw+QT9YcIdZvQepH/fLuKHPNJL3BPQ+uW6VHPE8zeeg6fd5SRYly
FIDhV4xV86xKyiQwbIU4+EzXIpYmqJ9fmjeAADST2/fI5SR7Acq6kQbi0xTjquy6
MRQr+6vhVr6EKNZQIKj8+JCjugp88CNiHayMgMChd7OiTbQa1dX9XSeUmuUVXyS9
RM/joadcUXw7+ot7utR/k5XRogbMtivbrPDg/nY0pr2UpYVmY/ftyBw1/KNcuFog
gnkOlRFC67fklFFwVunJNU5iQevocY2TKY+YCufdwx8UkxMdm740qS8gxo72SDkZ
lBpUjP2EeoY4frIzIiWKzhcaTgHvGFD7pXL3/mu5FoRCW59Bq/SB0IYMfHxxulYR
+U3PsxAONuA/drcfAAwCN38FIngjYux5daTkWzVenO5UcUw1WzQEthPW2OREF00P
4IMsjCAEE65jr7f6sCN/qZ1bRWEXOjhJBAa6BJ5lAPWQ0/urdgNy5DkgDP/pNLV3
9aHsnov11qAGy7pD5jjYiz43JUNhH58fVhLF2+upt3te7SZx8VF+TmWoWx8RZe/O
ZQu9iOJVc61DFGXtuNhLaBDExt9xoykUlrERV0oaWL0laBdj2mnEUoFpxcwphMbe
BN6miz6h+AZHO28zYyv6wu9ZFTHqlzRFBzFndaNKTCB82JrxXVK/lEwODgn2+h1l
B0dToh4q6+cX3Nl3cyYStdRbR0O6CieVsLNrw7gNXqzD1ru3gwCoVyuWV0RkxKq5
l4fvOk+Q/d1bkoaOZnYemDxLQ4dLTBTAQWqkKIJWqXVhmCC6IHkbcDL8MV7eF9KB
SZ1W3B5MkFvYHOBtWKRFids7ecTGbZQucJktiPvqVwEYge8gvYX4cyhXkDZ/u9Yw
Vxce79SDsZthU1Wu/W7zZCBKjDGxkJ0SjozhT21cTYZV0SJ/S4SdjEmsTxqXm6PU
fSSQblHyfPmzH0A4Es4FdA9KT+9f93G5mH5y5kxcuoATBtz6A2rEhgY5kK0f/Ge+
VPBDjI556oOZSmew73f390/XqHvBVaLLNBq0dBYpsRVnYdTmgx5DhEFYGHh/Nz/t
r8hzXsNK4HUwGHAYpnHl66L88y3zV/2qLQlAGONCjXTiZprUvYyPc6yqQ4fvsjgC
jy1WevakeKWd90WDxHiYtTWDqeot3nWPEvW0fpzGb7zm0blT67qEdT5Cfq9B6RPW
gc5h5eUAKwV2/cetAks9H7BrMTYMxF6DlY7ngEzAeHZQGBpMJYLE5te6OaptrCLz
a1wnqC/trBZHnrSALoz8GHL3iJo+HwABKloX5R3eB2J53yDymSfKm+d4SMRuioXZ
iRVQNS1xLcejYB/xLjqQWuAZ3MsDgFJWWKBCA45AEcVer0n/MdoaIk0lylfX74Qp
63I9EqkdSaNhnnHxSsYJW8vdCda6yb+is0FTJKFUmUE5VaPu5a8n1MjutmSMT5vC
ys0pHp/nSHa93glKXvrEGO90cWbyIx3gjRLuFfuxZbK1i1Rp0LkqKzseqbNAhYkW
Gb9g3WQKT8kk8SmaqnX8ie4iu1uFQUB/T1Z0hcU28cAFeTlfBnbRJVPtjjBuwRK9
kMRsxlIbXiHvXO7aidXlj75vRPU7jI9b1VspdDr79VnNy1ZSNYb39v3Qg6eJ83az
gZOTJqoNSM19QAR64JIKA64O9acS7BdISjP1J68K6yR14V2+h8+hSI5n5peq49dL
lVg4QlfKfQN5vaZcUNOh2mrKGWxw1kjlTi2B2wf6BsIBAwzo32e8cTMz08c8s/7d
hfdZcAz+Y+/KwwR8FvL3u9FZYMb+T4pR0q06gJh61ye9F6VleLV/RINMaY6X2mPk
LqpgGR68g/0QrCmiQTbWNPEUFMK4j/bR/YJwPr0Wy5qseTZqRq4npSeKNcquZJfn
8BRGMK2DQnOLZQNx9gEJqAuV3IHPUSLwp3V6Vd4X6G+8J6LtaTinLwpLugCBHH5K
E0g3FufosM14R5WTJiS4kmdQiKBjETWaOGW0Zast9N3xSyxAh1btsY8DI8ovvCJ7
ieBAT6KMnzdv4yqWnqSGK0zgthF7xVdGfdfbTl6Rw1rnu8w4OQkObOPwQqSUY32s
2Q2adkYzUk5PoIH+Uwl3T47cVbEQfIuST1KxCp3K2Mr36fBhkeFVJhKJ63ekOr6G
xcAvsPBBN7WNKDsuWD+1xZjVpRogxFqfNNa7UrvH5LVC+iF5x5q9qT87EkvZ/BvN
LCVxy6iY6Kq1IC+g6r44i1ez+aVD1Zi2X9YAemRVmR6qaUiBYq5oEHdlk/i4mRut
VvoPGvsyvou2Pf5PmJ10tKloaNnGdVbL1zlOXtITFCZN3y8wt1GLq5vFl+I17KDB
Kyyo8nJiLN/lYA4iYAKDFcrzDpochQxYtMzaum/85FBdFQlCIJjsHWbF4749ua12
hjukjg9w6fuTk6/9pTK/aFcrDDqSSTRFhgT59yLHd/GgsE0OKGq/SN5d8fLBjdyY
qFm+KV1Wp2iWz2hJDl15FqloedqmBAGuZ7ez5GAvO2+hF6rLWWu5L1rao/+AGlWU
d882QUaZ2wVjhebKbBXuZXwdVuBWujr6NBjf0bby2p8IAtL8apnA4XnX2XrvURvL
04SwLwkz2LVRgFxhX0KgCbrPKu/xbldW+dtdQkI6y1DkFLxGvLgSzObZiJLGTw32
7WRPAJo5ADf6sdiGM91LIqfIPJbqeRYZb1EoOzhvJj9ZRgzdkMDluBzxOKpdhfhY
rC1Bt4ckBO48cAQtN0bTXsjjBtELDIe5yJOxZT4nLoLh6giZkpGj4H3jAzAinFIO
CqOIviS0XShyC9e0pJujr5sJBwTpwXgp5cCwSk2pPd/wu1yzFmNh58iYi1LY9j+x
wjCuNI9ZNoRihvnKHSErbhxmfY/eNg9C8WBM8mwj+1ct8f6bif5JvuQuT+VZ6IXZ
sIK7+bvIdxqLuZpIIjfddVuf+CavaJu3B7x71sWMr2k8rsI6XoIk3gfdT7B1KEQO
U5JPBMlJdO2wOmpHQeePhCi2fF/lzTP4DKl9aIG03KRCS1jTxu4I+yryCBVHqNMu
vcNwRNJU2muTNCiGxIyNmOGCONROQODxA1sFM/gdgOJPtOIesFFy//wyurrj6k5Y
yOUesFNtICol9WFoo7kMioeyKr/wvLiqN2ysK4HtSmR9TzQXjCPhTexiCZJSbflR
t9XI0Umg/xeF4+IyslxzJDoXnPBqlsUa+BnbSCQjOtG2XyTZF+idmsu4GYFwhMHH
ePRRE7WvrvP3kWRemXcecErtQGr43O3FZUbVNN8O1vsk/6iwGbSZdwihcV+QtGZ9
mcchBkfSQUwPQVu2b9obtBAlHmf+Ww0XMXdKZhLrIvL8k1t6QGXYOPdukKbRob+3
mQDzMo33QPclegzrELYi3CdcnW0ZugfRP0/9/+W/d5LgWQqp8+AarfM5tZDShTus
EMHI0nHqZ/MnhYy3ixiRxkUn3di/FNTEaFD2hR7/xUn1+/n+Mu00HF3OLHrB2DA/
dlGVHP2klUpsyljwy+MytbfS8vEbkNm2SQTN+Anqf1t/w0fSK5uJgxH5p5Vl8h4l
knlkvzGF2fqYvyYSNenwRNYRKeXrDxDfOVXIjsIpt9KGPBPrRsxf1H8uQOdpyHc6
TIzYwGBqTtVXo6vH/AdyaYu6bUjvkoc4TiB2KPNyVzxcC2n1iu1SPSNlsDYSEGwR
PjstR8c3emukUV+gZrweUvtJNUhAURuanU9SRqb04u3qUUDgbbT2AekW23riDA17
bAWMrzteIO3XwEu2lNGHYOcjY9EpFH26SovZebLDFVIhiHlsrTZe6m/KB9ABkNB9
LGXpX7wtvq7cZxbW4lkq+1kYgfxU3NUJEauLVoGsQcNhPKulXUPdhuUL5sppDRtI
S175RgC2Ey6TJuswBQ3nF3eBl9vndz/kQRV7Jok4vZnphPLJPac/757V6FPPsiSm
5IGM2VKrostgIwwLCL2ggyYbwzcRVnnpYayus3oWIbtB++QSr9Nb2nHg/Vi/4JUn
RVeJsNrc9WS5GEiZxb3tW1KVR1cdCy+0TBGfBbv90c/Wf5Za7nzB4xpve33P+zxy
O7geRNUKdaehAUne18kG2+d1kAG0ciuS1u3Sc74rfvb0FljagcduPBtepcoNP/s4
Qd1okIwPoONQ0Pmc8qlVkMZuNaaLIU/GqzHlXOwlqR/+CvDr5cyodXB/4obxyYL2
/LqS51g986XKbyg5Gf3VtUzpRIAtpgop5bOJmwdDXTke36BvLeK6lKlM2yuwRBCW
YbEDpPk44U1ZeKCQ1XvZXpiK6lq4uXCVVoqg9E8qNnEKtwLgPnWSBa0Z8wBeS7+5
JHgbnMdNxzlwHstPMsWcLWKGVEAE7bjxY7Qt2K2CWOMpAa0Y9s5AqcDCM/0J7elv
1dOWb2MqQpxKoPA72LOiB2rmEMXq/2CtwMpqLMWbyzPEd1SpikgyAQfx4EjnDC1T
0JyNkLdT/qB45hkmELiikOtwuLPlvtzEJTae0WTQ+05e7nlK44tIe5urjHXu3/lU
Mblw/GCp9Jw+sq8NBxgK3FUZZHNdRaha2+Txad5lLPOGy1fO+4O9GY84b3gQ3E9j
3agFl5IT3luiPBNJDe9Lz3rDQX7eDmrdEzsGlhXZf3xaqjv7xNFE0hcLvBAE+d9D
ZgfVHoklpivsOhn3husIIdecCbxvSR+Sbzv9p5hR2DK03TWn6tso0yAvFd+7lnt4
FgzKjg3yvUr8SHPaNKtGZAyy4RuhDKOpZwiPYPyykLIyd/53aC/p0ooGyVUU7Iwu
L0GG5WQpSUKSkzptB2dyr17Ro9RMJCU/aSa/qpGvCQsfhViiClQf52Vj7lyApLvS
o0p9SPLood3ctqvSh/i8UgmZ8Z+e0tIU6TtLreWEX9WMNFS+teemBbCtYaSL9EA0
6/WPh9gIV9eDeeteTtdBEjAXZrHmxKKu6uAXAFgEK0zKdutl+IPIvGS8HQbp30vS
V8C6xW/HGqpzgtfrl33IA67qUCK8+2oHKz0yR5pkg2m+krZ89zNubWrbhKrzHQ9r
6qoWAudk5fI0TNWzQH+SZNWbYtY3NvXq4lqmNgQ1uV8uWYu8/jDJsVjgxDeHl5Kh
nuL/scVfPwMom04dC++RskWp2yQmMz8LIJ0kCrkKr54dIogIVOOf8/LA8t1L65yp
VE4iSpZyY5UizvSGBuxi7GFj65wShx5BBecmvaLRKs3KviQgmGifHP4zitiU/Z/Q
rXCgSyUofWV3E1I5vRTRgrr6v52HePhnZUQQEPp7R2GPSbj/MJ26/bzatKo+MF8J
lcgqKBvBaBndtKOD106x4LjYqZ6UJVyup0BGp8scv5yr/Os1Juy/c22c7A06baGV
cH4SxNcsYXCtFOpU1HLC+go78TQsR8fLgH3DRvkBWXdWyQ5h52bTseOp6Bm2cyBd
qmOECCw+smLY5H+V4SsZukmYL7id2vORau1So0/lxBo2Za5FwDxQSXT5Leg8YMTu
ntALghl/hlx/eVUR4WjhhFgQQoMwNCmDBeEdmmE+QiGt0hmeYmGtXtkrlEi8quy1
jwJFNyXYYkfRywnHpHxLvfMU7ky4ttr3Cs4jHIQ304QDM45SEIyz3vI7xr/E8xiA
tV4P8VPI4WXJJB7rN67MiyJgmVRX25ZsI87j7gNJyjyYg4Ckto8LDz0Vw5O48/ZF
T8hM7XWjzQGQz2zVPy+Jemj3kISJKmWCfnnHX+sAKGPTHgwsaItmBIED0UjVfc/B
10cBmx+Xhp5Cfa9l0sw3ShempgdF9oXsjFLRM4SRNVDAp4Bdmhcrwilo6EPzrsSS
zn3/Poya0f74sCyEx6RD0qtM1HsJU+vDbXIAvl4r8mST29lqGyuSItzMH98Cb0kc
VQMm4eyJ+CI5Jqc1IsAP1QcFJTHlvzb/xaSInPm9OM8g1r5qevsJ3ixd1EYMnyj6
kgKaNvqjwtIwozTeDbx+g4qMXTKO/pDb6D8jRiyZfw5hMK9HRbABt1x54cRfzdTL
iUIFTo8ru/56ricxoR8bEOn0bWBxGF2t9pc+E9sIlMJzId5gNaLqM66tPJQuskJG
disbZOUlIgisY+45FKB1tL2w7Wf0WMltk54ZEj7EQ/Z7MkBA5MQjW2VyqGLraXYD
cyr0xPMgk+U4kIwTjczKmcvmAk2wTJHFauLWfvEBUYn2TvYT45j5DRG/0KUFM/zp
taxpJBHi6KgoXoqibr9K+iPRAnAN2DOaaeLIPnXMiVY16uZjVUJ3SPMeFW/c6xQx
7PfGuAzCqpM6aTcCAa9LmRPVvc3KOnSy6YowoSejrEULbpHtdepUj0m+0af6YIZr
8xd1fkcg1ayAdSnYbkIeiaRfxvxwQdNr7s1P+pJyr3UNbl3NSpR9eZIJQPxe0pGY
Jl7P1KqyV9aKMHk5wisbJXB+dNwjL8V8cwbd4BFzFmR+KRmkExxyoe83Lr5iwIpJ
1GcC0LjfaI2/TyCx3i50ur2YQY3pF960vNHw7+DOxrnS98EzGBL2U5JUJ+aNXUY4
YemP4UuWCg4jqnEIqmfiH3LQ5nW3hDyCMDXzf7i0K5ht39tOeVhdLEWWPGgHm6J7
SkcXfZPuqmmq1EY+twAVo5jz7jbJ87svX5Wo8uOnGBET8PNOy9oI+dF0nmlymX/W
I2vq4fz90dOWm9yVgQDJSaIg/G1BN5HyOagWm8cLOU6WDH94RQWYPMqKS3hMuCsX
PhkbZcXsAmEL9uFPXe2/djicazfM4rF7megiJv5IwDHGvpYg9We/XFP6qP+tu9lq
wS1FDiKL8ZdRrUKIPTnOdRPWyDVDiyuDsHYknffTfQde4oMrPNs40sAEXN16eFZi
0GHXP4EswGWIg3GiOgBAYbax9TQNFrlQvHU3cSyYkbpVmHGA7zD10EOo6hhloz/r
KIR7+aZxUOiF/nq+KESRei48QmDRJpRXosuhKHC82+nVe/rLAaFdfqjVHl9Kbf/E
0PArqXlrjebint5iXQWMYwX7Re5Vn9S6V02wwxaeef+wJOshuVSQb0B26C6cbPw6
0i7tCVBGklQxhr9lgm1tUf30kyNwXDyXPjRLDM8GkNUhNxIKaIpcT8dIeDKa63N6
wDlJJ792LOtlCiHkjR56CSTEwLMpOkKQW6dyvjtzo6zNmgY4NsuFOSRL8G1FZ8x7
xRSO8alEbtgu96iCBmN+ZlzELw7jfmpZgk1MeijB12I+TohJbuL7SbtAiFRndhCw
KPirTSJFsfoSbDHeDq0R8CAn9UNocPXs6ohpeW+7U0pOuH5hKCXGfsVSBK+a3tsp
ikrFaOZ54UhoPmfJXv5j04ZTq4HilMYOuC+R8Ttt5i5EJVLLARdwaw2vXtvmbpNU
RA2hZpcCynfywXEvtFGR33/NdpR65M5v9H/eE3lpi1nIJ2OEJTvfaG77ZiSZ53LT
3v3NO3N707mZicw+YN8wP8VtgGbEGyD+h3fkglJeMuIBeOTwT9Hoe+NeCF2ORlKY
vNKckNcvjHsSeBheNedzHe/Tq5WT9CAaz9KBJhTJsU25Wpmsa0SFce/YCxa/owdF
RyN7ODotb5ZKyxo/KXjAJKnF6k/KZ9QhwXvCDyCly0+LASUfhPn8r6D5JezeemC6
o07A0PwhRsVN22n3AwMZOz3GnMX92YOIhP1qG9xU3uwtmzSZRXvZ0aN/kDIdPEZL
P9u9UhqRbtSxlZcbw+aGK8IRlZC+SY0YIVodLGm4d5Tyqvuk0rXx/i6CljOZDhcb
hr5AOxajFOgywFIA9KlWxKALLE7gUD2nYj2fU2N2hRYrgnGRmKO674EG0clqoHQZ
OgLN4t08SIkDbG10ytczW9jkH/9j0mcCrvTQngoChwJo/8kT4sJTL2uuCt4skwNQ
NQlBIk8vr2RtSfDIjkKOodMe4egfeRE2xs8vxfOkznA6sEUquUFs8I7LK3G/DxSz
sPzBG4f59JbfmMZi3p9JJZfF0HSGlsh9gWWOuy/2lo45A+MsLb+HehXz6mypRjEi
L6LHnyyfVSh5DGfZ3ZMcokTxC3sXThp8UGZ1ZElAwh8GHMViUvhAf73SVB3wLIJ9
t20L2gWa2Ts8d6ydYaSb9JTwVNoWE6oj/j7+MgtkFGTr7XHnJ0U0/MvVLinU8Sjb
ivR19bF7g4PSu/3W8SSmIjjEblKzgwlut2izey6AdARYCopUr7FaNCUuE24SNVoU
qib/Eht1Rlq4N0A8+WB8yLSjYTIFpQL7xYsneSr9tuFg4keWCTxvHFNgAuDUiXdF
Igsi61ximvs7gKed+6pN8Vp1Hqxk0GzDqHzKlYCvOhSXFbbnFdetq6KA5ZfiQSIa
4OJy/15kQbMuLEsSLXEhXQXj28rCCe9aqHStLn5c39dYA11ViZK03AOilqCpiN6g
Q5rKIa/S1Omi4Wy9uy8WG8evNPIP6gTByEpQ5aKmXRwV0uwvdM1fyjHbDE3nBkUx
6wtjcGroFKyTvl/Z22A1uTrtm/BpusOowM91snbZOXes1dbeH26wAUF5Wi8Qu/kH
aHK4JynaL9VXi34Gpa5KnBB7NHJmG00uJAzTsWeqt/kvWpGSrwnEOV8jx/VSaDqu
tcyB8qkf9G8cMh7krRNClZYCK3bzb/XcCeRDU54sab8KPKDolBHMz/XjgOfdcow/
0TjUrtoyxlaBQvLQlRbfsbAPgr1AoRWZV7fPRluMnU0rtSQlcI97ok800+g1mAQM
sGbhd20oDKre7/eyUyj74FapM7/ocU98g3d1lxDg66MGaZyp1vUZ+dG3KHcChvtS
2Wa/D/dh/hrEyIRge0/8bTaz2siT0UTiwwsnUnT1C4hhd2mI//4bkI0BKLWJgK5U
6yGzJgI1AF5zFqO9LprCcCPYivwtCzJp2s3ktoG2PMPWVQu9QIAg6B8kvV1GzTII
FIYq5WboqUSRv85Z2/JPzZDiJrvxC/y5PDchn20iBNIdWl/fKUIF0U15ng2kVt3m
5e3bnFWfSY+N3Wkz3/IyWxvCcB22ma0iHIzs1tQo8ejDLHwgFHcc7WWeZZl8ugeb
+S9GBJatEvaJHjCv8apl3/aeD9g7JWyK3/uc6HWP/6PWnkYQuMQbJhKOz5ty94W/
eVljrcvydlYbwtSYnTxZL4E9RXHdBwSfRZjIG3by959CSU8TgD70iiKHg1iHxFDs
4SBBuyKHmCzD4qjwmMp035rIZwE9lRwkx+OGWSc1vmnOYHizKTgpDII8eLQaKdFA
WozYscWziQis2zaL6btkWUutZVU8ZRDokBJwKEyrYWrR6vhY7ab6oj6j1kQ/tETV
kA6LvR/U0Bt1F82/nWgAr7pC/JITY2622QsLqONxTB7nvGhpJ8bXNRwavLbzt2eU
VxuG67GnFsoknzrVSwOcTBA8hdU1USckdOU5hnQ8B3zSnzEZRXQvJ/jE8Vy0Ufeo
aAVuoWo/FqN+aL4OBqzrmgLUysWT1EajvuY2zFWuZKqWfm0YB+xqVaYoBNNqkCIq
ztovSHMKwjruBHumZHXn63SrH2aQGMVy6jMBlx3W+PzFUVgyWKbyBDh0AJA3eRJj
DzeTkOa1lQoJE0HGLzI8K5aGeErjCFV1g/eUnNjuUoQNPA3sB6PGWoeQsILfKRQV
/xsmaJIUMe8WbUvQu4Cvpgm9XzvRA7YcILZlvE+4LXO0p+6NRW6ijZ4zo69QOfUr
7AGFf9A3TiR48eYKgztrnRY8j1qXosxD8VjPaCxtt2vnQID6L70Th7yg/U7K3ij2
uDqIBK6C5mvGHvZOHuzRwN6GALYa3c1iz/MfpJ7uF9+/FnYhxB0Yr5nm4XSiWjwJ
3QjH3hLBQM4wGlbUDpN5yoFzc67zpFQDKT5W6GtBshKNl/cZpYVK2AP5xfwc4czx
93O5tRZUQhC1/Kpov55jGjj6yBMqdjbmjGw4+X+NsDOu5gdeiZBn7BTPj9LDNKEH
0RP26XZkp623T+if7mNozwJCvQAm1L6undJ6YjRnN8awhRnPVyBo6ZIzsWz+RihG
AP0ppj6AxQsPfWf/MuuCPIYazsaB1Mzaall71FVWYXVfUh+XVPUgSzRUtJdShJm4
YSnEQKe6EX/kgWe/AsXgi7NMlfC/nj46bfvQzuUQgAv9f39WJnnBzChSXXZGyNgV
r+LXoqtFajsyBrd+UYV9qwDiNodRLT7Tv11xhLQxw6z2MXFz8Wh0mp4LADCq3XXB
/BPclidF6+qzTkO3IrR9LCpxXAcYDNRdpsgZftTUIpfqRhSQTeEfZEiEPyG/6AcP
IkyU+Jcg8MapB6n051XUHgVrMFUK7FWqzuTg/Jm6Taxu6NS03uc8KEPxWzvW+dD6
0WNNFu75dvagFeraR3yRUbIn1elp5GW/DsPkmCDpRgBbw39A3qbsthkUlUF7A2xO
/VuaJ0jckZEWIjwM1Of++zmKolMqWqbaBUMBY0YyY3N5DR9gK/Pc7zHCeDFnzRn9
jgEuQb3zr+lJjt8LMUM/261tcR/LGx0zj/TXq/e+1h7g7V/1uwfZFt8bQrNYhp3U
JKpYcjlR2kWaQyHwOM3clfYu9PifZ7leqMgxLeJEb9ZoPZCqbIsJxj//XH1s39Kv
jEASFD0JBsawIlVXV+DvPHPzLqc8OTA1B5DISmrRGU64oILzey8sEmm+dHdgQ12C
nOerg0Ta1CS+YZ4vJuIf7MGSUNgd6QQArROoOldhSyvQd6SCcccxVO8WW5KqdWyE
3j9izn1wRFqNnghxE9m7dTGND/zoVJPU+BhePJUmQ72OJOTfW7yX6WiAFiK03mx5
G6hF9EDqvp6Pukv2H4eGML5Mp8F5e5T/xbPm7OqyUEWYAk3Y94QNjhgOUrNPzi23
SD+sr88ORMiC0s1+raacUemLvQnkR3u56DKHcw+pvBzO2e2K45xMYWG6iUtUUlAY
VV7D2j6cvnP6VJCxR25l3tCejy6i1Yq55B+Cq1H7SnyahkZV+k41qcZdbGdKBCih
ptPtaF1q2C1Dja8JF00T3z+0v7cuegAikaIEImuc7rIDJUMR0xrI1pMd4r0q1cXJ
GzbvJWmFGjpzxs6p7E64zIb0r86rJkmJUdLysq/M+C9uDqRxCp6K6fJCTg58ZAFu
OBpZo+J02DmsB1ywt+DZC3Rdn3gQR496Bua/EeuOXQluSxQR7Vix1hJjUluhbpdG
0qzFUekT3i1FkueCEmWLnupm+xuEOZH+xvByudeb0+xGpOKRcRfRxFWOp/ER+l/s
nR9ks30F3X+WjkQ8aVo+ke4eCm7qLgy6/kEWoVbEKCiwo8NbWG9FsPM0ZqNBAtuP
VRpFtREv6P4GRqGhk8nEHkBVkYBYgerYPTVKs4TlJ5kXRaHuBS9ujDDT9u+udtnU
uFhivssCp36/VxP612tT/3i3VZnWgnHTQSEQFpr4tamvy2W1rn/BbBCG9vwy5Nhj
Ux87DTxNLLSKpK7THo/1O6F8b6VkJ+CIdYCeoqALnSwx6z9/Ws0eTi4SWJw3T4WX
NhnNdEHrZYaueMe8t9Bcr77/wHkDaQ3izz9qGOyZGhD9pP/DzzHJ0x3jJVJaQf8e
lW+ll9/zoDZ6ywVh9qfEsItK6YFzLvP/VwSWlCTVsLfxQQhbpcFDwyBYexWslj1/
YGJAiAdx244Edc8LW7mViJ10WGZQckZ2UrBZKzgu2YTvRlJHkTPraJOSf1iur8bR
AcKqxxWloye4V1mje9WYm5v4U5O/czZQ7ivnVSgLHeSIXkVj3nkDF/hL+glkRfJD
VeQuJnXgjK2bAhPTTa9bPqR/SM5La2poLypofaB4Psh6/a/YM4IVt7RoN63LHQfL
ohhxndUU0uApEVqw9ek+ZQhlKZpvesn7K+ztYtkN0wFAmwiYNkUmg2TDxEBEybDo
fMF50dbvBTyyimw53g2pxdbJ4EjCHQewbu0JQBXcXo+i90YfeJafYpLkA3JuL65F
4/uJ3Fb+Ch/QPMaCZJFhsXEq6boVtoECbl6QuC+w44bxAYLBKwR0TbNBjF9GQQ9j
Z2ZISTqTUDc8o+Ci5ngQJtyC4JIKU2oKjbpEhXgppz8T+gGlQTXvtD4pEJil6K7r
tVjHBQNwqOWTUaIGwtzA9dj7ZL5TZu4vfmK+GOmpaC3C7kM6zt3L5bnqAiaRsNpe
WmmmmLivONDAFSLKwxzBrf3rNvalWXnouWIpsUZmgPxm26OfRlZKLfkLPndrIBPp
AwcD7xsvFflOqoTpN9v2nVik19ziLNHyk80K0vumKCEBxlgB1IyoYrtZrl6X0cpv
EXA+2IfrT0cXZWt+HDm1lHDNpjYZGWv2gbhchGQKw1S0+Iz+JoUT/qytuYjIj1IZ
Q/ftBFrzuxSVDlE2j0swc024kP2A/nbrytVwZdfOzgEAscV+i/EV+KSFYITGRcJQ
pi5LtQNxPDOEHt8VOBCJiMt6nscrMPk4Tyf5uA0vSBZteZS8kHXYSkKJ+CqYAim8
t3DgmFOpud9bzVp16D8hY9TaD1M/lsrhH5lnhAMzl6jaA2gfxItwZ+bGNuL9s1Rg
x+CUzr0Y4wIMcnrqG09Bh3f14XyFEaB6nUvLRU+psL7Awd3LUF/gKb627ZCUVYpy
sFM2eqglOdoQwk3WM/dnI5pdOExDFHtYUhkFQ9kvt0yc7Y8zWRdeabuXEQnMou0Q
V/v3/NR3JCzxK/lwNtwTRQ1mP7iNxR27xAU4SVQ74HD6V+C2jPaUhEeTM3fNhJc1
VkAdbVO9sO27h3xbTC/KF2hrw54uwmN9x1zdjX+LZtiqnPXtNWm59hz8M45HOPne
wrN9hQ8sQyl3VI9NFvqkft3Bw405+qnMG0opjYkgl38K3NZUrpMOQhutikkAlNUs
BVziYEBO5f12eJjuD1EL65FGpB75vkm+raua/Sw5naMjwadrW5ynqSOTWGX6AjGM
G7dcvAsDMax2qklVMUlc89NFaA2uD4lPh7cXpbaw1y3nNQQ6AgC9Pp+SggoMWDOm
gqcoytN5M6vTLFZ3sgWai0YX8naDWohRpSAi+7w0OLzAfHaPQqbT2YLWeAR7SoT7
t2nWpVuqJIMczWKiU/Fi+28Av88lTFR/FXjiMZN/nTv19eIvxxAZw3T/UZyGp/AV
e6oPhGM5DAkAF8fJ3oayJsAH+mF4/J/XI0BqZ1/1t889ohfzfrZ15io8Lskx/2XI
2lo3tAfQqT0RuI5tUbxADfVGHaVYzr6jQQIhh0WtWHVAsfWLHJv3VPpppXEFnqRJ
d1o6XsjVxwDDY+78Gea13CBfe/B+wRM7aJLwhQRJXizITA+wDRYJh7fdhz4e8u5Z
BIyC+121YIWwBB+CV1j5paztV+31BzLXfH4/FFN/g0AAl0IO1rWdnPjgbcnvhXLe
DZyzKI2zqq0zaFUeabQRfzOW3O0E13fXmc8zJ9BHh2Z093tlcEb0jVhXgLfbjDv5
Ys8eYfjL5mgmEQtzjcgJhwb51WwDlHyN4HGKPLMulEGCptfx0krmiFLeKCuIrkEV
rRJW40TXDJSBy2IcT40M3xgWnreYzLIsXDjIYGrZQTfJCzCIOk9/J3Rbfh5NpvIe
4Xl9yOJLXt02o2xKIPLnBeMZLIlVSfA0xy2TwXl8fRUulJCdu+1RWaVri9JMsikD
83Prd3eaKaRTtiKLeWJdrn/KLyxIB/5SuOTMdOe6pE5RM0+8zRMSVdhdzm+FOL6S
x7P6zM0AKMvJAhvDfCG21Ccsp/4jsYT5ogSaSn9mcSFWLZ4zCDzuFh0+h3XtkQip
schv+WUNihLP2kYPwEf+18JUM+SLQW/hcq3ZYi/xT+F5TN6aFrmmKmS9rd8DlnW/
+071jwkLkIUo7UTmnrbRJT1XBiiz7uXeMaKqueCmi/e8E3n874cDBQtqu2okC8WS
iuV1XYVEC4Q9mqrwS9qdjXkbqBVGtgrdJfpMqdyFY1851WTNo40DZlX2WMmx13I5
u2MUVy/T1skUJmrVM339jz/eqetYksKeQBfmuomB6799O+/KVRoArEkYH/vY0RjL
B4df6uHIA6UnUO/G6DcZFoH3isw1urk92B2DogYOP8B9kWAJAXB3kqj8NYXHG3Jm
4M3p2QSJbXUvIBjtmmRCdtWepp2kU08G3yy3R03XZ/vvWFI+r0TxWP1Uj1rzEEIp
XgTv35L6xf7EA9qmOiswAih6x55hqzPnTV/08szIDdO2SxlFDN317oYUdFqCpYpx
AM+NIYmisd2BRx2NboDpPPXhKKzDMJKcJOmRghKEdW3IoVPfULK/pzcUZCNiJ+1R
gAqBQSCY4o9yaHH+tD9UkYeaNwVHbgtXDMKujA8kxaPMBlsf5f6/rPxlAWRWaPMR
cbIjVhCi/rvTRsvSN6G53DOIi5Dh8rMhFsG4lDfVC9/xpVVZESc41Gap6WDcq0WR
7dPVuHk7jU0R2vzLOUaargdJF8LhjcOQLb28EQrM3r+a74bD7XOzD1Ll43ulofi2
M6F0KyaIPs7eZyHBCmMbcPgnGnXFzStfOs/N5mxjG+D4CnekRoHbxrwfJBMNNYts
H6Z+P+wMlnGZJ1mKThBWjdnV1st+45CEN/Tv3YDdsZBweNfFdUg8/bIDrwcrGrb5
OGnVoA5LgEv2jM1G6JBq3sTyAJAmL7ZT+jK7id1LwAevGQN6mraiVnhcellQuawS
1SCASlYhJ9f34cfIKqctDg6Oq/xAfswC2rTw3JUKgrOTZZ51sPHpnkIYArCH4XTy
9Qwm71MyFA7PtVTkswxd2C5MrDPs6KOIBLilXnl3K1/+eLkINCab/Uxyp5YRzTP/
YBcdWIo9l2sqDJrYS/fPohNKxNC8V7NEQya537fVlGCjVNaGHuIELzyz9p2s1ost
EtFfdZObdsWzR/wIHbxCqVn3a1PV+HA38GPWxORtrUIwZrbPblDSIjcIIjIH+oUR
KimAT4MvoHjttcQv06bOHrx9K8y7dATBP3tKWGglY53C3c/yDLTAlj5nyx7h3Znq
zaJHPAA1a3whycyteIt9qVQH3RuIAK7ZXwqSsjh70JrPJPPq26VRIiq2tBqWw9e+
28m5OduJGOSjojJuHbbBY/P6qQCjuOQl/o8pNel+bft+2NR5Gc+MHLoBKzgd61SS
5d8cc7nJIhCpLUkE57ROU9K6XN6y3QpSca1pq9MUhB/TzwkoZ7nIB/BirL8ya7Py
WKV24jDvx7ds7jCghV2ZvfUApFBz++w2/KoTVKnslv9IEd71aeOQHOUkzdYbq/B/
2+vS7ouJGHBrMV3b2c3c2Zwzj4dZSVXvBjwHhr3bKp6KVKN3yOfy/9vQJMEfSgdQ
jFJpS2LwF9sBaN+5e3f8e7pYmhKrGdZ872pBM+3G+KgzjrJ21cyFZvSXmUcxK0y7
FIc+pq++HX3+wHmP8qe8IIZx1agZBvBnPZZZrhLNBZ4ehOubMsF0pUuQRAobjr4o
2i2zQVB4SXwLVMynvcbeFOCa7hiIQWo2+TGsXhG0bzNlgiaeF2FaZJtMmW2mNE1D
JfzhWlMl0+dJWiznAqlyTcK1MlwbK7V6QgkcStWtHzc5cfDTsYlus6pQJvDrERPE
r1Ni71houyB+JWCbnK3aMpPEIRVEDzJLEgze+6LzjfuawuPOTGeNBMVI8EGZf5Lx
hpCRVkM9xM6ZmKzAiYGLe82vbGTpBlAcdpTQ4cc4HfOXb/WWS9+xhlPBzz+uc63v
sYrijuHI84KvQ9ENCxdWGFEL9TS6X94SitxI94UbC/OeCpifKKHs3UaIbqDjshsD
0QVMX95qedN5xSY+zycdG9RMbYtDim8YDeAF1VUa6Wy4q99B8moRDBptYVbiBJYK
PThyE8xjTh0wXkZNaezpI8+hnItT59oX6itZLrsgMArL/Mtx7VDDOgna0XHhSEcT
TWND2ZO7LUs3c5wJgG5Z48uhwBMJbgxQpKu13zMwidddCLVUykISjT89/HoJ5pnI
7DAbFUC5Jlv44jx9kaW6XOrAoMGQ9Px0UbzPi0TZF0UDWd145wiWaLVqJHK9D1Hm
sdC/00l2SJo4K3yTsQlDoDAY8X3E/6yO2OP+H+rNByx1DQYHxjM3kxAUWscMF7Um
56v6SREyspMhM9mGAWyN5b6+LIh5tHo5Xuoe8cqWmnivwiG4aqhfDPn4Ev+VjYO/
bIPE7in2gsH9aFWlBnGCOSbWpFj8MLzGEbyvDaKvwBYWZ0LYHhfp7asZ6YKqJ/x4
vkCJLGVzZhVsVDf+riuVHzDnMCFMbbeI1GRmAU2z0hfYTvKAaPqVIP/ufb4Grm3l
5ZuxeddlrlnfPHuZEUZ3dLEzfWDoaOar8H0ZTKvtq8jfHG82DHZRJRGijw69tg8u
j8P2nrDgg8761vGFySO2/B1T0W3qmZTPdAgTh1b+t0WsMPRtwnnV/XDAGJ76olT4
Y0AFeHY5CS9s0TxEG/8zOg4ctMOmwJ46u3O9FFEotNAhJmnYwGOCUEDbhQVp+Ohr
Pf5tFtL8BfV/cesaqIDARscEAX+6zPOcoFfgUIPdhJYZoTo50ncpPVAKKYZhGV3Z
nEjnjWddb+pbmVVZPYRuSOaEE/+zK1xrLTJNzEhSwfUVoR1Muf7oy1+OuPSRSy1H
u4p4PMhPJEkt/mJPQyw8CmV33Z3dJEIGmtD5jMnpHO50e8DLr4nVfySCaJ09DYC8
GW2vQZAoUNLrU+nudmpnzyL+/eqfqr/vWkRLsck1u7nR1eU92IDDJCCdA1ECR+04
nyUbx7ST5Q3bZe+EsAX9zhdul7AS7b9HN0lxhLsmHwMdRU+rGQgYdD+kjjoeEPrF
oA8bTeop7ogTLT8/5icaFSbNVqk6uXWUw2UORFG/oRGg/7MXWDagci1qLPejD7/4
7TILSGQofLafMvP0kL34++g2ig1fisf0oO+hKqutF3b3gs/z2sBEwO0kZiHWiSlC
InlGegubXkSwTwRmCgaH4clw5EDpxDMk8W6udAxht6ZzSIK7u1IdjInB5n1tjkTD
SiVzwXErXuBzxIpTThXXXT+GVnxCSjOH/yRSX8XSXVWBNFcujZ65l2euZgC7D6q1
X+a10ItWARFFLhzXji4qX0wWCN6zfoYy0O/K/skpgP6wpCPYMFVQpDuNd8E9s258
9C7P7J6kbYSddB44wRv5pQuioHEqcG6MO7c/WsKc+Nqvhl3OE9cSUKR4zelaQk7K
Q20orFOFfLx4AgmONQ7RR94fuF90Adnreoj5TvntgeQ8N/ohJwuXE7Is4QG65WHX
QNBQvCuTWE7/AWw5Ta9sQFIH24UA2j2kZ9afEzqfI9q1RiniJm5t0EJnIFJ73B98
QsMCHwa1m3Secjz0Wk8HObIHXWkegM6xuOluFaxR/rCqLZmKcG0N9xhVjEK4r2FD
bkdSg53iCbyHWQecvs+tO2B125sD7cC/80pTz+82pokWjynAQcj8xh3liK83KeAb
YkwKMiBWOesoujH8XT9gyCfl460pys+/TObw0tE5yd/FLijeLvIdZRfswUleHrDb
Aj2zKCQNncvmG6RADug/sami2FnmAUYCgFD0JfNiF7HhqsFUjtQvuYnrL6jyaCXw
FUBRd7M+wSNR98GzlXglpy1DJTXjmCXSnk78/KMVdE3c1PvcC3jNli98CgA1VHU6
UXUrdzBz80TVaVUiD1ozWS6qcG5js2E/c5bERZbWHc0mIIUUu+e+t78LSu9UroSh
eEj3m1yHyMYkel5H6D7C7X4eE1RKv6WpHDZCijPWs7y82z+oEB4CAq3mcDFrXtER
4ZgOEVvz/BrofMd28icW4EYEa3roj7j/HaSltxvNLzgrYjNtcmW/de+R3j1Bs5hY
4liqp/4BXCTvzaH2sr9/9+RH9lJ/OPciiJKwO5tX5aCLwdb5WMSsDh5930YEDM5G
xn8W81e5eOjqdgxi2arapurmWJ/Gzx4h3EsyvJNwGmKTn6YJIB5ZW5ImnnKQz9WP
DWv+jLYdPOCOZIUYJcRAoW0joGMd+An/AylOxLefJUtuCHUOMzEnTdouWci/mvN1
tWEqB9b3HcFeeORCqkkvo1ogPR/7j3KZ3JRhEWUUiLK1k5uOT4naWO+ceUSp/Dyf
dteYQJxag2140wkWeUnEHC+qBQ7GCKDcqJZ02/1MbV6m5f5VjQVjHw950z0W602+
TqBd+LC8k2lvhIj6/o5M2IPl+33/jsLRpPdHY/oVfJQhzEdwleMeYakoSnyADpO3
yfjLtYJW1RRg8XDGNzCeaSooKq0CRY2cWCxgOY2pnSetYcab1i088r0pE3XurPEp
0cR7vURLkZkMGUnn1DFldZ/nJ8hCMqeB1HPbLuJGRw7BE6j09Y2gj5LDnYjybra9
RT4svTikINIh0O2qTHG/3ztFhtdr5huMdXHxKOgcRsFOF6vIsKWVJ+pJpenuHTXB
hE3dRd9v5tHQSVLCVKsG2OpN9T/N+RYyt7I6m4mVvXYM6sd5rwnC056eAtfFb81b
eUqcQWyKK2ihrmgSlF3u2FeLn1UGYWUHtfvEX5twDAa/mXQ3KrI+bMCldmKh8o2o
mfsrXK8dSXXEpUhQ7UcRMzbzH4eQ45zJZoQ5oq2QHc1qsApHSDx1F7y+8bWcI1DO
ov7u8icjzbZPe+U0DotntGbDYQ1RrB31PRdbKrbIOigE4FHIRUBhW8iLR8kccH4R
lPN8L8s8s8QwNd+Nl60T7INGVDfPJaCDzQRj7gxZHJd4+HVVZkkaBrVP5183MUy5
dU5ueMjzLdwu8KlUmE5bW777BilbmbOo3oRrBetUtDYCQwdW7F70lsA/CxPgM5Ih
nErvFmtc8xdBzn7ZiJiqi/L2AxZrBcEUMz/mGfshVefnIiEFSJ2QZbc2oZ5v2kRd
KHZccPwEzqA5st833ka4hM9oA0NZBeoa9M2WpW7kJt0nEdwOmZsSzF4ab5Tc0yCY
SGgHc0nZ8oqGnAW8PEM7/+fOPHKdX/VjAAFEWdIJm8xjgaK/dyqLrkmQlchcSXpS
nJk+3v2fQVTuWMPNiwAwWZvrAYZo26E2i2EEw/gTNQW1Pws8AgxWpWFwp4da9Udh
2UxlWWPa0NKoMo12ZGfbgteAdOWnDwMe6xYqFvoXThGDH2Tz7Y81iCyEak3eRZ1b
dls8Gtcc2WOJif+YHtxV8e5wFnI5wz98VKv4e4ao1O3soMHSRA03rq0qAAtL086F
B8vJDgzUSsv9QLdke2/uiU/bqSpRq+g4OzlBtGD05qkcfK0hDxaCl/Fy81msPljr
SlTJd9Rj0wAqMrJjGSegPD0tiGAi8O2GMz2mc21/ztBW2brJ4w8PESThfL1HZUeP
adglApYxeQWsZXO6poEJx3oTSVZeJBJ/z18jcHbB93UZGLO1fpewZfX7lVZ4aPO/
pBikIGxg4FezjHP8BQG0G10GtKFdKQ/cJG55+6LPM+UiwXAo+mjyy/M3Z8KEAvXK
iy5q9rZ6cSSc7kCzBG3iY0Wje2dsnGep18Ez5mHz4dBp0olOZit7pA9pUxJu3qvS
JXj9ulpTtgXVMNZpZiSkqxBstpwE08kkLlzwBl7tYRtalgQTK+O+Sd5odj9ra0pv
3JVKcP4STwRjZzaee9W0il5tNzBxJSTgt9B0BaC201cdV+XRf+/iliqdNmk9vfbt
IzwKZUi6mC4nEGIEuLEv9C3G+1jkU0fqWfJyKsILJTgwpvbffswOWrLmuw6NhnUo
VtlsnNq4lcPfZtUJiiDFo1racpJBbUBVFLGYwWQCqQ6NqUDDXstBLM+WJRcczdXN
eySYiDr6U4ymIcR2YXhdjIpR6J6XTTSQRhTOWUhSrbKPVTCqhGn/2hrMmkuZbovn
/nPvlHKw/WMHQXTgcosn7bnBw+IncRUoabOV5TX2GVNFvtQWCxQD8L52nea1Zfb6
qqqPoakmHALYDej4oJxuB0JGoX0fUb1+QkEZBO+ZXOORW11F9EqYo9XCEhQNBuVD
dkDFUw256nmIXSNSfiqGwTpS39Ew7+R3MZEIUZxKNW9k92CVDo8O+epbxRktR2Fq
qc4pCup81HhrcfjqvYNXlJb6GWy4cgkpZAalyCJKE9K5azWrrDdhkLBRDMYSEzPk
XhUiJz+JkLBzSzekDgL3qo6U8fXK+VQT9Cf9QmvIznPOPGKP7Vkn9tsyIO53T8Mv
cMQg5MBMTnViO0G4WXmZ5ecY0kTdCKG0EnXLRgqn712zEZIO/vOhAeY/a14nrjSc
eYeOAu8gdkxKS5Jx1+Slhx6DchOmWfBJ6I8wlipBXYzC/qwX8jmuOWpaldKN7M7/
ZLYKnbZ6OIjq5JNm6MhSfsw2qeGLBuueBkl0b8WLswY5RszTVURFIgqpgKQu0TcF
hM/PEivDZL2tztQni6KkV+vA62avkY/BSYAtpM2U05WNSXkp0KwtotRa2bkF6Xzi
yPL+nLKX4Y1GjxcW4vexsK7KM/gWWzP96poHO5S30KsHAOhLiTrYtXsDRnpjxh37
2Qp59DkpFEMNAqw4XUd+O71wjaT5gAVdprl+JAhucrY/9ZHPhYqwrI3Edxvpxm//
dHqXYAIdoH8UOxyhZ+ksNpGnQ40FVcpxjfcgNjfGo05osQqsQRTUPq/Y3r/sewJg
lFGWg4goo+NaOWGA/ctYwJffIPxEldgnFrnwWp/OVMG5aIlmfgNzc0DQfjO8CNlU
7JYV633Proy6mLgDmjp6NccRDMPTWp5EJV42GIxeTFS71WFHx5BwxA2TZi082glo
P+thPPmy82Q2sFmdFUqndUWnUQo7theLFqTfKKI3sxrQT4m+iePxxA9UklF5/AJo
uI8eiUGGaDW2O5Zn0NJ639cq40rWYtNBkcyAl+9pz4nODTv+86MwCQFWqGZRqvik
IAyH1NLHGbjhEarQBlisBtxdAtucU1C35XORVIMTaqoWhR3BPEQjt7qt8LPIiuXc
98oU+zhoWXBcevzokNfJ9ppj872nqv0pwctJHxrN1a74eiGPCjKsfjZdN7VK3IRM
F+yzV147NUDdoA23WKknY8g0Rhao0oGfxI/YQS0zYPIFjD5ML6NK31deIieiwzUP
VKAck899GX29k0A5fbPE1IWONYKy7l6/dRpWbOK3PasB63zjs9uMU6f7YmgYqWJI
gZbrFSQJ5sjLYlD/57kx05ywmQq9mmHFbylldZgY38wxekXsZuB/HZgjkMdnvyz2
VtpyHDZ3tFIxStd+970SLizH4u6k2Q5+Kx2NUgQQJ3thYJKdYcMwJT59mFB0IZkN
5g2VeLBqyqeUMUFWKMvtyd/sTgud7xWNJf5eEbtZ3URZwziQHoD0NusjkseH7m3o
2GhnC/Uve9tX77J6IRYVsmA5qdQ9+pYioFmO9igxvGawSOg4lNYDkVEn3ysy7tDh
Xp+zJadG1612GGgCpzDfWMd6kBiBN9bE29f56ICJhjAe/bCqcEVNrBCZ51IPHco+
m0mmE0+z7sQpEVO9tr9sQ9LMftLLXupHLKcVdeu0D6+jhdaBfMjZKUnQ8xrZBSQN
fLTeDmQPrIgEiAgOXuQhIGWIHCwLqZIYU2IIi65LSZagKX5lLq9rd5Hg+nX6c6cB
3Hvy0XrjmnQZvdNZOX83jhLGR5jX0D8reFKlhVMQlI7Q73nrIo9EuxnwZC8IPTXo
lewzsVDiMyAKZ8+g1AW1OPnZZXwaVUgXYHuk/pRp1M8+JjuAzBo5zgExqt38V5FT
KuumUCZ6mE1YtjINIkI7uluqFb/p7KYu1l4To+04fab5N/fzU+uo3N4LLuKD6OID
xhYJ2z/SStRi8O9/VlblVoXJbtulTdmCFGVi89oHpH+6VbY61nIl34cQJVYkH6St
BZ0tWtjerA9APuw/n4K53jfbKy9JptMJIa+3NcQd6VngpWpL29oYuZHJcu/Vv5tG
eJ3QLohx4fwX1gzdhrYJ9zMkw9Z1aipURiZwh9teezAoYarAVQGAVa0DHi/3Eau1
SyWXKUV4Ln2jmm7ZMRoviNVGbuA5+g5vE7b2oizk6XsuMOiGB51MG0ZroVu117Rz
mU/+f7N4PU76yAzVuDFa0F217sXeZ8C92GTKSx23WdZvdVutM2v9A5U+qyN453ag
mPWDHeOpKz914XQAnDObCr984cd36y9Pg5/0SxeYLq+cMBGmRR8yt+FPcoYqFv6k
d4ZtIvkCR4pd2xf5LM/MttJ9kmkd90XCxpm2TowzvHZUmwD30lq0ccRUs/hmPCeo
9gdpLSRh9WuY0eyTZVpvvK1ozFILLv/rcItBZBXXqOWp98vE2gEfiSocx0/BBJnT
Vq4P+j99GMs8SruNTBJdnyrBo5OslxmIURZaQHZgRAF05Jtm2e3EpJOJGdRyB4aB
OY3aOKjId0RutPJr4j+qwnb+tmzA6MkPRdqeauOXYXqKBLWJr4+M/TB7K9WNKdHf
jLrcb9unVMzLz1g/Z+iIdQlAUvALticeOPrKnE3qhssTHbwd/RGZPUok/nvc2HGk
O9b6+PjLQ/iSt1B+S51/hoZnrw07KlXdW9S+UrIlaQeS7om75nk+mOOsLqCEd96V
XjAYyEQmfPrqo8zB7Q7WXmUULbfJ09T4aV3ZwtsEu8PMaYgFWvHdFfFppRdBzkFl
D1Q7ZGS00493fBJeWBx7BILnM0jLvd0bI1Yc9VenWVTI8vJ7I5IznfG8hQCs9xB1
TPiqe6IzX+Was/QO24ZHXnwXLTn4E6yC7ZDFc6aNF3rA2RdQBPL7hVvunmyqnANo
NLHLpkV2H5odIvUiXwjhSs337hjRPq3j6OTVZVbItl3ySXx+TlKFieKRMfuZozbY
6dTuBnc3j2NzZQ3yvpTJX9YbYxeLxMwUhsu0gjKs9PYk5CDFTz1uvTrRTREJoX8Y
iiydDRxKFbSUGsjM14xOrpQbGTqfbJ5CoC70WPTMlMzqT4AE7oOjV8CH73CMBly2
VTtXW5oDc+0OMVyzFSiSe8VK7tbh+flUZ9AXLo2sfAKHhbYPLwTbWB2VP6vFlJmk
bYQ8tw2Ol9ys+LkyFrcll1zaEYtjI5eJLzYenza+S/Rr0r4b1C0iiTUW0TAeRoBG
T3cRcT9wHEcsVIH6e0qYjVcjPf/c1jBDiomVIofXk3daJZrYcOLh59DhbSq42hcG
sMgBC9FKYVHVZo1yG1EWloNxYNsmqLSe46a84Xw6Ey1YCC9QYVzV7XIe2b1UufUC
BNxnyZH+ImN0RwzRXXafeSHLmsTt5bcwhHgA8U9LReSWG+WL73mv77dIkYVqzPw4
zEEz2uNIsfQgX9jr7GeWYyjaCmi9y6kLi7zbZim2NHAr2eDGAxnZpasckwTYHd2M
c1DBXQZTGcFiaVCTyhTjlYDiXFgF78XvtWgK4LXAi1zpiXZ02PTFQ3PXUFDkmGCM
/uTp3KZGiQ+o13zDcZ3ue5rQVew2CxtPcbr9W6lhH5grXPDKpQPBnO5m8IL+RT8a
5klcqFa1t9ClsZywU8dwfHiy6dvLx8yAB3oxvtR24LBPpTfe3f5HM4GF0Fjkrhtp
Dl6+bLr2+pHhOqN2ZCUUZ8uOxXs/v6BmbKKUnf7R/bCtRkEnwM3M1jWSJysUQpS7
rP0k0Q2Uf6YfW0gd/DgRMYCQ2nQQZ6qaB/6453BBVG1ukuROszb7cyFbAm0+HtGT
kHZ2iXztYngAVX+aHLCBijo/JtyZOBE/pM4KdBCsPPCbx1FoMbcfldvbSnqisUn9
Ej9nzPcdXgDnEsXOkv+F1Eb4Jb4yPiJNHcTR8DFfAYH8MZZdsw6VsO+9z2KI0M5H
E0siu38AoNpqRnj1j77r9ZWKAfEp+5qNiF0PkVjN7CZ4iJaY/b9nshCqVK+Oe5Ea
WyP0x2LXIJkcsO6tM8RrFbnmw8v27WeLPXj7U89bO1DF/vXG6st49m0qux33P9yx
UUToSBYnjLng3QIn6FaTWIzLY0reKO7/6fuvhjPgJfio2PP/Nx5p0zVVTMaqomic
2aRrG0Bzq7td73sglOSeuTKsnDX2rAAcSCB36NesvArNro7v+ZB5WoEGtI7r89hf
oPAThaQdzGkkYUYnuEELkycsO//M15b2WVykLCiuGBxwuZsdAN9sO5EJU5MiU/Le
KaDC3MaJL94WSN/qTykzVw1JFyL0cWy1NDbW5DEl8VR5zHtTkfIakI6KVf3wKilv
MNf6dhQqq8TSMjuKOVhAZ68wkKLU2qcmnnUIjECx/uOkZQxwnf+Hemsz42W6rVtM
XxK+c4kAKXz5O/xqXIahhrFoZxyHYSM0SxfMf3ANbteC223QA8yF+5r5ydJ1qqT7
7OgFqaYAvNGiKkYdyXzjYnn6w9GVbc4K4Cy+y/I02OlZnpLYoyXJXb+sNFV7AMbI
63Q1WL5NUilzHT1at6WXf9iMUGI8QHqUzByzA/iskW5e4hdbQnZDv4AnRJz6cms0
sdijEtvNEHALATk69XTrJhbOkrH2S1yH4LBlMIngVc+bDq+NXgDyyUvI4pjuqcX5
k5stq7JDyri4VIXiQQnQ7xr2sLpnboxW2TWidXIXH766h+3ZHaMcuRswUtv4yTk9
3UJplwgRHBa0Po5NHOczdHErErtBUGNtXo/XfOQjI1SW36hodX8Oso3uWQSaWKg7
D82+lYzjp+DJ3KpBe+6okEZ+dNCrMy7bzvxHKjQ5WVEzeuIldbN0StHjg7LjdPeJ
/mxdbGAnmj1p1Kk8yCvgKRQlfX4Dv8pNsbUQXOwfCELqgyPY8NhlwQv/uSSBkxXq
OEGxN/GVYvjWxMQxX3cGEx7grgU27fpHQGuJq3KrmX2AkkF7agqaDgxTEwrTGtzJ
0dRAeXHj6jYKW06x8PRJfgPwvWs/G2UiLfGhiN7Au7X3k/BZYpT6g2NEhdEsf6VV
cNeUtLSWnCAziYrSIXEmqEBzVaCrZhoNLwRxl14TZsDfWVeEzbCvqQdz1EjzmaAd
sKq0Z9MNZnySWZRMnstN4ci0G1O/lz33sFs+YdB2Czr3exsWMyHKWq4eu3WZdYlb
rCutFyGnMj2F2lgfGKYFDADpx7J4UP+BXREzjjydehLr3leXLXyJq784FqC8whoP
6HkEdVw3iy1258dJgeD4Qj9diFBgvNh3du9+X/7xME4t2EFFSOPXe+4Slmm1hxlY
TAFFTnIbEECiiX0+nNjx021Cof93a/lOtRInl651KoaCFutucsXC2E1Y1/kCd9bS
mmGI45XnnWeKxCUdSUckf1EezDbm2SSm2ZhXRhKkvW/GqaG5d5ol9wZ7wX90Ty60
3g7HhL4IAjx8gGgmpPPI0wV2BWUEpcZ0QsLhH0rFrGw5q7X6hiT941XoXXZGapUW
HriD3QrpAcvn/uPwteIeTBhquNqspxgOWL21IZRlDSil012853Au5x1Ym9uB236a
W1OTvO4PfzyPm25V59GRgFYB4lS9xUW96GHOamffc1A3NxbBFK5xtfK884UaoLac
RDRAsK4TH+ER61Py7OTPg96wwIvy+azRo+KiJfx8V7aaAwffd4vMy97HM6RuJDT+
F6HvGA0XsiGqEg9Y1XXIO2aBrsAkyM5b6jRoW/3bxCm6HckvsnJB95K5ed+CtArb
k908BOE5AAmQWUl/H64N87GTM2Owzkndq13Ky7sUEdDmpEIEnSn81PTp81LmzTvm
0xwxMsiBV8dhipHyI4ERq3UDdOBYUp2ZRV3pYomhQ9VhE5C4VwXK2yt1jyJYYwg3
Vy7gQ3qXjVN85LR7alyisnwRUXzOZimM13OexnCaP7YsDdVEJSJyvVjgny7jkf3Z
yQimWs0KuAwGExxo1XUSYUUj8MoUbNAYYYvEVKgzJMfvRvN46WnnZO/i7fpyl5wG
O2jgjNiMHGJwcPlRs3fVuTqC2Z7rLwNs/AcEUpn/1ZXAUWUiO+0KHxPX/d1s/JFg
B0QHksGngBwKMZC6ROAzNLghDuUsX/ovatE2tLfft5JDz439NCBMYq2dek2nLoG5
ycil50qr2H4ntOUM5QenNmGrdA7uwU8UBn2PhZVmVmSh/5sDdu41fkb4FsdbbsOn
3J1ecjjKBKAf2mXjj9PTDe84HL2KBs8xQy2oft2ZHbvI7MjOWa/BVw0JGeSz0S2M
VYCHstQ4EjwZ/Fdzaq54m5k+iHw/bVN4eKnYHf4mxXvuQxz1GcC/SKDEBYiXDUAK
5LlDj0o848swo6RLsoQfcD5h3tvW8OAyZ4q0G8OY4RnRwZ0YDNx02JI4cbMmANYy
V5r/PfGvBErHjwcNbqvn2rhFBs3+KCwYVaUQqFuABcAg7x43vUaTVf9R1XUqC0mt
wjOsyc0RWI7ufRGfmO7bpvyCuTHPdeCLczAxyezXJR8GY02Z4mSL3RHwKDqcYWuF
QQMehs5q2B4mdpdFQNloPUCBuRYeHpu0rPCBLTY4yDIuVaF+LZOqDVpNjE6v8PhF
Xp+ETnqF4ggn69McZq1OgjjFJ6SR+tL4yiKWH/jTJgRZy+ZUUE3ieUrtKLD8SN2B
0IHRMjQrYNK8puEd9EM5Cg/CkD16jOP4LDDZ0qhcJc2VTzCcvPa5O/HSlSCyJInj
yrbKVyOCZCHEIYpYHYmwp7pAw5yZhEy7W+vXyeelBE8DCXBy7RHCMw6AANjR+MSf
T0fFQLoW3En5Qw/hqBRH6VZSBNm2aeYgbAt8tY1N+2iOl7iU1MLJIWVRSqENVi/c
MAaiBJEcj6sA/baCISZqm0huOiyhU4Ozo6ocsOFgRZKyoxOi3SRGShAROIMl3d5D
OEBGd82ea+iZOmPKnGYMCxb7EhEyahlMH+SuZSuq5MVYxR8rvX4iqT0fLfI5Yoxq
A84E0GLK64lRh9vYQNf8oYIsDP0N1vJa5ldbTUrX/5U5s6SLmo/12sGMgIjokzNn
R6flGURnEdeDGKk810Bm20MQV345ZcNxtOA/6MdU3z129KWpZOP3kTUuxyMiuEtt
jZZyeaMSnqWC/82wXXYKQaBVq5hbX2449m86jnD98DN7gw5DUAbRtinSY1HNM7Xo
pGEGPnHFf9LdywYNy//pSepkhatUpBktxJM+QR98l7Dw2qQEPdxn6/s8GhxZyX+Z
kLxpr5Bnkbex3XRF/ooQamj+i+h746K6H61iHkjUjVNCz60RlyQ6vvBptVCtrHoY
shIb/Vh3QIRgzaJlDIpkorgm3iJosyuVVl//ZKzBD0RZzRv0dp6ho88PfYSWVQd/
+VP5n/EdGZ1IQce3zRQ/dHd90sgq9mIJ933A8Gw5tpKVf/F7u8nom7wMLe3T+iO4
Th87MwtlDvuxAV1oWhgb8ELB6O4ZkfoXrqvh626oGn9CjBeCdpRqK6w0+bnZk5tI
lx0bHVA0QE3sNeywTzoE9C1kohjuyj4AzBlVdylMnEqwjmStH73jHf1nmhBI1syo
ZvetG6MtvV7mVY4/82gv6P/Jn4eATct0emRrv9VY1k9otcrUOA/wgjUFP5Plsi0u
r2O9TnLsmxFJyEa4gpW16pC5L+GWfAF9kyYxcSjMbDlhVjbHLDJ9bGGoqQphB4jf
QQKRrmei1ZuSF02t6gYbxpxI3EqNnqrNl6p9nltJegzTLXHNfOT7pmngBtFUv8jo
ea8XXApbTh0hAD0GKGpbPDIotoFdV81fIMIdndFkCeNVqwsUp+5V6W77EidGr+lf
0AQEfjc0lC43qEIb1e3jmnQdacj5yLTnHBpvZYFHHgzSp3MyEAGWvG0pdIkaojII
GooFUkLc65RhanB1/2dFgsP8WX80Yk/Du7NUkl6UyeSt6OciADFfVgp7Tg7rmbPJ
D0nGkLCzxpgREhI0VL8Xwd1OcE5aag5mJlUNab/Zcw4sXTReiFF9ZtHXHtNx0y6w
fxMI5XovrvXVJHT+xT0ZixiknPVGuZbqzfx8EKN7YSwS3NqJzKOrx6ZietXT3Dfb
3Jx6u/IKIGrof2wp7tpTt5NXxDyoXJFbdI+1SjVCRmZhrEtDi+fwV5LnQZQk+LZY
MjCoXqg9h/KHEGfI6br1mN19FlLIA/I9dxyPu/T8LsxM348SjyV/zLkpoGzWvUe5
8zbHZ1L4zFyAtH7hOZIus0rCzVAXEpT5tOA9T0WZNDBd5+ykA9qPD3lPcW1CZA1u
GBXJ+GdY7rs4DmV7lAfaLoiYeXbcWdfwibaIrXF08cyx8FIOnfSWiLtvgpr80V0V
I7YlP0Yju/y1fDSkIzD5qFi03yp0/jX4KvtaajDl/LrdeMi7iMYK/ZaZP4kXGif8
SPUjQRtA38OsXRUeBXO24KSzEWwqDzSF4PYbOTsxtkjG4L42ysBn41UpDVeC43zJ
871EIZbIVp6mGsq/91NWPVLSLsHHrMC9/aFQ+DfkR3yJ5S+8SA32dswS96Xmi401
/AKYL5v2lwpsQbsQIr0hU1iMAKs3SQ0LWCLF1rkPoBrHeVXUhhWHdwdMP9VihmmW
vaxSNTtPPfDseYb2yCZd6IWQTN31m6eon8ZAEJH7kMEQIPHmkpp9B/RwFpK08beY
bXrEnbte3EHwt1pmW84MGoUN27OU2SByp9pWh/uHtty8MLuLiuWBP4fQJ0ywEm25
OWB8EORWudVCDUusFehhAVuSq/4yt43xIw+lSTLkiyfjxJZT/9ZL51oCIkL9qe45
ZvwaA+qGrs/HEewe9uQSsYUbJccPR9C9j/zlQH7mkFaRIXOkoVMVdXdpLZU28QD4
Q9aHstfGpk3HBc7od6KG1JJ2wWg3qYoVtBRUikLAj5bdhljpis/jiHV+KoAVapZ4
LPt9AP9Li5pyVi9PzjTBmsx08wa2eRyOIDx5yCD6YBEA3qDxacxF6VepaxjrAIAB
xD32Seocwn49JL3d2LkjzptyOzTJtMLfUCzmgF+uk7XvdtzyZDbD5nRBgcBglmUf
nK2vR7HT3aDbAYMb0u1e7u5WyazE6Mohqh9qNZpsV6Z9fFlIGVX6yCwsSXk/CVw5
/tZ8oTTvwuEHi2ExkkN1k+bbqRwSoXWJ51J5kM9CLFkRL5eCZkC10zVu688rEd46
ws2070/zY1y4o1ytgddqckKx/NnviNrZgx1e+kUSwkaRsG+V72Nz7Vx8tnZnNfe3
ft5x31WQh1WCDzQ9c2cZch7ltnwcGkezo9E8HwiDTPdhX38zKiYmAi5ZcO2j7WCM
yr7T5YuE7a1jMdw64nKpP5dEcQhS2WcOh04wpaBGgJD5HMYHI+znegGdwTCm/iC1
83N9lKnw1J+u16f0FcK4tOlVM8uaApHTYLOyYm1/GwvRReddkkPtbEk93ax0Wz4v
2E8lFQ3sdz8acRo3pB/SOoSpvU/Ops6vnZ/wItZ9f+B9+eqXYoAEA5ubjXtmU16s
Jk8vub+cRWpCsPLG1xY8vo+xI+jxpzdvPrC/fVb99hxwQw9vyYLY/kj4W1CHhPY+
zNixKBAZ98tU+PUj5cy7fOPZcs5H27WOvbW/V9+SCenUpzyhtqozEs+VwfAMX9d4
VaeIqK1c6x9Ld3k5oAwQYC04sGSYMVaxREK2al7U4O4vxHf8dVtEoenKnzAlVVRC
5pWBzqw0CpbzV/jcngftYVxP++RC07un3OChdS/DYkq+agJ7HXbD2wt7Aw8SbONj
78gvz1YbkFpNTzR8lQi/Hg5f/wFNN0i7RiBExljXwB0aHVnFO2p6NXLWtw6AtVX6
QSJak1LZ77su02aqqUfLVj6VfO4KC7y3yWV65xf8k7XT1tm7fT7/EyBYYp9DFDT5
0CQfXbJvfJF+EF0zpyYrhW2ztz9dU62EBU0MvCjoypxmE83d0i/a6Vw6Tu6S7Ckk
AM8GHke5kdi8NvQBOBBHwFYocGTMNR26/oMWZ+c4G8p51lpCShardz+nrULDZJt6
RFxI+Wnx2T95umXkxgKZ3L+CFaBnVh06reQFaQbaJ/1d+CduOUXorRJtZNaRK74A
ecZdJ0y1R83VixCqnjLNT3pWRVVMVDqyrqO5itfPlpauzSFxe8qmE4kuyexe9Epq
z/XQIdzS9Bkwvko12ShXWHiFiI7zuGpPyXBSm+5UH5AKwSrtz3ikDbKbNKC8hR62
x/fTkR5pPtsfb0JNpKlgTCatZlszkA0cy/00FnOWiOTCj1bFeY8Nxsn/RrJSaqvH
jxnvMYpd2+V+SyqN0Vvmw6XRqL6cJAkdlMCd/Eqo4NfvP1QuV0b41/8zLDXsojVV
3RARAr42RV0HUE+iEGoATCFtGNC83LRFhLLyxuQswL2NI/ajyVCEEXqz5MOa8B5x
qJ3lYAuyaAO3x3PS38QF8YNBcUhY8xXlvQ8LU0dQJYwllniKPQfmpirSd//3TRcK
csw3qo0rtpBmQwi8iCKzO9RESbuhQVlOLMod2p+xHMMpcLDEv4sO2fxBmq7PXOM/
k8zFLspgtjoOiIMZMSo+BVPgnKyzL1/6OtGdR1v53ncAXHm8cX9T3J6geuSE/UCp
ABN1HxiHe370bnbnLeuYudV4g691z2YY+Gr4Yyf68oDIpuLuSbXtZYF8g3FDnhI3
5knmcad03a4CErosrk8nDZvfjWskp9ONOdlXwVhBUrGCbgWSfa2KBWZS9aRdUErP
8XkW8nog/YFAKKH+dScyESbIRubeu32sCJJOOZm1Uj4hKp1XrcSOuJ1BF4R+i8D8
10uSuGt6HtKmskvYWy2FJgE1rzwsD/t0TfrFr0cFAHgW+LOIYXYnMHIqUhgYZ33T
RIMrT8BxpvIM/cXqiFW6F32UgzBgeAuCAixMOASHb11WDIX1K+Egw1eT9IJO4KdV
0tQzq1FmKpEfhs2P9cSEPGpKieROABuLgXDgeYRgkkfxcxQZADfxAFEO72W+p+Ba
HIm8BUujxuZKfNiPvCIkOZxcdRfTPKCwRpnUN54IoIy7AdxAfEwuTN97H3a94KJg
200Zh9fArt00vqmXL0//lkFhfaIWpZ46h24Zlg2DPHaW4NzJUId6yxkOgOdQ/uMR
7POaNQV9otQB3UlmXWkf07zvxJ1L2y80c6vO8OZswC/YuKeCc9IgSZDiTJMeRu6T
sP+1q0StxUAXvz+4vuER/XtPfXyFgYNbAxoQ08uW3CMsTX8R3SgZa7J6JPyaFzu3
iGn1aUikbsfd82+QD+cVHlv330sW1d4NUEutAqQ0TYoNH+z64OEP5zKhX2QeOTd7
kLcnSQ260jCrkf82DTvPd1OuAMeJu0x7wmH8XJoyOb9Z0aoeTLnU4zQl/wjJ5wHm
ovDLEVdwtxKd7nmucigG4w6AqF5XtrHyabYUXl8AoH/mmJlsoYzLf8QKbTsUOF5/
L5eDyw+gGJQzU7QR4e9cxWWv6E0UJ2DBh99P1COVddIbAg8ZrNZLnXN13XezJd13
HjYi8YuyWrOgdDwaUYYlt0TYNM4Orh3dp/vNQ92ENmikWzR31X7G3M0e6kHYWfmH
wFZNTyGz1cZT0eVqiX/P/D2wF/1RirK4BUPVKmB151/iIoiXpR6MoHOdQhf2bqSJ
Ucayt9gWwJXG91VAFQDbbMi7lFqnN5WkF24StQG5IW+sQLwoX3VhjIQuIBy9uz8p
lSw+JL+EVEVfhHVG5ozTSEuH9yTohAfXavGmJgV8/tvOyOBRUNj8g9Jt3bs4nPz/
Tz3ZmfYQ8EfVkVO+VFM48CmoDv2CLNxx6N3ov6qgTQshpeugBbZc0Uc6c0rwPI2N
krwZPrGcnRl43yz6il3l6CXs++74lcFLbvH7hWdxaBMNVsNfxOfFHlkMZD1vl4lj
Kx22yPwZ5p4V+Y1I/lRpaKKJHYCiocIIGs152pdZM8/QGxiFxD4crLFk3yLH6ZJg
ZopmXbIX7uFjv02hbkI9PiZ1ey+hkefX0ZW29QyrwdTzubSGXXV9TUj/+7MafjbS
yBXHrQvvLLDpW2+TMBiGCAfPGmCXHVOmR8nS66x4YzMyB6CqEf5XMuaeiLZG3VT7
iW4hBMi5heqg/m/v4O8FYIIgyDlC8GzfkALmod1HsFWLHHlCvZLmCInPHhpx+rP5
JHY2B8kJqc+pq8E9kdGR6ULiU49tTYn/alPSsMP8zbjmSw9ztu2dfQlRQtZXnUVX
1SiwQhztnqUdfpaFaxza9P7kgThNw3PdEh3Gg98LLx2TUyyJHGgCFPsJF/jk5d8O
u5Tk2GMTrC1WzobLfSBLFpVKVhBnHawoPymi8PG/pmh9HpJwpKp1ifLDAYsLf9NL
WrjYLgDN/zA+DklYFT8OtG988BdHOVRw6ZFliEmEFJaIg6zXReJzC1JDwesH1FLV
u6//PVboF9jNPXEsJcqN364oGIxssvkN2f2fXslluWv+wfCUumCXrIMfP0gFjVd9
fnw2tBqZaRnudwK4r5XnpPjBVtTKEwrgazUMTZ3Jil72BHMuuDDc6H6DdxOocKWL
9Sz1JOtqgaX3zY3HYsOmjLnLnPRppR3u8npX56adG1ljeEpErV+6J2HFdBaAI89n
qaM3ffGVtzi/zCnb/WtnIzLiWbStmQJ61J4BJEQzJYjFzpkmaQzC7ravqHzNSv0d
RymFbTtxQX9nDkOGwGcl35QPe7MtQznD4BKgr7TwUCMaP/GH+VHJu7Llig0UApg8
aU15SkWxydStwzm+FBQA3OtpHLEALlTkOn8/7sRunIWFiITSAuwtm/0yTz9IkQ75
vOqQUqvYmXYj8yY/8vLWlNCZ9yGvvzCLgC4FmuHYv6ZYX9js2/a7hjn2hOFlUxGB
DwoXCV2+/fwDsplplqA2O1Dzxg0Z9pr6hXCjaaMiu04iTGoC1/uSJadPcpxOugK9
iS35+Qze4WpE0Wj0+ghB5vkPdH7938VwbGrMwnzoii2ELSYcr7fKgIQ71b5nCZt8
CqSx39XaDchn1ixZswzOcjVf9QMHKSpdbMViCut5DgJXoS7r+DdGqZ0x/6nme/63
e03aGcsSWFMS9ZXPSzNHmJadGwQlTyZ46/qXykZwtEGIH8A/69E1cld6YXu/I+XK
wpaCrJEHaqDdCkOOdoGojYtE+D6QMJLflTFVsRcUQ6Jx/hcEroaaAa7Y372JTPH3
Y0OU4PpUIGz7HK0zL2CYTP5/RtlNethOWmYcM8maTXPdgjv44lI8bO+ibN7Jdk52
5b5WTyQ7fi+q4HTNtv8eJTtfYdvsCIR2rBUShnDkgQ0gncO6mTwDyHBzZg7RsTVr
Oee2Jm069sDVadxNemEVcczAh0avsk5Wp2X9yit5cMcOdIe8ktMIPLRwrIwaYyle
Pk6Tr/CNhWa5SxdUuVtNVzuLCkfHQSTShXg+gg3Ku6070w2aJiuCB83/8KQEQ5mg
rug1e00JDkyX4yyh8+Eot3bJfAzyXeqlARYIyvb2mC4BgVAA68IVYJg8JTsaDnyX
Q8KwjYY+7/L1nyGjzionN1tLhxdUPh0dMLBmzM/NS1Wd8hdgA0SEcvSyxMUJYR58
1hpy/6r7j4sISUSd+Dl1iinTPg0BK7m2M7Vbmz62LaD6sF1skzUgjo60XRf7olaI
1FtDGfq+CNftgrr9XgCFiTAphEqLgZ2Db9eRNbt3BH6rFEsvHE4y5joSylmE76SX
lSzg2IOdsqrBKy1mKbIW1Vcz32mB0rqGc/N+WNzSxIsXNBlZP0jabOCaTBfjNAGb
DN9POhrpAY9J/u5WUVK3uXEuhDlzeJrlgQ/WIAKpSR0kO8N5xaWZSyoVQQG9ixUH
OOEQiVkN2gsMMuqkeqO8Mt/Hlx7o1nal84hx52oFZ0u5XDx6yAVdZpkJsEtDc027
f0IHou3ryNE2Ip92T9gJypHdshYim38CvwDZGjDeiu2vF6cDIY4/+E1iTLNDg+Le
/EwEyQ93PpuXbJmpmpSMCEU10ZFo6wOiE85qIExXlMiGdEWte9EyYtoDNV9BYm2F
DRp41WYTAx0rUpJX3Lo2G1F6hqpeu1LKEXEqr+0fnfMYrv3y2Oo8iqqhigzDypID
/m3qWZUuhpgeC001VpTMX3il+p3LioDWAz7hdFR0f60dl/sjE2sOma9bUXobMFTr
hEyBN4wHErPJ5RuXh0qtYmXnuUn8PWKqUIU16zv+goESFBpj6wos+blSgVPwkSTg
mzN8NqroVLFDdGJDpN1zzybbnrVR/EjCmOwcBaJ1NYkHLh/T7QBq4ww2nG1jTM+Q
iD4H4aDZ+9CP9LsaQxR2KNvf0LqXgU6dHuMi6cqFtxrIQB0oExsAd5gJRqrVBtZ2
Jf8JuUjWM46/idbZ/1jBviU7XEx4qZpfj0hreiNwlIa1ec7Gp3kWTZSIK6KAA7FH
FyrIXDVZK16HPezFwMlO6NUNFzbPtY73wpIrSWCkW8QrNUiCORuVUtUjVZ477+Wn
bJ2unQqytCVUSIoor97KdmORlfvz16swIw+87zlvLawO6F8Jq44eykTTIQQfCV7M
ZX3j/bn1RjJI6GFxyszN+qUnkmtndMY/K1SdPIzLy5KXpW5Oup56/0MNZdzvwTw+
2iQHMUlGGoAYGS6jnOcjkdInwbGM/6qwX5UtnXDI7RnElxkeCc4Op6j47uvdiXfn
RpTA4mfAEXvjz11c8Dq7fuEDoeG/8BLSUoOKJx0NdFcd3iDGu+kErr+jmDhhhs6X
jVzJlhneTjeXgzMUiSWmRgjW/estD/65FQnWFsoNqRYNojkWKPpA425ZEuecUsGX
RFlfJ5aZXwL9RN+Bej2m5cINX4SVhvYGy8aVIJpW50U81eb2qVNWmOL46QtyCjX+
Me9xxokUz/TCmTjlZEXgmjLK/TNpcby9ReRV9n5r1VFHcnt2wYqo+QEAlgWtSQw0
70DRTjbFQZVRUcxEg1OQNvulAg/tTpvdE89w0O9U2cUelt6qzvvR6OGaX19tHW1s
5sJOOzKggrn8xRexddWzxluFVCRW6oD2xafwOmmb7h7qaeqh07RwBAonDfYr40A8
PJp3dWSAEXcEeT6TRR4aCKD2FHBQG0QNkL3Vmb6jwsTDeu6FfUahIU+CHn1OWlMR
Y+BaiIhOOIkF4vX12HxOgMG1oQS4g+mwQ9G3tIwmArfrNZVW9Qjim4dSG6ZmcevN
eMX1ohVz8CSgRZ1s7fggF5Yuvgbr7Fun3ydidfWBJ4ogjB7v5TL7YZDGCrqSSkEY
l9//uDVGu/Hmx/XEOSeEi4xf2KR5BbU/qF6/00+FAL6GQa5Oz3R8Wu/G6X2y9Bhp
att/hLUpFga6uoLhSnTXCfCZg1h3cl+tHUkBB/fpYO0T5A2V/Vh4Tt6PxANPyuHc
8Wds4foqwXDSXJScqSeyNfXfWhV4sPzXt5cjILa1hTSdrsW+JPCvR4wbl1T7D5cI
gGYRkgyFhuUflpdkBHy+/Tvt7ZO96dOzBg+xnMzb/A7lOfgr9kurkkYnVorIh8eD
ntqWPz7ZitJpn2x590ldlVOmm50e3fMRvelQi9G+/w/4NPUJPweY5XZ59w9s+2/O
oROtQF/96hq250o8BFUy4vxBz9eqZt6gS4yKmviOCmP7MgGIVClDrloH3nnHOzJ0
5cqZ1jA5KgJPR0qKHKMfCGEoESLBnISDmr72z7LB5OkLW3s8sNLVmPrnSlMsNwQQ
yZ2hBi0Q18Ig2fI+2pCeKE9sZnz0JnT8nijdrvgjNlK8p6dUTD+Tn7NkxEWHClrF
WS3FHLkjP1YpOF0ittFi0q62/1+8r4rCW2f5+CTTnQ9cKlJVPzhqJJS3C/x9hmmn
pGSG1ypBdXu2unwzjslwPDLRJzZw/tzie2I0euTg/xoKkZXU9X3LYOMjhMXiYjwV
LSyJJT30T0mJp8blFN56NcfRaoMV2nRh8LpfCVZgVaRrGDpqOcobwbcMS6krjiik
aEUey1yJKdyvcWN8LE0qCWmoZYte5+kaDvqurPOcPzsp8NNhf+OQFTkRfsbwUGSB
MiOiUiqi1Q59PxSzm84T70TuPF6mOlsgl5HBVCZ7rEJxTUgWRI4sY7JoJ/odwAJZ
WLIiP7MrKglq8GBHIMrJD9jUG/Z4NitudzvqpWqnV3fCoqOJ1ZtbJnts34bXbz2u
fAW0orQgj21Vkzuz+5jKRh2VQ1O+PqosTPP1/FfggRWaAKRDiH3P/+iJIrm7XZa5
DcQGZafUhflw28GbnVurD5u5Hjb6BTEnWNtI+XIsdvScWo4jxP1dZtrrRBH6K30s
9p+aFa1ala9UxvA+TjbOfqMl6weqx7aV4ezSfSFBRp/9+LRUov7i6MdSM7hAxe/5
cQYO7KR+PueBCi16jO+5L8U/nnS9feIwcAEms1Jb9bN/hEWb7zuNoMhSFQpzFvOU
0SRr3Wv+T0rfepoOq+585TTRDJF+Ve3WLxLhMsw6p86hl49LfbabRFFBg3hy/f2/
4Mf9M53bYTKqTY0yldgC7nLKTZWrxFAv57YOJWZSF+1LTzInGK8u+zswtIiY5vB5
TpRuGrfjUJm0P5uUzavK+x3vU4wucpxcBLd3QxVBH3U915BaDvBGxMM50yaB3CcJ
KhziujDoCMGsIlbyizqr/mZtFmoSr3yU2HFMxNsW3UlFVHTTnzlu8eQmVYvwqUxA
w4Em+EB+x3Z8G3L5k/NARwId6oO1QgZA7U0OlKsiZ6vxQPmukJXr1OQY3r2Kplxk
FiOaAmBGi0q1ESARabIQJDvucGm34c2dxztZjjkKay0l/+QKw9eHyDhLGABeAzb0
zycLTmMOmP7kAyx1iSF26kc3Wo+TvrX6nZtblT1oUI7W5/gs5w4yXh0IFjPgESkY
f8t5eURGxWrOx3874XENkiCTSniTXUTsgYCJkAOVY9Om2zo20hOoQD7x2XK3gNSz
8NlNbFM3ibWqa4Qrzb3XIJmqhDO6sbOx31dN8gcTpUhGfgs/g6wI6wf7obCMn0lJ
b96yib3a/xi7UJQPheM6+5LQoHqO44PSBbsgZvZF6TYP0GtLvbQg083cIfaXaS1z
450QugkS21bpBZn9Z74HrpAVaBGno9VUCFFxHuCkK1KWw08TrKZJE+vq0a/mhbF+
Ix+KJs+ZqBlSTsfG6a7TSreFEqz8KFHGwBoobj7H+N/CLYT6poMPqrOi9fgDze03
tRFVs48OJMDXqgtQ71eH3f/6c3BuNffRXuz4Y5rNkqrIz52vGVDkSm5RUXfrW4Xp
YonDVXK18pLEQq+iCjgWMtzOsDpRQi+IBWv8PLLSaXAkB6W6D3arBq8DG+CMdRGw
0g0st5/lezdXOo3GOQ4astQHTwRWMnOoPlOSEuWlvVnRqpoxvj5Z0PgWf2hISqxM
8agkaxDdRKLjulve602SnBHWw/RkPTMzpoSzuG4Z3hlSNT5A0E7a3jypeXXU8yb7
47PsW9LOwCtPE/JupsMWwQJUshtfk4ptA4X7GfoFI0G16uU0ZnZHhefBU/4SQ3n0
N53XmGngoqHhk+e+ZClM52i8cgQlw8btIGxW22875xv8mEPARG1FINrQDOQeidcg
UrGzaoo150TLmg2A9NJnYaMRAw6vnyiWdPHbOWNVAUK6p4xVRDSNzeFDLrV4Ngtq
iooNiv3mlVSBpCU/87I0F7MUsgUhKmXqpHfc9IAnfGXnRABDwsIQeoLwoFBe0HdQ
5+6Nz2kkq5+ibBwTW1Ukn0bJ+hIgpRLTr27yefYp3O5yWi9kzFM8pWHKYxhO7Rxq
2gPAMHeSmB8/sWWxPzgKk1i4HKLs7zXVDAsBBoLA1jIU8by/7bvrtZq69mkaoTuc
15+nDF1rB0kWhn4QMM4QM1mBw9qaGro8yVo5wFi6820KM5De4FPEgUDduIFnWReO
M0OBR/YsC+jrGlTAXWywN/0weyskmhk76Wpk2Vm8Nyjb0DapfnQaMyaM4rqRhQSz
NBmuFWzCyQIUZlBFrAX+pkNlQL8Nr1nGP5VWOFEf2kpvgwvyTX+TXASzd4SCnN4g
1/MOwBtOibbo7LppktCgxUr4IIcoXoXjH4QCf76DsUZ4saTKrrHHVmdZcc8EwcOx
AFDj7EzE9hlKVW3ZIjcvvdayCSlArIrKQGIlYovoOJGoCKY6Yy4/Tr6zp3RB1N2o
GB62irRccIa1pDTjHaqcG+Rfy5gUYeLpUC3quqTKPDYKJeJm0t4aMX1/0LEnz1Ub
Pe7cf1tDaxJH/BvTb/C+/+8wzGh6IvTsiPmWuaWY2fCSZ+TxyNzrqchcBi1hBYzt
yhUea1lDtylLq4PtZQlQergIUA25SQR2c8OIHFzrSvsJhM2C2NPmJCtEH4BOZLb0
9KWgrpQJyak3H/54CRAvUbD7Zbq8hINfn2weBn5xELdJICPeyrH4ddU6SbX7QtgI
G2UOBRbpXbaay63wC25lNBwJGxbwL1i/n8ZnqDkL2SJRAjkVyaD9VVMT0WTqlNnd
/qm4AaEEqnFguFmnIS4t/cQlwNeDFu8TFjtdzpvE4jjwdSF0Cx99CiqxdJ3o/YX0
N1YOrviR+WGIpfrQm00lVZzWCIIacs2t4MIhbSGLuGjrgcr4+TGkFdpzqgLdGLT+
l4dVLkBQ0GjcJ1E+IWreuimIaZEFgvJS6GkzinADS809GbyiVx12afUuHCkhz8M1
PUjf/S1tifos3WcW4MLWM5hGL0QbkXSguVE1nxKrQhcFrJogB9ZhVdfzUwMi/hy9
zGEc5aj+PW55NfpFvMSNIKAEddFKToVstK2zdF7MZIFX3n+0aCBYqQjk47RzrEZH
7wGs53gI+TUk8nmxpO+fh2YfODBiS7sxPj0UG4o6FmaHRHefHtsNrIusrc4aErHH
1CzpACb1Of9YSVmnysctsZTvU7zQrBLckVqxDYPqao/2usLiK76yztBYg5ezXWjT
aPogh6wDhyZ/XiHLHGmODVXWpv4RtoQ3cZYeEFgXqQ9SdG7V7nQRpLdVmlYl0A+o
a8+XRZXCb3rcIqyMP0d5YGQ3gDbo0/qjHq54m3X4cdyAclDKmhP0QLiWI8ALe2IK
wo6kX/w235dSMk9eWhwiUzIhllhgAuw10KXfnDvPzMngTnmDr7AMbbIbvz57W7FM
3/u0eO7yajqoHzpaIwXPIQJ4JItaeoqpt2zQbbdmjfY6hGGmIltuc5yf7c2GjD+T
CRgkvd5fpyO4TfDJ+6C0JEq72H85wbBgc8axgXeGt2g/JLI1QLc60YJ5f6LYbzCA
eEY7GhK/f39V4PCoshi/iB4W5lLCMu6LpFMnkIuVdDW5DTM6/gxGtflz96mqBs3r
BSIUOqGMNTtPx0s3NltqEbqsX/HO9zqS4ogS7FSZC5gNA4U/hSwTAml3RPmbWtA2
ulMVFWd3rMND7jTHIBOGXf0BAen+nNS5bA6iOqsb9cjFzdqc9nMZeWWwQCCK706s
WJuBPdRs6VOo5gwQQQtGB7nhF1TM1tVGLO9Gip2Bt/50mZdTIGPGs+nz+X6J/CqR
MBKFEMu0xgb5rqaHrbo7wVh0mSBfKpoJFtZQF3wWKogetEejQDhQ4iyaxYav40Af
iJ5ltc0udHDRyhvhni19g4jSh839v1tIKq42npJ0TQ5vnlO6sf5VFvKlNDdrItRK
i2KgyqS+ZXHSj/kiKqW+ooKZc3DXmaV2EOoZNx9Zh2xxPqfcJb4PnXwy7ptXlUVS
6AUUF9O04W58jiRdbSTXtaKE4kdFDL0STEIX0Ui//aktQcnfESWGxkDrfOKqG3PR
W8uco/c7adEjF6eIKnejNnU4931I+NW0zdTcceyoFZrzh91ZFjG7Gq9Tsc+RN/+/
+lTjtEqu7972J2qzFNsnXFIZnYD487AxxScz/CXcteMI5uMI36TeIYzSeoL+uKrl
ayoIb5jzQIm2VZBBe79mGijh/30wmJIiQoqrGE0932PGPntwPQjEw18OFV62rQTa
ax37E3j/kjwgMjOxCXOIlhHt/DR1UeOBSk/dsWTuSxol21XJnEiqFGDn5LP/XFek
ZvKRiMQXV1RQr1sDcMze/vkz9pPYEz+vHhikdvs+UxFQ1xiRVY5n0XfslLmNJ6B4
NwbLTyAu6EYcisZO2Cgbi//zbHL3QNtNPNg09PaX3qHxiNZnAL45vp8Xn89LV/y3
+bAmT9DbNccclR9TSuEGBLESlT3wYTI5WO/SkB7MAVEiMaA2CDlytVcQyQfMyeIt
tFKbjyp99Dy/K7jnxoUWTuqe/uftn/Ju2mG2bIJG1pBnitgOOUvDxTjn/oNXg3LA
EkjkeH0Xrjhqzt8Uhy7Wd2l0JHTtzqjpAD3Uia9iEIuYpsAV9+tyfeD7vprhN6UL
/dVChMxBA/MLa9NpkxmwqL+R5Y4/PlUCUPkwG4LfuD9MF8aljY/acxafpWIJfQ+G
4WtTseG+YqI73/d4JWqDnTcaCCl5yK0LuiAFp2B4zmWNJPhNayh4nsl3lnJuoR2Q
HerbZChJMs3H7bZgo+OSa+pi09u0EnVSO3R9x5I9XLMJciqH1DTnQhCgJDrvGVD2
vlflue960eoMKimBmP4XOXhWZ9SaNOGDlu1/+HJey7HG5560wXd3sVgFrXDvmRv4
acQ3Ck7MP/ME0lOE80DE+JBm+Pw0dL9VsJsGCrDwvZe71bh4kdPpKQXXo1xdEfUz
5DNgGN9Usp2H44uRD2NQlCScRzeQWRujX3H1urVnSfUmjfBffcxMuiN2rHL/x4l+
i/nOE6Va+kJF2TZx3rgvhVtk14GauCoTmUAG4aJu+OvlA0HjORZS7k1HGZ0L/Ad+
DPi+9GA+aVFpJ2Z1eUI/Aaf+Zj8e4vH2c5PPkxqkGw4C1cKonTWZrufnFkk3Ihp+
SSuUBwo0UwQ1Xqog6p+o5ayviTbFgrH/MyIhdvKcTeoQuDl1s9sj17IzvW9HT9QM
nWbuGL7vz44D/Tyb9S/HhsCLPVYELjk0/j0mBauWLJHFncgJFd+6mIoavde0xvgj
OpB6k4Ag0+gbkvBXniLfn/mkBituaTDimf8usWp7Fz9xHiF826xgjVAHluiLRtLj
d2RRwwqc+lEmdUQgPB6OkEDJGgvJCxcd/q82DhuLSFknd7IkOISIxNuZgBwT/tzs
Xcp6kgLxFmyvq+zx0JZCSRe5PHavtqj074Mn04CCIpRrrYlxSDfQJf/oICbXJ2Vn
UWG3L/knkNY/fOmK4IrURxD/2Pnqk3FiYk4Nxu3qlqFWWtHu8C+HB8gdSgTOuhs0
CEJReYn8CgJClpEs9K1sBZ9FWWY3uhDap5rkZmQeOpEIjTzrN8LbJH9eqdkIcLDh
eqD6TJh8ybsBJqxTLuRrgyU5yn9hCuToRbT4iOpRqoGomuwUIGsEE0uMUK/NVsoq
hqrJ3ZD6PmqzDbXln8qnY+ZmTWejX3oGb+R2rrhzBbQDKBM+MinzT0Qa4bqxIwwk
y5AT3IvuvWHn026TK3ZEAeQO0vfdDd6p1/fwobqxrgaDYZhRZbmZGHALdX3Jpgca
gcfl+CL3QGb4aMDJRHOrOA7pZMyf33IHZAyPHdo6g2pxUollWYB6w+H4qeyV6+m5
Fl1BxnlYzChq9keSz4tdpP2TwGw0/N5SYD2e//gaYsxA1Q73SafgpD6F+cvHK7C7
UZN1YmgIVuxdmjFTVyoRK9fEc2iXg0JavOxno2erBmxDDmeL24wV3IySKzJLohYP
oTkEn/WGish3Etdy/gZvSZnp1aHES4SZ1ZUUL4DyVtHRrow4AdEbdMTTa208/mCw
giv+g6rdG55UQqruTECi6dIBcOsKA4BfLkcSffMDpQ+dg0iXTQvYJbZcCSdT5gUO
GZXFEgJmJnvuALIuROlRv1fWL4/VfY5nJZTf7y1BXiiZHF+Q/F9itWC9V+194XPe
UkW80iBJuImyicWqhYqh6fvPA539jj3DZ9r3HGk8e7pJ74wb+9cuOiBprvkBl6fy
6uesnetDJxtvcvok6tecw6/0tFb8geDbb8+T/Qf5+eR/X4wrRhVSVSanvx4ggwfK
xuZRG60HENcsZs0RIqhddr4YgFLz7DAPsnEGoRtDFTuLYK9xVGXxPT72vmkf6VD2
KnBP86s52bMA4vONEEykE8EBfMcfm3SZ8KQcqaGkyITuT2DkskuirAw+sNp5rUWD
Zy/FTclq5lgRNYnCtc75XfZX1qkl2xrFqZCassHU8qQdZPavFKOsEF+oVz91FETS
ggfl5p3DMACKaKez0SWXh8aN6Y8VZBq3pwSuR1iF0Y1l74rBZKzDtOViXBPX8p28
IwT47av731t8QgKfeMdOqR3ARQZ/uJy2A/3wvx9UVSUFRSvwPgI4dv8wGZaVfB3J
pQV4EuJ0/TRg8T8/CeK1HkWdRIGxrFrc1HJwyakZ8OvY4+WnUCP0SCJUJAL5RF+R
ZoVH2NnILnSaWUtJ2Vc8JmhbmtbP1Y+6e2GduGjmcl0xaLYZAVxxxKhlfuUUqyKb
VaaZcnYf4U0sR0HRp+yHqcCZnZdV4mWWVBFlt6nUUVC1GW7CPLrC2eh6KE+BhGg6
Hi7fmMu2sdwOzohEC7NrEzthm7VEiot0ihWqQwVfeCkb2DDKK0Y/Q1LHMJ4slkQj
e0snk23w0hyYN0NEz+6Lhv+REYBxqgIZy29HS+FS6/Ex8O10JUccSNY1490ee7EE
smirlDNpQQn4WJ2jc9YnPYt3uDBHk2o2zi56Di0okq05ZHDbH4wY50d5gTvkEffw
QXWDXtsPdlW5BhT3OuoHYYHgN46yXS+O1VQKis6qlVMbwmZExIa605ay2rQVqYHv
Tgwm/EgKaF1FKe+0BlfjGouvyghS8wkbvhxpRRmrwBPjG6Jrk8DfTP2WPxsnK6FQ
POGhTf9atjraOMugB6mGr06pip90OFzfFavp2ZAXjtfgjwgpNJTmHaekVavFlkXr
ToStNAekXtBxtXzH9xtadxcCBRYwAlbTk5urutVm0tvTePM++UyKSrLNO0qgLSXt
cs6HG3OHA5e5cMmW2CRtdrTGOilrgUWfE9+ZyFWj34dKvpV1e8zk9kTBHK/sefjr
I9fHPZ4oVPloUIn3mURChTVW0r5GKlmaC2u/Qh1REWRMehqJBafgg4kEKObdHM1T
/PGiFtSZdzvLfwQYjwgTnFCOm41/WqB+lM5o3WrU8BjiqpQRg6XrVijMASYTT5zt
ETaDTvWRPnNiB0+iiuNIE3XVvGN2xesWFNAh9WdpRNBqpDMPQy9dUPAOtozaEtIS
Lfboqa9HRu0E7xX/2/cYxguLG/RBVEXp7HSIHLqCAPrT2djJy85rCFEu5EydDd71
homlB5ifCnbPFQ1zleZP4gMFVMYPqxhOcDAvDZOG4ZVbr51+5z7akz4xZhBdipna
npFrKeO8m/vwSAynxBwE+VnSQ5EnT+IqxlcmMBwPcKFr+FtaEhY8Re9nSgCjk/DT
1qc0nSVIduXZaE08745o1KWfyyw04IKuAn6+nDbdnlLov/oz9YjaTVgkOQepZO+n
Yazh1QlQiFcwS92hjig5DAmIY4aAZ7x9AHbXt60sI2G5TXsUwEyKLMfPGEWaUaxE
zScbqswk0q7W4fC2piVtDRFVe0dxUu8qUiVsOL9GCyIOIxkIS1/SGyT+kn+Czeri
PURr4o8hE7Fd24nPhdv2/TWLwsCCpq/zoEzNVbsQ0EfsDv5ofJMGLqXZiQAxzv5c
jZDcX2IOwwGs670Ky7QxOF0tHBkdVNAKrpX8jMOTOBLEFEC7+Kq6m/ni966T3WvM
YuxtyuUM3Mdo3629Si4xBZvlkSOUxImY/ncuPku6i/ThM2W4SpV1q9j/xgx87ZFk
WVN6T+JD8sK2QqeEUcwAlLgly2cprLpzRD49H18LUYOP9w4U1pBC3gbEKqhlWVUX
wA8td8SuNohdpD4Zm9dPAN7wO0vGw0FK9t+2/wsLwbbdE8AUGLiM7xXVtu8cO0WO
4ZdGw0FYuHUXirGmxTXNLylx4bJfQ187hgOM3px2OFD60qt6VIyAmWoEoseVr81x
DIxXxd05P+5J1CgDoL46tAPTH439V73mAoqcm2cf37nXUcnbchynR0Eu31hctfWc
I5Tlvavs3PJPZF7MlEDZ353AzWA6HS2pJTZ1hQ5xXeSFjY+spWbEVP9z89YuUcyC
wBuMIjLe62tw+bhBJcqRKisx9s2w9/yDF+OOL/Jj9UMYXbetp49lGCP+7PEhrDJl
oS+k+VWWtdzgSNnkQAEuUmXd0jfQnQD7ZZOMSgh8TuDNNtzVUeGf1RuEZNwm1hla
BqV7GeFqTt4RwaGsc3iBB+hVecFosm/+T98WsI8qJ0BpAPNaTOgUmEMLRsjGzPMl
nGvvKHnx5NxTwScFmQKbcKqRL1CEWsv6y9wJd3xWm0Fl+r8T5PcrsS0OaouOfWK8
ETdKUJp/ZnJfqIje4dc+YJXEsmxlrkoq3+Hct4zi0KJMny869ohlBbKr97RefQPY
KIv8gK6ArRvJz+u8dcf/i08j82KMy06WfK2VRdLcMq9KhoXv4DuhiJf8LcnReOC8
2MZKXDx75R8gk4R+ggOPAuvf1GesQZAmyFlJjerkBxoNVRlz5gP9PfSup76o86f6
L+HuVDMDE1qseIW/IArT7lzPaXTtKUuhHIeQOZPGMDGyUx/BBeR56s8wmkNxA0MC
kZ5D5q9Mh/ilvGnylpCZWzilrpdRKIO42hC/34kGo1iPGK9MrlYexwO7/nVYASTZ
l9K3HqTbTvxew+WYtMgsEi1VYQxA2zSNv/khc51hZY9Ig6/B2nzrF2RPZuv0mgNT
6ZAR5ZghFgjmlVZ1s4efEoZBUh7EpKYaFCGLJtR0YlwVFpuId2gdYpO1qyuH7pVg
EIPOU8jyF/SQiZBuJiH6vvRSMooDWez+xu4XJGs8O6D7624n8hKros8fYk0ZVBC8
0c64AyMz2666jEiGKClwvMEImVjHOaoj/QnaIN5aHxEiuUESfJhzHC/w1hjC7LIa
JNCeN3JlROKcxsk+YK2rYv0pytvSuuDe7B/nzhbJl1rbAxc1IBGxFhNyfAqDNfEu
4BIjrqgBfN5W9BfFoCCwPe3ia/nm6JlZBcMawjP1I91ZfvenOZdqaqKtqsPfFNWB
kXzilMTlGgwr0zyJ/jbCd6QvKYEhI+2hjcZO49nQsrf+N8UDFW+qHJVLwRdfLXFW
tYAwPm1xCaUDDEWVMdbIshVwGQz2/roeKDjDQtFEjMOAE9tyHVd/xE6vZPX1PdIb
KgTQ6/D72yaDbQi9m1yl+CokyEPvgDwqMPMTT/VVTNc4YBnWnCdPiyX2PCrhQiR7
FlZZ56rSQ0tco1FTc0UN2MDKi5FXBJJEZSTYtbN+BOeT9Y9RR7JusVLcRddlI74M
ouvsDbAb0CJUdRCOtF6KXOFzUBHODe4cD6IpoRXU6r6BbqexHFfc95VfPBWltOBS
bOOyNu9y31xJa1cpxS+3O6xPC3rDbAfqX7WPepKAVVA6TVlPXFjbdLpTcG6rJfC1
TrlIdZwVH8OehIvAJ4tgwS0GBn3LUYA8InE5i/52Bjjk7SQmZRDUKiQWnOyHjEAh
098U0Mdmvefmh/fRcV3JhLNnLr/ZE/qo2RWSsTzViMaATSHLbu9btrOd9NwTbDLI
/MB5t9s0KYf1YbNBOExH1rTuBiqClqwfd+KCrDry9+cfdap1nvyANCaTipDpM0yN
bbyeJy/PybDUxuHEEDdOj1ge8bej78+BxVY95gJ/RLWahM4KtFgVHqmdQ+XSt4vG
hlhEfnBN74RFlRHPY/Pkcp0velsURcpXhT1CoapMVvmNdYzXGJeNmlVAtbsTHQyp
bNaX0Pm3BWsbJiZUERvEuwC3Je6RAZkA99BoUJLYV4oJncgfkN5m1ZNEK2BPqwvb
btN7pUvjvyFeGeq0IwpbO+IkqqwaIU+J/flsp2pxeyGvDyxl190HO8nzxeMI4du7
nxray6kv4wmb7N0q5wV6AMaGhh/jWAkFb5NctAcpUHy7HDHsLL+X6Nol394RQZQK
7hgxtAAuj2h1wZmf5qWFn2peHf6O6JsbynOUMeBrNQC4cM10VWLHTXCJl/lPJG54
oTb8B2v5o+P3O9d1BOp90mE/yPjALqZF5NB0pNdzlbq0iMF19tGnuxrZ1DpEQMvu
0nBil2LcIVxig7852+htKhe7dmencFifOyIQ1nMaTZmWW3ozg4Sw3AYz44P1UW+4
T6vDqmAxcRni/EqarCJXAa/yOsPbpqYbF1djMtiUxe962HP/vhmXNPZc6X95f8BN
OUk6KKv9ivmJzBor8DF4tDuzowLxDqhN+KFz3wwGZztvS6hLdF76IvaygXLqIO3d
451r1qKZr1wsSZOWTpgA7m/6nJYEdtA7QITPrDq/R9swA/KOXWgZEYo7cFUj4jtj
TJgWJjxj3vTmcGmA94C6RiNeI+rAUq+/91yIC4cbfNM4HTZ1c1GIqvot5hhT9A3l
tU+yXelaVMXurKXcDNUOroUHBjdbObwZmCAze6neg84c5WIqaKZvwXIlGpdETm3S
u3Zjcx49Xk8dCr+v3IBL6I3C9LS2oaSX8K/XG0V7kKip5rEnZPr+KG+fsgMEF052
tYMbr4pOEIQ3CKcPsptGhQBY56fk7xae/5vVSsdOiXCaYfKZi9VwddhIqVs48mGG
EpL46pqYQYdKBH1IAFSP/MBkJnfxKRcp7YcWMY32eVfogRHBXlcdsGxTQ1HylxJX
UB1KmMZpfGHLAlMCOsq/V1zFn17DwI4ry+UMp3JorbEhHEszkPwI2L71qcNuxjcH
rDiIZvSOgRbFszYXzPpTtFWa1iWrFCBOfskUxFzJdpq/mx2gQNjZkhQD4VvsLLlJ
/8B2OiAvL397o3kH4KC1xBaelKH4mLWiN5iPYnbONh9qKqX2B5fOo+1gCiqtHMlt
pqwKoU1FotlJVipXvE6dNV04aC7slWbzFaNMKh6xvJg10gbtqMAcyaLEXiO1pEzU
3o2fQOY3O6lNvRZohCLZ84l9P4ivHxadUZ3ir5Ku1rYxtjD/IwLbpNlGXQ9l4ue6
5UPKGgcs/atKrWUsKqZX9vuu1Rnc5Rs5a7rDlqr8pUJ6LXcU3YdB8tRTzpT0QixU
ztDpOa9v3ki2FmNnmLHZUimXuPM9M1Y5oYI+dIHZLGiaEmfN6F3O41nqcBkBdRyF
SypZjfKqTyBc17XO3wfPE4TqcwAVfr+RgBeRI17UggmSaYeuGdADZtzdnCV8nh2x
uBj4Si9MjqqXV8soiTmmTRuNx1FiZlZjgshijiuHnJzdeinl4ZJe9bTrEMSHCpDw
hsGxQtKK91gO9w5EJF4uzyOAbfu+jTla1/d24JLUHcKUcnZkXU1gV7tdUedQt2EA
QcnXfSksBmCGEOL+EBUhm8/SyNfYGSybdOvw7ZLinLbSKwaabS1dyUIYdAYqe61V
5+UZuEGwWA0UnUZlvy5imjdNFeUokk9wsLUMNA0aX+z0aAtp1BzvAfmMndv7/RcW
dBWgs+0L39FCCkNhZBpKR7s0pxChqxdfQ4o2H1Cx7k5DNX/eoKNCYIQOYhmMrOmH
FG389O1Uzd5iJL8d6JKIJbp1jtDQvFq8Z6rSOHEcRWJCyGyop3B1bVEqglinag5L
RmWL2CJUT5G9wp/0B0qidyMwmVKJ0mkmWnGyT2xvCSwell2XT/GWk+kM0tU2VH0F
wnXLuicpIV9qks9QJm1LFxQBM2sKHWlQwV8X3Exa68F1n7KYSWt6z1m5cHf4Y/6L
hqPYhCqPOqTt/7t3TSaNdwYaK31zQPt3uJo/ZBzkKhhUtFNc3Lyvvv3gyKSpUFZG
nQoD0B82/TKthTASPyT2opAmtfRPld7v2GMfANT9ybZPQsV0/ufPGlx82aOq8uvw
wnlBgtS/+AUf8fEiS1WZewYYExr2VjfL/6q2mR7YC9EsmNyyPHnxpSLwcJuDdJV7
XH2kBmGZFwL70psLSDagoKbDGvHlfN8DyLQI9G5bSECgYgoAwHgHQKRx64vepxoN
PT8XRNHNM0//Cxfc64LU5ovXYzZyVsOlf/wTwOFS3gg7vithvXc1t6jGDbDTHrPA
9XjpoiFwDwVcFjuG/hD0lrDxS6wjn9n1T3nGvv93+SVnNca+o5ueWD3An5XFakVW
xCJOttcbeDR+9Jc0/zXAHCWlpqcrmvxcwS8U67IAHA5elNjAqPwIR4plD9BxcUYa
kLwhPelQOoBS9qrvLlm14Tsraz7HFiiphax7Gn9g7W7kUS1vU7QsZ2fj+Zv9tt0G
eQpp4aeWu3xd7fgWBFXGYmduY+EAjINyC1gVV182/yZc2NWGjXNB+uIsU07DQX/L
nL3xYs2BKvSNkpJPNP0JO3oSy/sFVBPVM9ZdANNpS5UjZwxLYKfqHFbcR29tCYDK
dWWIJLLXgLlWAPsv3u0KCwEhdx162KpkNSXIs7frQauPhZXR4XDzcuAixonqj+0K
6x7BnwgFDiW/AylDDxghnoSMjZmOFrE8neaglcwkajWtZL0uQ5Uyf0tuX9caAkWI
9oz1KDdhx41ZoxN6ehMz2QV5BeOR7mUtoay1v5a6qxUFOf7jYE5/wjG4O0l/Dl9H
Q8zdwB/AN136dzVWgKh9MpJO1f58eqnZKxCyY4vCzfOFIQqSGvttPRxvVWYhnUpx
toHOqyftk8KZux+DlOT3+Uwd2v3+0/zIilVNuMjmctKL0PDgs3ILUaEKSkVYTuRy
PWUo9NpUqvUjDrEHux8f/W5qfa4ptLPO3vSytKm1gEcFlh8Vn7rIgJmz6AUkm8Xm
zDHxxQ1lIDE43KKx64TZUfkt3sQOUhFhMuZDvLX0tv2EBKOJqjyrKq/EKWZvt5f3
HTPpMFKe3RjCu9iN+xsUIjvhGnteCsK/LG1Lb+MxcBJSl4efAQzm3+d8pRZceaJ6
04MperJN/RvVf5tAeGHfqVgbcYhfzFdSwNsxdeXm1fPPMurPFiYNsHlpOqeRKN7z
H+HzYZQcv0nqQZEPURzolaB8I2bRugArjw/u1t3j8xZ0788CeC58EW1yeQeoUBIs
NyIjMZyRtnykzfQiRGLYPfFEouiNRQ56MjU0he986EYF58a3z5qAFGKCn/z+CnoE
5QyhTqZ8liM+bOpmWywwjCDt4mjqE28GWsPJ4/Eqi3H3laulnM3EMkdiqmLeW0a1
7V57JSRVbF1dG0lDI4hXYNSd5pemXNkwWUU6EgZhZkLRewkjYgW5rlueqq1VMv0/
ThaCvZffXh+UjMrTRv287VfjNKZRU3MwjnfzvY8+vCCyaHf5wBGY6rlqAG/u+ZT5
ryIbWTSiZTwpdSkB0OzzFHXJdnZLMoDOFLIhIKtbX1TwNHlymRxeBLseOKO+e2wj
I3F7XJDl8Xa3jxjpfLejnZimWBQ7SwbBiXW18G1hbYIEkg+ksnPS8QZGm56xuIal
H99AaSDteOJEgLuRtecindV3CyVVVukYrTq+LqV0KKXcwtPAa/3WuIs1aXHhTJvy
i+AiXtEVPsDFgVUrzY+rqBhm//PdZr4VqU7RC/yHOilQvwCAVWIG1ISjmz3Be9nU
1ieOIIiB3fciIjRILmhLemVf1f74XACMmL0Ox8wr9LPVUMHWHUAAwiTbsud4gQ0z
XF7bkI/cx4aU4d/9zJ+77+1mv3eIx0rQgj9TJdK7MrvuxYeAWtgC/WzsSwgEmW7l
tmVBusJpduUFNmb0t+wkpp1OpgA86MZz57mXJQd7ImurTN5eF+eJPUrP1t7HQ3xl
JRYD9cvWSiL4pLP0u+jIg3ejS3Z46abnWheTg1xx+ucO/TiKF1vSfHypt18efU85
biCVrfC0Sgh/wB8n0PLCnqZ9u31TMUhEf03EbUXQnY+zuS6yeAiSDMyhLsR5tOUb
oqLR4XC8nzOmFP9C5Vw4L2WpGg5uYtx1W63TLNZ6yu8Exe2jDvES4B/Na+H+ED/c
5Wi3X9GsKceDP4BY54aJMNyHM6Emk/cYAJQ813uu19iQAtOouzIVvc1fRgfqEcUt
oqLPSQO1B1n4fj01pnEjBWZzozsDP6CPfFsHWolWNs5rE1iNgJK5zioYdoBF5yNT
VxEQRQDrf2FFhLCusfIVKVZJcWsuIthptuwmUbLYLUqzWK6c+SHzN+baoeTEOXWM
7pZuzu36YS0UbZVkCyC5bayfDNsv5YOhFyzF6wN7oE0Qm+/kpJZTbwiKWPizQEjx
/4kGTU72ZJ/DHVYAV1GQeaNQ9PZl5vCkLVuJO/JQ1JUsXfxxSj8zp9iE3arEK2cf
TvX87FuRXWbFACN4KK8PT2fOpUGUdKld0XYI6hEbRFxxC/4E81pV4YcUNJQfUlJs
/6+syh+7jfT4WUD6fIbaKDlFcqY5QMxK6cimrNA0c9aIMNt0Hh0T47u/pvKCVb3Z
NYWAYfp2XkejErRYyqRXihSaOWQ6jBMzX1WU3DsDzfsRjxuXCqwm8c+AVQ0S5L/C
djUu5TleEHhJTOefrQGWrhhencJN1c+krGtvpJm4e0TILVIqrFrUj3yMiEnyQEtu
yzq4fxCgUqZTCpv0er+MQu/DzWmftBzwS31LE9gLrjTnx3ComwMSJlLnJ+jpIihx
jPtlm7Y2XMWNB1ff35rpXRd652XNpd/NRreXKYtkCqqVI0DKzV2irn7ibtmGo279
uADqLU+YjioKN6VBqk3tinGJSGF7TdkzVGdXaicGvP85N/EMgGlSpF+nPe+KJ4nx
CQmYhCpLA3wpWlBzQufFN/FlWgt2eELO883wgAUitG5jkxDrFEVKL7NV1KAV7V+7
EmzIQI27ueovGS1Nckidwr4f3cpJNhwsxQbGF7mvvytpA067x9NsrbnHAnpqYKvx
7AyqdbfKx0yngTrLuUnH5r+khhhI7BIX1/9qupqKKQp2f7ZYL65mfxGKLJdXitDK
B/G3f6EqGJFE7C6CA0QjyaiMewlkNaFtRgzqHpFB4Qlh5nUvPrFIIQQOZOlMAN+t
f77xkfpyaIB9o0Ff027qT8n0dyfRwiZj404TxGZ9i/Uho8yOGS3KevyZuO4p+xdT
YklcD6e1Oy5yuf1PBUbXIoR7ExbiWY/hrlLOAdcgCT8x8pcyU4EtHMo/mHeWCXi9
5WVTHTipUtCAiC6GVW/TkLDszlGqg92vcEcQZS5tFuwnqlV9+EAC3j0kaPBiup16
o5yJLDOqj0RZSmtQlU4tMrd7XztsT4zz/cZ8HJWiSb29Ux73QeVWM+Os9oef9jv8
Sx4mFjkcav8nVpuPsbxa3a5mM15gez+vJa5sGRx6u+tTJCMdpaPeGHyPhsZhIebx
epYZ/ja6QR5FSKy/gSPYmutki49xTM794KSg9qp7gaBjV3bi9LafLZciuII8OumT
teIHyXFl0bU/MWlKTAGdpnO5/1mHa+YbuVB98mVQQcfCC6trzRGhrCHe5/ttxWkn
szBzkQnDO9xdTTA+qWM+oXK+igZG2PQIeqQ00XTQ1iOcVozYc1mi13IZdhPHUDRP
Q1dnr6mGGyHUONVz5IJJHWvY0RVakW/K3O1EezaD0+v1J0HBZhGms0WYvV1kVtEo
oudxN2ivec/vEvdakldj8jFUoSnRaJY/bTRp1Hl8dEGSgA6g1/KuaAPTalAE5DrS
ENez/SCKKcPMtq7lEUaHK1I83K1MLayouxI00sjBB3hQefkZUdH8+17Ds9D4Jja8
hZ2/51lilK5sv+Km+z1GyyH74KE8a5jkZW3JITKjY1Ou1gDzSs33mvEW5+y0xwDT
aD3g8dvNXfjVwvZdDxvpzhL5yagFR1f0npDkgSG5GZBbVOZl1GdUN22LP+/vcVpp
m+/r2nCIRcwlAVTuwh9EWiMoLnbZE1MM68G+AcAS36AyWaOYeQ8Dk0Ad7CLnnjOu
4NE26IwPwMp6bfEI1LURwYBKgwCmRDnpcKgFVCiYA9RMyS6ZJ7jEOl0ng0NgfRaT
C0z6/y2GFT1hfEY0GtcRMN29xb3D50VDoe00tEyQgXJKnuhG/JBErTAkgml82zPf
KPv6ZZlJyjEAz5krcxruyK9v9wdfirbvcFeTBPUNW3SwZ+hamQGR6NSbXr5Mg+VJ
KNSkC7CAaIfZhfAcWpmU2BrgHVrfnMgdnpt3dZJ9+s7R95rhzY46i8I7pnWDO6Pv
Rhv3B5iN9c9o0NmVWJ4c7fWu7pZTatL27W7dvFGQJMLvdnyr8YJhpAN0uUcOhyIR
056LGzOUAWJtXoH+I/qy4vfHaBeDOXMdTt6+TUq8QqpKtgPOHe6XSZHu/MjP+RDn
GM5Zot+XHAbvjZWG+KzJx71YyqBmGWVZV0+siMLQxvz8yvnT5ZpVZuO7HkLzQY4T
B6dPyybHaJiZcn7uTbzYyivBC45gpwnypM4+1GUbgw8MjTaoGZHxzFxcKZ5A2gza
vXvfjNxggoGiRAWBdpMmHutxfK7xyavwyvOF2mcR1hF5KITb73Gc09YWDFpryEQI
/9bqcJRlQiXbefm1d8X7jlzYpf3Qa0DUhVJ6mC/jJZu2vK+Is7TDeBnuODrKhpuU
M8VjwnAB8c9j0Hr6PSVgpWT+W8KC0AHn/KxJk0ECf1uuMr5rWPlMLhE9xmRrCTSi
+uTurV3sDYVQ5GAyDHAYlG7OzWfKCyJfeFlc+nmv1xvkz3VPKJS5WwOY5C81+P9g
0osEaQN8sDcQMehxqpgCTOmALaAKt6hMIgP5ymtR++wtKI9RITwD9ephpS4xUbYJ
pXRhwBb5Dm2Y2Vk7MK8tvsc/x1NSWAVuWvnul+YorXLGOHKly8kMgwl+kEde9WCU
k9THqwlvjMOeEn9KX4qcjgeaV7p5zDTMhquN/ducnXvoP/GmPi60FzOid3rF52Xw
jE85ktRq3z2UNCQNh4YfLTC0crziHLauAFy9MWbx2P36pJKGMk09gymvAJ4y6S7Y
iUZ3SdJf+8BcVxaqBepk8nEwc14IFF1ynpghPCsNfIZD42VqpKndLTcnEwZTmrys
loTiS947gY8I8JCI0AtqXTk2Kz61ntRqHK7PqUcLkqO1uFcl9spOIww4PjBS5h6E
Ytio27r/8/YVGAqmNeYx0Wvb+61zENiST1Kx04+4zfMrfVUUvSALOx/slPf5Z0yF
9Yw7mTOJVgOmm3euu/dyPYyKTmRywURVApn4eE3/PbZHrPuGuLRlsUwnD7ewOsTg
zu3sV+WbeZzKX+si4qHK60UqEkzpvVKfEgKK+P+5hxrOriJfweIQ8u0wnl5nnSME
jDNLl7EKIblL0mN0bRVkvI8W+CPQNgq+Be7G80k4LwNBxphVf21Y59e+WLvEPd3u
SzGkZ6FL2KFvGCUo1PnoUenuMioRSt9t6gmpkCFaAa8nTEGnX6c9TuPfXsydHD0f
pOwV23hK4WRPo02g2kAd8j43nvPr929ucQZHvjc5Gh5f42KnsFFz3xvGgOG9e0Wf
zG4xxGWFrBqrXcNgmfqpxWKgiXV2YM3j6x8ka/DHgzyzBn7G++uZ4kRp9yxNOLEJ
hH0lSt/IXnMEpM9HJsRXtaWY9/+bNZX6+frypcKo3espnKOnxcHix5b4GDXzvIac
UMeMpv8roaQ6WTg8qbTaEXnel3IdLbBoxl1hIA0l52b3LE+uc3nd1ISWHeLjgebz
xy6XwJgxElqfKPwkKiFoTAkkCL8+hHrAt0giPwHOL6Alit9XJI1qTv884xNP4LAe
EJMuE6odZ6jbx4Umm5OhbgbnVQnhSyW4khBLAIvvXxl56m8rVSX3YKsUXCj53RcF
IfzkH+rH9jW9+U2sRq/bjOCX5Ef8phUeZgcX0iybqb1/LLQeRjPRtKHEYd+QYVnQ
XaBmRilDrWtw8KNMeroJ6t1RohXNjhzchC+nw9D8aUGvB0hTNBJpbWk7eiQpZWku
ZVJv1Exo1GDWC1XcqX90S5dfkUKR7ynf3LEnZKug/ZGlT538kAlh+7kxltQLt/p/
ELTh4mTMEjxY0QFJh2OrTrk/KuVO1TeRMTMuCVxHlUhqROr4S0bRxJ+7DmX6vMv+
xP1+xrg1/gKh1PTbYEC3pEv0/WmWBhjPRVV3roHBQznOKx57eu62CRWqNPhduHmR
cFD8UXM+O63gK5Fb9quMmw==
`protect END_PROTECTED
