`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9g7UnZqWzUfydhOOjgyQBIOPJo6Hb+6GfIbKtlmB92Pugww8jKTCrcKBB8xhTNae
ZVCPLoRiabMfNcenBbL9BQq/SIjujsthYPH+fJ7Wv+NQXSq/YM7Hi36s94JdrXi7
9BxfohedHjVG+Je/Ftgouh99GMnwQBdlFHW7B8g4RG9LJ9GkqpfK43scSbmu4L7Z
z1iO0gab3goOTumBs9VDPqcDB6wH08hU+vO44rj7INA+tXUvZZ/LeSPHo2gEHdd2
bXGLd60575p2B8gPcQmbTpts4AKJIAL8ahTe4ppLwQSptnuwvTuy2Xiiv6jgzUJt
g0M5rAZeznVuarxWheOXgA==
`protect END_PROTECTED
