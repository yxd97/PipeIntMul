`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mt6tKW2y4Wf/3dGxqWFOlsf//Kt6uTl+9M4ZURbrsES3HSaOqVlEHyvPgH9MzEln
7oNYO2s32pk95txWgg+GhJ7c3FL9f+aC+Irggd8UllR/2adJZr4iC5ru7qcENs10
1MO92Y0FmAzBg+ClTGjyWn8qUxJoJ9Ta6r1yaPVu8C7CqXxoDXFIe3fn2tHb02Mq
PMiR79izvjh1xueWDzDu1/FC+ja/nNPHnCHY79FsJ54z8n09oJ6OJWEq1HN2xnND
7BlVDH6KJKSypmavASNjfhsK3s0B9QVwDVQ+6ng7r9XNzxnAUZFaSm+2XC149hpu
C6/SsGzTHSZPhuYWu7djdGcbTGGmIuDB1/TVPN3IGSzR6DeGThY51U2QX8+9stWV
dB+w+8Dtbza9YSGuJGep6EHFrlydSbDJH7cf7dPUkdL2O+O8fE6egpn0BKLjJ4nr
VbDOhqGNaAHGKfahA0BeergdoPNPoKVw5FoRHzOcNG3++hcC3Fa6twjV6BJ6rrIv
zTF1v9rUAMYXu9c3dC+t/lDD85+EbaaOAuO9EfyL855B9xl4W6XLOuNJErCBuJWI
qJ91Ba8h5rx80QeoBWMcJCZJgpIjSzgw1eReeVKBjpDR605IzJxjQ4PpKVCO9jaM
`protect END_PROTECTED
