library verilog;
use verilog.vl_types.all;
entity OBUF_LVCMOS15_F_6 is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end OBUF_LVCMOS15_F_6;
