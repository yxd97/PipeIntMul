`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hcad4aN3ULASiA2ut9gFYmRDfFNTvhccI7cuBRw+CL5LELAThJgPQxuW0o+z3B2m
gCJ2gv7KHLwm6xF4AWzL1ziKjP19uJ0eH8nW90oIAmRSIUBbAaIGZlsw4n9f7LfU
W17D9dTZw9SJFhEl6dF9LLLG3OXZaMI7jrqnOAApZZ6Q2UBir4X0z8dJSJb5IsCA
1docXmHMeR1GSLD3RjhMeM75E9oV87wLrPwpom0aG1VzVwSTs9S4cIEQN1R6dGq4
wIpo4KbSjzgxVFBTYMrv2pyMynujltF2KTSQDxAxQTiIdce5v5D9Y2lQyHJGQpuT
/hupBjFyjvocybvc/bXdylgGfWXeElD74ofkgRnzbEA3jY/eaqPG+QnAgORsMoLr
ihbbZyPnES+5CAIhvBO8/tMx7uyvNpmX63xDlcU0k+E=
`protect END_PROTECTED
