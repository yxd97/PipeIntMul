`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9D74TJWGGF7p/bFkEG261OlOwWVa++VpVsz0a32Xwrehqp42d6JxEAXB5dRx+hV
mfoELxCe84KOGCq/wOgSS67vXQhoN/UqeHjmNJH26zosipDyzGV6R9vaC+q18z5o
18mVMOQ1QYNtgVKt7r+eHYjLFRyhsjuA6qQgfYU1My5JojaDRHufDKrRXmOHYTGZ
NnN4eTbFEYr1Mr6ysnhdpA7AXv8rlXt2/aPZc+noEAzeb5DRpsKKHhRuRMPtrHdw
9LdObWGJYmbqdahCb3lad6sfx8qgMU7HyWOfbQPbW1/o/ROZ+mvSC24lsV1RPCr0
35RW93yW+hBtTQAZOjIIwd0JoXMXc6R3ceWtYVU53d15UOz6NCBM9QT7Uh3qsqYT
xe+9gdja3rTZO4jZ2L6P3nkIDch014HNTn96wckYFoqwJ0M9N268HQp2cw+RBdpe
jrX7IMUnUbdpfZ6T4zzWn1Qwz+jFRWsa2nudHaG8rjM7Eh/xXg6mQ4kL7XYTsDfN
hAmIUXkTq58O55mhY4d+kRH1a2Vokz4wpR7ypuPl8kTKtcqUeU22LThB0acOkc7x
dFnqIbyqvZJgiT7PxvLXLMotRTPlwLIBjz2OoO0zW9ddmYdAFR9BDjIbeQ+ivKMk
L8V/SfdVT4w7fVADxHA8mg==
`protect END_PROTECTED
