`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hDs4jljjz26Qh/RwTfDQmg4BvJADRgvi+GWk0kMBcsKe1hYA00AGJdw/JC9xh+g3
iDlQ73jGu85pJZkRH/EzgAb1AMPqTwRECL+fx0RZDUxihogw3tCGO5gMwlawOLzu
ZdQ3vi6yX+XCjsJu5/wfFcc++TNNXHG/0drgkVnp+VQ1S37WNVxeuH+daRDSjtbF
ex8yXJS1/WUOXFJ00NOofs5f2pGzC2Rjs0kVZFQiFaG0DGuVf2JjDY14ESWHfEIW
83iLCpOMR/ifzuhRdoJRHWyLawTkvZR5WK3RGuMuwmYrx33QIXjD91nwcQT7YDIz
hf1aJXM45rf37D0Ot4BF/U5r3O9qFHlK7bGIsUvnGGY6znS1CZ1O5zmPdT6NFWDL
deeYOvEcfcQNgwrlQRcVs0/DncrpXI1TOMp72dxaLYM1gHMZkvt9vR0KHdmiTU57
Pc1vFUyKosKAJpBe0AS+fl94tQdooAHC0h6pvuIXGTGaOnKyu1fCNMnCoNRNPETm
jyCEygPpuHUMQKzni6KpETswzEyn+6b+zQfDSFeOcL2PywX37JRr+h3MMFyVTkbn
F5WQ0DpF2to2zhN7T5RVkAy4elJqGYgjmWaX07BZAJ82WW4qUywHbeUKVunBSmCW
3hUu6bYnO+sFxG+yyxkAx6Q71AnLmXpUvbICNodZxG4zhuARb/E1yOv6y8TiXCZe
rverBS+4LyyYID3DPcSFRzretV1pfYfjHXceC0gmHh7ikSTwc+Z481ThWYce0J6y
Ry5Cty62+S/c9IOL0b3AlZH73WuVs3dwfvwbeOSxzIndpc1+Ly5aksJIbcGOmJ4K
eX+OESbDA/LITF3D9udRo8TwkJj7zct/ZfvIk0z4iFsg9NnMsiaQY4N7nzpacoiK
D04CliOLBJZaX+yh5WENfATLX/uot1RfPJb4w0ESCvir2+h7tvgpJUqxmZgHFMf1
/VopR1GkyHPIgD7mMMeF/5fSUSHzXJR1UZNxfcsqrshEwvJ9SBFK+ycgh1M737Fc
oLW3N8pj7EaUqoAdpduqaBGOWArTb0JxQCKlf5i1Mx9Q8l2Ca4oLhAmG3xw1fahI
k46PKYAiNcdCvZWqodF01H6D2+dYH9EJGzwG1KBasxeY772IWkSiyV3pOfesqagg
LZT8MKLVMsbV7N1YXTxg4GYKJEaF9vD6UXRjDqmcwCEFCztXQpEj+pPiyFU2X3Dg
/gnTdhGYT01NCZyUJOIlp18NSV3bUgydvK+Dox/6ln+K8b1HFLIDZYqofkiqutjO
TUlCLBAyJhzpEoCncyQtdK+02HyC0Ec+NJpN6Y19dgI57fKNJoFIM2WT83SdFmaE
Ql9icg2BNUraAHo8wwkV5jd+0NM8KzAAfXgVfwvtOBlQh7rhNtZ1F+/1Jme/HZuI
XRnzbv6MDHCiNVCL3RN+9SAQjly5+jSHGDSZzPqYVCG8JFNnkIWiwg5bR3og6gH8
/1ZHNzMlF4oejg+2imYgLjqYVZfWW22tFU01xQ7MuQDKJVUNpc0rcbibIIpxOKKk
gRbaddib3uVFEZZNiEq6m+jqYtUAZkB8dxLy9mo5hatMtgAA9FtAEq7VsITYKYgd
Q1qMOQY/+q+hlo0J6I0tcDdHb5Znlvj3g3Cw5IeOrK0YQpfSrrdaHbH+9BxRLZYx
cV92Fhf7OdbCslsTSAsDWODfMY4IUy9KAX8hs3yIvB5eoZ3TNbI0EE6+5CY5Lkyz
Bv/5gC9P7cSdEVZs1Ig33XqPawHe8mEesdO3JZfOXcvVof7vCtYEBNj+SdwqzDst
HVbQ4HfX/7vKSlqbqEfon9gb90zbnQx4q5YpDJamSweV8DASd5FJ0lY83THZQQny
qhcWN6CkjDuDw8aAQ+cJehqUR/4u8USAtD+Tw5/Ao2bialoiwp1t25o0UgYhTxNm
pFSkZPAPOS2NOBIoVMy1GiZj2H962VJznNO6QSBVjMB7QpQEe637SANefDmb4bmi
9H4Rsy+u9X8Gq750+BpSrO6dXv761fLO3Tf5z32DSthMmB5mFERuYKWtP4TA0R76
Bu4gxBJlC+R+LKxFjzlnNzMHTCkWFuzMp0g92Fay1P3sdcP6SfTHgYK2kF8Ar6dL
blYRXhob7rIJnGnxQQ8tD2SV1DZMsY8TPkaWFMemRMppmVOUTq7R+KccfHeubk7u
XHtI/vsqXFGPRmBYhO/4/FJJ1PYwbvA1gsbT+ZiMQEZ9ywCUQGuKzN3+ad5LLmlW
jInmO+b/8nDbFz4zAgWHC3Rlx081TH3Khi+OvW4dmpagDE+zIUUODy02OJfTx1yD
u8+FJMW3Rxl/Uavea5dr+RIC4xHsVmWVYKLnNhaGwCM8scEdFsLnGqQNwm9VS7Ds
Nh5t2ECPZdDbUw0jvNmwjsQ7gjhwh+Yk82skY5NAIwDx5CqGVdtniojqiJqzSGBS
xgobTeWkpa5U3Y5UN1gFpcWx7nYMYwn5ut8BDo/N6K2PCzJUkoTRI4CAQyHUZ7CW
PyYk8QWhbBJukjGLyz5Mp8yfItLsick+CUVkbCOusKS7Op79Xc5A/11vbXadMas6
MmZHmONR1mm0isoF9Xg7sYJi1eDgugBeyE4w5cgGXj/SXoe0scGrDLXZKKANuDhk
drZAgrYgXqy45IjQWw88VF/TVuCCHSfYwvQlp4AujI2O389+Ljr+z/d9S4MpGwGj
rY1ekg6IrEji9yHA573Mv6gcCkZBZT2EuakIGU4AIbr/hVn/2lIH4b9/AKxaEmvt
viCG/P5h/JOz/4O01HVhg2nMO8Uz2Yh4C9g+ojplrGhxXciv/c1FwrWTki3YQ0ht
2hYVtHD50SPbg+WbBSPxDQC0CnmT2SWZ+xAXo8NdWXYk0zOUOLexb4M9Op/0KmRb
rDcGMlqS32zGrBWpBFH3bkXIzI1uOUlxrwr0tPC/wSOJxupMHQI0933u8zXoQY+u
nlvfucwm39pIRBHeF8ORSqCA+D2hLGztlIyCBzUY5F4Z5MtR06axlJOXRE1g21wT
imqoWpCV2SXiOmViHwrxWmfu4PR9+m881RLWF2Wjc5+jLlhj7uVEHqAGqojZpmwE
Njzg7w63TwCDam336E45vemJrZBiCLqaWQK0AtGCAVzGNog9rf4XtO0XU5CuhPLT
hsBEtBhER2RRky2rgFjM/hoZHuN8yQV6kyYvMZHxSXkQ6mpOCA3Zn3O8X/DNIv5x
LHBO/wq3BdzLGRymYOwUm6eLKg1+57rsPIoxOFXCqTVw6e9LotKgKz4fXpCG3Fmz
YZk5Xtd5OFEMRQysC6pwIXM/dp9ZImXI9UQj+aGaGDSeA8LgVhEZS9GqN0g1hkwx
VvtCUq4mPt2tkHYES81OuTKSoeJ55TpFQBYImqvSf5Twibw0brhvEb/Kzun4/0pU
2N5xvHMYfbmgNEVqmQslSg==
`protect END_PROTECTED
