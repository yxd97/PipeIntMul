`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3zXEU4IQibQc68o4aWgSBK9z6tBQkNv3o2JyneE1XimjsUgp29zLSVkd7fcNJBe
1mAoyRF9hn8aCy/qULVmv2/WH9BN53XyziaIRyp3HlgpqGZWXP4jgHGgU7Zmwmuu
K9otqc7TpKdyn67ChpUBWiKtt1nwf4gRoaAe+j5Jvo9uOzlSZ4EKSLTK1xlKh/vu
YOgwKhYhIRD+D7JkLkvJ7bNjPL/DBaPfwJv8xMJf4/1MzR4dRPUHqIqClx+RQ188
mgMV+ZqeA9KS2ZvN5urfG23IZas7vC8i3GKK7nIFYKfqc9GM12VzdjxSQ8kmz+3k
KiUum1xlEZVJMsgxAnfHoA==
`protect END_PROTECTED
