`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SFQlTYSuvKtSscBGpotl8XFe0Wc9HEksFGhUTtXVOA2DtZdOj2cVQlMuy+MTQLDN
DBJQ3FUBUxOv6Z1kUcjoKglGlmyHoS0Wl2YeIYSkKS/3sJ+NOrXFcS3IUu98iknd
0/JQycF4IRkxZOOY7oRBgrgWKa0rcahItfdjKjQG4OKZM2/7aY7iTBLYHC9fi6BT
6NktzYCgG4O0481cEPVNjW11AUKuPDNcbljw98wPNMkonRkQ13BXJ+GcTbhJa+zQ
FIxEl7igdq/64nP7ZrG/jj0BT7oTWhTdzsuHEfGUdve/HKQanAOEO2+dXsKnQEdi
9TOyyfmBXBNOiOjU1zUWuWaqf5DXc33yaBIDoRzSYLK+bVO0lNGSjOSdB8nU+UUw
aavbNKa1h71W9kAXcB3DMAchDzmbzzLvnuHnkta8G01JZfElYUN7CjVcl39Vk2MW
vyjp7CYUwOT2E8fc3FfCN1qg04OUfnkSbo5dq/MBGmFJLTvFWkGA5HlGgO44zyQG
+ZkBVhZ9e/0hUjLeRfaKDOMGr3n6PpwDiXTe3dtWRYQiHl+nNB+exof4RrtCxGmk
/s/iH7M0QNgiFQ8kv0aMafZxaNCA5zr6g87iUMeUWkWHuryT1T4lKMoT9gTHg1Ab
zMDW2+O/quNMO7C31Ks01RFKxekcDh5HEQgkYVWF0GOshb82bxxeH3V/vNu4weLH
5+/5vhFOXJ4pyDRaOhwM7kXsWW2SocQ4eXBhI2GEWPGv2gVLIw5ZP0VkhGnnBxTz
b+lDG5xPSgEvlEzYM1XRNq8vLz/a3YqbSTL51BDf8NCTZJ3ORIP35PNmxCm3MlRO
vORlgTHUiPGADSVUwFSXstcSCz6geiqRKxm3kIo99wqH2CGZ4gEXuFvG0G7/ue02
6D8PksLS9y5AmYGNbjKgmqs4cS7uaYPxSMEEqfSYTmUXelQsK4zNNux5yGihmqq1
zXzJxP0OGrx0ZbEj2g/EcpPWm1afRf4tj0uWkZo5Vo6mCx6WlCtybBTM7Yf9Gciu
pTzFtKBjhuYxI+p3kAeDYZnuTiQ8BF+cjonD+qfCtPy10NRy54nyp8AJ0HT22CNF
nLzgEPUEZhq/TPfd6QUhdA2nNTQDPTtK26gkoK8L8/yupLizUsG8v9TGaX4mLgJp
P9kctzdp/YToJalOwY/8U/d4NIAWgYowKW0+QVd3dcqxJQPGZHTEQ0FA+SCmpr+E
Oiii99VQVJH4bdqfi72hLvtRnUkWk8+7Hmy0gponM2xwav3X+XS5LHxZj9FHrJWM
sfd/RtaaJnvkSR6DUnRiP6XtWvQeoOR/oOb+x8foNogJeeQNj7tHslru8+5Ln/gA
b4Kyi4Nw4MR23J8oXyOOP6U3hypt9Ch0R4NmCdrGnb4AYq6eHxY33lAc2jz/GqfV
sNy0aQEHpBu9LiJrTIrn2RHByrbmb6T9qdUvkE/e5nYdIQtnw4Xdgl+wHM09vJFR
Uo0FqfH1cPAOpp2YCo6SSca1mXCos2c7XLVVRgnmTFsKPr95UDWrGSIZsVJ/As6S
2TJae/VSQ2klEaWebMZAFWeCIp6Pk7CvgJTfpGyHoeMp/WDfcm5sqeSPyMGelfP0
ECsxAHi7RYnhpWGYQ+nx1jt/u+Df0XqeUOPCkV0lbd6at2n1nbysGqX9Zq6qLHYv
kYX8S/porRx9TNE2xbkvvt83ZxqWygwa8Whi666WMdNJywm28yLpI3l0/bDQMDYr
IhXcQXMk8+9BzPvfg4vtDOIPf58L1DKr4hC10Gh2D3ncLF1H0UG7EazBQ5m8BodW
Y3Yo2cIoBwxAAV66613ZN+4W6HOe86IAhOfK3oa+PACxxQln6FjMGHt8Zsp+656K
oHTrrSNuRFJRfNwqo5cT7N8aJgIsQ/P5n2WDfGZPgho1sQbYQO4T9HeUp8JMb8um
0fg3u89P+DRyywEiaoDNv3IMQv+hRmisNM6hB4r2zZTbA1SWaFk/4q6jglrGJmVP
0u/SspC80jPvX7Liyc265H5BA2x+5D+2iPBLC1WYhVUTDg1U0tUo8pbXM2YC9L3o
Ul8WpCzFz1COhKcB94imxWwVRuQTn2r2XEyaeFNefXJY6cXMzTMqdp4sa4TQzUeK
k8SALJTjYa5QNt1X1otUKpDbs35e7irdpfA38DQYBM9BoACLZKB5itU63qzC2uqd
vanMzvpnzaZjNk70BNljHR/Gt9Kh6u25Yf3VcC20rmmixlWUCCQ81yVByxO0CxSB
wkd7yg1Ny7xYx+PGsh7MdbIAvDowL5hYm2iyueJE8k+KRKRgorjuKwV6lkQrVkPt
yk36/QYmpLSA2vmimNt06EO6gsfTnHXnFVNND4bgmYeiDkY8MLscTxE7eNMFbHA7
NuJbMD+KvXVEMJF/GipfoGEj1kdGFplv/Qe5/406f6k1ihcqghFiHEEGKPm/vgeT
XfPdKjrqEb0afRIK7AnNEY2g8jFNrz6gt9NbIM2dB16SB1iP4u+qG4ifAjqX5asQ
38jCCGBbWIISoSemUXTbiPnodfQQb5+H9q7yxoKqAUjZcyIrLquQ+cgsA/blEfDx
ea+oogjltjxqctkJD+vL43r9pxi4Ya27/I+0ODmetRq86KQo8XXqcsBUJGnIMPq2
uaoDugItZ7Zse97LgdMsLjKdVnoBaFrt8qKQXiWOlc157LxmkUGE9JtVney4D237
pwjsJuLWrtlH9ZjRZMYywImOaCxx2orM3CD9Y4jMCin9IMn6A4yc4DNJC7V/2LV0
BI/lYb7BDWbqPtmOR0xEog5fVdoVAxXka//Z69IDfxM/AOSQyMZ42ebS2mYqXA5e
wVQZYYRM5hxAvYt1gowzCu6u5E3QtSyXQsD+OE77FZFD3GQkv4peZ9u+abvzrigK
nDrxxHCtLgc3CyJTO8TZmGBddIYz0s23BtMq8btS9so0ah6H5h5kn96BdmuyYtOD
n6woystnJokN1cQG/3m7bdQtjmWf70Xl3RYDQlgS9u+8tVuDAln8tzXL3aJMk59F
c8swxSljrIV8GSnFnL7YyQ8y+DNAC3TXEStTp5OO6CJ4L6Q5jKSObUMl0ks7fO5C
1Pon8YkJ3sUB+pjbLAgrwqwTmNlw9o/sJzThMMPLYcsTeAq+I8F78EQsIlMOzsv7
ODj+a9SL1dzwcB3f9k3i4HtusRrUFYQetlwc66NGRLw9wU2R5MGoAFpanMKuPc+d
mvGAi9DDvlkqWt/JzCTBqsafB+P1RZGRQDvwjBjL9yTH+dxH2wLlzxJ7tySUBrWC
g3U5I+uP4dskPLZbhakzR5b39oDCEQbGvW8HMzkLW3uO3zxAecLjvtx3rF5rtI8o
FK7t2/Cmi5wFVinj7ae1DHHbnmXY++qW+yJ11sWsRcxvFp0r4yLXkHLUvjXwoTK+
Ed8GjLqixW6dzupRU/Oukm2N8sjn98QjTMoSsW6wDK+uvg4fXesPilxMNubxe7f2
Sigy4A6UG/yPZKmRRvdZwpcNFGZlFhD/K/NpuSRsjsbNNcck648lQESQdtl/jOZ8
esl5NI6ZAkn1zd2FLtqy0Tf6wqK9mOY+tfq3Te2EV0L+0BO6Dj0/D+vsexJvwpJi
M4L/bjPP9e/wjtGL2BK2OgjoOIc/4PMAIu76gjuE4GBzv7dF60nGccYkxmJRd0Wt
muYZonVbyLrGYLITtTOj5aOpisLVW0k2XXrbsPwHUaZefVUApudaMyjjiYKreJNe
04C4D0XAaXtQZqbmg3gbNOfihXL46/Xrb7Jxjg5AsI1xbii71spzGxwncaOq59Zr
Ed2TdU2Rq0/VGa7RjzY+/1a7G+B0MIj4oQQaHF/enMlkJq+tacD9ezy6KzkGLL8n
kITUq3M0GZVfMpGLddnYjze79+gJSV3Guxku1nqIf+X4baw5XDEWwgD0TqwJC6g6
ixLXYTbz+qzh3D5zwhll1gjqXz/3x2Crka3SfqltTSGwA6rZJm2Zts5vkbnIwJCg
tCpB0QhZku0ASpl8cR5G9a71BjvlaZ47nOgF8/Wva755m/FxrUOWmaEhFwa9P496
PRhNkHFSFendRjwe4jk2sIvC4JBVkNvUK64Rs13Js/txIzbtk254nFF5z7Yafw5l
VdUydeOmx3K59hqEpsKHdKVd4cOwp6PTzh/EmtwQjw1GPU+Moz9rImRaYfGWtzKQ
ndtPjP0tXNCzlRC/C/6DzerXO/kfv2yGuSgC1ERe9tWFdGQp8SEwQDmsDHttcs+c
JyBI1jx+A0Q929IeasIQEvzV1oprb8hQGSNRuJw6ykmB1ZEDdOIZECeec93EuWcj
odNcCk52hDnkrpSrjawx6PvS1AmCX/Vmrf5IjeNiYjndYCDCQbvJ2si4l1nPy+Xm
jNDtrys8J1WoCyaSyz7mQUhLIrjSSG8ItCoDLZLMy7LpOguqUT/einKAzTu5GxGh
QO/zDUcchzPgFxDC5IlZvdj2NaMG4ozZVYSo4N34lBYYWDQek/UJBixEpTTvR0hd
G8eO4CVeeQE9NUACb2NWXwXdD9mLtxHW22dZVYp/lYE=
`protect END_PROTECTED
