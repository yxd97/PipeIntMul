`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nTnQz8x86C86A0BbRfn3z7uhPEXeXTitYcPwHIDzgX6Kc32eAbjndiRKeGvh+kJi
v/i8AQ39Lc55Sjvde5rJ4I32Sx9iPa2bI5JWs6z+DLGWLPLtxoMvKcYqszZ2rhhQ
xUDqkNqEP0dhVH185PLTXFiOqpoW1QiB2lEc86vTS9w9ws0KG6uN53FsvegkM5IX
aMBiJ1QVLP1Nr9xBxSOzr4S+HUKwACoJvxn+OwdyyqpOKnwVKrltXS2lSKxYeWj2
THga1qgGRf96E0eUVCyhiIfosAnOGynzjqwJcqc0y6ovhzDUwBcH4m8BCHK0lBrB
hN8Mtyqwvyxun8rW6/FmJBXZNY1Xbk43zWvxQrq/IMqwrQ3PII8QFd7+ycIi/51k
D3YyejIjIprivP4CQl+NIk7EJx20KeAKf+lq1/Oh5PZjEk1GTS2isPRQu1+vOrdK
w852le2KY5YnRcS3E/71WlBshWqnVi10KfAEanfHTvDQFEePT93LHoEv9UWJRa2l
fEqdLGFnIe+bNPHCNnRCI8NmqCgQo7lJeQQHdYsSJFJnjZc/5qzTp53sLpQ28JWu
ibMPLqdMCdu0Cf3Pr9l6oMbXeYsg98GJUE4r9Ki9d2JwL4MWs3pKHxKVoF+lbbvL
bRoMxFc52uorO/npGjeHmwoof85LDc7hZaxSuKLhyXVRFl9kOHXpj1eTydOHo/p5
Fha81Id7Y2/huMQ03y2MsOTe3eduU7qx4QKr4m3bWQw5lsGjJ03X8+/Rg0p4pxB6
mdEfcShWM20hw+NEg3nmay0t2OeJsf1xg9J0x8L7LyBjk/ZS2rSTvfgmB53ns/Ws
ixA40uiT0Dk9XbM/uZScJdPKvdI6/NRDQ+KPhBhMZm8ByTadXk/2abn2/5lpp0ue
F58+IFOeYKfX6V7rPFpd/uBWqAjbvFyNGRFwajP9RBabzplcvh5kLcwmrUV6Ihp7
IWnfS0iN7jwterWpgnTbOt2LdZ0Hl5xjHapY3hXesVygPS8t08ATqlugbQZ+vqkE
we4NxQi8bFVb/6u0EnZz6OL4uBRqCJrYHjMx117nyYbyR6UZzesDEwqC17UWHb6o
oXP9o7X4KrJ/K1REia/sfcVcdFfY5RnI747T3Bibh3l+ydvHwdIReP9TzxUacCbI
k/Laj5GfnVu0ypvxqkH8UsCr37JKMZ0CjnhskPtKsFUphOP1YImYln1aTgzuiOg2
emsK2uHibABOb1494FsSxOJoLbtX6Ilc0hJ/0rIo+N8cxa92i7nHm4PVijzQQj3u
1TgwascMHgDsduO/9iGWlNOnxREA9sxWmq9Rkyfm18wtfTl7ogZo+9PyGNRUG8Ts
ve7VqL9e1hP8q1RZtwTz9ZyTp9YVaQdycR4pY6Qe2wW4UV7XKSvsm+kj1dzhS62f
LifA5mjpDRXYp2mUPFC0/M5VlHyl89vjV30K3OWmSGY2YGoJ+dZxBb/Y2n3pfcYn
ETTpboE3KnspUjT0Q2ZpjJA3w8zpD7oo9bFcNFH4LRjbLtQYFX9et5jqhdB1qtTa
yuVpjnA6sR60Ht0Y6O5jW7Kpmk+4Tsj4+WzXsIZSnQu76NP1sQ+na13TXXzfFDb1
QfEoIjGSDjFW4HLCSJU3yK/NJVuwCuhpfyBZdJIzWV28LPdvveDjOFkVN33xHhAm
A4/o5mnfdKeI/isVmUU2dph3qNPogNl+uPqD6BznSidE8Zs1HLcv81KMLXRmlkcZ
ENvYa5RFcXuMBb5XWLnzuJHi98ocWPBz/b2kRtDlXKmfRe9ANt7O6jBxpWHwgmL4
ocsUJvNaXsOXmJLDac0lBlA+ywIPDAtx4b8hxFyu7l8zUq+3JEnZYisLZNSERl0A
YGnXv9IyQ73iktojZOaEpAOXeuRaaFtQcukaU65C52lIICv7EQ/GKe6Fm3x6bvxW
HrlOtYhs7iIIQjqvCn/OdwFCmVA3Ob9NWLPCtRkd2yLD9RElmsMh0+9/GUWsT5xM
4xeR5D25ezYZtHyPSsxjsQl3pjVhJVUG0d6XzOQM+WhnaKnoQomHFvgs5r1aHo5r
sOxrW1p2mCVRub9ox3hEzuoAezcX9QfpBoJ4KIWpJbPp41Q6ZvJk5EtH9JptcVwq
/kbvIljiPmMCbouNqanzoU13IDmFamnsSOaMyLB9OQtwuEh8VEjVOTx2ezlurb6V
R4ERq4VVuA4+Tem5kuaBEegFJBGYaG1sZDCvZ7A/94sgVV4k4kX1cvP7SRLf9sUm
Ip4YqJn1864V7etnjdkOYpgnCoZc0GtegW21ZOxw4pma1KILhHkTl+A8T3UDekTA
zJYlU2TR5QKGqmw5Y0KO8Q6T4eq4wzGh6IUNWqPxYSOr9g8mPoSVq2kSHTlEAmsp
KIzPZ8sXyW+xEOBmpthDUR5zkIKeObmUcSXFf9i5CRld8awJKjWcZNdNdJz04n3F
+4r/0lOWPtTinA+rB8vxIeO/+TWcR6k7YQrdk6TjuroGzmAGiqZa8bX2+tSiO/hP
H8IeOMYGpfYKfxq8QqQg3ZLPwAhOAEZ4S0mO+VI+LkcTt83W1BLvRsOt4/8Cj7M6
Cl6kk8q1fYwv/4KTGGaC24kU2vSZbtypm5eLKAuSkbgAK+zvTofnW+1tpC+1NGGe
OtgIi+NIcfmn/l1DZn5dHHq4gbPeoF0ppbOUdZ4IZiwDVsYfipYYkYykkZbVD/RR
r6ozLE3KylvwzEdyUDgar+ReXLG2L+Wbhff0lI+CuWdS4MJtvwYADOJsgHkWHa1m
trMfD82dCWpPi0AOdj5T80O3Na7DG48flAPL45DleMj26uDH6MYlJf8P3wFcL2HG
bstOrO/sSfUY8VBtcbAvcqtC8Pr4Ckik7FRTiAB0Hd07fTooJ+xRbAmOp6xh97ZM
1RXA9YKg4GpI+8tgWZUV76mjMm+IK4Li/KYyQm5/+B+VisMWe8OhMTk2+kcYf2dc
yX4Z9CvXg7jRCGueWkPkFmW/uZ+u6HqEogSBln7K6U8+QdxFz4XcTyOz+sxUs1ux
sV4p1KkIBlI7NZijrntOe7ffb7+2XbupIkZhgUVX7dlzEs2HT60DBv0NtR5Xfi0v
9ibiIzjVxA3xpZcgrteGU4UR3RgzPW1mUAEjjPvGWExgQbMQ4WQ9gpXB4vrusZ51
yt3K75TEibIHS21YWUeAvG9M8P2cEAfWgb+YSauKntwE7faD8aJdn5jPqrFdpza3
8tVHy8zj15bLl1cCIQHJaIvfqsSpoSWU5IseQToMPlEAUW1d03eMBabeDPGGNikQ
fV+JrJ2Ka778pPouWIUcD3DeUANBBQEneij1R8brWn77a8cInuX8AeWNqhs0tsoZ
aBw5ey/rAH8CBXN6WX6a7Zi+dCfebQnqaAz3rlYnd1tUPacVQbqYT3NceBf89cXM
XFbLabJM5XTPL6bez86bjxu1LXI+xNCpzqvJLmwE2WqDReUOI75Gc5jQ3X3wRukh
72fzLMybOBwrZ1ptIzXv2in7zNQdvIqoy12ULey7ke65VKEKJWTVC8rUC/1POb6J
+msuYXOMMrmrzRZOba8LSMJhVTTdiZGwzt5OQcYVVyCd5NF8qV6ByiHTbEpxDVvB
30xYyscu4TWOM3/uzKWmFYR35v2MBPS4Pd2uHwst8d2qbfFWMr293JwgWwzZ28xT
po5y0YTFiT+L9t0U8ILZb7ZH86t4tT7ke8XH1Qgtfx2XjzHzPP7Nacy0fjFeAj6Y
5pQESCVDNQLx5PGzDI73OoNZjpFjHG8zQI+EyEqAxefqaqOPvjULNVjoE8z0jeNc
7GvQVJlwUifnAjmFtxTfDfY9rnamQ7VWhC0JGD28NeoWzly6iaQ3EUL84t+yNjWV
4z7OBujDL8C/MX+/iAyAfU96ggY07KiGMxAeJ5TzaxEz58yjGgDi3xqqgQa2brL/
whQlQKnDgZWRY5HOrzq6blzIuWR7GAEQ211VM3x+GTBt2HzLZZC/jsBwI/I5lCmY
IVDTHjuipA37PC+Sosn2QhSJdBhHLSEtjdPftjG2iEEcbU1RVZNqueM0iTAV79RG
X/B5GdmDAzhRP5tAcSzA3MmrhDnJ94DU9oR4Gxs+01DKtJHn4aBfw2AiS3Kve4Pa
r49vq3w3bIgazBblZGSVdB6H9fhOpQT87kZzHWQA/3vwV0T0wP6D4ptF/YWpzss6
RqgUm3TiKIdkBQGUyuytdt09tVWzLzE92oGeE6nCFln0zl260g5hqmKtCvQmFQRB
z6MkjivrwguCa/kSQFNdlqDwOirYxkHz2u10bzuWMMkk7HDDCWvgYkREnvBrvbXV
P1sIQ0r9JINqN5fVG2sob4Wx6FMVyS+ngRToK1FGBmaQj2gxkEpwIziRiDOrzvRV
zHV5Nx2ZBJWlS72C6pR3XEdRe9LI6WYRmiV1bfBa9KJXBUsn1QWImAzH+AJZHyNP
S0jdW2bDrp6ssGchD7iRqbzPlfS1dDZL4PLvePZBPvaKZl5Zsu47gR35imDYXW7l
8klMTKNra7VrmmtK6RHOlBsNO6qXOVg56SW98rmwLLy0xdU0wX4R/LZnQ9QVAIrl
ZYrswOu1hU20PE6t5hRZcTL0s/ebPuueuwmAIjvUYMdqtozh6UC69fmq8IoL+XYZ
hD/Sx5ruRjrEYjiZZ5eOOwDgbuNhbgFGEzcndYeKitygfEAbULqxOdhZrZX4x4Of
7DPIuFrrHU9IP4TByoIK+tx7uBv2SuDHvpMaodBAnWE9KM1Y69HfrnlfPCVwsRwe
t7nJG7G3M3XUocJgv86RMCvfnfEDERWfCg+Ych8q5oPbSPAfyEaGIP3vJ1knvlfu
tDaNNSg9QbnIMjposa7rey5b8WwirbLEBeAWroVzJ8Pu9DEUPS9l2LaIM11rS2rQ
XkpPRwDhd6fPLT61uoFWcQ==
`protect END_PROTECTED
