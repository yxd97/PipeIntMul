`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBA6APmRYSfwILM0zbTeRIFv21UhQ4cvEH1P9XdUtLapGMUrCyzTWEDIA3wlGSjJ
9QzEmFH8r5toX/NOmzhZpZYMbbGevQ2pB1Q5z13UvDiU9u5UucSp3tly5D7VjyBy
veFgcLD0SyHHf68sAmEeLd8J4wct+NWLEHTm/2VdF9nMJzfDJ0NHmDsokOQHTLxa
g/3Qq7iah3h7tJNvb01QZMQuJy+ngE5zbjRk1cWsfUtkl3Fie5wUobH5s7CCxqeN
jhvkZdl3AxcQOP6jnUDtAQu7xYnKqkXfLxRl90bIvTX/NxmIPfzgspk8JLmHZgdN
DYRaOKzbPg2gGuSTtnxLeOjFyhV5JDPc/N4UdELYE0DcdARzxlfAhy31BeXRjese
NxZjGzfw8CXZykuJvOzkGhUXcN0lWs2HZHA1kB1DmMzL13uENed3/lHqwIrdYK29
Dov/USASmbQcNByRe6CMw22P4LIHVaQn4UkFr7HbQh0=
`protect END_PROTECTED
