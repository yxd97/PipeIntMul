`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BeQEwvlaQ87fsIdpdAzQlJUVj1mhS1oqT1DsiOxUBdp/dh8Aab+s3uxEdzD+M+ag
JVHkcPZP5/YrgWvJ/92gvqpofQ9ajs/j5o8U7qlJ0ycVwmALDQCzZOGKszEMJlV2
inGUqxz7xCyzgCgRWCA8HDe8pUSA2bQNDDP1lIWWCmT9YMyWCOLb/tKF7mQ+MDaj
WHXY0krymlRo3isdGUoMOqvivblFnwBjgnTqDsqUEBhaTDkM52DccshwHJ4OHNI2
0aTCdianzub40hlxRf7iFO0Hx+2jYYepaefcZnHHsxDmlFRgY85qKgPS4hs4PNKM
2OITfJZEBZ4S7Tu/gVlEeGLEAAej6R+a+qKcOZ2Tng5Fh+o7FzCTdBr3GyjoLSye
c+Juq4f45gTAMlKB4GRR+DV6BH8ZMjZbWjh2L802hTdhP/MdaCBiReVsYsLSil2u
zoJzuPvZNeWEwFag9Aj76l0EbKB9D40L+ECy3z3NmDRTSYuPSz3PWQgy3qf1PVH8
Okz1PhY5GMNxSzdb2zpgzGAnnNhtDchD8+7aygKQGSGQt8XaczJFFqj0G1Jaq22M
wMOfp5ckvASYMDIj52ui8cmNe+aQOFRN2fjQ4Jjwd0drbHfvazrDbjyIag+MNzIA
BdZtBvbjZBFwTkBxwNJxH+tde63J1vry2gKYuaxQPABzdy4YPQa4+b0qb6tXwV66
/gfupgzGG42lNmOqOzsc33dD4qOxgKVbqLVa04geCII5HzApQSWDG72I1Jqk4B8j
rA2nKJ47ai/oFHrFngB06DJcN0vxYy8k83qt2jfrkA+WM38iG5VJjoQqxU+T5bV+
8SzjypqlaWu1c79940i0ruq2smo88q5cyH8Vl/I1c157rAJOkSrpyV4L8XJRUi8/
sbpbD74DakAnggVAKD+dWw0BzFVzuEfeF8a9ESokTqJlKSaEDZ4+ZwfEzY4Gdywr
/xu8NSmLgJCxyhLkBXcn2m6IPwcMACb/xUPIrkzFTAIjW3oMMDZnms58xEGgXRaN
pZHPFQnOFKtu5ck9ZqZYIUAH/6zNUEuoD+6BX+ar7LrACUIvptj0q31LZQrcPPAy
+wwRpmWNvV9wPNuoQJlVjgLB4VvX3gcNSh/4Rvby8tqBHvI0cjjzqATfYy16ZTL5
R0zAizXRH5ZQbZZHYK60NBjFXiocdeEnre27vJcy1wDiLk6KVQ2rpPLpwcLUJX3H
lAynnA27MNfPptFiE/BnSSGXbecIleBAeubL7Z6W66jn9kjLUZRT61XD50pxqjLT
W5ar5uFRFXs4m5GN5YXePn+KzqOmtOB6kAExkZNoBOyrDvDKBiMUGRfSEWhKcrcU
iT4+HUSzDsmGUR3BF2shs0fXk4YtckJs2jdkg4yNHTbP9WbM2XEZ1C6o3iw3MpRn
ZEHBbkUU4vxPRQXgmVgcTlDNEFCyqeX5ydd+b4DfVQohr2Y4kIBJ5IgytBDx09CY
Mn6DZ2YkO5lFdmWnTHI7zv8hMZTFnaBNBX7kySiIu+JCqTqDbDD6DflTAbs5oetk
m3E5skoc1MZYHhvzSrntX40/zHFz2HkGq9cLSRNdekBtMcmxWthfzxAsLnAenM4z
axmLGc/o39D978s9uI/NwHLFGaDbzk5rNdT/0vHK/l6tKEu0lEFL29pCO/KIjAhB
RQAUMJ8f+PRi3qwCxyUggtTmxlqlSsazZejyXlvQkj+p9DOrmZfbZd8nBJ6BKGB6
CZ0M9zuRv9+VyWcap40sOx101mRUtyq9ra4vDh7+02KvkEszqNf8XVrMO82mZDlP
C6Cc0w5jwKJzRbOSU03eufa8N71nf2uMXmcy9S6gXG29B8ojPuM1zECM6yTZdaR+
E8tJO1UUfoA34E0D574D0xkN0GEB9KSZEWSLfDi0ygbgiKlK8DXUAn8WJbQE7YHt
pKracb337ktftjcucdlsBH0Q/8N/wkvFXfMQ/vfOZQF07Vg0KA4NqoeLB5iwsIIa
unujQiHtpjQfv1l9XScvL31Kq/a+XWuinEJpMYhDFItmOpLmoqPyydFY8dNd68hO
cGbn0EaEAov1U6ymS5mBNnoOJG78KJ+zr8Zo9ne7Tw8RClPeetXSqQtREVWIa06D
M1yu3zCJzuZczRZ3n5iDoEpexNH/7A/yQvIvVzDpAZqDVj03JnrQe1p1hw2HEkY1
JRgswCbonkjD3740M9I/ca3lh9/F/6Hev9kHHmcAQa5/eccD+/cpLcs07RJla8i6
CbjGEjyQ/psD1E4Fs6mMw/efA9J86gSpAscuI5xwXsioxf7x+43FV6ncqGrvxeJP
4wTajQDgRPH+CkUG6jGGQFg2hUOqlcxzCxFPjUWnHslMdCYA+B9sSlJgZmaIzes/
UFp32LrDbAbUogN3qjiHGRSS3e6KlnYGsEP9QSoItMXZop22ItktA3r2ZEPgpYni
VJphYSpk+wJXqy3znNynCFA/AD0wbWqmkOAhgjzZvh8JRvJUeeoOqwTuKpPl9w3t
1qXuXzAjaLNfWL8/fO7vjQPGaTzZyeC5LjXlTV/Mj9LFHNFT4/RPEevKNhsCkp4d
u5uZ6oiOZrMSoWAQhTXE0NMagCmyvgpMfD68ELVi4wlwOwtQVDlU4MeW/olMMNl2
Gdsde6nE65Uvh0fig3zDbzzOw3u6B9C/Gqdk7FoQ7K+1bC6Ic0+OiVrFIUU3VHph
ke27hQENLhtnGuGzP/d5b5aOO8nM84skoo7B38hE14SzsVI+H+GJfIFrXTNbeBFV
rPiD3BTXJEjSDWnR2DOPaeZhZqN88pIqac5qVFdDVVbmo/cjGsHIhaqs/YpEBDJa
PYS61VRspyX4Wxad+9ZncE5q2+uP3lwVR/qb22hGHi5ENrRvnGbqvigTL6tkoxGx
csrZMNoE62OWzVIrhM8Saropqaksrt8nUgqVffSP+7H8HqN/IYEVFXHx/FHihd9S
Ira4Au6q5nAhztfpIZemHNYxkPMSVxFm1UMJdQ7DVTnWWGLvGP45EBPfx7avHYMu
Virv4PYhFqAidVshzL8zHx13nfPH9ljrYoGlbLes71Kf2Fd/cXPkXaYCn7kHqUPN
c3Hs1JUu/N5WPjbgh1aXgNfKqKT1Yk9DKBhTR9TS/+CQtHRyH+w2nSGoJyQm/U9l
FT0fojLZYgpPXDCIn3TVyxBzydlPV3quFCDwAynwaZH909gMFlDRGI/5zt22IjIM
7qkIPW2IdO0kj/NayPuOVwzlHTHx4XqZCuzBzlDMMm9kPufzd00b0BGueJr8kGCI
x3AdqOYwXXoR+PCaBPwD3s1Xdwblak+gACDYs4SVkzNVbvExrUCb9ure7pXx/Tvm
IoQ0LnSDs7mHtasyYBVQSe/r1VaxRhJBxOmXtUHlxRUwbZOCRLn+3JWK4O7SOF+7
OXhbCJy+EF5Nl4dDBoHk1Ud6/ggJadHdbO1WlfMylck+cwTuwoD9qDEzRMcvYVa0
UsVEMz8DgbIRf+kVnleQY6yWsGaz0h7/aZY9MmdpW3lDA+0/RiSYeQRmogzF/jxl
Bnoix7X6NnRwB6jWvlS1yTgKWf1tmJB5fkr77u9VhtvIeLvO8bW55wYe6a99iDLr
yBU6UhiRQpDs8qN+EQrMupxyxRXYVhr8oG2UYPwS6EHQibJ2UrYXItVVEqeaA5Cq
EFsMaug1Q6rF7BCXncFL1uwKiLAXa/g5lbMLoUVyx2DKeGaR106B2zz5665UaeWz
dH5GN+H/meOgtlUga8o2HY8+XE3qtGvBVEnc++eQ4p4AW2AsZgA+8F7hzk491224
t1wlv8SUF4FiHydEqbKX7ETqj+6TfakW+oZrHTrX+5PLDpOgkJzrpTvCf+Mv7h0a
YY3abQ4uzZO4s8dsXtUXI292ySrVViN3a19+qWrJ4pGtnfE/WgbUPVZyL3Du8Oin
IWVxSg04HXRYvj7ZnSK9V0z44TSIqxiVXphlDVrKzYUxLTCEoVKg2yC4l7DMUpqy
Mq2V4ExeqgJ14O3bkiXJIP6VfDeIZUZUrDfrx2KKP8IMzKCCAA2bH7VyDruNFz25
kiDKQhrkZITaPQPzy97REbYdEoQyUBw+NfbOgc8e7qrBCjV1Ia+S2XzmV6/63LLb
rUil9iCunWV4+QsnY8JpqyjthEgX8iEsmftxPw+CYvlkIXdTqFRH56Q6RE/jpOJm
126ymy6/GTvKwiup+1PAdLpgFyoRM5RjjTeWv5UpjXW+K00gkudDUMvVCfWT5xJc
jpgH81CiQZyLsKJ1F0qcD1soRHxIydNi0rDW/TMmmHy9Wzp7LrQFsrVk9npveaMT
iY48wc0HYlV1dtN+qmmIUj7LgA5TPv5OSBgXAfmZdFU57VACUwISqSBAUw2H/4TA
gYUzqPfJGs38Fm0GcgUNxTcxQxyxDLBJ6oSWNkhTHq5r9q4lJZ4nm7lGGoM0j4Gt
5X9f1pMF8x7Oa7ZDF9ifkbExeCIRlfc9P+JtnG+9DEE93p6af22T4mXgRIr6X2zw
3aTvkdsQinCDJNXpHg+vdYTMax9iJiJBHWT9i9tE22YlKFE04J7Bf+rJom44d8gX
NohRG33tpYD97WLuqcDmhLmcy09B0gk+CnQepL3BrBQkHFtgzcYitoP0nG3eY15+
rVZ2zE7DeF1bcsTn/aXT6ETJclYtwi957txVGRmGzpbCef+RFR/6yrihYCOhaVhZ
/sijQ34eQhg4/XNO9KRato77iMDTX5Xyhe7hQiRSlOv7nqHRwuNJ9Mbotkw0+KOj
QOnv9EtZTn9l8YVGA6iu+CAYu3ZfuAtVr0227bJkh9lwGco3pHyPpG5Y4nZCE0lH
GO43yOueBQxDy/ymAf7RyqMOLJYTgNMxCCvcBZdqEZma88Y+oPbaHf6uuLkTa1SP
yDecdc22J8tO1PH0LI2Je0rX6oS/KvkSNzs6YcSWIWCc8VBwSpa70t4AGFQ8nmsb
Nt0ZH3uEhYOkoagqSX7norQ0rYUPzifHVj2n9Dk57sAH2xtL7khywJ5/Cngscwd8
0vHl+5l8GHzc9AZM+YLWgw4flY0tv4aS/vhX0xX3VS4kSkyCRH7HCq1ErBBXSJE6
ph3v67ObOquqoG2D2cMDJxfjk5VWsHYIO3z04ANa4Qc7qMnutkYkAuzL2q8Hq++3
BM4heb1QAzmm00Vmyxr3kgIXQb3uocsE2Vit60pmPsBuxMrkhNdwydC8OpJdNbUA
7Sm/IxLlZFoJe0tUId0XEgfp5KVa4Ij6zMiEcTibBYyVtW69iWWlaILuO2kDe5vr
mAF8/UIbvY930G54z3AvRmtZm22A84OtsA1In+aqCMeW0StJ5eJxxGp9lR5o69h4
GGKT9y9w2G2CnZQ6PWbsyy0dzXva77ib8OSkIh0AbsLhb+7UprymWKzQA+2JPFdR
C8eLDBtYd4Y33NYKrVB7r80dUkRZsFo8lie4cnCJ3DR2OuND977o9+6ul0ynw+d4
NkO+a7HyyT9XtIcn6A3kkcYD6haYcejUf7YhLCF8yDpkn+9coJBy0aksctvzVm76
L1R3Z706nmDmRRa++pyAB/uzkWhjpmTs/wtdijKAOxcf8xQKw/19pZ691sHWJ4fw
diEDNmyYDcop0YW17f06y/Nw1qBA00J6tkI3bzK+clBWj7AyUtf28ovm+GfYLy2v
UF2E009z832nm3qV5fecAbHekkcWKuYdd//QsMekiXch2wbCXUlrr49O5fXAh5qJ
KjCh9UDBTk6yCNVUkFbqwP/MspzQjVlGjMwcYGneG+Tp7Hbv0NLKBxAjyENIsm7C
hUPrqrFwDVDSqaFDEDlcsD4cveDkPAT8hRg568CEPvFOOiUV+mHg5k8xvRMF6WAb
mAGlIsuVKVbvS4u64wOuXXrNqTCYTNxo305hwNnaMCU1+Pvzpk8e6OhmDeL1Phyh
jtJ6iK89EdEdJln+CnJ5M0SPmh5PQvlFb78/lD0St7eQ+QYJ5HO9UPgdnCMIICHM
oMpuccFKmQZKcxUNuUbqBm+pcc5CZxzgXdn3TknE/gOzfcToakq2wVCNzl02dNWT
G2EjeW5kmRNhI8LPwSTdmUNx2grgRkgAav1wtJsUuvouK+UdLnbzVd5HguOLU7+g
YlPHC2lObNHM33MD2/FS1Q2txFneCPiuYo8z+IM7AT8GIm/JQZxwOGsrpqWRRA1u
teafbcfc0vtWnNu5Mk6Pg9rm18G5XhbL216zT1zFSE7kbeVghpmb/eYprTMKHvld
bs6CpOZY1qSlIKnN8qqQvCcbxqQAB4vzEqHBSzIuP+nk+FxC0DE4xerY9+H+PIaJ
RLcoXQlI4ylGL60nYgHp6/Y2Qi1CYIEwdvyF7SASvrZKHfkwEw3bs6xcHhA5w1YF
FxInb1BsJV1YuPodQACYVwmDrx9haGWM4EISbOKkbws=
`protect END_PROTECTED
