`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OfUjYP/7OkxPvNMclWFFx6aWPugtoWkTfy+trqGI7ht42QY1uCfjKEAEuz1rRKHl
uB0x4PmC0vawJzkrUflaVivk3/gVCc7MrFS7PIHXGrCvmrTGHQP48/SRqqvOOkB5
nJHD5j7NF2tAYXq3U2XpUmvXe5Pun7Hk8ZcSII7IXhQWb95aa3IyLWICFuqHu22g
0ecZQX2xJyq5Vyfl3jOEIzbmQPWElo7T99JPd6+XrzcziAGwBmyxoiw4QlYEbRl7
1/iT7XnlDy6yRl9eosRimnJPg3126aadtssQWLuag51s+eNHE+jJWtpjq7H99z78
aVhRs1yxe2FU4zxiJbVXhLMdyRa57ELUoidOiF3n8VUZDSr7G6cO0+KTgXIiQEgw
8Amsyj4SO6V7ONCo+jGoYw==
`protect END_PROTECTED
