`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ttKyt4+fCJHCayfTE2kubzdfsGKrQ9Cns2P3oBa3KBme6kWcb7fU3a1kAFrdU3yZ
aE451tL8Ho+gbFZLQZNxz8aNalAzVruzV+W09+JR/yW3NrBQpUrm2e7yvZFcQhcT
lWUtSw0FppbXPJy3gVDHVQQi1YksyL+BvAsOhKkqqu8rBYTADBYXyPS9INhWYYNK
2H+Dm3dd+eQabSgkTm2DEw5ZsFoNZscozi/+IoPEyt54VazpEBi46SltVhMzYKOc
xbKYji0GcIY5pVwu2vRETB5JKhXlbDFEst5IYcNGNAgE22x0wymb1EH/huZpxsvA
S2/4wLagDe5lF1FtU6/zrvk29z51cmPUadWTOikqDmLLEyukho09jYO/HOLrmr2Y
Np/f1z0ehka7oGQq46Iie0HQUxQgS3KgteQM6SgM/6Cqtd1+prI5AieYuYrOC07p
7dYjClgmtS31s2/6wzJFuxhg8niEXz4GZ8lsBssbDXMhaxZKVlkoIS0Hq7OQb2Ux
QGeuVCRFskTUzuhSkTxFFZkol1UmllGZU+RdyJNCW4lG58HbhU5hj3QWF/hiOU8n
Tife0e/KgRUzvxcCUUG79g==
`protect END_PROTECTED
