`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9FpaFv7GvSDzrd4ImAbD1GVB13uuaKb6+IXjyPk+EiPoEs01JKph91GLYAJwTUp0
BkMk3COK+k4VgqIAuJkcT+lkfFgZ+v9nrP5mloeyLmeLm1sVS20MERuSIhdVtAHV
cmr11FwrTWcrFe15rC5eUND2x18uUBxrG7ZQ4dJbq82OTSMhvVFotGP2eqmgrgv1
6+6fQtl2lEcNwGTEmiJbvq7AedXoM7USmiLiq4MHJoiO8Y58m1aA4mtBTMGAzx7m
W9nx6eKQdt3+bGR1o9oXJPwkWcWdsAVWYOMedX/mPYgZfgStesfNVBzil3UWl0j+
9obLzQv9auO3Bdy2G7/IPwpwP2AcF2y0K0mS004HnObzYLRRLE/Yb1lVefh/rCv8
JfqMnQohwGtG0s0veWg/iELe/c78cPJHQvJGVRasdoqlZOREAMh32DJdG0zBfJKA
rDIiGS1w6/Qp/XXEJPyOBd1vEVEhKRqfGA9iGuwDNgDo7m0/1HvdVkoFwov8O5T6
b8hMbbgsAGCNncHiqCNeCyCC4mu23M0fobH1S7U3WhxRjsRCt88w3i6Wh4QxRkhV
MBv0MQeHRkcyE0g1P2oTpN3LosQ+8I/TnxSprBVo4jYMd1BEMBc5F2bqtPytVc3S
9uhHhQQ+IyNLnYLhQM3hfzDLk9ZIM7ffkAJNCUgRTpk=
`protect END_PROTECTED
