`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2bqP+SvVjTSHWtzRvndqmpaTyEFmqM7m1qijSZmNS+9A61PN2gw+orl4gYA79ABh
eXX2q2L7GcEPoK8zWnBXriL/CQCiBTo0TOpPnfqrlnLN5ZX8VtBn0oxfJrDbg8xk
mJXza3c5EMUw8st5b7F+VRlQGTFCy9TYaYuErzxGIY0m41Eek5TLibu7FBxlZwbm
23w2obOyvMTs6hTRIHXBl8lP15UD8mtER+tfJrctMQeJF58oL4536eTqCtpJ4lSA
bT9dTw8Sr7SLgqEvXy6QiroL0ubC3n7yNezFu2e+DfOdeZl0+ay09uZPZNkk1JTS
pqN/p8q2w2WU/7wC5yzr/00T+Uk9oa0iOdQe976HzDrddF7lXbB9dEkU8JFyxbPL
s7XnURi2X1kJ2jIRVvp/NBSEPFX0yUb6DKUEfpKshZZB6Aw/Hc1hfzb/mi+xn5GV
5CJSvoj/W9rTjMmosJV/7hKRLu1JSzEoDYiJ/HGihv2EUo6Cgphd1XBtdb2LmiK1
`protect END_PROTECTED
