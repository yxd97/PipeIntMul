`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vMi328bTT45mntYrKOpuKjZSLQgRZRa/OdEQSDO9Mi97H8aug1z3kz8pagDJkQil
bPlzxmuBDWYJuxHwAQSvIedOkDnoigLZiXqr6c6NWJwAr4H6fQ7ZAidE8ixutlIl
2WLMaQlAzejsfBPnz5fro1A/HuoUBMqWXg4u6RoaFbHCp17YT0k9gXMjZ1Fk2SiF
rQvcNFzvkNR/wBGoWsKnnMYwNy/NAbHyzBK67dxUpPKkgP2kX7JAmR6xR0Yc7pgi
91EqZEKAyaKj0+wnWwhU0wVSOZO8cfJO8o+sDeJdP0e7iaLglquPaa6WtZ85G/Q5
WPEhsJYOqhYcTMRk3vZhm0hGymbnITpqTr4uxy9exWJtUK5ixOaY61jL91aQq/gZ
0ZX2d5uDtFCe3nZ+fxaYrXa9eSCLwhxA8CPebwi0e1GLzGOx8wSM5cvU3RRFrqpt
l0X9JGDMwIRrly2xspugrEvUvg+0YoCGAhmsojV+fAO9jq+fshNeyo9+YjjUMKUW
1FZP1BXtEmHv66FRHuE2Ys9dkqulva0JFtx4F7tR54HCeWI6NNUS6o7Fua47/MpQ
IdkACGzusRTTtoRXi9F/Gw3Ts7F3ou+PuvTzyqJq4nPaGtMt4W0+zOFhFhggzHOr
YLo5o5g+jZQ5/WC1FWL2gHl33yB8tfr6AYifniUuIYxn6xh194eVKdJeoc0EmlhH
zWJc1pwhExAcSyGAPXmKABtiJl2CNb2CwM3R5f18oxi6rVJlIZk2AB0pzXJ8pj1v
YmPkwOdfZ4mFqyNhlc+OF9FgP8Yn0AMkQGC+oHqjVPQT/OZ8BqkF/eELeef/CiGD
pYkVjMLYI8wEuxvPLdyTMc6aEzrzcZWUHyjwY3RE1jnMRkWeyfAwi3cJyh80/Pd6
WpLYcjqA8wdTO9BAZxNFTGlrA/2pZT/jkdzvAAQwoxoctHIk3PNglJqeh9tDTTcZ
Q85TIDzS7dZoLVcV3D38OKuXjEU6Z/wM2z8KOqg0ebdk0CzWYcUN2rsuiFTRwO3y
zjEiX6TAtzieyvRFed42QPB+0Q8L64Ztuai8lVOU189co2P7CC6/vDKJFdK8HcEw
+9OxDtxIjyZ0eWch2diDu6i/8p15uBnubzKbxRcBJsPIx+1VJ5kHBLYXoRl9b13V
a+32ujogOuwnorpOEI6cV6M6nDY7NWBRZL1dcJgnlEwC/KJ4yCb1sL0LO5FXcFHo
Xdpj/+8mMltarwIy+3v9Ipnj0f707jYaw0ZmkJ+SgglKsy1EmO0E5hGlFB/SdDUT
sgsH0lKOgwwImnlBnNYBS5ThdVgdx10cRQ8iSUg5x3iVyMtaYKZyn2Q9mRvLDRkA
7ZHnO9KX5FT9/ySuwNHFC58YMtGTLyfxyBWXSZZHjN9u1EuN4l6i29h+QG/o8N47
74pnBthRAEve3+mqxG+SSw/o5nTrqd8W6251V18OBl5k3G0881+UvJ3F13pdv8+9
dODF0AzcZ6hSiRvZgaftU5+QXQMSMemY0V0VFO9DW7VogkOYrm/givYbLgx4TLkK
HGsasaGQi2u/YWoaWEr80+pJyfQXfBly0+8EcwRmIj/j1ZzyCmzuFTEbutARQsBB
6fFOENWOJLIKbyd75+PPSfXH5L9LrYs+84asgCs4MbwVLnTEIr4VTvUveE48Cmf4
3wYSTDWjrU0DI5Xx+YBCNilxwjHJ1fvrLxq/P2tH8SA8pnNih8n01s5ZPfsQhPUB
pU/81MvGQap1+JbxK4k496JmHKSiS/woKo1WH8uad59HV+m7rwJd3A0Lv2gca443
eezfVcl91crD7hOq1Xi+gU/b8rVNnV2pAuJTUSFZ+lUvXltCuvkOb+Ub8+BBRGsm
fhsPgIqXNWdjJOGHeV8X/zlcK8dKkzcJJA8kTPcnBKit4V2e9A8WyI1A3hOmXQQw
KzkKlWHr0SWnanJEBSNnE7BZd5yWxkq1bO0/nT9v/9RS/20KL2rRynD+KYcL2t2T
ZyjsP4N6nYwLmLCllTaIYI9KPZuN1BDtKL54yV34fBQCOb4a7Jw+Dva/1bUd0TTQ
QsAce/eRD7f1X6BkpeWbfdOcAGbMSqpgg6a7v32pFYRYso9Sii4Mkh4ATflCWnoZ
bzybxGVbkslHrV3YQ5yN3mnjjFqUciHQiEpBI9XyVIKO+NK5gsHUCDXZRYYqi/8l
hOeNFSkepS5YlcZ0ZLX7peo8Pz4eN4JkowlUYeZPLUpjxTtFO2yMfr8zh18sNWZW
N6Vm8fG2QgA319i0zF4iTg==
`protect END_PROTECTED
