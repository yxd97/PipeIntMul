`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KDexTnMlWrcpc03SRrJNR9I8DFLQEGaqBLzbd5OrAR6k+Y9nFpJUrmOjSZr9fK4H
CpIe/D8olXLt/tqTYC1DW5RLo0I8dl3idgovVN4lVm73Zo0MsSTis6Q1vAQh4+IK
E1pUOQyofLnpRsRAodb3PBKYhSObzm1HnyZ8IitTQtTqtlaoNPArwj0bMSZ44VPz
tFYmGOY8BtHdAmrlCdD7LykqK0MPSTljmCN+rCW49W5GexXpxjslpMYWpWh+Vx0H
X0pkksKR9wQekhZLJ1asE+1nK/lyQZ/Td3Zg18jyf49ak15Mv6a3hDz+QPyWuLta
`protect END_PROTECTED
