`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXiQRlOWAvdmFeg70Z130xYkKp9wgIbcKNsPQQvB3GrRQ309tqaE+HvE0AaH2fBA
kLZ0os8tM1Bjh2bIPKfsWzURWA5sQG4iwl559DiH7KiONu2gbjBjVxRK9dMUzNOK
fyNj+SzmiAWVu6/kxhn62PjiaXYN7rP+NlzBt8hYnb/h7uWoMIKTKOKF2QjVUD3Z
BkIwQLoh9Thx+y0T5x0Mufj0UEPfQWDLIeHePLQ7Odj84O/pYciXLgUCXY7Gbnnk
JYon7YpFHaOmR/bp595PIPHQiOlwl+VJ627hnyhW5uNAVuosgcqwRXxmb26nMRDw
bkHj4CONFucMSWbZmEwRWNqbJsqIVnU4s/bNUxKKazAF5xcDSs9J+JxPKQkQySo5
+P/DJNphqcspl7o0EMPWRLo56Q+Ai/mUS62vfPV4ZYxLPHqvhwih8yLjngEsLzl5
dJjH6fWvu8GSuMeksfinwdRaWU4WRvTufbMgZY5W/QmxtJ7Q++b5pg2urT8S8sy6
A/msaYe5EIX0T+zsOgdHPC0bHTGKn5GvWzi2H+9nfR8=
`protect END_PROTECTED
