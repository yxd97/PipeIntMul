`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
omUxapVZBm3YNJyWITiXDjWWt58tUMZDNpbSnQEVY5+DzHdHzd+nydI72dI+/z/4
Ty5eWVqroqzMXbnz2B6wZYiAhbvJjy7X7A1MOFMTx/nCf8BdI//DL1L61Ce2g2yN
evIwMENgQTUb7D5XK2FqhHZI9g68GM4Ajtf541Bim9ZSSzlsg/f3pfbhhPlaNKuL
fqWbRnXmklzIdBHXbtiGBBI8WQgZO5hwBgxI/HsduY4tZWhlQMN4cVqB4sqwxn1U
3juW9JbST2BHiub95XT5BhbGFouGkCqfqMb6ctuq+9MpoZH3oevsy9SMNNX55Ua0
uvLcFu3BOc8tmdXbbvc7bzGHOcYVWE2gPQOpBAfPmVJLYsL54ziK8ADMlF4gWj9r
Gy+kK0d7kzQVuKtY6iQ3pygo30eiyP4LI/s5PwI8pBKR5EXs0KimYa8uhJ6uya9+
6ZLsL5kAm42baqRrJCV4LtMlaslMrW2Va+Nbu1knFfggTheQYqombngny3g/stlV
fNHZDA5TndPIm5Rcot56KqWxQJqqjw3Fi4RjBtR/iGw5N64p/8jIwm4neuqvfX7Q
JFNqYb5hEJH7lQ2dWggcAByxwhBx4Gnjv0k+ogGgQ2Ob5/VB7MiG1QiSjauuosFu
It9GN0TtIkvdOQYJmnsAeZq81QYH1LMSIfWzU2RqMo7PBB7QOMllks19LOxD590d
Nu9nnMXAhL2ikn7m//JDcuvqqab+lII+/ed29N48nfhV8XEIDXakB+WYvcZhQZWF
tppRuslllA7EnUkic6tVwfaf9huJgSiJw9Z+gJj4LE9oFHctxxv80zI51KsHtX0r
qyrG0fcVbithhAjeZNyp60ievVw/0K5qA9z44iAJVxvSIf3FlW10hnzCrb31zAxB
JC/49DIomOUPKN8L1teZGIOiVG3glENgnHj7I7lOvRNjkdPZop6usAeaTYNQflxQ
Lg1R7W1hCPbl+EGnniDYeWHiTxDg7NE05x/QAMbOgTMDqeIgoQHu0gzGyQCDv6Mq
L6obdaBJXdjL3hguEiXCc4FWAjLtPy0oW89N2+972W5ZIWI2PH7hMZpjPUf3je9p
MzPPydqjxAzYv08WWoMiCQr9teOXMdKtrbJ6TzjKIbuZkmJAB+HmWwx+4/igJSc0
CKlDFFCMk1MhJbsvuzTxpXOfnktoTmSisf35r0uPpskp9rxZoRDHv62mGEZrZS+r
8CLz1BgPFUfi5xKYrXfejzSz7j2BWcWhVaME6wuS5Upg8DoRd4RPH2pfpa1AJXId
eqfz3DVtZFHaMLWQv/I4p68ARjVYyje+v5S4zTmevRYkIZ5nEZrpv+pkOsUFJkdL
Qtf5Ir/8ldCa9PRI/wQ0er8DH9uSTHNU7v8LPHDkiZrOg1/79gcs2HWLEtwZE/b7
`protect END_PROTECTED
