`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LPCJIuei0Rdmt5Zi+50LSbdtjSz7hAfDVFcgw5FJM0u8cIUCrqp+9xLrKnmK5YK
roKdN6yEHp3mTE4If7ae/AbFlMG0sYj7VXPqlCknlVOExTos/7otTZBp8PzUPYJI
xzkJtDmF54HIsnPxcuAXaoXJ3V5o9ewltT2+ZtmCyN6XCaJy2qey167iX+g4BwjV
otrsyfuApBp9aHKefjm2/TStixEfM1xn7Q7WgoaWMLceJlPyHDtm/JFh/P7PQfQA
EBxKc/Vj3xEzMDlXcovhzlUMccIYNmYAnDaA0kaq1Gc=
`protect END_PROTECTED
