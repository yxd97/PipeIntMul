`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uGigjoCOeycszPgW+haciUBmWEBlV864jaso0hXiXrtXK1xZewSH8fPbq7JKDewp
0O8CBLGDv2HQuWUze5N93JO+6QeYLEYZbmwi3jBaqNlS8dhZBbosO3wVWrCLX59X
WXL+FUjg9d3kJTW3HqQwqb9DQLSAWW+w7qunFc2e4T5qPS08Y6CJZX2QF0/rxoX8
UAWxiIw7chiDpWjPCQgPuxLtZiMwFwachy2x8klWndjmhHp3EzJ1K7QO77L9jI+2
6fTEBEXtnCOpzjsAYayVMyQJwKUQrei1NAa0J7cy+cI=
`protect END_PROTECTED
