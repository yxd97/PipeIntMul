`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c8Hmlf4uBHPlbOtx3kgrphJJZ3qksW7fr5vCck01oq+O8KHL/yHxGuTosURz9Wqd
C3KXKmfDYD030bIoFL+sDkt1oFiOYcsUtpypc2SpZxLJWK3oXR/kNZIhogTFj6F6
3JiSI0rM9zWZYbeTtjPUYTAYC85uuQT/aDNLcfCWELu4OX2N6RMIhmU+0dHdabyH
fOMnO1m1Ts4+6DC3cS93Wwu9hD1pOYCukXoH1tJ+nm6GbGwgdvG6uiSawDsGb0tO
TsTVbqyGVJQzNdecZwKfITpTNWMnncniNVrWJELNCH2VbeVgj3MMC4g2JyDbwKyB
PBkU9mVB9KATETzNMVQQw0eGJdW4Q7BeUyDvuHc40ixGWJyBCfg7A8VPEVhwwRIK
dlbbDMWtpjLNaedxbDX2z7FMRr20vI76/wjcWc0RBYcjlpmQn5r/rofihFl8GTNl
O00g1TYRIXqAbIWC5u3s8QSoy1qsuV1Az9Rz7qE2SmizhFrTqW9AwW4CwXJYFfyd
8ClKJArV/WjmoOyIxomT+544bOZ89XNYj4AoI3qS7TtrMi7Bj2U7LqDzyvE7PxMF
kd5tE+Kf3LZn1yNE/NnaUMYDPOjRfEvPrR6mkxbLwiPp+l3c0lbBFzjGNeQspysh
OOqoyf6WRF6LqyPZV5ceEySRly/6u1rnD99VwxbluS8k76sOBuE1uB7vQOA2gZzN
Z+QrIPz5+HUV4QGIdDJ6lz3u+duu3WHTBPe/19lgJtE8EhEplcKN6swzz/XUVDHY
Jec0ImocZhb/mnKIWihMQLE2KvAeAj+/xh4FM5uJDfJhdG0Rlp1a2Orayv96kttO
9Sn+MidC2zeeKsXNTX7p6u5cBsHf+7UPvoF8Ty41h2GET4SYgqGC6dsGkFeCoxKe
z3A3YDJqmhwnLYe1saa+rIAbcJl5fexbmqtVoQtnAn0dcZ9GGckeBBP1l9GlFl0g
BWujVZ173f7B6i3g5RCOw1MQkM4wCn4LiiWU16jSc0aBiXnuGU/dOypBY9SwijPV
JIS7nMRkFyGZ1tt7x6rl13H/Y6UImuM1ARcgVth0YSHvGlARyqlaz0yfKinFu7BM
vR9WRkdwFxVAN5DxlJVVCpC1Qb4FaBtznetPAgO3rCrEoRaK+YR5n6iEli4lti7d
gseNjpw+6vxWPeVqI0Oq6bTTyhiI0VF/wbPZsZuCx3cV3L7ewrPhHnF11fUBHwmo
xQ0cVfozObQv2EgIOCTa2DGLXbdtp4I/oKUTKNoONDID0nws00lnZQEMN82dAHz0
DjKDdw1gR5GKnxtZPTFUrGLVMRNE0xRX6fq959Hrnq1SFNMdBzOfwTq0h8VGxv3Y
6KYwHc2P/VDUba0NFJlfdsYE1PINf9xA/uh6NRH/qfe4UdsB+TFL30X2sOuAGy+x
b++pIBGj9OVnkvKe4mwFoTznQJeB97Lqv3HIp/BIRnq3x0h922ArMiGCWiv232cr
UBDFj+t+sp1umwJx3q2QvIaqdqkTtMG1Mqe41ZUk0x4=
`protect END_PROTECTED
