`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eDC5fQo84D11571s+MDiUipAqK5RE9Mrp/RBufiMWL/s3H4lgI25q3z8C3mx6+0h
RD4bKrYuLLf+h2v6Sd6GTlkNApFjRMvMMC2aczdWf5AzWcFyVR91OpFwMMxZLybv
WZQaulBE/bmAZ3M7JF4IWNU/aWrom3xHZI/af/yqMd42fHNBzgHGv42ls2VSIHeb
hapV2n6FeXIAx+fg/tHCvetG9DgdNW0UEcXl+HecmJzd/2e2FoOiN/7d+NdtLzEc
N7rrz39I35gMMA0K2wWw3n73xFbSwKnpQGS5xDG3K08f03gk4m7NaoqR9BTBkMUZ
TZpajQyMk2bVbtST7gCUs6Uef/ArZOhb8bsaAAzW06yZT64JO2AX8riF9BG6zRYm
`protect END_PROTECTED
