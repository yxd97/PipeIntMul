`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1yJ941qhTVIVWoWNdGJrhpd7hhfS4PaF1hq4wVVEdXRxXm3fQnbKEeKt/WJ0AT4f
ao9Z7oa3yVuNbxZO+YYvzx/XdamB9YEjVeCOQlfQD8TAw7L/yFuZLnrI0KaIpz2N
cUATRAa3rRoxvZWUKsmz5OSK5UCJpBu8I6sKkVpoqXtqQOU9T6TIpdz4DmBzsCDf
P+flvnH42uz/60clllM0xkTXCANR2C5FK9vSFoZK2mxVISxc2WH25OX+6WUuaoC3
p/rYGSK6DVBvemjv1P3RdxHd9UoecmI0jixeNg3n2dUUO8WefWxxiKaTB/WuZCsZ
8B2ljouGLzVddqFzwpywVBPpk7maJK7JTCj7ctE4QtN1YOXq8ZcYDLchSxGx4yju
kZX1gJwu80KSBMalMRNniQJoAPrniEnOH8i2gxx16V9zaHeXe3dTQoZX/iUSr12i
BfGgnzWWwQqPxXQ2ljJio5A3cT9PEiKu8wadhFYvz+uJ9huEbdWj/DNDSMJgxSL8
QrcSaDa1qTn5wr/qYV5LVy6GhFCNsgvcVIG4XMkeU+cnE74PA5tM1JrEvN1rTRYs
vJ80LocSMqJ8RbHDL1hxGyGQlBXx6IvYaKu4/zkUyZfbA6q8FQLZCRIWhjoaNe5q
nvIG5yQ2o6euoeIDxP00oUZsMzJTrq9FdAtG85zWzTof+BdEKDi+3n715ycIhSmi
nf9dzgafiE3tdYPOZaEh3GwyFAznOoXRo6pdjlpVx89+B3P/78wOeQCau+kXBrxY
mWoNWyMRMHrB7MTBE/0yT65O6o4fWti1P5bQmpLy3jDXig0CKUR3OgT+tB2epDmX
rFjdvTsaaUSd+cCFJfNFgQ9Azo5THXp4la+1PojSHddXL94ESWCsfwWgKYaVUCBU
7u6nXvSblvZq6RZRnEiuabsWN5ByC15agHXsDr3t5ML9xSY8OC/1F5Ah42JMBjVS
QD2LL3FZNB2TWfODkTHfTwXYwvjRqqKHQGk53U2Ad2kgxNM8Fa8KeBMDHqwzewi8
ygo2Kuui0LCu7YDwdN3f0pDOoyb1w79EQwyE0pvwLgMcwil2+S8pryGMC+HZEjHR
0KJXXBUyWzROylKSFNkkxH4YIsRqbAfqDJGyHxj/A0Tm3ZEvlmExNlhBxRHdRUKu
zv4WcUrZh2DIsIzl3avD764VtNJ72zLqoWMiXqmI1OMV9bD+tOkuS+Uq+XvikzSM
s2hEr6obpkBm9foeI1FTwfwaTbUvEE4tHAiKWRJf8LR1s8UOexlgw0hFrtkrv21H
TIZRDeJeLHUXS4jZ4TcbKid7ThPJZf7UNczUEYrBfVrJv8ny2trgTRjOHnvizSPI
3MsdMyL9NrgO4zjt5YbnDZkUf6Ob/Wgv5fzdiZNU8dLE+rFJUfdf03degfdk5jRg
ESS98TWbRotu7PVWIp0XaW/CMmyiEs3eVfT2/4zU+tNeP6CPd8bwznnV4gbTNYdo
00AqYV9ZkQDKqN27F0fkHb6/fa7BCpaMaBk9IJtYXfhewsIl9fIM/irmCSuC0BZ2
KuSCJ+YNOalGtnPSmbaEvKtEvQsgZ1n/Jk2OA+9Qjr687s1lVegkWEZnQ4REn01K
NYjKMP/Hthe4d4KJHjy8oOsh4qJxAajL1Szn3H8ykDc/lrvfC7/wr8onJtaR4e2E
QkiFGAtkyTDz84+7patCDvBtt8VIxVFYNrDW6fe4Mn+nptzQQlEkniGIBpifqDDI
ErQ+YndvrRk2fUSNyVq/HXZg6SaZ3ZpavaFRYmV8wQ+6LYabUnEuI2FK+g6P8lBK
yoN9wv8Rv26RJFjvNjKZzL2kfxb98LH8Vf+nJPrSp8cFAHsBC7IZd6KZ6D5+Svb9
knucSIAhJQWlJPQpUkn0P72FZeEjsS9iEbm0KChl7JU+CWkSIM71BcUGDcFFV6JV
ecTiQ4Mo9qHwkPjEIChrgwN5KGtHQl2TuOolkiF2BNQrfxM/dRtSCFmWuTY7CAHw
Uc6w0U7TywoQhzHOlmYuSC9X7c+SHRe6NF0ZFXSkfEdSGBkfe9TKtGi/dCcwxVeK
cYGdoloUlFBAsEYZH/X2TqK0aLh3cWXZHOJ4YDobxlyPWeWS7fISLjaI6DsbNEQN
aGlVCEAm/Nb6Hjcr31VNaL8cQkYK/95vX9Z1e2akkNSuWk5hjZXrisHvTtHlCyuv
fNOtbURa4Hs4FMU+nJFYSm0WUivTtnSrUEjlXP8qTH8quGb3GlZGKfV+3qXN8GFC
/D6kTLIOwosXZAoYLQAYH27LF0K66n7D2dVDsMilRmVbW37FJWqsN9HBgNTJHV3m
7OxQKyrBgLGhw04K84GKxIGjmpNwhYjRdNPWKjzbfTvttt8OWKRkBMHIH61xzwGH
hNFRotnewzgxRMQwnl93X0XFqQHdgxpogvzajT6AwE6AIuF2cnNfd8rhCQZJbi1V
I7kYBmHIMFVKNCsBODNrw2JmusKM4j04WgpPHLGQRa8cdOrqA4tRG7hz+L2DZsmc
HrSZhfN3jBGe8UmomZltkY4b3n3H9r5uYEmmx2vLIoyCVBLHHOz7rWDiDb5zBpEx
zp3i1+u/AD//VWlcjLV9jFihcSs6R1rC3msyApn4nYcJTlT0eZrWhVYbGhC2GZ/t
NhbH8afEjUBVuyjQyZTOP0eQnjDfRwpOCUOrrO6bAAcb+Lof67moj8Gh/t0Z3skw
cNDol3tae4fINV6gYY25iLAf64ionmJI2kwOmhqlov2Ir2s12iWiY/S0Dm7VP/A8
h5lxw+POBWtDxssKg1JoCJOOJedgouasdaFu05Dq/CrXnL8QJUIHIqQRBp4eEgmT
set5alZ7VNxWLt1szggFczfOVV1Ku+8ZGrRYW1btVL/fbWDMhwjRvS4g4fXZwrjX
qecwKRWk5YLIgWjP+wxDRZrjtD6fkchLmcJa2xG/YV9L1RiRJQMa1qQdZ/XXy8BG
6VADmKtm5nYa7JWJNdaHPj2E7w7zWjHuSFxloccsNKKKVphFwMgEAUP6cPDqSUZZ
I9Bspx1/vXlj34TT1j47Yf2+fbeOXykN/El+9+ONT/EpbC6GsCB4mNdzd7qwM//m
m8obfiFyCptYd+klXT6+2/SoL24eyB0Ck9dihDdD9Q2K522KQ6FSJDRMutP+3pri
PtrKWMshd7pYbR/zQZPxTcp0tyX6fwnHUtIJiKQ2J1hIFBCT6IFWUuS76GTfZ3D0
fj62VuZZr2uV5fzaS8nkF0/4imEYRJVfjTmQHxjvWE2EzjnbofIcdfs944W06OMk
sukhD/DpV18SY3w9SBNQkyPBOY8W8DyebditEvICcrIcxzWh+BcmnnqPs/WE8+cX
Sm6Ve/KreX07yYY/pEp9z2hYQHbDG/MPxvg99+jCLPOS0jqlO2LVSAvyK+9Vmlvp
FtlgiNrLPFB+ND6jL30oRkv9kKKdax5R9pAAwJru4IcHgbT3LEtFsJvgcvPjHaeZ
ymax7/PehqdA5SUvJDM4i75EZheuRKJbzfevau9lQJyHKIsi/ZutRcGzI+2qWz6W
LsMKh/1il7EhFCtcYlVMVnOeJbWt6UHUrvVCqOKp9ZTzj5+J97zEFqSb9CVoPdP3
AhfK7f+I2ftqz0M55yos/MXYsvPSemBkdwCIc54RUKLAG0PvtelMlg9Fst5lEbcR
Qag75wJOYKcsSOZRg2SRglvQK8ZShBaQ9si8oqmNqYD+U1PYit30qVDMbGqOOOn3
QbMbL+4ZpJxukc1jxrpI7WpMX3p/vG0zzG4eauqZhdteYxbhHYxHQ6W1dTg6l3v0
oxxqlQlra3L+UTDFevHi+tH4f58kwL7TYQSlp08QDjHZB+rHaEpJu3C4mZfowtaq
W+JXyOtUDBMEdVcztsQXM5EOBrNrq0ieQ8okRr1Wwpu7WwULPneQLJgAn2ASMYDl
WLB9FPvCUY6yYIePu1VMgSpey13ELiF3prcN4rB11r8rmm8ZtzCUYmagwB47ItFE
uEYJleDspjoLDKn2Lutz7sFw0jaiB9aMl1u8QM0StFP2gT5Gs00DSDeKAcwoAwZl
xjmNFwfYayF1oxtGJBq9emnBV5P0d4LW/K+1tczzzK+/KHxG4N+BqL/lXYrND8wm
LfCCguJa7EBtQZudiUnGmj+YPP34VZHpX/jaQJo/9bxDVycM4lymFfbEI/GMJ7v5
CbWEsGRB5PLQpLA/efsBm8WA2q74WzZJjhC0RHIwJCk3IxUb7tIpg7DoUKrJG9UL
A17h+w5A+daQZRI7GL41NlZ1A3txYaxI0C6lebEtwj2J9JTNgdZQkiK7xLNlxeEb
L683I+1qj3u2yRNfgWUZfFkZUgFae7jQueFhfyWuShiYXVHZ/gTG5fgtvnqIhNnW
n2rgP/ncdTzT0uYFp4Ipfzvhmcfx1YqqMIed4I7nW3sHDmP2vqw0rAoY4DRoz5D9
E/cbv16jBBQtEwc2GT7kDEZNiVEs6sHjer0ek034f4CZobbPF/ne9yY5x6/93H9N
j0gE5RY2otLiyQAmf/vaAhySmZxXphrABTtKAnhTTCI9tV9t031X/QlWWHBI6MOp
If6PuAn27qh6uBB/tX4wkuolp7DmiGrrRGEBx3eWvAcBRhOjo9G7brPqaAyTksTm
W59FGmrviHzZfWQCjY1wCtWwG0OicvcyO3EZ+yXPNuWG6Kr0XElMXv/6xglTMKay
nAml4ZR1hIhz87Fry8VujzR5EotOQqsHOwDp03yS9u37jj4RIUjxVr/2DTC/ZaFB
Q7muSMC9JZ+OORyTHVMWfu086ZohdjSFBGYUGW6BXHraC3SuqBN5Wdxw8yVQj7fp
uas9ibxfuMvrxHn0+Z3TliZ4jcI+ww0Mg2XRNFT8yKttEYBOxIK5k4sCfWdcLNBN
jAAX5jSg7sWCipg2bGUloizYTqE2lL5PfpqcE0wTweSQiN1+u7293gplq7gVcPHw
YZxbRschYCAixm7BbA0rkzYX36YoqNZ9rCZ/Pe2A6vWKOqVNo+btbwhDEdtb4frJ
olBxeJ2SukGoJqhyXhVcFRnPwluE5xlhL5jI/9vcSUanbUEPhMkARgGt8A3UMUIB
+XrP2ELM7DrYzFuvnroqxnoBJpUZi+h/I0tAmUObeGFxRNVHlznLaEJOPys4WEk+
y9Wd3DHQgKdhnt9rx0iCeZV9TLJV33EkT5iRK3HwHgpA7MpWPgBQzi7ZsgVKWBMw
8ntSISTOZSpFkBG8epyTnJUbCnYwCjPII1C9zrf0nIXdmRRPaFTPoHD6bOS0pIj0
o4+nFMzSTqCmDspNZQNxUYKXLOyh0Z9tz71GwAjBmjkXsYSRvYT/LheQRu72V3Bs
Q7b9rzyY3+Z8a29FiSmwGs1vNoKAob/K1jlGYk/xHhJ63+aFTJHttvuqEtR6KF7U
R17Rsd+k3kZ4k17oQX5M/XEmiDp80uZIoOv9oaXY1+CwdEA2fcKWP0/U34l2upIo
57KDqxSijAFsXiAroz/unaOJnGO4Znx7HAa4/LQY2XUtBmQkc1e5UJ/XQpEwUUzy
IZqR2R+9mfZqQF1TRiCE+SO6slJFLDawlCMhMNK5gfgdfsSjSp4QosBebXZSclJC
x0ljgZDiMNYKRTLGQKa56mGVjOMooLR+Z6IO6+EbjbzxvnNh8bixYvFKqEd0xwgh
K6CUnQMMIaR43iXptXYoCfzHG+UH8VHfX0PnO6F3K1MYr2IUU9aemHXlAVaRDFJY
nyt1E/0NWgeos3Kt1x1twTA5wyYvg7bY5C7oatmf07S5XgLky3T0d6REFnvEhZfY
7e2rpnZbtilzEziT0CSiPk4L+tb+VIINZejIM5Jn3rQFBPBIglqnVyTERDYVWx7n
EGIMj7e6rjMpUbsbLwankMVXbUOJvnhE6DCPfjWA/SH+ZGd0rm83q+CK6daRvmuF
HReLVlPM3Qm8XrL8CG8HJstKFmEMCKjlG3Cz655SoWjdqLpuDd96D/i/C/kuJY5B
QpUOoUoh8l1ANqyRdRw+iCPhM23HBpW30OCnqt5RxK473+pdE3mWRloHEgtzUyW1
NptVHll75hhd09VsU4NY2q3BcBPWgMg6OtqqAVHRwpKrg48/E8fnaYub+eLW2HAZ
3HYUl9S8gHSnKs1WefehneHRixtfuLGCgeL8F1T3NeAlN6I2IRg/fgMqAsAgAVkv
2vFetqqIyoOKutMdXqFxA79fF49psPm+MGcjUHL5JyjtvRnx1f3ZWGAgk2OxsH6j
injYR5r5FqpBAgp+6XmgCQpmAeNwHgbb1rLZrwnvfycmyWIt1Qm/vO29986rvQnM
NccOytHQKptI3KBFkrKoETajt9vWdhuSyYO8KL6y5x4BXW/aKO5IhCrR8sjkyH0E
31VmmaXf56nJTT3zzm1y4n1e/wphUKOGzlciJzNClzWPpRn0jTfYahzI1unGJSer
ikF45BoK7Eq21LAqBZMMYemUjNJ/KP/Qf4FZZAHxLT77uZAJahrlwPh4sNlPvfnu
7TIoXNOzOIiwv9rCAvZ2i+xPLX6puJl2WM9n5AibhAjepwVBRV/uUbJoRhIddWwa
OF0bHaBVcEf+0NpYcKGIjW4gumBSlWAqQwWlSdMfA4yRuQzShi0ub4dK+utyy4RE
4HXOjI5zV6ArG6OBi+ZxgKkYfLPBmNgECry6gC7ItEyh3qjTvxKBf7r1A4jKyHyp
Z9dUNM6niptFA3Dw7EMr7ig09HAiEMSNbgCkv3cIMrnYIFT7BDYWCyEzgihMKMpt
I3Pee41oXiQhIzb8x+4JbKg+5FshQiF4/WNCmd6VDao60vair79Zarp/K6cwmLYW
lS39ZOyle1rgizZDCFsLPQR0ZKV//bix+5OtCVmsqnM4XQXei62IV1Hf8PEkkokz
OTp/dm05NtfpctJR80SxalHgXh//eUTAY7fskULNTjOkYHOOmhW/njgNdysuVOQm
2Lp7uYXzxCkFN6r075nsfhblm1GacLpYZxivKShzfJJ0rHMbYxam/avGA5RcAhaT
alyYcNkmfxvJe2Zk952c10PPxbaIvbn2tvFGJt9hCGa+H8wpkgNyqPcgXHkbjzKw
yKKerSeI0i+5JKVJfDJoq6r/pbEiwRfTKN0OaGF2ihm3gn2OTYe3XYPudd1MTT6L
enecCdQOJ3hpuvPC2qLgPzycYEV1cVdAKWlSDs85511IPy7HGOsLXKjlktw2+LoX
ePgObZGJZJ/4UmzCOTNKqSnO5mUkoKQK5GQ/34icVXux55tUSkL6f3P8UILBLszC
ff7b0TUCJkdabNU10doxGDLIROblRRx31VktTT1h3F2/WRQaEvyQ+dA+Iw7lP7KI
bJ7n+Daw5vwVuWSs1rGDC4IlfEdFQ7/Ns4yZB0FtlvN4NWhSp4HfETFcO3+Lt9lP
xEhpZQeuXZcTmAtp99lCqb8Yd3qGNk2CAU5EhgsvQSJiDTGR7PLOgPhI4mvryZNJ
m8hEPa6tFdr5xBodrwreIs5Lth2tNJysPLika46ZC2VI7trxns17a4RbLqtWJs9K
++lIBOdFI8P1P4oemrgQOxqlpBq+08GOjTFnc1YcxPohBWP9HsN0Z/zxiCBFpvbJ
4EyQEXDs3RIt5tnNooWE0gAbPn+whj8nnnh3JO41PIanmKQ90a5vcZTgHxSoTPGo
wdHIxrfadhmEKJpZle2PCBIqQu8zyAVZs5Ihz3Zhv/fvET5TDE/bo9AEvgsur+BU
YEzQ/XVRslWJVnoVzz48cNC6uQAyuDs2oRNxc6q6Ewo+GT3dBxlOhBf9yWP9lGqN
T1k8Id0kMlB/4r210i2aPTA67+UUHXLRfzNx0jxacIGPdAnbgFaL4bur9Jk2zKhl
XptSO1KDmINOxLACSUbA95KVVbLSHtYLoOjN/DZTtCalOHOrA6SUowNw7B68Zb+u
uoWHKgb8eem/vy2QlF6DJKE3gljW5jxp23IbstoJ8zn9L0rKl1femm+XOptyiJ0+
sB6qE/cNColLAYCuNfYnsF74Y5tzTsEWWvHm6tiPm3Nhf4dBo8bp7IxYMyTkOsxV
I6+utZnH3l3xMNhgw38jJzzSJJUc+TaISbqZjFxwKZ0Nyj3f5uFvnQHFkV2xqQv7
yy485izAL5B8JvPWOvbOBweqPdcju3ZzKed6todyqf2H6NIgli8pjr46dfLjEmD6
dkjKHGge7CxyIEJHkw39LbiCXIMWvFehzZONnkiKKzG+/gZ8Rr2+3Qa5gL85RIMj
8KUdso2iVd6EY9Q6lnSKdMYtx6tR1qWcY4AqEWKVfWYcapTYFuu7rXG3/Ppa1Nkc
7A8j27dBp3iUziWyp2lL05je6uze1feF5tRcFjmzot5a14l2/OKT4VPYZXVH2+VA
zRpPRFF9/K7Yei6Gymnxt6Vs91cvZQGvwt+xA1GlxRpOoxobNevlpwes2asRM50j
GGZKVgO7oWOSmy4O4cK5y9Y7ZfutrxBqz2RoOpgBHNh+T3EW3+jULfqVDUBSBEIq
ymQ+DadTGpb2K+ZeqP7eM6JH4G4FKJQlv5YM0c1VLJw/iv6ySXPcSWZhccgd+Gti
7nxT3GM0WtYczVQ/yteddhMxah7me/aYXn3ISS9i5cDMV6hKdb/ykKVDZ/BSWqji
M5UbxB4qq/M+biejUSRy7bIDCZuCVE5DkCzGuFLeyNbvNfFnraRm30CNhLYDuvTa
PILI8laOT2fpPYk7mg7/4OpCbUrrMesaJVJc8/kKvu+Qs3a5bJyr0B7nPn9zKRrG
bzEM/XEhTk5xaB8MgqRMDvT4CXhJO5sn7M1xXNenUPlZZgftZj78ITsflzzP4jSL
OoBvtZednvieljBBrr4mVYoJetHK4q4g9EbUjHEAIVKiRIgweEUF/DjVooYbar4H
3liswkBq0KssimH4yg4b+gmFd4FT2bDIQFCDnRNObbW3I20tcLo7oDnFWJ0VK6LP
fGbbGMvl48aEEq1HhJktFSJ+PjQIapaSNvCDXyjEEQsY4YHr0UfyPDRX6N+UCDwS
DWceLbNWKV/3zxAEpb+Dk2pCqVw4EwJu+z/3uv4DxQ2Nu7CsPOj7OP7niM4EaiL0
rR6s5YJFWDpZ3mjfS5eDFzbjO9LRBEPJiswaueeDfkcBSHHcfx2Z2jQbOyoNf2mG
RnoCOSD9ReoKZOv17vYXflt5lV9ZdDYrdTqnRR33sqVaASF9+q6GINXk4/ssppQX
kNWE1+KU+lkIGSOetyuucz/KT2lLA9+FYatZ+5KVXtlTfvF2slCw82wJvy984qUH
O1Xd84F6jDe7A5JUb7zW5B7MrHskPvYAvpvAYPwDyKP9xrzZfUbGmttWxx3S1MMC
pj0ubsw8CJxWp21BZOUUuiVIOv8V0PSekEzn81O5j52/4VcJcGmSGpSSz3nR4feQ
jkRw9HniZcBVu0g5GN2lM3y5kC0ez9z+pEJG8n+FMCO/Npe3kHOLcub/ybteaDCv
x+amwCr5D1v6LMOiXiwHXRM9rRMygZukt0j0m4jfHp9ECIdgKT3yxHYWh4iHiikq
NmKNxLpjWr9TTtygHV+oEtHjQktkIRuiX6N8C+3McdB10VRCkzv51xbIQ34qzjwA
JvZgBjxSlc3/WNqd25GTgoM1mUHXHpSBMxT0hZIxStQYnAemxFNC0T7BylToz8kl
MNPOabFXnvx6R2IItrAGuNUL9NdhtdD9pcd01Z8oZkBR67vxh8ruPIJOTrXTDG20
bBIp64bQOaYpDXZa7OQyxbyeTQ3AwtvPyDVL4AOFH6o4m7L4rIN7DifNnf9NHQyj
ZoWfmi5sFa9nNwPQN6A3xebryMczPox/r/DBaP7WWufzowIzzHUj5mk3M2F1RnuR
91BeCun4aCZBtUEWvwv++apJD+76f6QlV5RbrIZ2S4fdBfUq1CXX4Ikw4p6G/o97
0+qi33/V5hPZkanm8BOHZQKsu5cl6uwJA9WtzCimBQ3EThXlFoZCOAhNfyphg/xO
Y+64aWk1x9pvdRm2SQ5GD/PCuvccbeKS53jSwK5wad2falBgH2tLP/EFKdpdP/Pq
le3pYn4BmL8iNGO1XrG/YTRFxCagSdBA0E2xH/QcNhuNg+PyVwx8fWsfJl1CxCuT
WpxqdQVuan1bIUY8oil3eeaqCz2oHzWNb8ooSx/1wGfC6JgapEIFCIlamcmLnWkl
mP9JYxn7To1mBmBz1N6sVUsHP5sQjwkd2wwyaS8OG1zwi6E7fg7b7p566bgd2vd6
9Lp4kN4NWN+aIT3PeagKpWz0fIgN4EkW3QS3QdLJCM3Qun/UeCD2oaGm6eK8ZSUB
CSB7m0r7sfNRztJ6tEKpCFnyxGjHGX0Al5GDaxEDSrjK1e3D4q4fqlIlt9TKeGCR
U0esvtExwOwYuf3GfeSb1KkfUtPLM6ubgzF2VA4Rm+PjT6LrV9yg7KTKXJ+2U/D+
cQNVsJKC7XmAspTSnZ+Ea64jq7yzwV49CX/4n7exPQnRcgbAiF9RTFMIKaPh73rn
BP8TmHzGHF5qjw9Uim3OMCGJZ6Erz4z6qiOx8YIQnh8Bex2xdtxh4mH6UY/2AbwG
r/qztYHfwLf4GgBONxBgdnqpDmbO17KQaDVWqZLPYzEY/JgN1yNAHWzETvJMlrEN
ARPMecPmszXrzuVOiTi95kOAnyd9FcYahy+jDkhNbA/lTvZwlF8CUBggpUUxpETM
HFJBU5KnCjt6xOddVrQ18QT1TdoB8EWre61HHejumcZZQTXyJgPLMokVCVFjkKb8
eBlD1KUUoBFhGM0ldJvMKNWjcuuOzMJjGNrUa733S+0btf2b84vWDHcdLMZhjFxg
Ypv3O/t4o+V22Do0+HC6wr+7rBmH3xdPRVADb2H+X/02vLL8J4P5w5SaWegPV2Zc
T0OtqdFeAA9jsvUqUYGyv7WyqWH7BXbCpQG87Tq1S6w9f/iB4ieMU0OAQzuSab/a
eq3S8aXeaxNXw0M7zTKGR5WxeaLTEh8BjfagZ7bLccaM1BvnHUxxWx6mS3w9vI51
Z8AMoh1dpmWmdcnwiUrupMeuY4bLqI1UopSmALsuXxMwP39xvhoQVbmfhjdGHBbJ
c07RTx8KGdAfFLz1M44abxY/9YBjJq4ZwENhNcuDYYHPWeNqVrHihtqB0+sfd5pj
/Po2zKBX3aVppoGPSWZoRW4uqkf0ERxSl0RsgN1D4THcqecvfspuyHMh7ENyiyGz
DFCeF8jyTLxT0fX2PxRa2yjWPHlVcBk7QEqTlpfzGk5wYiVmaI3iuyz7oWxKwbXQ
ASLHc/Aj37cKo38/XgmaZkwBjqweb+1NvRlS0k1GkfGCdG6sE4jnPPcp1U3ilZzt
UDtaZDDrs1nJ5FE4L5CGZ4JuNvk8LeZ0Y2DGmuQT8rS7Rjv+zj6mU/cQhAorSS/A
b0nML+2jFS3V5QAiqH75o3Cnuy7Pau+vQoTfOfgUQDhmRL38fgdOm39i9pBUYZq6
8Y9WIHhck+piyEkdxtDXM690CMGgmandVo2fqrG+L22/R0c1g0cvQ1gQ+q9T6M9M
bMF62FlajFWFcC17dvrc69XOrnuaBHB3cD4YZvLCc/Ic4SnOkczFHSc2r2dUynFU
oWzmv57iHPR/DtYSLAMoFIu6lfhwSIxOwsFd5A5nCchrRTY4skiu2l5ephJHxtIW
LwzVuJ5NlgW38SuqG6+S8mVtLiXP26NhQiDEYcLd+BuESPBD2rTrWRxRtYdmZgpJ
aqIXWBkqdpvVzgjTLWOyUNoFZJPU0C1bBP3fvU+pGqknWmnLROyxI1nA3oB/Y/Jz
demEYtCu8VPF7QDynr9BDHa0Ioaw57gfG8Rt2ySYljjfJentZb4N34BsGEFUQHmo
ypjQsqGzvC7XahFa/bagX1W026NceGE3jo2iRfPHxTQJ624y4sbW+zqBAGaw1+6C
cSJ9FsRJ7igbl2f+hbnYiElvNMZ8CWnqReSSg/4GmpWWwuR3GMNpzyjzfOqVZgL1
SdSD/Gdf44sQaZyH3VEtTMpQHzl7X85lnxvS77BijKM029e+caRVsG9Smm+Z/gT0
6EYRixcU786obdZohHTycoUcRNbTTaXAW4GxTb7SAvSEGrbhIZOQmFkDwwZXxdBw
+MNOoSMWdyuOwyTDK/Bn62n0q7OUzyX2nl/v4qBHDu6qvdsoukE8qVk/g4Nbf7JZ
P2s+TTrxCaaU8sQakf3dApM3vjFBkucL0KNiVvX4EoBLlPa6c1aBVahk2I+bNwg1
Rig4dURNcN3qR0StzPfVKV7odV2l2ZnPsI1sHYTh5FR/E1IVuXDjvNitqpZUlb+Y
ZGmSh+vJxNbojWIn6jTg3cZB9qeTLiEFQhl/oeoC17yIfGuFRhPelz//FJBvmVub
/G0AzY3YSDbsQsKW4XHxR18G5idkg0ufTfy1eaBUjT1Ia/a6cHA3npa9DxaIY0B8
F4SRYjPUb/TQzUt7ChOK1iB/CJvoqHhFoFTAQUKFQopg2Sx3SzYFmXAPg0+jGu+0
m70Nzo7z5BM954vunly598A5VmB0SgvrfNJOKX4cNUfxhxSkTIfEyUvlMpDBpsp9
QLV9FsJmr5JYD3SbgYRUEO/W4u57yGjArzy411KMn9tbcEWun0hXknv+Q7NES2Fb
5phYonBQIzqt7ZOErGEaQWzL8ooUa64qM7UgaVtKitxrmUDtcEXoq0vbjqHB3o/y
IRFYP5+l3bzLWsOM0Tn85LmVV2WdUP/PThXjb/KREcDN0JxTTfMqvm+TU+TsvvEJ
IDR+CZbzQDiZfTLtzYiL+RWlX7/vWnrE/ioUHuuo9fBNM07MM0eFlf4ySTqzC+eR
ba/6pTSry0stgMV9w1ivK6YVhos3ahPTLUcSjXHu0TaVFFGTAXcAzKhcr9GCRUzY
FwxsmdwX5PbycegEIh8bTSIdMllnqAHOI9rmNIpKMGQG00oMAEeGM+V7SGTNXhnH
os0DdrhrXeVRkFjsfSNp4HhNEGALPv+4VCHzsKNPgGjTaBugdFJugMz3kCj47kjE
w0i+PTodPnGIALko7JhwR7z02i+N/JpiP3EdQbLZ0OIaJMtSDU/nc4Zs7OgEJeQs
vLrCty7v+0fA1G+FN26twgRr2UwDCAA7hfX/rVcY5wJUM/gr0SaSmNApAmUPXd0R
1doP+Gm5lDYlqyKpdszqOXDwHY+XwdiUJ/Ip/UYRTGoL37trnyLe44zYJO2oE7hY
4wp+yKhbLrtWC7/dd+vTHSyWE0Y3aZBXp3v353SNJcP9IqP7n++k8y9ZQ01qMFu8
PZRGvBj7SMQ7rwHh2VCbE9kVDtKB+sncE+8Vui3djPtO1nywf34502WixF7fKWuZ
LImARM3D91TTYg+t87Ko/OkoApBRzpSwNSfV0lWSAGavN85LmRvMA95LkU8EDrkD
2urSBYMJfYUTUcoBEymqJU/sdhh65syUgC9356Tm5T/QwkvlQeCRm26yu88S9nBV
dHTSPqync/JpQMDAJLI7QDlWiOwDvcbKrEwXAh76uxPMjppUhgx7hGBMo5suULSb
3XQAllstIUOPRrJnsLMAvbteS4bO6DseShSOf916Q0Tmxlg1HizU3djQfKd94qPT
cosT+Lu9uypWbxvJmCaLjmrZ/gfmZf/EgOmolvVz3ipAxhKmSP1RaIMiICOSvzyg
r6gOr/Uf2KtlmotRaen6jNZe8Fz/JMQXtuoB00vUiayZ5WDvMXHe9/QIBbta2FPK
CphJg7+TYE3b2jkumGgBlmnraBKTU0SX92sZ3HHgiS+ZxyewVzU64ra4i9BVO3QG
Vt7bObl6A0RvZEG3ntKTtH0LEi7Gd82iJrrQL6zyDzoVQCerQtO5JMZug+zF+9SI
fDc52R4Ey2yDbDqLs/bma9RWhN4diUHU/50DstUPXk+Vy7InuXRJOlhOoOSvd+wk
OtxB3cP1k/cfd6eRTcCgBgXkU8OHlIk4IdivqeIHhVLH+iodbfbW7NCZgHeTjaPM
lhU7SrsAz/iZwO0pbjcorH9HGILlUbRrnI9qXZF0hAn0mQ/GYgoD2uEeB9LRQMhr
vQwggfbuEZQHosuk2O2JJOzf+jDMIJU3HPItRE95dyvjqG+oK9wqpwdSXpz3cRFj
cJVddGBNSWxpQl2kOFtL1rsQuv6zUinlvq9XlsNe43kKH+Jfov9E9bfC9AbgvnL+
huUx4Wuee3F9BuevkOld+UyxmmUkBumocDSFsO0eOzEh/Nqgn3ZfXOh4yHonthXh
gHYzATltHEXJK5JJdO6+LDZaqKx9Qx3T8kzTUP4yahC7bKecbHP4dEkw68fGp/w5
P4j4xXmpdcZjQQ54Tuf0rapVb2KaiMYkYt5Ir1NWbgC8/0g7zsmou9wnguCS2RjU
j9atTLDzMpjCOiwc/Q1FK0LSvEn+0vG/YmLw0+IlTyaZjx1EXNRweBxlxUnkgBB/
y1Kez82bBinJUi3gzRJkt9tKz45tOGn2pAxmwR775eg6cnjIitQz0R3Rre9FGRJy
N65ESgmuEdHNg1f1YRB0IFMZNlpHZVWseHiUMJqsjjyaOkJPMpVl1/+qBvL8WlvJ
KP2o+FT8sBmWl77Q3aZku/dt2prg9hn6OLsep8GoaqiTPqRnOw77Cbis0IE8c4j1
QtpTjHOe5ZfaHVR5I1d5weXQ+WVuDLVQZc+VfzWWDa2x07hWG3YxQ7hieWAqAjpB
/gh1fPh4C/bPP2+u8+ZNweQEYKwoo2DubMjUyceAlpQ75TKLuYfworNrMoEWYbyI
LtCAKdNI72joiGiRRexf8cc6K4iwDPBbCLFa3tQ5li5A+XT3zLXsW/iULY8080TU
fNJWMOcT8fVhfaQ9EUosewb1ZMOAToSlMs6xDg7Rf/IGtiNyG/Ymuxjd39Ibcd8u
haAA24y7l1DxXZkPEj4Sg0XMr8eH/5IthONA/h5WE9N7xtW03fQUinw6ASTjEqrg
3w855yJLN14sdjpLAvBafBPKQ7XRxQ3z1sLxdW00I2DKen7r6gQzS/8mW2RWNj6x
FHFk78XNWfGSelHoQPF+ROU89YI0VwFnIM5TPYqTWv30tDSk2XDYOXWMA+llGUpN
47zY6KcbRigf2tcXx7ziVGQ5pslnIiaonxClrcrKmC9ol/0u9+cYWlb4JhbFXUVP
2xdbmPtuhT5ggANnmpo5nZX3KaVBNoqsBSj67OZ6EcoyCRrZjcqKeX4VY7sV2lPd
4+8E5cv+Dp71Ak1en3Q2+M4O5SjCjJTSZylEHjRiPWWQS928HdOvE1M5CQbU/MMZ
QtuJ6T4pAOH27CcqggHjfYmdkGF/lomJD//W+DFXtfN/SI/7LUrVFc4AJvpx9YeN
/CHb8OA67j9HoptmGzXUl4jejVPUHpkG0sGh2HMFfv8YZDkEryJN9lWm5jDDaOuc
xJcysnMd59qjI3BIMxA5CW6NIgf0kNYNDdTaXCDKQNvl1wSkDNLI+Ud3wkzHtG0D
2ONM+o4ygJYFupLgwpGIHGKqjY8HGP10wzaCcdlC020NK4vuMROkhiNyykcmSybH
bKJ4EeLAKtNVtVRTeXOFSV4eHgvt8RRKmIrRMI7bOFWElI+s+ITUMLk3l+/nlEJe
AtaSSmIlzAkeJQE91Mf4puxfuW0wPaSxBVU/0Np9F685Hc+JejVf9h1s/T36+rVm
Bky5BXIvbtI1cQQGDA3Zi0UoKcVx3bWFwJBHzpw4OZ2WWd/+3OPpRtbuT2CY8mWQ
SPe5asW8+BJnQQr24FUCObR4qXBSxi1QzXe+f80lhXaRH4fcKeU+vY001Y8r+OKR
1hEx9xXlqH1x3aecgMV7ieIdr1Jd+hVHppGDJksCVtLEjNW5Tc6jqf2heZKFHdp+
NeOTuAt/yyJhCU/Pucvy9yFTJRkHEh0kTB/4r+Iju6vm4/hhkb1TBfj9GUgJV6Oa
qEAM7TfJFHkz15VIsEsYp7Z4ovZ0y945C017zRX32nNxRaZWRzcl3PEZY9REuLIB
xzqX0+Av5071m/25Gb8bS8RebUDV54f70pz1H0h1b7CjCxCgT0jVb1r6u4oAoXiX
DhRnwkswVSsCqvpiAbE4qwZtK+PByM0V2QJVwMVqpRkEmcWluO6v6uW4A/iXXLwr
hbhCQONhVX49o6ClQrdOitFNteoJf9kje8NrixIVzxamY5jkm0QyMslHUr1mN17G
+gR28enR0VuVs8DxlPO5T7NYHcfu7+wa3cy0STIbuvIgzjF3ZNYKmV61rqMLhgQ1
tQ8PMUe40NXAcdkJCRqTEBsUlSAiaATSgnA/zrGWbSoTaVVUpoXhCy1EZEFu1KMo
je9f2ma9J4tKczWtWu5kMjfHQt2+5HQ9s0jZuJuKRrnhMJ08YNxoQBUe8wiceziw
Vexi7KRcnmaF9Cgd1+pEh7ql6lybcmHSmUc5wyREfQxAQyy1Xpixf0vu0mAeeNyM
9+itEv2bQRx4a5gTtavIqG28o3p8d/TNGorDviIndYFKBpjBKTV1Q1VL7Vg9pSzi
G4tul7twNZlk4TozZwqc0jttIe7o4p0z0BEX9fP1k/l3kAezMJIfgs6NJ6PSk444
badjBpre5Iegw5/38JYlYJafvnWyu6KetQOKUl8894jmnANSWJdUdXgQ33JzuQMS
KkWmIqOEuR7ffw/EDs+u1BixAkB29jShW1IIQ4O1gfI4SjDekKcbHCaWhvUecC0l
AYasU20pJuKkYG2PiSQfzpkoG2LFaoSEotSwHFJSXL1QOJr0/XGM0/WAaNuvmECp
wPQIyk0Ys8wPVSo471/iTI2DQRTz0MJBJjkBxsbQFJ9YedxjNVgL59AKaK5UUwty
q2zjfNyPHCNUSSF/SuQfvUDF1Uw243DscYvtXWi/j7M=
`protect END_PROTECTED
