`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8XL9zXtNKUS5Bl9929Fx6mRhjdOTiLzx3zsUdv14wfeEaYB4MbyCEoi0A6u/EBO
c7EdhSicj+PBLMeGnPS88O0HioeAYocJyCRzKarK/xQ0T3OEKUTkA+3pduEAEPCb
hx7/Q0y7RZBT/ZYdqBt+98pVJAaxXXwk5AjTrsxWxlENEXABsgXHWCIeICgqgeyQ
sTaLdXXiYb4FazXKYeQdD3Fbdp5pyg01fzg/jOidq1F7CtlDcxtFK5zO152/b6OJ
Djrcc6dwXrcZphTVizRlPnyF80YcNc7ynGY+IpyezVpsmHwoUDfzBLO+jjgw7t6V
Dq4kmKYyDWqUfv7+HjZIrI68bnXu7DkCGd6Z8bYdXqykAxFtAkQRPEsBzWdfj7NF
n1BfDH3v/aH0sE9TkeHWZpn3ih1KdnLBAkj6jI5fBHWMmtpZtVRyRA/nRUAQMHMn
inELMSWPXcLeYTSWFnouz+Pvf5fjJcnIbC+EbLxtH7F+eP3KJx82merYJVemLvWh
ODBhrYrRMJeWjEBJGp3K/a7WixZ0kndopYyDhpi4j23RKlJEr5rn89I7bDLKqO3L
MM0/3+B8PEUjj9x/aStuyPIrXb+AjmTrcN38seAr3yo=
`protect END_PROTECTED
