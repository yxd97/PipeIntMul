`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDh3H9d/WAD1cjb4dGI+rh3BdGg7Edk6YHZtebFK9TBFT4ZEHhldauYaFMnI8tlR
PvnT4mbZvxSqEmXOTC1EzozdCLhup8LQwMTyE9qhdSwhTJlJ1DtmiU+2DNTkTXeu
0zxka5YMKfYPQ/ibiuE8R+K/9d/aN+2ROk7YEx+Rrgwgfk/jE3XdnbQMmmcNIT1n
CBMRLkOFaGlDCh9Oo7kD4aFjKn/4Zczj/q3GJ6ebqmqZ4tyqAu8VY2ML0xnyU5eg
8Ut6PI389jb56ogMS5cdPghK7Mq06MIlOWi/7F3MUUH1XNWmeeJ0bKj5L/GPb9BU
31swgbtHYSOFaHQanqJ6WABH6VZ0QLomszI6fAV61tmNhXyYsRBM4eOy6L/OFlpN
EbYt2vgOHhlEwdw42WpArm5fPytblNgf6EagNaJyraMlXsFAnyNxw40Snz73NFES
eEUKK5XNdPVQTiynI7Zk0deNgqIE9XGtGukCHF9+M91eG3RprWqCxwANCZntujRR
n62MoHFucOickh57g+F3j26SnFiXrdT2ucHZ1O5FOr7Mj3DWddLb/l/pgFYXOqPd
`protect END_PROTECTED
