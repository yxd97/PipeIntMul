`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1d156Z6nTKoMZjYESnwPJdwqfv0Jf80Th9DbZi9cRaNjTzz7vPUUav2GWaXOEd1
axT9rz3BeljPfTnArSfeZKsJTZFRCroHT8PzZ4EzL7jafrn44rJ6rUs27DzkxaJo
bjMLMA8vnmJF4XTKcdB2X5US7IQc7s3bCSLsxRKdR1L3hBIKAU61jd4mdjrzawtU
qmRNU+GljsVUmE8JMbl1ejptRPgJr1M10bMgIGjbw5RrTyTKmyuOxDMxdql8Ylyx
EiUbGNLQVPYTxy0TTe+TuGhbkMY8y2FLKaFQCFeLeMseqjitCa6X3CqoQEyDMmCE
fbsM+ESK5mmIBOR8Z4vCdPsX5JvX+LfftznwDsmPyxJOUTN28O+nCSIgxM+XBTjc
8tL32gjF3a/Hc0PFhrdGeK/4rG3jVnDnaPgEUPDBqwHZlqZ0Pa/jxDrLNMab3SrZ
G6/p4CCwiEAv8nydMl0wkdiPkOwCyqlzQNtNf5elnyy7q/sFEo1mTniNIKp5Y2Xs
/p5Tvl/yGukPeB8uUjx1fuRA9RbY8dC1koCuSV0Ub6eLbheQgKB/6KKpnG6PI10V
1HSQ/XhvB1FETwuVnFEcgnpK9LedEtSt07mEjqLZvr2Um/q+bvmV7vI/V8fbvLIq
w5mmBKPls5ruNI6iAIukCtKyKEh9xRqVu+3tUsnDsDruj5mL58wT2xcDRbJb22KT
FUDkIc/6KuNzTveFl7Ue+NKsddqszPVjT3PN5fcL9MKqHX24EEelfrUp3b7rUhsc
a4Qnwl1M7LA/gdFMVVpxjEgahCMxNFo01WKeQM0QAYU8+ymuxEqRf+iHe6Uwq97R
zw5P613+Lxcmx1eig4HAm74twzccDVt5P8/Y3+t6Vs1CnbweEPg17m3YfNNbBSDQ
SVVTfXaRJGvS4cf/Wj83+bb8YA5976d03FaDkZ8t1nfJIEFV/cFHFNilutbYWwUR
cD9v7pVa3/IvuaAAyyvB7U1ka9c68u464xYoOYWNnkpLOeVN9GtyTqDsHiChR8ps
rLC/EnhsX15vFgJYT92YCCDK/IbAx0I0VLSlm3kC1v9JcGiLbiUKsaBsD3u5iepc
/6A5VFAgHhTSFhheHRx0ZyVvMDmUQvGVehfMKEYKm52TlSK5MYoXq1vytAO0QC/M
mqvyU39AJjdZn48LEz6dEtMiglKgjRheImrU3guH4PuDVavGp9mVak0biH3kGfCk
mXjp8XdGBuTYMEuLyFpfjfzgcB6h/zuT5oyIFZtdOKPWBW8IdqIQbXpN+uo92Ubj
dS9nfXoRR5CTPzbgolW7/6TOmEt5XCJmPbAuze7029x5hSaHNHSJ7vLu+5DyBiWU
LaJuW+TsKvGacCxxFjmGfF4NAsm4wBXk9VWrCEATnE7GLwWCwWsdNcqOvJdDLaOU
lhutPz+Itd6mJu+qzLdSmtUb2sfPJkJeBnuPLXiz2OHRif96WuwulAl0MTqNiDrz
9I4SsylML8Ypv6QmHj+3SS2Uhey1IgR3SD7piE8cHIGUEDLZQI2q8n9dwIaOoIQB
7h3+qQLWn7J3hfex87QnZdRhRoJKkbZTV/kZJ6co/NYr3lfIJZIHRLLa4RuC8qQg
bnwInf1Wmatbs2m5pTGyNKFPjoYk5k7WCpz01IwMm1vC4StiPUBO6uyChWEdxa/4
wnNYQRjznUUgusQrQEgLztgT41l13CCTFxx/dTArkPbO8vheF+j2m2GF9ajtUeaF
yofMXIdfYV329XQ1fIG/FGN3rPqsdI36z3sDJ0us2sgsldfmBJ6UpxkJSK4j3Kgl
z7CymB5fN6gHQR9o9KZFpFSXi39Q/tr3VqtHNB6dVH57MO6TestZrX6iApSlWThY
M9Z44FlLnKy53oD8L5P/rtubLidcFRpoUFEqpZ9C7N7EWfETKz+Ro+hHnA9DQODy
p07RvWkeuXbpCbx+pmm5QbPp/tlF+YB9RqjKEnsJk6Tf3s2JT2LJv3wjand/ugtr
TGKaj08SpCb/363qQfBxHcvK13YyYCewI6JmEBE11iLcNMTT6JfGLl+DCpDaxBY3
8b9HEISP0Drs/4wSM4FzFb3KyDKvEcIYFZzH7ch3bPvn13H6njvMmrOv4XHw/xCJ
9VKdTYFs8cc30z9NVRCI0YWawhg64lvaJRnktXfWip8LqWwS/WpJ3RiW+ABxlaDZ
meRCmMGdMp65JxrAjudVC4mJnG4I8Q1lLQS6FLtiaWbqvKQYJumNDnEGmYswJpJ6
IAxiOwV8sYAFN/1mLKO8xlsskivVYWNX5krtVR/DD0+V1KHlHSQnZLur833jErY8
zM1oi2xXT9ETaj0oLbnat1nH2V4YLvsMyzElopghTqO1u4X3snzuqDi+RvsocOd+
BUYE4LvlPZmZSOx/P5wxoA216+/0Ne7SUfOH1MKWNVK/6WDy5BMmbo1YuCBOik5m
NVYalLLHMM2ik3h0+ePjUdeijNVEEyLKjD4cHnQKO1T3k340sJjgsPbUob6X7nAN
JmUc+O2AYxwLqvyUsaMDoqOfnVAfjJfPo68NGmbiYkZbNwF6KE4ltE0C+VwYDn2X
JlgqF9LQ2YwNm84fH4ZGj/cQ1ue095/U3nbKhEYan/9TffX/IUDikLEHTNFGzQAx
Tu8HVMNMSlN+3x0asc8MDTk00Xd2elYe517SFA4d3+vIfsNg0hlZrnlS26PIs3rZ
v5OqryLgaT17cg9E33axsKyry6WjmaKjPM0OAdXL6s1soOiFTvIAo06OFrE/i1b2
kg0uBLy6/vT6WICF9ifVhr6Qc23g/nwum4TMuek9DkQ4yy16cNwOizTP/eJdp6b/
x+ofCXE825e4P2sagwsFOsFNxHR/h+i1Axh20D0HE0KY8Q69T8FUnNLM7kozvNJ2
JfXUBIuaabkZjUvQL9VFjCEXA/qiMLTg1cCW2dokoKRriXLKs6aeW2mInQracfoT
93H0Uwf8KvYHOtYn6hosZb2tVwh0Yrvz1QOhycnWs/CjU8hVpGQEWhkApHoCqtGS
UwtV2/q000z339vFJHSLg0qXXlAhoyfOETg5Ed+Ad3w=
`protect END_PROTECTED
