`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ez5LSciwdrEeIjNGKHpDkkdMtlLyePD4+fkzN2HbeZEq5i0Sp0RhknXAcM0e1amb
RywWy5gd+QlRZFy3ZWuTon88CtVdL+5rEIb7CGY7pkx7ZDlUmHZqG0GzfFBptB1B
ZQ/TEKwMgq9wIcXJnQwyNNqyEbRdWLISL04gMITIMyD/nB+EvAdsW292jobSBDGP
fygahOSocTopF6xHmRC1UOhOaelmHBL9rePZ7JlXG54vtfPSdiZaBOlwoHpkCCmW
s9mJzVr+11rYx/QyfHYzdYGK7xgU6sifuC0taABJF23J30xXud7JPZPpPzvT/1Di
1O+J8VE0LsKPwQDi/MOa5U2G9xZifcjt36zNMGMqPhW+9bG64U0BS5e0eywKpk2k
h3oJXCvCEetDUb8gj0GT0Q/jWcAuag0EosSjqLbOq1/WCqpqo95siKjvkBkDo/HT
iKRJYBBr76zVzaghmZFVnlUj1wj/w22SHoj9n51tmIKUgTyGiqwj8MoF8oGy600o
zXVEBIb19By0eLdXu3qPHhY4rN2Qszb05XTuIWNBb5vFwfNLHPS39p2wmPION6CL
VLmBs63BdJMIykP520cVnQSPQ7EIwLcOc4zWyrae9WAITFwoDag6lWNesHqzXRtg
BGoMOUMGuoXR0RPnwqqzGJNzei/fQSSPIGP4tJbhpzjsU5Fhgi8V4zO6rrh68MBR
/kXtvZMxi1FMR/7CWl7oDtqmYH3XtfnsyZCpg0Zl6h4DLPyiHqO4X8WDvPE89RBQ
Aj8z/A8f0zuPhBdwiEB6jOoP5lVe9hW1MUPtkJi0Hy+7R4EWU2TST05mpw+FCjR9
1Vd0uinYXRP3b8ntWDq5Iizq2TgF6yAU/WauPgPD3nkHhZAyLXT2LBtpgW85+5F1
OQTh6ronUtQz2QW2jCGXwipleC/2vF1fy4eEZwOe9ZvwZ1kYXlc9voijdgAJF2n0
jOQ3+pdLReWh8WAixnCUKOb9LRh96WFxfLNTF/mG+T+mjivTE52l2NNno7PE1s5r
u3Dnyhu7KpigXGY0JJDjlb7+zKJwcWGRTD+2rB7+m9wy7aR1FnYNAXHC6Plut6pi
W7FnjwfvWxTyyxD6wBpsNHHcNrJpYwgYV+fhC1FAFpOKrYHxSwMIh95gB+LBn75U
+adx2eXJPPNYvYzmbfXzYE3okWJtbwR5hg8Y5oVoKhPTQ9oq7BwbLp+20zuw6PVB
P48PeC9TXiMJBd+65OrwvkbF5MVYStziEl9loTQxz/VRdJfwPLl3TpGT9mMxVVOq
ol6catJ74DoGFYYJAuUH4BcsIX156WPvqXQMXX3iJi0Nm4jX/MZ9NZih7pYaOcKH
rIw17Lbk45cwQcXlLCvsO9EsgxKbQt2udcW3EZjus2ofb2JYylYpwCrHTQAwlI/4
VNNo7S18QiWe2SzZ/4uOgYHDPNDqi9H8x7biVjtAJm71b42kvHLfsfIq0VJu0dHA
8qn7aWkPLImTd5OdzlOaUjbYACysUca0vYsKqq2KSm33XjrsQaRziDW+CVANcQO2
zA4J+NQOz2Ze+LWeVyRqNpDvBEEgsodPBU62XPNWLkMzU7OUlOzbcox6RzF8q7Eo
fQwmeNUuRD6FbL6FWF64GNMQUusF6qgrz1PKXQxN8AjzNFTYuQvD0nQsV/8SSFvS
sX4iNBVWfzRtezxA9hA4kDq8GvlHKVwYj5ZD+u4azAI9xpaV27b7BKl+GiznEuZF
ixV74mdin45muZBH6L6lSIQAXMoxm6hNE/pi1TILer9yCXyrxrS4uiv1TZy2p+Hb
gWrL0GAka0ArJTAqZMbTHuL4hTajs40v/vfCRHt0VakfeRrD4+w4bNRoANclzFV5
1LcZdh2Ggb1KB+hC8Cd22h8LSv6rC6SSjh1CgJH9hCiHeNB9fvaWGJ6rixzwDof/
NG/3LwAajsQ7oNg3wc9uqJQJ7tyjFw8bgiJDrf9ZrLo+HxIn8CSRKdZpxCPpFxIG
JQ7fs0b29vx9mmmaQ5ij6duO5/IJe9qIL0ynFdeSKU/HxZR3ooRoBoy+hvSlLCmN
LW6F9BXCgYH/MHJgWN+IsjK16Lyc7rkgFDCwqlQIXJAVjodrJ6ZgFdve+K2P+0cc
bQiXfxyPh9vgdXpVLDpSDVUMafi7et/g9PzBeY6WFSpi5sF0FMoHg/ysxgEDb9w4
aW69/jkMytw2eLt7lbBAZbqiAmadFQ82Jl4ZMFsrW5sGUQsWzZ4+CZvFP4IfqME0
YpQMC0JzHInZCnx1i2w5zCXgQCNontbfTZaBZ9PYd3PEjglKN+/07Wb4NyKeeJ3v
uXrlRP6I7ahH5uyXI9AWMGsifRo32M03KWIncuJSm+tUcKAhPZBJ0KD05tlJVNMA
ZwAVXKCbc410yBauAgZRjt12J3B0G/v+BXUbypX4hKqTruq6S4Cfvb4V+/aa9dMC
ThbO2nwSzqAjisHtBTwLrPAkzpuT6mtp/gbWKzpIJV6SWaHRo0tZ/JkIDoIxOzS9
PJZFS1qweCJPcKLwPldc6Xl39TTw9LllnnszpXhbyYPMvop3A//Y2h4sQ3iB5s2v
mJbIdQoOKGngGgPa/+tzXEzQkcQ04oslz6LRBdbwfuSppAVEC6hRC5Xxgh0HGHsa
ZxqDz8PxOR/ChHM3bvA4XjGg00vyFomBDtEqcEgp5aS+gxcns9XiLwRw6UD9Rdkm
`protect END_PROTECTED
