`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MD1InHjrI0+iyTxdtQSv0ZHNUnLRk+Svnb39pyI1xyY6F/f2ztvjnWw+SF14Oyzm
/T9nS8if5u1bGmnQdmVHIp1uin+yLfcXG9CURU86mnAfSdLG2SyAHVTGasFZ9En7
JjbSWgCOPNdcxjJHR9gwP8Y39e6QxLHTHecK+3KtZ0qozIqm3FQYbs/WrdlPGYvC
4TeM7KF3Q+kLIWvzLMVuyaz3nY0qHpa7zmVkDG3vgqVL4/uyAWILJpq/uVqQlrVK
ZWsO1z/MtPGTwkpfiGxcvXn1q24mcsniZ445LRkRl+4=
`protect END_PROTECTED
