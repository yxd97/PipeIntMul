`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IoigNCYxZeWYer82YrStxBvnLyKs9KkiGz5h8/Go4DoFAp9wIfwq5CyuwI36G1P9
aIH53JD7ThkeXLoXxVMHgDalXaaU/NsRM72W7UdLDGrXG9lJfl9iugTg6gQcNR2v
rYFlucqMl0xZTeS+desLjD/1bXh1QOxTv2KzpAwea+YTXu8u0iXBBhZ8we/llXl8
ntRzoTrXvwhAlBE1EcG1/XIPHtESSB74713JXRmwTqw37205JKrEO6ZquHgmf9p7
xf9b30fO+kw7WBliBmZ0bepYdyfC1sRAy9hZBK34bqeaRtWZER80hEXZipcQ8FJS
tPHd56cYCrRQKY2OqLNhS8XtASYIav5VictOxO09nGUqt036kP44r1fwOVmw9MsS
vVBYOmn0ktJ9Y2I2JKeea4Dfx20FR/3PQCSmeD/XONhF0R2xoKfFHdTMoTpl6QoX
NvB/rzhJanpK7xjOTajT9VioKJjOSLuxguVeBOBl2sbaFRsLfr5fj4uDU/ai3s5H
2EAg74Hm2mlQmLdcytgMIQ==
`protect END_PROTECTED
