`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ro39vIG8Ra9LCrG/6v5hBGuXdeNgSEjt27uob+1CWosR4ZKsBQuPLznnskR48Nfw
lrw8WChHpzGtOYMBkXjzpXkeZ3nSclRQeaw3XF0CZKxtDXn2WQDt5uQ+G3zJtlcU
AXDQ7zcadVczgzhn0PtWaZAGBR8A1MfQJFHtEi4787PVMLvil6HlZ5E4m69IbGIU
aC5ps5XbMZfvA+8uBM17C9+9Q9/iYLWW9o2mAfdbEcgjDLutulT/AB0ZUSUXbkR5
QycQRyO4L8Uud8vG96Wnd/CknQKnAbb1awh9qLqkDbEaOJvdd5y8oE5fTTs2BhQX
dewpUgrX0ZXyQisIvEbEgkIjs3fZgodql2PNUqiylF+kjsy3FGErpgcqU7sRw6ir
iLeBCpQIL83Ht31zxTqpE91FUYcwk18rgjR9OgMRFsCI72G1EqFDmqFYa5bwfKlw
nZOiNApQqE17uVU0sK3cQda5uzJxA1gVwR9H4owGYCfZcLNWgCyxyUbnCeP3sWzF
ehj1WM8GzCxZFiFjRQSNV9+IoyEM2ES7iVT8QW4BwvRlDgjaWcdY64jJhJw//okl
VPegQAKbG1JFR9Ox1mUCBgLYhIk3ZK2RHeYFxM+OwmLoZBspObYy6VlYBAkytEmV
ZRWzWbj9zbRb6wiXhQwl7ZTE7wPAYnqE/M2TWWrzDUSbey6sxIZ2GoPnhXRsF2m3
8JrnJPuktXjUIoNkIAS88Q==
`protect END_PROTECTED
