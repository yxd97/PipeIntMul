`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
92mzinEjXk+zqzFom3Zn2h7ox96SUYWpLM2Qvs37eH4RyzagVeIClB+y64qUf/o9
oSRolPKpePIapc0zLi+bZXFhvYSLj8Fg8qCmG/yNOynGV5F3DibkNd0ouNHP9lQQ
CNDt2CMw04uHPYqrmZg+CGF53NR+h6aQrA6GtETgSKi1YAxquv7k75H4aX9bQ78o
MfQm0VAxlrSMtPrWzTPcqgq9SAcD7SyaYgoUtO9+LY+wFXjIZkG1lNmB75843m+u
NvrZbtAmTXjofr+rMRK9t0Cwiz28T5w5ave+D8g9cF+cOclrZ7GQrl6XxpLFr7FT
dxB9q96jM1B/3XrmjF0Nlh/Dj4gcw7ThGaoF5a93st52tQcnulomgE/GDJtpv3LA
3oipCMMZCfRuBEI1xyapgKwDRLG0F0VXDjXckBLTQEcyTNHsr1YTj6tyi4ECdhhE
yHWNpjwBwyG+1ufwvgXeYXZZTG2frMaw4/dFwAe+QpU0/CMrRID+TDTtc56CAnuG
tU2f9h+rJ45qi28SDm3izCtVp6PDCxxIDq1SlnUaBWkEVF1j4Bd3Hu4wbTQSFGMT
fTtrH6e1zbCnSpvkHLCOzWMyO3inyQfgeF0aYN8bJ4jsgKexvYAQcE1gK06qLc9S
3Gm1n8yqfvmvjx67Q8bfcLlF1aCWfZNWppc5Xz3xYhDkGju54hbv33BjdOcVG2WT
TcD76fO3NJ0d57jmq26DpKbb2kaKK4n6tZNfMmDR+wA50dZg3k980VrFBHdxf2gm
PvV4Jn90NHCNduLriy8xpHtG3GBrnliQRNnmADJvQxlF3jWTs4PX/2+g6dsNoIhM
GcMuBM/UZ/Xvn0mHBGawOuwwpQEoca0QFC+YGlwF0DDTOQoJtdzaWkqlfL0JmUaW
nh6+XTuM5ZiqWtenuMCLm/FGQyscSzWmJjdPl+/DRjEkHacr5p7iJWcQib+DTmD6
EsjVn6CVtdsEfOQOOoGd83MkrMjtD5/TxRFy9nT//F3VKC4fnb7Z5YsW/p9HzQHc
dcX+hcOS+7wuXSOx97Pm7BVNneIJDlYbJxMm85zmpV9CllqRkwyMZOsrvP4/vCVk
wrT8xd7KJhkrMDImkAvs0Q==
`protect END_PROTECTED
