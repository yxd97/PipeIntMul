`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4duZRKsWER7BXofJtVdFDdemvS/8wy5F76UPK2cE7fiNiL20B1lKJyNKO9I1+DVt
q07KygMgajiVDeZTuDqE1M9zWY3nGA1+VPV8aXX62JfnUEOhc4OfT6DLTjy1Z+7v
DxlmlAiE9i28G63UJgaa8tmeY5ji6+VOmXvoh2e4GB+hLmMtraz6J3HTMSvrnVh1
MJ8XciDtkJBPYorX5hvHY6R7ts8OJguGNniJWb7C+UKqgucdykrkgx+GdYv8j++V
WHA6Jr4Ke1MR5hqYe12QJ+pPmqFyXl3v2D7lj8DEGN+qVX0crs0971A7uoITN9zP
5oKnoLeopOvToxVFeLd1qp6X1uj4/pihPnGY0+NFsyP1Vwz10sibULNRSx0/tyPw
wzfYIi7MYOIsOBilyzluD9zc4Jyuf1L7ICFDrCTrq8xoyXVzEXI839OJ1kDwDzrS
pLBbtbSLJmRznNn3YkMAaOCBSPYXqhFPzwednDOkBCToH68/8X+HYCbdAoulDf/E
PuapIERI0aRNptvoNIxPK0jUydjcOEkHv7Jwrb2v3u8XacIC+zswGIC2/V63kVBJ
D7MZgub3X9Yae5aAOOQ8varHbzqszUHpIn9/NIaA3gcZo3UiMi8W9A63GuOQdgtQ
lvyTwviDNDYkuR/W41lAo4p8KjI+ag2P6spLa+nJmmx0Waskczc/9pt+nTYeAiaB
zcsTlVk9Nuo5RIZhdJ0E8wyqXikRDCctqh3zb6m3rO3rjdtBSnOzIe+9xw89hQ+2
pg3Z2fp5W5aIVgyLW2kQYRhx1HTNyETysm27h44DzJ9ZX1dVvm4YbEaw0MgS/RsS
+87UryrY5lcpXduJJHCuVQRI2Zskr1JhH+1rR61fUsJdH0dX4s1EtkisZePyyKkX
ryyPh0Jvdt6MnUTcMxHO1tgzdNGoYSLBC877zFKpvX3XQz0lDvB1C6mi+saC93EJ
8yckGezn+KGihQuxjJQukDevvan5xhY8TOYcQka5Wck=
`protect END_PROTECTED
