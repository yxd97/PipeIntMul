`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qf1ib55yoDx06IOWIPezRfGhLS/CzECMe5hnJgN6Whv8IKNUJBDUVV9TMij9M44X
Lh5peVNBZSjPA1DEW+APIgfD4nCVydevJBKgxUTBp93lgXXYJGt9uHgGO71mfrJC
dPqER9zrucSyx13KwUrLX5olrt3JKB3XpNCe1V9pnX75DHUHfNgVZqO1HFy146xH
91ePv30PHzORkGZzE3+8Nln40NnKANrIQIj7ldAGPw3S7i5kn8i0sD6OrtCnOVfc
4moglBkkyXptji5GnXkyKLu2zT9CEu3nxwXCSe6XhHKLh60q6ioJGyWVdy1Sw8Rw
/hWtuRn35VKFQrcBtaCv4wcj11hRMlBOxqz/xAL1wyiAwzv4YNj3VNSpAXGDpC2m
WmW6F0CKgJ6qGfHIV4lAkbR1t39q34zke1E0ImzUcnONY/3SrQFFnsKF7cg4H6sf
5XfCtpkLhmx2wnTNhfcYIMVygJ06BzvwXcomGFtEQRKswl5RcTYxg0an6bbFVvBG
gZ2sfHh7QfykDV6y3onxvimmEk/qTnNofnAghsnNCZlEZkUjEra6utKtWuIn3JIU
r2R1hNQ5bVm3N1e2SyOxa3su28+gMhtvwm511xp/LQ4rEm6UzqdAOSvOYNnwaFmI
x4Qj5lsG/h0wSqxe0M94EwvCvDFHOMcxcPkuxy9FSckcpKXxVK+WhKXUyMOTmDmw
QJvqDCG8BIJnHPxJocjrqBwXamd8uhejj810KCmsjOAkBTGvqsw6VlVjLHcGf4po
PN1C/BoeAESmqs34Z3DM1l3wWs97TtS1SMcJLDYnwJtNbc220nWaejf/6OyAsXT2
0aud62cvfRZzQkAdup2LNaj//bqZHgdnLwbbQkWBwAwwAzJ7DytP5G2bA+ut87eI
FHb+BhBWJnsMg6tt/2tJEQ95KAn/1OMcBbMIwcCUQEUzn45a8ZFH3J5wAsxQxrsT
`protect END_PROTECTED
