`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I18ygZ1DAlw89HkYahk+lnuCzfWFCMQHmKTOpvEHdzf5RFRXNy+1C1YDmjZY/q5v
1pariicYEChg8EmkmgErR0fJvHF0hyA9B2rLY32ZZ+FM97vPM9aI4NDsJ/8qyBif
GPaOPmUdnRLP5onLNlkPTMGgTqegSKPb/aP4phxoOq7YB2Kg3ZLRBrq7OfHeNzBc
Zw19uWS9oq7ELW6m9cmja4YiFGwPyyNV+1kaK0jMEUhEugbLcTLv9jDxyRg2Ifti
`protect END_PROTECTED
