`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Z4HCGDiSQfPCMtVTFQt9zxvyD2NrLypA8dLY3gXgKs1IOhrlkLKm0d7lRpp4U5H
C56PyGep77J8Vebtvtl6sKFWc1gD5af6/kiI4PfEvdcExbIWHefP21m0y+mr2tVh
nNdyE5/MWSQJ0OEG6uqd1R5DbEA5MEeU3EKaZWbwCucEH/Ykte2n9o+n4SzpA8tS
tiT0M1H+0Xi4VB6HUbo1lcOsa+QhjRySGauKkizZn4YWBV4ZDnEHj5aPKQkeGj7J
Qra/U+AKEOFycEerhn0NYXsgNq1whsksO+MIfwFThq86dDccTmwtp+vmU7kzSO4d
lU8H5a/nJF55KJA1GmGZts9sQ9F8WUsgep2Fxc7emFIIDzpoGaROC2AMoz+9D99j
8tdqq4ZLkAoH388JXsGi+Qe6aAPvwLQdxn7JAt5yuVeozBbd7DGEsxIeeNFMhMJx
Rmg8QvKk4XsKTWYWyQqrPIESWhH7EqK106/VpV1lGLzhLNEW8yUMDqCf+Hcupw8O
7dyfUcSyZTSipQQtHpFWBthA52wHfJNO1E1vHBpYvdZGL227n7VsTJs3TN2Q/Zs9
4+9rwo7iNx//QsYWTYxWtlxwRplogL3mRdlt1YZ2dxp00gYAkj1XMJhXt1u2soyZ
phs/qzP/4Jw6hQKZqEIIT1hEvfpY8I48vB4kvJeXBGqrQySJpsg2QBZmD/reqVKG
MIalKlfvlD2barKrFEHqAeOH3YluRlbf2WjUwW5mh6Ex/vCWw8yVCmXVh2IKeu4L
ukRLHblHBap83bZHrIMWfZG1e3fsSlzmglGOeYh3BvbD3W88XCf/TXWBa3PMMf1X
W9CkXzDn8eSpq1Gb3bmm3BJxSgD0b1x10CQLxseHZrhVA2FtvpVZ5P1DXrhGaFw0
n8WFIwuEEe6W51Edtwjg0PtlAhPALlOaLGqAdCBbPdWc8lJirmFtwVeIor1tFOJR
uwxfQaHZ5721aDM6RtyZR0CFaCN5bGvM7J84mnSmheHw4FJkqpFJ7oE7cyEWfDzy
i//7GkGtCKmKoCSHXMUaejLlgkeaDAc9MC98ObdCUNwOZR6JUhyvqVCRxCti7uhQ
HpJvpXM6BgJB12WYejdgpbrZYZ6imFQJfUAHYl7vKM53+GP0vSs+k04+HQelGGxE
3s6zh38QsLYib0A5p8yCqZFAdmYFFOnt4+PhUUfdPyNmLYEhR+FnD6+l8tZlIFLC
kiiQEOc2HfLEEVzOzTxJYYHqVnmAHb1GL+nwvm5GQBZUYFBB6+ai+f7nKdnYebQa
GqFX/NhIU/Ts1O/U0JQyKBC2lyerQ19lxzK8W58+tUoxEZ4ejTQmLg3PxUDAciDZ
IJPtEKJKLKoSHHeycbt8MdqqiezdSHfqTu2nmb9sdwSrlBZ2XurQh29b6PmU2sYt
Yi7WE5iDAd12swleD6sdXgZ8h9Bdx83VAVdCbtduqoF3sODREVrDbx95qIfs9wAv
xKVMt5m4YJvX83oMrK+7EV2AN+bBbTBzZwB+KPiCBtHawHnB0LlxgfOMzUrFQ7Cw
9XLoW7/SJrfFobPvEFEz1ZgxHnS2OZBxPuh+/TgFHipjMfJ1bXnrvWXqZWNQGUrJ
6e9oKnEhfrSb/yijtHbjocq3Js3dZTm19jGhvVs8Un6GW8U2q567f3PEZ8LTug1a
TEuPk9og6SYFKMQ1Y7rtQu6OUdzeWixfbBwlalDA8LKP+Dzba3V5on/Yz52a8sdu
pv5CI/cVNPQU6U92N0XzD2M3KN8/S0hKnygsy2Z+00Nxbg6v8QvNqtGrggha3lrY
6bpJXgMGewoa8eA8llxrCtmxSCoVKz4GGnrXoF7n1W7AHte1lyV4Xpo3k26ohCUm
xPKbk0XdqqDEnF/9afX0efLjSr3h4f8gHzdfn3F9sLL8ZoOXsHpw0+Xw01/Q8Yck
EQNNv5Fv1cSbZ3tCpICfdYeNUaIB90d9iEvGFUcd6KP3QU5dbw/sQqfFO0bYknIw
Q7tXBbwyJpnLiYgCkih4CL4uka9mGB1PItxcX1PFeh0j+84JotS7zG1vbgzUSMSb
V8OSKmLJRoEM8yO2vJh1I8F2mjAnVk8/vLJPDSFmN3rage6sVf2wKRLTQDZ35LH4
w7IsxnsfeU/2V+nsWz1lahG2SSsJfINzF6UGWN2vL9LFHtLgc7NfgiwQur0phMhF
GhTr2RlYVoRaUhU/NMvT9tRKgzzgC9iK9eYijYENdPg=
`protect END_PROTECTED
