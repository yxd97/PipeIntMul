`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8c1akME/lmzpIiuhvlM8/6bks8wgFWBpnoi2QtGBZ2SW48/5ioO8QVwTOS7A7uPa
bZ/0rH/6FgqJ1/BxNEFAD1U2c6EaZ6xsRhrHLD/11s0WWjvK4n8rTRo/17GFzK5m
ipANesCp+W4VLrjIqm/CUM5toqq/zYiYkxAdsdMp0gOkTqswl9eowrn8nXsciokQ
uddzC+H0KyJ3KCDkJSG5AK/QufUFbXLZR3D84GGQCoWORdR4F53r2wY0K0en8/sV
WnC6e+qHs6lX179J02jETTl7ZDydf5Zv17Dkj3vuOHxG41Xmvcg5hC0pBxBgIr5M
f5wIKzRvdMTDtBKIuIXUQE4riLyYt92ztlLWWpAKILIA0NEQEJruxEURDOXSaYSv
14v99e5aoRDycZbG/+vwMMG6sjYRS/tXrR6Ji5P0C8Dp7CCrPHNMhGtNzftdIU75
/2NZitL5o7tUY6ZzoJ7EFTrvbHwgYIr+e8+G+OvQBdbuy4RiKGjQArEc5KKQmOKL
fAQ9JLpKpKqlpNAFMuvPvdkQFF+tyZowifS2YJ1mPT8M73kZm7RsnV2rr/QbbGgb
rMtKISLUweFR6mS1G0ji73bqUnDVFha4ThauH/mALItmf/U6aK2wJRzmN02qEkQu
EYl2bcFWRKgGAYg6nSAUNOpFuzhlcuWLplFBTGodvx7xG0cMBVEO87nI5QFFlLM3
ZrIHpQlku0kiTIw+sxmuekMZtcJ/bhYcPOzjy0inPZejb9NwpMDHNqm7EtyycLg8
i3hA0SGTW6ha9Ip7LDikhuwWrqNtCX0Np/OgWGu9pMyAKwkfeZovj4/HWDUMHNgh
6epPyXWAyP2qr4MXxfYOUMPuPVWXRMyvb1Y/twHM5yxdh/gBaILJ7QEzrT/FmgT0
ZzNDayOARoFfrLaQ6CRwxudgFAB28DGo27DCoW9Nunwx9GfaefrrmWuIq8Sq0El9
9EYXLu7Q7iJRjerdyXpm7UiCqWfpcDAOzxAAbkgIU1EZZkzx9ldEXbcFkiN2F6NT
bmovN1UODH9VFqzRxRHGJpGr31CBG3DWuhYa1/7AxQIDSebFM2xQuFHNbUmSIOzO
ZQu5cueA4CUAGrUhmKiXGoDwRfaMTvrHvPd3cyIzSFS1Yu25ZoleeAYqb4N1qGiH
fRYBmQsoMooQfgRMTn4gWIqgJ80FQdHpZl+tPpkXuOZlVVsSY9kwLhmXv3ec7X+q
kpDZoprKiei4mC6NArjl9/RuuU2n66ic9AlMS5VSDkHjx1evtDg8Mceerkb+uHW+
q2++DOc7PTXQd59mVCCTJC2RnCmhzTgJEVcVT3Xy1Xzw8grE4VzscJrzVtZ+YBdo
4cvDpvwiSgxNtiyIZn12x8Co6cDGmS8VOTnKHrRwrbZM+bZfZfnbtFjEAr3nwG5W
YQtUcFQAqnLSr3D5rQAV3EZyoFe75wIev9rWnYVLu4r9IfwSsaPEPrZt2bz3LSWV
s0aeBf/Jpkb7xM/UHjqklcVADYHnHBw17JtTagc1Tg8xPd93IL7FpS7vGtY0kvoj
pYIYxW65g7ksZDvtAuFXo6bVq2tqj9Tmd3Az6WHJGYOmXGxqOHsiKSoX9i0nl5VA
35xXXjhoPCjG05e9+ZETqxyJLhfJp/1omniXcTwu5HRYbjAQM4AfyiuCHcM0dEQw
yElFkApQZHOzs5yovXXLWq8wkqUn6+uXbgHn0dzdpAJqyfcJqZQuQ2fCGF3MGKPW
2d0RHePs/T+9LEpGA99qN20b/dkPwSQHFIk7dn/souScBbgmxLTKK1MfoJYXOqs3
qyy+Go+gtRNx5M5t2cv5+leOSMHi+fZkY7ixhtOmitIeRp/mk6B9NhDqNXiTMxg2
xqt//AoHJ9cB7WVDifjfGqDge6xJup4Y8lB5KwtBE8gaqroDyO9a9i+vPpz/9xRB
i3htOXaEXWPl8wvA5PBvuT9+R9PGwwxea5qr3RLW4ZGDexuKaK2LRoF34R6VnzQe
5bAIht2sJR+6tQeaPc9EHKt8ecd923OmEeBUamCHXUQJcptkhb3A+MTBOHv+4sSl
p1/+Q2xp7JE0IIgDgakZTfAgrpyRLttInsY6IPkCNyRSF77JPDJVnhGDU5IdGnvF
qtl7CN8j/cumPsTDycA8qJF0jVzfIK30ViHHJpXY9m0kMG+60B9pw/eJv+03Mmla
der+zfRAO6IZ7dA7rBvxE4NLu1kNu7OAQYS4HxZpZQBCNGkvYtw6M6cPvOR8Vn4f
t5LrWHeD00zqfz3bm3woMoPb8hZQ/1c0flfyFC3jo0P/fH/RsVINbuwt5MdrklL9
Ws80rOpuVTFue1xM9AajRkrwkPyucYZEPwKeftbpwA6z/zLijnBrGBfgdt/l2VM3
1ilRVy8ZK55/y/zjLABRnOH7MVfZT6uwsxcTdTTfI8qEGRCjUx2oKFz0HTuKOa7v
mmLo2Hd0ZTY0Sf/pSm5DcO51KUrnvz5o24tgxnvndzhayhOGxugUufTg9EXMkcVd
8ahG43KumAeMsGJzAYOzFJCO1ciZWsr/Ki3NRRF/p8OBfohd7XThj1FpuRs5c9Ay
T0iSGT2sQtb9naB4ZiyiVOz2KyiiZpMUw9//Y5ek/50eJ/m0trHIDT+L+YUYDaQq
0mCD6wlrjLh6TmAxmfRsyjliQPDwuDWb+XSMTYukjw46CEbVZ0gWxW9sXPGBSnCk
KSEKNkQ9Gg9jHz4+hzvxu7fjaoxlodnrYQ3fbI8lDPB8rBOgwX/SezeuEZ56Nslm
ql+EwB7xJbzzkMtMxiSyIVXRlVwIVf89C37OuZAcIURYz77wyFXQ+/kBNp2fhVwx
jvu8W5JIniXlS2fPnNvzPd7MIzxHegLaWzSxas3uRIIhvNpE6X3zxQOdvegnBDnV
cl/LrFsywdzTy00ChfoGWR/anD6Utei4koBxPsYA9Qq0SvXZ1HqMbZI6aKUFaAt3
LcJAasmbiOdXCyqiYKJzLoZEAcZtRxIOVYH7PDmxF+NAYZ2cli6wEDIWIVNkMTAP
SLPcY0+r2cYgUVLBq2rW3gtkawHmBr8fBKwkO7E1MlkKkRO8j3EbZgGQ5WYOBz3i
LrVsFkLHBfBUuj+Vn+rrEq56hLGQQMNtAwQ9X7lIfkjqrouPu7bvu3RX0y8wfcLU
fZHOy8txagqLtHGnbwC1rwQPk+vbQRGOvZSWzJtlNLt4E0E9+1FzSociigrV1ss8
uz/sWNGDa8lCDv9yXPbDdwiE9X9JiHU963nDuvTuBaJJiex827Ulth/JXWsRXrXY
NkmRDNtceoQLMZTu+GdFsWNg911Htp40lzls0FBQ3kz4AYVW5X362WmS67RX7mFC
IOaQspObirF+qpL4FBmYYFQ4ckwUTEVThIUTmvHaMcct48yMo7zkcieI6FeXeVVh
87wmJlq5xbZfOUu3+wc4HkgDM+pW3ytuziddIQl0WIBJkmjZYZ70lRPNvRxWr4MF
YGsH/LVEneJt3Lyzcj4VXtxtkOCFpDjoei6CdZxVI2LwtQ5yMlZAJlOTjjTPa9mz
V0qVTeF+eLfAhmKDAR9BRtvI9SiSCDcmcxOFGFzC+7S56dh5MlPr7oWJISPBddRa
lWm/XfJymZ953MWJrvf9BKB/neGmm5Ol7SXn9eoOkchODWIc7NHSTUWgRzYyZbut
SKmdRPulLoolQJolNUCOV1CZjcGKrLUmnkUusKO/CqGsZa9YzNED8YY8Zzxzn5h1
yKWRldO4s4Z0TYNnA/y/z4jXAm0pEgW9wWZXFcdUMVhZExmT+R6aZfVSHMlwODQE
K/R2GV58vmndZu2PWG49rW6C9NQXrymSwdjYqr+9BlLvYmCSrt3cEug+yHXhnFs8
nEBPgL16i3UvMyHwXvF0KH/aihl3r7qh9qzqLTjuAC2xdIw6J1r5uASvLdc2OVXA
BF8dQu4iZu0v6hCJxjwTatqXipIsxFnkWLr9k7g/4yMs1mTkEn/XDMVfCxP8tXDb
rWe/DnjCOtPQvp3qnp5JY56H4psVXBxBWfsgxYwP9606lcFdpisveuvK/3AntgVj
3xpEErA93+JPRs+0/Lx0NPUCoGLG4AC8+JEFnxBZQ2TS1E7rM6jJ8BDzE5PZqFXN
Xg5SXycFDXnoOvWvhcobR7Z5bktcDu9TxeyMd40wjWCqNSKAYtZcS2CRQzQmUY2h
r6Gz8qARPzs0yAaiUyphdtcRaW0M8bFWx/mXT74IIxKpW4YBj4MSRLVTlyRWZUvB
ryl+yeO2YJ2BZndIR6fQFKE22WC0b6PmZIX9q4C2cR6y1qq7Yizr9MIMAZJq3Ily
VdBxFZlmyl76DUMdoAsNQ749yLtr/GJK66iUX4jCTpYN6s/oUFqlNDGTZEYKa0Z7
mpR1hYZi2YhdMIn9WVq0AUfkU/cUDQJdCbaYGJ89CDhFjm7c0Q5rpJ3b/MS3VkDw
V2/EBNVjduSeKvNIPpmN6h1ctKPquxsUWL2MwZRJDH2rS6fdGwkDHb0P5BgJ9EQU
egjY+JpVIHBKtPN8ROV9lIJR1wPTTls5owZj96SHn8Ae+41eaYafxiqxNkIegNo3
gSm8NkMitEYCEELNHZDSr67LtJjEw6vDofc9YiLpkC0nWPBSo504OSR5KCWbs5E+
T38fCnOLJcWftEa6eRxt+IJMapVFNJfBb2vvDj3FA+t8yqZjBh1gvTEfwV4Qs7FX
k53SiAwL7qgeJe/hphhxG4Ilp3OCFtO75kTyZFKzQBhFmJDZsdMPyma+7rCUUsn7
P1fKY2ddU1CpXpnhekaGP0kS6Kl7t0Faen5fg1AVb1xa5iGsYsE6kggXg4y2Sm66
edehFqDWMY6Gf5vfnsLGOiEMzwyYEqlVgOvICGl6ytBRB3VUtcUVL7U+Y6indf/y
rjxy8eb8r8DvWWBJPEAPUVLK89PGE6UqmtMqQC+8xn+qra0Mn7QDCBcKOjtPjiHF
DyzxIffKiiWKXpvp3OTnyHVYgBD3mugXvVtOb5dDYnCsF3nLXbPo+TlHXH4xms8A
iV67+JCVTAvZW7Mbq+iQfHVhr7r2Vbpc5waRwPpCVmbgjsc2+QhEjzldfyb9EAPH
2ZJyohQdYk5sWjRl960/xXXlCUpBbfLfOnGIoZ+0Eiz5+p+pLhK3JfLJU/+diIYK
X5hpsXsDzyt1r1RlcV5QylWAFGs9AFYjYtwkepvgQOgVXaEtnwRQakiA+oUpRxX8
z19YOTCqdvAufw1Win5c+TPztEWaqpjWAP8/Nw6aEth3Ajm9G7+sUVMwQjrwEeH3
v+nDxve1Q5pgBm+nZQB236lFWJHNWss1Fj9rgZjxDhvDFd4t4OLCU62E6pp2Rjn3
GYjS229eHtUffv3oj/1A00/kVpdhLpwueu9mRO8eFKdtGjcGhNvVYJPwATBgj7CW
PEayXMCyZbF0tqbeGfXTPfXNNQvFOAU8XQDO8Lojw+nCX449btQaA7aBMeTRUWJi
hRHUhVsGLcJOLHND4UthRRTygFn/LY8TBH2klNrdGyFNqlZXw1CGVCFS/VPQt/xp
hsJbc3ZjitCEQ24kUjW5/KoKihSenGKwwNHaHKNl5xrNLQKyCGV+0LZCGCcRIz8E
YrUJIu6TuNGLspFinbdo31nbB5TAcpqJrksIcfGfpd6e5rkhFleNwiddSp/Z/8Fg
JzpXabe25UM7o5W06yiyPlJKsVMUoo5gL9B/SvJIbtcrfYzGSGag0IHL8zlW6Fvw
SW7sOr8+XRhqvmAFjDMzNcFgfyiUp0iMK4RMFg2653GmbB+fR+GFeAgpA7d9+46Z
nckQMdx/ciVmrVH9sLdWcs8MqHdbbZXkL3c8FlCiCJDBPv5n9m4t9Nz36kkSpOM4
bLt+YacaiEnz0S11bys5SlANkSJ/KhR9x6aj5ekts6n1bgW1VuZ2bj5o0hANFeyR
arGnLZaGl08jGRWEU4J8KDBv5bSmJa9K4K14sr9XkBCWGmu8QV8T3Al65x8P1CF6
26LerAI1gOSKBr6AQW7H7clQVnzvgP+2ydOAn2cY2l1SE/yiXC68keaFRmbG2gVW
1+vR9H+MZEOgjtb8WC85pyxbCV4hdmSZIlplSSiZ1ipVHTtQcXGqIBy26edmTNQS
SqGkWUVdRLNu4ProvWe0J/Hd/KzRwU7nyN+Ez7HNd3CS52RF0JP+u8EAq3Ji3Ri0
2ekTjyc6RFhbClhTD7Z4b5oaAC7L8HS1gjENzycVlnjqNK9tqIY5zAza22SSl9uh
YYssiLUF2B9FGjB9sSsXHZMUK8Ky8JYINV6tlKem3zJHa3k7BS+ctbbF1qyocnie
OeIF89srUDCc4Pwp9W6JRv1rEHNcJo+ZNKmMAwjilK73fiZp4bzLzfXyJqnDDQOk
1MQ7GFzReSSFXvvziM4d7t/z2Je9s4G/MhES6x39dM/jgiIonhu6CKaKV1l21BVx
AjLrmljT0OwadoH2VzgnV8p0F5eS4W/gcovms1ARSk2cIFbkVxqPf1IDhRnXgtc2
4eUT9AW+BxUBvfQRk5cM5kh+gowL/WFtrzRHyHxIqakPOH2ztU3KL10eRJGv/ewk
ndIn/gwOz4ZTmGCm4NL+Fjt6mJUVf/78mMN6gqHiROt7ASEUHHbzthTwOdxd9cv4
PRvTFiWdLvL12Y33MgRp8YrqfQ6O5gB3LOLTv3Evkq8KUikkVg0BQHFCbSnlrLvP
dXio7t4zn1zu9wZL+rq+3Y6x1TGiq+2uQAzIAGuRgUhPHHPrtsOi0nygZB7eOkE2
nhr8xvY6WiCK2qglfPNGjFyA3Uz6dx3GrzYvHxp/3oM4RD2QnTLVc9lnAbhXpgPK
v1Ol2mW030+/wf20rOVeeBsW7gC69Yig3K37fH1y1gO/9NNkGmcaES4775PolmQ6
f6t8X4tcL5BzX7dSsIDs64GsDCtr1HMHOSzJYW5Eey1yKgcJpVA++cyii10Kff7X
OMosSTaL9MaHxmwf2BevMRdZKiINvHn+TfmKprWuBTl3968prALxC4ZWslacRLv0
qSlWlHSs5p7i8+y0v9+RTeohihmn7oYBZ8DIw3fQRSSdya8EdWLI9bSvP/kNHR/D
ivh1d8UMBdx9eVqPk8lKaqf0fWbFmvpjtYLkMoSAMXRC+BDBz2TfcGM7+TftVcxo
X/bSnDc6uONE7DPnMG+uMSB2XMXz3ZXZp65RhQWL7/pvD0Rw+ILTCbRmGtiUu2AI
JVAy/G5LPgv70p31vToWm7hMPZzW0QSJMcqQ677WMVYdfssOYxZOA8eNVQPpNnFq
xzWSnrGePXBSZRjS+FUBixnDPoNWLKO4NVC3shtr5Ob3TaQMgvjTIC03NorOLP03
QRnXw1WEzoXm4/M5NsZM8tV4wwkIs5c12ODOMIYmzYa247yLIGegvc2Fdo+qauk7
2/kBIndDoT5cZr4GyVwmrIxNXPLQpZ6c2dFRjCsotUr164aW8Kjmb2FyD/Oobm7s
/PTNN4dlVDbvurq572dS5QpJCIoP37oTCmFZjVB0swMGDptFHytcSgXNMgicwVcH
7z9g9DRNmrecmK1aXfNbFz+Itk4+7y2lSAxrZmVS09NEC+9V/W3lh+ml0wDiDQHh
FRz4Da/HqAVsBWTTwq2yx9Wa7h4ClcVAbgGUqJ8E9ts3+3K/iP3aMV1ERgaIMbl8
0ask7Z5WDmR4asBj6Aboz8FTnQFtJiQhEokhoNINvg8BPxCg8auJg/Du7FIO/h64
4IMMEM6/FlE1A7r/U1NUqFeIGgNxcOTk3nA+OlsuceJ0e3m//YObXbrgudVIWrX1
6QSBhyDWY9m6vI1JH1vyWNUB8UdOHVcyiP/YTT4hu2/iFVl58r7QdCLnjCL0bZ3E
LQbCioKwNfxsjDOGJta83zY3EjzEnRCIPGCXda5oFnyy5p5tLBp97++nfQf7gqYC
ybew5mDJbhxY6G8M/PjTlv94P0ouwiZc2/ylzviW9rfgQ4LHAU8DTII27RwA5DhU
e/0+lfFZhjNljaJywPeyjVghtFnS9fwLOaWXU/pOmcmrP6mAdoeJB3pq0RunP1Q9
1wmkEptWpb7LXFgGZ5xtFJZ1DMkgnk9IPce8CyDKuyf0VC/drvNIxxWlLC7MMHXY
+Eibs6jC+BTtcGZUpVWqrUnv1aPePIQPTM9VT460vqtQayG97eoG6Yp/+HY/smnD
6K2UD1PvfH+AQ8sdSvRla70GpQrH9LXDUpmwUHIm/VfDk9Z6i6JwkOsHKZHtsGSY
7U6Jxkbsc1Epudvr/Zla1NJeWRt5sWBpf6GM7CmpxzIrpKoQUkNXc/v7iwSYQ7rn
wIqDlreRe0XehBifeSZ3SxXjb2IXxgtsIGgXJR/XimkXvSxwl6/39ia+WXzyoBvA
xXI4oTWnxzzAS1fcHjwjNtIAWaRpMgPhHlV40bI0Nb0x02TVd1A5TpratyLpKlxl
89Fe0fkiOO8O1jAmW7mjaQXaZ3PTZLNn5zL5JmNxl0cV2/WqC/KGNudy40IeCk6f
S/tJvZDvDEvGD28or2w2Irup1vjUFdhUg/FEFWGpoyFLigBfvkeKVKGk2zgxuUBj
TWouUFgcJGJ1UKD8ojgVzyuxTA7hznTxxpxnQy2mKrF4SibD6Am0sSw1LRogblVQ
DLwp/2mJQwRxF9Z/L2gJM+6rtXzkCFFWENk0izSNQe5xfKKNOVXw/CDGCvU+CMJ+
Y5F1efETSlcfe8JQsFm7GCfwQ0ENUwmQhon1WeR4r9/1QRFA7kFrltamKW4VCB2P
AtL1NvTgcK0be1DCR54xh9oaOB252X/koQj8IgfDF3N8ltps5WLskg3WLt6VZTaj
geLOTCGs8Atc+zvstMQa17qFUPilYEPObqB1Q2GNyip15nVu9rUc7nQfq4r5bCB4
iYKdNTOeuuYlrurIA+EvovjwdzrkTUxYhuNU2EdYfmwhZ65aGYHB798KZNegkBtC
zFytKPe8af870vbkOL/MNcBsh1VSgAnJ6IN+HVjM1zlQcd9wyC3EzvhWYJr1nzaW
5HNal1zUBGrg1gQ1T/HA+QczioeiEkMkdcqPRglkfV9dLlUPwfA33m22guJHEL6I
l7jxOCRPBAWRX92SNS3jdHbye4Jt+Hw+Okark6lYiE5Z8/eYg/Owy+Jxc3Xz3AXY
ia3S2XXDPCVRm07WPSa+mF3RqQVvHAHKRhZNp/wzHsJ9xlJCPQc8gkBjQ/HbUi+/
b2/48VFTQncM84C/vCsd9q84Jdhyo+/nvJrECkFpgxxTFkRdbkKMbyIs4ZcwrOls
Ygjj2pHGw8y+jPeLBtSewtALsWSHB9vF0W6t6a+ldleoWpc8Bd15HxQuU5PLEI7d
vjqAWZPqbzup9gM4R4dfh4tRFSION4cYvJ3JUjTEH92i/M6TZLyQBpVBJEKj4LL0
rAN/EmjT5eCjADXDtwP4t8NEIapZLy5rMiyc2y9UhEezgUxJ/q8Wr2S30+S+OkUp
297j84ayRfFpmjIth+9XlrXWnm+dfm0yHCzMuVTAEP/SPeJrdU5+rro1DaW9MLpZ
hTNdNj5t+LZ7VWIw/ZYDPJBit8K0JS7oJzvhRNqrfCTtPXZVKF6/otXz3pSbz+YM
L1NG71o0eKJOoAjuv1VQtKkS55bcjHaxsdXOgmWQZVmjfbaI4d01z+8qJqNCDH7u
HEe7SbZwebJNP06n1JLH+7hwkzSk6xhr5zB1noIAr+jGiT6otKElsitpItL7Vdlp
qo8u235b92nG3qb27akHc3Jo/WD3C9yr5Crt+WW+QOgpd892D+YAWCgFagHh7xd+
MtR5olmOesB3LEQUaldeiLt0a9+h+8kj+MroR3mMBNFY5vb0fMu18aAHOkTAQo9q
Xa0J64uEIY+PVxwadZPwWNQQxycVIDXKBW0wMF8zfbNmZItpNdhebh5c74S0bB0B
4urfNJjhOjt+teu6jtkeWmrzmOj5vA0W30LsJ58iegUPhF2QwZSSSyKhqUhnJfcO
QtaRNW6gfk+iYAThrcnlymr68yVZGCQZXlufugXeYxvLkm0C3T7d97dCVdVMnLXo
mnPSutL3VdSFjVuIV0gj9kDW5Rz2PV5sQEdJVu+r4fI5YHQIhNmlYelJ7o2zcLmM
9HX6DPe6Pn3ptIJ87xXb6aVtNxEoicNd3lnq6llzfNJNPpAcltT6hcS4t+2J3zFw
HzXSohz6Kh9pGrqSG1AULwhtJbQLfhZ+DtXEpLYlLGcbMte41NBvkjPjniMaML57
PuhaefbVkFJRl8NhZO7/Si0DGcHnuar6v//R/NwWek4Dpcf0W9ax8mF8/rmANgwo
2ERLRe8c2uGT1S4WluM+Dv+WcjQfrKomFBz1QwvdpvSrKJgPOmHCI74C+LEea34L
FPByQbhm+5brisAK9v5E3/wPxlhqE8iZYHExBksWlQXc6efACEZApiIk8Mccc+U8
6imAUK1len4i6GvpiIvStFpW2ZV17Vqhr3r1Q2c7/2eznbfrEtUyORMxtKJSf6KG
6Ey8kV1bMpyUPddXXWZYw6lc3XZYWgnCAduXmMy4yPYVqSWZYspIzC6ng77yipVG
UIrWuyHplomPTXi44m2TegNbd4HLr6VOIX2m7y1YPg1Q0ka94apks0I25PhCbc+H
6sSI/0qkeyRa3AarOqDonHwGezg7YWrv8915X3IL+in8nhon1LR74qVW6gj8kleE
EpRD3tBQOyulurGcdwf++5H7j8GhTCfx06Zjh0Hox40yeUpKpZHIjd56MOBjDfDR
MBdOV+abrlrdpcQB6OPZD5owTeQSVmeqDgL9iyGHgtnkNY9R3X8MBQ4Jpr6zFpD6
456/sd2aggI3OkoEbYYYsBKWTLtEE+d5uQ7bHu+gW8w0gK2t7Hy/TKiarpQc4raM
Plp9NZyQMLvkB9jEm6WZ9UQdZw000fCG8Ub8O7nOLiidVy7HjhrIf3+HsUNCiqnd
DqBd9hkGBVmlvDjxOKM/BjSG8AYHfzpjnV5uc1j/oX5MrnnG7UHYKvOAsJBku5Pg
8SR9uBpGvEVXYh64v5YGA5fBayrGGRavpWBV8JYOSe6G1A+mYkpN16hxRlpGTlSj
1iquPD/kOp+dJQnnuCgJrpPzZIT14qfJugjMxLs6DMMgI+GXy7Z7gy91whfUCF9v
QG7HSg7UfuKZXGmxZqfJs4bw2G6lQ5AnXJE4lnncIN8gpFkWyCL1nvxOZ2SzqezS
1WFUawEsTBC9TOFdXuEUybwoy45Eqcg4a2kZPfEybai/qf/zTkwRXWCSQ6XdeHLH
TO0so9wyig7C9WL4kJjMRmnJffkOIfw8LmGRLc0blaHYUtggq7l2FMH55R0cWKKN
Yw2jogDmCSNBQ4f9K4WDwkV0PCc9zJ0o79JfdKBkYmY9vQvBkybZ9j6CY/deUcWv
Ni8RT+OnB89k+lZggOkFR4YzRzwkF094qWsbwSgNfdYHx5X6frKD1iDeLys4ZUtj
T2uHV6/5QvRrHo21ISXIu2qG/ezAeRAQnD5V8IseB5JzQ0OZfZ2QEct2bETy49RW
0i9LvyZ1nmWCe7/61o+R//hG180sy9i9fv2mvp1bARGHQtAdg+5+yX03PTM7E/Oc
W/4XTvaVeXxzsEG//6VRIZiQ8v6vhonZvYlnzFfg7P7g4/byluFZbm12VRV4DBeG
w4MiXTfFIjQr1Hd59ArBKWSQie43R2i4nnxm9Q80Dpy3Ev/zjw/jpD0ZvfkKzhi8
2kZLninXEwSaNqUhzmTXs5ugC/ALWrky8/olpujKF9EkX17EppEx22EmaZ1PC1u2
mjN22aIUJOuE7sHxA5IpfOYa7LMM2Oy9w/UvHVy3EdOG3T+Vy2i5taN4sXyDasBI
2AJ7nZELjeX2B7Jj8mII80bpP2aT/lI1Aorv5TMSUQf8c1eTBylPOnAki4lTI9ij
VRK3ex7NzDfGI4/QPg/fOqxnk0aG6E0xx9UeyP6gkpgHtI3kXoxzKQ/d6vEmR38W
nQlROvgKlTBv9nVzqfFW0PBkBuGbp3+6Bo5dhNC9A7k=
`protect END_PROTECTED
