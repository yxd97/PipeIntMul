`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8nNhdLISz6JnLWXXWtVRg5jMjezQ4tgvxtG2o3wpDFxH3KY8U26XvdQGFUjY7RzD
jBGuX8Dm7l+mKCEcPMm6irGsJjIUN1I0//qt5G7oXQc6B5/ya7okAL8qQ18es+Rd
e4e1l6jx/MtDIqw8cvBBSTjOkoYftPp4Rd+WUw8E1KW5tMl7YHrvW6+0ssQjOF0z
3BTtwioyai0qhrAooCCZ+/phwgUmDJiL9EYVTwYTlwmuBNZzkjC4SIDEnGL0xt8O
1Pv3qEmxCgG8ivZSD/ZKaA/nT8oe4/OV2ClsjF1v8LII3X7jKyZoqRyZCF2SuCbk
CkRLYYBRvk3GzJx0eleEdBdqIwdbesh5qBWujlgUUdpMzkBcd9eqBogjT9QT/OfT
8hRrHD64UmBoqlYDFRs8SD6rLjd4yI84X3JyQc7Nw4ZF22ecZ4hmse4A6Leyyoa7
2N1Di8N2y9s6Gn+Bj9a9jQ==
`protect END_PROTECTED
