`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UyUCBAm6/HHfkde6mqcPbTllF8+w+gVSumNbZukkioPb2WY7I2K06t3I2jJtLqnn
sskEoCKIJg/Q6zFjxumAStjieG95GiPXHA/CF6CmAueYCcmTWZw68LRohSoInDwh
4cp0E3HChyy8/dJKr9ExqTlPczMDNB8yPNQXLBFbsV96b0G8RORIdB9NFRn5Omd5
F5MKNxn01ukx53Fg0UUO9giIuv/VcF4k56NwDzXjTJ5nJnFHBD3mUSNdrUJ5/V4p
yK4Bl3ZyJaIzW95NR8NjbsiQr0Fopzj6NznY9aNKEB7mwPmZS/ZxNlGU7MHGJTul
N/Ph34/R4NY8nadsF8ZTdwEwUHXcffvCvY6agc8OAqwoq6VPDWUmXoyrgAkLJmzj
p3bmptxbLbR4Z84Ca6yMLJXK6hfgBk1U849GO4GmyljHQ2bDvUaINizYbp36AqLD
+wnBWqKz/ewxFFSsaVVcR+4Q0dC57tbzYPDUZpoXkQNsYbM2EuNUHwVOdAJJSBnu
`protect END_PROTECTED
