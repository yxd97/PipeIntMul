`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xFbTAL5lQHxzeRxQMbMyq8VX0RN7qZkeSSGB5jmQ7aHpUEdUaEhSvlXVTJjCtJ+0
IrIe/7PCeTtgCMmRL4HcI0q5Q5TgNR/SAhuPVk41b8a1YR9EjO8H+VkyjGm87vbC
+DKgpoWWa/h7qTTb7Oqgc9cFb2BEdOgxq0g2uSCfc0YjUh1IISJXJBDbCHVMRqbo
A6owT231+0ZWXw3oaVefTpC/uo01n1aeUt0fWJ65z0gRYd/8aHbL9FoeYrduVpkn
NH5LpV3nRsoerx9vcaBRRzrFn3qrwucViKvs5ar2v9mCfW1cIPOea0+uAt/XDv/o
9kNa7wqeZ0sN0ZYBoF9T81mMKywohSliVD6mCEV70fEdsWXQtGc0C8WC850E69V5
qS1P/lIH4Ecy5MVGDPVrroW6p1kgGKvPGPcspTvAwVWP5td+HFT9KSj0/4DrZXqK
lljiAgTwghSFJNq/ALbPvAsLSaUp4463MwHg+MWW0L960cEcRuC5WVS+xorGQnLZ
oWj3ikOB0Xx7GIt5aeU/aW9KwAp6koZlUoT8ZSnQKTZFlkCdHXIi2fKiebT9wx/A
8QRc8R8E3XYliTfOLdF0aKAwSAiKgYkRFEWEpLTTyhvnhsbvcsiHkJ4kby7aQoVz
xRkn0LQ7f2DT7Vs5oSrZSqKciFydqhBxJLeJGZ27qx8fqQeNStY9Zk/8JLyoNkq5
zDgJ/Jq8Ko+3ZX1liz+4rjLIK8cgwqFK5qfoqNLmec8z7uNGuNYUCJE8QNvqLjze
z0YLNAm9f3wmOcI0xpG1VhOUqnyl9oJwJfGWMucUPfLEVGHTvggMnKc8Eg3z2fEp
26IfiFGZwnI0qDC9G/KqdthG8luoYXZ9B5Ft4jPSmwo9JiFdbPSPT4ASocH10ixL
9Gntw5Mn1CNNqJ7Z++BAiLa4lcDKrHuUfCLC14ui6yAXj1ckuhamRSh4hR86nC39
Rvt3Sp2zUzAdQKb5lugUZCFcFpA0dBFWgKgJ0Atay7s=
`protect END_PROTECTED
