`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bC/m9jFFGNC2XM4F3NK0aR/kG6/b51rTMgcxdzIO2u7NbXHEFN60JLADyshR89G/
tqPg62z1i2SAOUMyF8G9S3XsYdMmny2wjBH3HYoqthshpRXRpKJemofekvv1fb+6
FMKUa0g6Qk8fZ3MUhkMBxnqIpx1pRX4ZgaUZKQJtodOZjJV0725AWy3vsFoxTC/l
jRlLfOh3EwoefkT1tCJ3ivwtL0hoyLP7otZ1UMPPQ3v640GQe18HBMysQWkxMlYj
SXetaZ2/DeAYKqEGCyblcrr4MD3+N1opJYKmcRMzIBgqXU/hUMzjbyvma4luMIXV
YB2Vc5CUug+15ZQfR7lfhy/5KYyQBnUcp457NlGskvkV9A782TnoSNJaManx2NKB
i9J+QjQcbw7XZda1pl1r/2jNYhEV2pm7ZrN6y19lvxXyrz8HF+W846nwtdCOwDhw
4ljGCCiDk7gsF18Tn7YOhm0iMUQflwjevhGoAfh2Dif41hWIiCdSLqrKLzOhz6Fs
pQqVLiNnirxndwqQ4aZDuiVKSG9DZNaQCURNOpfqNw72tlNecwT6evkHZsqxv7RV
UjQC02AITX3SRttKfYoz9PQeo8Ow7xKkipRL+qL3CRTOLUmyO+fDoxQnetF1luAI
UoCb/weXEMBax3XYSiOZwrRDaE6hBQCkR6e8nW6ML+s2IbSxq3Wzh4iUeeQ3k3Nh
+RNFxfik9A0bOzvR09+G0+bZLnVreXkBLLt41j5sAdrVTxG9bAtfRe49CmDTTLp+
jBbMQ8SvE9yDNEtsIIqJ6nttP7E3PHJZotjqw9PxGUlzmVUq0A5oMBCH99xXCshL
y60CY1b/nfOVvBjsu9mwxagifqHVn1hbEvozlacSyQBYUE8ow8VBLhEUEVdmEeRZ
fFkZCQDTOP+Nxs9J1yewWggkr2Dgvv9UzyIOPTLYsUTSHgmcJwA9buONNoXK4lmM
cbVrib2hKKX2CHR2SoJI9z7wnalsGhkd6VoQdAxtvPIyh4Lfc1DjmfHVOefX8ASw
x/T6/ou1YJcyqU6BkX5r9RDeLYmK89iLjQKSdyiTCKbR1wc9yLchW3ybkyNMyETx
NoH0tuFZuiTMehoC6QbgonhpETfq5HIQzu6fpHaK8m3S7cEhJxNwgJE5eqani/Kt
wIA2jx9eco1CESX3NWbm2SaDZ7aNu1i8bIawSYoLXzxQZx9MNutjOINo/MFfVMeR
NaeHQOo6KjCvU49xLdC13OlXZ0d8tCSGvgZOlNqq71vM8Wy+GEU6eKLdEe+iEYSn
nqTX0iGwVZ9kj7FZcw0M6BtBlmIe/XjCgBxOTUCW8fH9EMA7A/42y2hhtI1vRFS6
nhaAc1c9Vi2fH9rTSHOnhmUqPhJrI6x1av5oGrOhiGSL4MKdoYgy9Aertlhvi+M6
Io9NYgdX5jcy3W0h/5A0losI0DwEFB3fsJK/OdY8zGOIaf8prKa1/z4eFwjKzp0y
oNuySZ46hq5Tg3FiHY0g5CJ8SRwANNGSZS/fkNp8Tn811kuGMmOCuJPIorBv+2j6
//4I5kpVe7Yc/mxKNQWe4xR20zkcfiqdnoHVs+60RRZ74K0nQO3SqZdGJ2jh17TO
`protect END_PROTECTED
