`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h3Zal1kXI/+iNXUtnSF4pOU3Zwo7C6+RVvBAouOvLoc8XxLSpUrgtSF4ojSLqi7D
xJW8/yVOyjjsQrxw3nyxbEHlQliNfuf1uCpRsxiJtqWThgxnwdfm5RjIERsNPYxW
7rJSRaVRjHvZkickaxrAbWEY9r+oO018DtshXkcrF7yHv6zB9uZSQJorHct/eZC/
UCqiJHQ47afl2RO34a+vnbf3NISlko7pvuO/ds+z18DXsehnXEz04aaR4pV1QNvl
DK5kwHSyP0uhQ9iZX+ciLAe9So1KDd8gFPS0/yEBTd9ccOiDaTDUrEsHZ4ZBXchm
TmWqO5zCWlwaYLMMdgM6pSM2vwbifYWEos1l5OvJzAJX7gbt5nxEC7onQ6OOB8qy
CrdeUKs1y/5dMJld4Pf2kyFySJnOI3P+p1AIFJHdJT/3dDyRGwxn3lvrq33wDyUv
lSBj36YQfIc4Ka9vFxLhA0nLml9zlOtkubrar7enpkgpQS3iXE34ifMXhGQzWoSJ
WY7WbabvhkY3Cy4sl4D9LTn95+YrxYTleYgi9mkU+bvDCZf+pEFeSXHBgshmQZB0
`protect END_PROTECTED
