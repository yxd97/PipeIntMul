`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IAs3jhDYyg5pL/VrkSdOAp4zPvZBluw6ScQIY38TGJYLzkU/7lk+QiYIFoR/i4Q3
05ODommMHDBI1I/IVpOsm0L9x6mzVxRjRsuK/bKjHtTKPcShFlazHQ/hL5xWeFok
Xv0+qSwgLxptu77Hqx4Xcttzj4b4V5seRBaeQKLhAec=
`protect END_PROTECTED
