`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lc0icbtFuVTn//a1g9NDXVKav1dxzcbmdRk34psm8O/Gl/od8x/AJgb//irWQMUz
lBYf0anWrMmE7Pj+C2+5uqdEzmXXV6dSoNhrs3gqWZ3PlDyls/lB7xXuiKSP/JqW
fcWp4fq/Yd3vTxncq4F3Ei9Fre+AeYJcRr2U6pUwksed7q8/OVga8h+Rp3PVeH0U
HVNOnvnHd/KjfO3hLBgmMyQhpbmkG8Qy+NupUeFTObAQUeZN326HI9lnJCj0QnK7
`protect END_PROTECTED
