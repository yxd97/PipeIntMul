`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GODwC3IeZcZGRvL8junC1coiFesXjEhMpw0Duh0lgFife39F65N9FOn8m6Cxn8rx
QdM5/CSo28GAH014iG/lfrLDzCm+gT14wvVLIO3e+P2KSWWmEOikCpnCFB0oEFYG
Qre3mUtu/rp/DiLqLcD2obYtypypOsEQFSQ6OaFTBWUgnnFGeZXwiET8LwmN/L2G
mF/cHsoWKlpxTm3mJfQRrwlJUC+0g3zarX5yWGcjw0T1jHN3SDuKJ8JEm5/dkJ/3
vY60I82Yl8Bd8sWbHspkW4FyTV9MBzzGyHGW2kfJIuB+nyU50LjzZuEadc42xrzM
dZ1TufSiKMb9KM1vjf5TCNwH9AoOx5OwM5kDcWByzadxtyfgVovQFF+ZMSrlQgzC
j/kWQvsqRnPznc67nj5yNvSjDdHcCnNtrywBIW//tw0QZI+LmqfdqFlSX6dXO9XJ
UZFidQQj4XPn1lplCi20wdI6IQLuPdSvs4q4lgahPCsCbF7RmBKcjs1r5DyTPqw5
48B7E9meisZmwnwTHJVJaUEp6x4PlrxAHJAH5E1L1wFY04l8ljnVn7FF1eseA5Yr
F2xDvRVkTz677qrMScTjZj7G7bzMnhkE02pLyN5UUgh/A9oJCS82XHLcMRVCz+a5
epxNuUqmvAdUDvxuphnQP3bli2I687gcoAlbvaIRIDiCux5Mbcc4kTpVHPWySZ83
68QM2hz2N+ynxmy8+Dmy5POr+wrcHaTYrHMrLuTyh1nZOAxXRfWiMQkLnX2iZ688
e7qvJglndeHEnGIkeoP90mbzz8j107Dogz13zWf0bLs1kxFDZR/uy6Nuj5ZxoAWl
mr2lb58mbfUdYqZaipICLX78TVBTq+ti0WKkU7ovB+YHkvEAcXTb9mGqoDwfC15M
OxxU68mtVreJGu2AwvVV0rKfBhxGAD0oSjzcempPI9xB7O6YxnoqxqrnZwAM3g4e
lVzAQgcCcdov7HaAzl1u5aMTBxPtiuYYXyhhESde1aSFD/3rq07u2rcR+XeL+KYU
mHqj0hl/bAkm5z/poZYvkdsDjb/Hv07DcJPcUU4ZMWYW8RVhplq3Et4OIEiTRwSG
PVUdpuNHpKikRDG64ooIbvhi+tquFHz2OUIU8pBFkJ/Pt05ygM47LMWyE1Xv5pPo
Gr7aUn358Vyepog2FXV+KtpjTjp2OFamsR26ckIsa52KZn3qn+cX+yD9hSQokZ+M
YQS15wz4d3yyt4R6S9YgdOg0aqkNFAEvxMQwmfj/H1AR3xaGt9cwIm0LDSjxiYnX
`protect END_PROTECTED
