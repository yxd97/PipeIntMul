`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Z9ymTysrsr0PCUeID09Cxhm4V12UKBzagF8S+WWZ6XCEA4lt0zD4dHBA4vL2J3R
TWrcpeZqRkg4LYXfBPwNFhVVe0skKS8HDFL1Mo2gnkLNiIF0QtYnWsAhOyHcZDpN
HPKDbkyX/mCNwEKtxYqVYCR0TuiLSlqP0fNgs9xl/CSVFltu9hA9rqeFGfyUvtJS
Yo4HZrWlbqXwvOExTyNZjSGLC7BsODiYtf60we3E0arEWbtdeGKhammn4iZCkW7R
0d2//mJWCWsq7slUJXqKC4wNON7nh3IVJDJDYQ/jO1GDKRHGALuTzfQkcZrVFavA
KDHGJwJptr2QmRoWmdVbWsWS2LpZqHoOvci7QWPxDLhzLTG47Iag1suJaqAnky8e
TA461L4SStC3BcipYpDAVnmitj4J3iwW5TsCDH6ssXv2fmIpr9P48xGblRrx3z37
`protect END_PROTECTED
