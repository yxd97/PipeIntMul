`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6GNLiuMFMUwAfTPUIPd46JhK6FzdypDVazMuEV2Lk9dHIcT3aVkHSXOKuvP7aNg
BSAtzcBe0dPs0+xVH3OzFog6ZJszLzUFekEebhTbkPXG6fT/uadXphRrM6aRQzsc
ZYPLe6giJLG3C1DeyyW5rx5yMEZm4Dwjm9Rs99W2+k/wUYOmgRk4KJOycIfMbGVp
DhMG0vyAYikSljEFGKRAdv/xa9hReDsSpW18veTHJlWm4bwytb7q2FZro5nNtG9j
0XXsITmLn4R17t0LSAPWUuaO2G3DTM0UnqpMD+T5wBeIMdbZ6nFalmO2uyMYCQ21
SHHu8AvvFEup6UfU4SywveUIkchATpSvg8kIYJJhwOqqfukMd339z5o1nT1ZT71O
vqF8FLuJTXnBjG00LJ6pj77EVtQ2rsxe19XhISctTkOiWJ5O2HS1E/dnTRHgSP0I
qTnUbtbj594O+UIOYZpE4Lzpi4dGV/+D43MnMGXwaEQ=
`protect END_PROTECTED
