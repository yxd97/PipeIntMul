`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4N3d2MJay4rI3J7vTzkNZ+7p0uxNw7dAF+z38t5BSv+9S8gB21BpjKXs8I/ocYBG
Bc0KLKshAlh5EK+MtYc9XbA1NDrtpypR/lSHjANtg3nbNU5Ry/MnxuGG0ESyt2TO
2z9puUnq9ZIvzLLGeI0V27uQmCbnC7zKD/7QO9LxwfRUlV8oqYDV30DlHOaQ8PQk
03OnX0Gm4HEB6ZaglRaOHxRG60GjoiCutn6hfZkJv2VvJcGjPdR5CN6fVUV7stxm
fL9F1j/1YmANDBzj4lxtXs+dqkINHfmSuR9Vo5a+41EHwr7t0CVoBhqAId2Q4QpT
GquQTpmNaz4dezgya56SWmxXrQK8Aj7fI+hkEgpsLLD8IAcNhTX71olt4NNtnyZ7
d10BsXLBEDM0dfAYYMOJW3piZ6UW+T0N5kcMZ/2LV4q9pXB8YysjJajna758xQ+J
yVkKaUPB0ogtoHHeVfsj/k3sD+ZjxESL2Y3nmi1iBavIoJGCCUe05hJBsxS6Y28A
irxMeauEqCz/49Kojbv5O/3X6rC/QIO9GrPA/ofhidVIQV0y8ixurpoAwZY36Wvi
9fpxdE5JzUsEtKEPJMGWdJoeA6ice22/JQlXwBmVApNahG6iNJK4W3weaT245pQ+
P02AUQ3iHiGqNO2KvTLYwQ==
`protect END_PROTECTED
