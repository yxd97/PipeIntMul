`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8K2YH+ENzb9O57DDjIBIxCJWFGu+KibPLQyQ1lRR0XSfJq1syEGeGgdzw7vePGu
73EqeSjYmK+BbvpNCMUM+y8raeo8N9Ji4ASit8cSXe77Hw2EUe5JG31Nv6OCJ2S2
NG6szWQfaRxn0YdArmqoap/idgjHxhcwZMQRXbYsDdkDMSXZ0BPIo86C18PL4I8/
iUCvK5BbunPxpJbOB4URp69Tr6e0bbVNIZVoCspBO9OxVtE92P4W6EWnbPO+Qt3R
2PJPoY+RJ/hNhlZOSkvycHB/x7iLrSYHELWCUXWhngw5z0hweiUcZXKSyEBns+V4
LtDEYMgAhCAG5XPuSjCidPvzI8PWSmxS9SUvUUKv0U5khr+IqALQbHf7wi92mA//
DQT/KzsVnBbc7eyFVrik3Q==
`protect END_PROTECTED
