`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pfSsuiTu8Ks1wvB2MIGr10fxvvCPzOlpIEBECRagPuvwhlSbHR2jXpTwC6eJHwR2
LaGcm1q0GSaiUU7WCCd92SZE/ojwRle+nI8rKI2p998o0twgS+cU2b3xLgiv+TmW
374Ajva7BO7czkMIsHMg3RZm3iecGn0ZfjkpTZKOVAhn24I0QhTD6utPbOILsBrp
JAakT0g2jLlY1xcUZBVv2H1t0hs6GiA3izuD/DsjaLUlTDR0I41kZ/5/Yv0B0JeZ
EfomzB14lwXYwfk0WXOj2oHcMNo4YhJPmUS8ShrdBev3ppkodwNg2NCRlLafrnha
K5MFzk1jWZ3jYzQE+mwIcVstas2mI8ShwtcHKdQf8Sg=
`protect END_PROTECTED
