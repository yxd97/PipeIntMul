`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2hRKGuxz0ce2RN5FPkJzLhiZ3ey1qWn8JHPK1CYhJmPWNaoSV4qKMrJBKfcaSHh
TBKuRy55tpqtUu3c/AMWf9Dijvvri61rJ/wM28nvDcU5yL4iVn8bbAq/nVydwooq
0TA+ZSKAwu8uyiWaD6efg1MwD3LGLOel0urWkWver3FblT1bahj3C8aXvoW+ZllL
2MKlXFo0sQzIbOK3mXiZ2/MUscoozGBm4LgAB32En1OCxCvzvxMiu3AMRZFFPGrp
1jib/7we7TQ/OZvvCdKixCXNAMz8f0PHqCx4ursLUrYMRMDFp/xJIMnk7+H7Avx5
aF7HYcDB0E2neJyBftTFFkwk5LKq/Pm00CO3aN3gKFmUq0OSIdCgVqsmAKy0rOPI
frIooVPuMbO9QMdzQBsYkoJajPCGHI+xvY/RbgWjqzScHoWL+AnQPLueL9VC5jkb
YJlz1F5gnRUFuWmQpPZxxNYdpA2NF/acf+GAyKVRHgqHXngQ7adBkCMZ84duqiFe
6GoWZKHJdkJG5rRzPYrRdhRmcRK+Aplojr5xQCSEgrdefMeS2bCMpK+hFUfjnBse
fPXecI7Xq2muDL69NdEgzd+HYQN4zESeIGQ6wXtY/AETmZML7S5WMYqXDjGMh7+1
0CEAxHKuDK/RgiRug3/HYZsM065PVrwvbNDgvHZFjdHtUHo+3RVgDX4X+ljINQvW
IFcwyPf2iV4Lvn5+0CgIqJ077lUlW47jLk3X7DTqwrmmHdbGZR/T9A4we3ZFZTd1
SKwEwE77aNag4VjaM9H0h0KeXsDwgqslNrT5elUhgfufZzzQAfxGFAPaC40ps8Na
qQEkvuT83kf8wz7/a3cLAc20t6yG/Ay3SlX0GjgNSuNdJVYEyHPjjrcjK6IsURB8
VUlvNKVBxs0y+nLJa1c626/t9QlKxXFzf1sgPKRbAB7JD6YMjgU2LhLi/B8o8gDR
wOEPlJvGFWelfmXyA2GEto+sEVBqudPQWnMo+WLUu3bKo72f1pbmCmgouEQF2saK
iabtPzUHkoIiYTiJlZqmxgmQKUnNs50oIu/2sW0TxtoOOWUITAaXy6Mq3ItFtww7
M9oi4pYq1ecfOJvNnIxsa+T02ZFvGAKObs4QgJ2D0zfx2CnCbj49gebFJs8LpUmz
qp27+TuGqEB+GFDr3Gdb5sLNe06JmxclP1qiIZXgF7Y7x8hIpBU1N7UCG9I85knJ
2Ahzgt5JUp2VOSBE+NBoJCFWFNgvOmsskJ00XBIcIrBf+xQOYqRWDbnfzfOo7VRF
ZVLmmxPSxb+U5OpgWDq6P8EVmIQnm/hlFOysW5N9o+p4BikgfkOw7voxSaVl4V6s
3NgWzJ37lum1TjBfIHC8UG71NnIz+jjABr/WPH4VIGIIa+DyrJH1XU+G7fHiqCB1
oLtGj2hLNvfaLUpUNsCrFWHw8sshJEGnkRUGi8mp9e7rM8+H9jYf1dMB0nUHedFS
+38RMBBNbVsD0l0up22l9BpNIR6wXU4Kn/iPa266Yn4csVhwts/S7nKT+/Zn3Y9k
qXQUOHV9L8Kq74sz3XWyZz80ulFionlY2v6h9oRm/BstamgIg++RVQ7RvS1OSS8P
5jIr8PQG1/oSLbIBPjORoPXDaz+0l4YE50WGxdaq6vjSWQpSN8kByS2tb7on8O+n
bouZeBQyb471EtJPQUF9Ng3i8A0Vr6hzroI/g7XQ+rVGvCM4cgRrDn0aS3YURMTp
/y9Un2tRWrmfrWXNkN0tx9QAvKbSMTMS+QuB5h1UbK15qnzHnswt6C8OuRssSPtC
Pd+v3J8khRKlc7EBQCMbW8Ma+DvNosrmbkRRnE3fYoWRULxb11NWdVJ7yV90ctmA
lW9JLX/rkMkKbJbRzPGYfc8Npu+i8AaiWfWM3VzSq19KH3oTrbIKQmCeVYloinjJ
g+k8rm+qhBHGHd1iPn31zpcz81cA0lyNgsMgH3F0oruUQVe3/QDnwe6R94+ScGQ7
ZwiZOiiglM+JCFNV5VQomwkKaHHQOi6wO+RdUYAsUE6vO2z7rfpBzWPLjKNq6atn
fDP7n2u9H2qwPgNjNLH79EyFTTmPlEpmkS9sN7aY8KBwCsxqCshOdLqX46qPA4G1
AhEwoa5Eq8EC44q34YHDbd2xH3N/dpUgAeLy/g21VBSVh9WOhXjfQVS2YHaxATKk
e36WfHYYRRJpFhGJcJnqEBYdM+KPa73yv1hncYjQ1GvoBg7fB/jrAj2vR5vlJUZM
MGvr4HXvfdj+y8QrD3mI7Hqu9SAqo11qaLrukFfYzrjWqqdkZFr+RQ9FufylmKYH
UPQRTOzA/mOS3Xoo7FgHtbr0Wo7nEkR6zqeluOblan2G/JIHLFtMxHHc4BGHqGLz
1zkOi8glqX18n0adLXR+HaYmmEg1gDWOTyOKt+nxcEJB9nb4iuTl2Qvtjz8u9VZ4
FUOrHhm1VJZKpZlASOPBF73ALWN1aAI88O19jlTiQKLQzgYLXiRRk5BZPJJStuP0
Oj02CLdx4/0cN7i2RLsKYbaeozP6JW+xgT6wwnpulS7NB+y+4UnwFgyfdpUy+ynd
ge7ufOrxlntk7c/h+EwHrtYkyL2FEjk2PG8Oy2NXBgwzbT3cwWlTObbZoQ4v/nXR
gjzBnJrOdCHgr/sJrlr1OMKzUoYuPqr+qm4Z4dzXNoKmdhGaSwjqYYG66sSAmw81
XOmKouWtblBw2eu27c2WVIs6cOvxojJLiGUlO8a2kF2fMIMxRae4lSTz1K7EbOKZ
8u3QOFFN1oy0UFos3lwfGH5cmVNXwbsWooGOhL9agKJIdVXtbCJ7cNuRZJcjLJtS
/aN/3fjZx5jVMyx0Gzeq8VZRIsNucC8GiPnizszaWa0ir00LbnIm4g2d4jo+tDWz
lvN8iD4i1huxp/E6qoRWKAyhFwbEYaohxVQAixJQwAtsPH29u1zRhhdYzD2KTo2v
/QL8BI/swxn0QhP29iH8hnQvyslu4O0jKYREgJgj/GtzWMlXJ1s3eNzZCIZcGhSK
9RF6dl02vvjQuiSeo3/rqjSNibBs4kDWVNt4DFEOqjnYS9kSoK1HLf3JwQTeAbl+
pXq05znYtrdN/F4D1PQPg7T8IFdLeNMB6CbfmexpQHPdKiDMeK+W/ValMZ+vFgxN
Ml7qb+OWMbgTq0KlpTzSI8HJuvGc77WAgw8Mq0+WJXys2/2Nj3F9cQqqzy6mvcxd
SYBKYMqaXw/0XwmCbDA/sVM6aE8+jmR75HtakEZkkSuQ4d5rJGr7AhzlWJ/xcK/F
z4+eSbDbLUZCWgAhvT7NbU8a6vRG4IozUTIAzvWWCZPeDn+nQu5Cg2ch5I/h1WHT
yoDE5dlxtd7/D6TwuxQgnmf4lZiYQoNmeKaYRfNow7uivQHI6FX8IE/YnfeD27Kw
P61N8RpWqefl/4sISxWKVS7wfOiEq0C1LCFXRzPIKi5hzs0t7xUpCGihKzg66oSd
Vkc+5DqBQsan4UqC3NkB0h8In1S/oJjsv4Fz8UNtD+N/06CAzeAIH/ldaQBwz9Gf
8Lz1o177BP0P0LghCQGkp9qz+sIepVZB3qkkhJ1Vy+gpRo4mQs++p0fIEmumzD6y
yy3aItelnUP3KIFnmDJidIq6vfp/Yw+iYP3z/qbSm202XRWLy9B+3bJONcUOXx0S
859EZjpXT7tfXgpJLRp53YxQQwzNOX0IitFgLUKF3PDEpk39FSyZDVWUqV2Z2Rc7
+Cx4JHETjxdQYh1A/mTOkTsANmTkroJhVRMaMjMiq+QDNUmU37Vwl27Pr+56wq6i
1v7NaYyv0KYwomoGQ028D9hZva1U3yLEpZVybcPUWlFFV7mPgzgMM2t6qDscmPrp
rUmkM/u/BIWHukBPUQNSeEXOS7LHNrOcYLzcZdf8W/nutQetVYv8Z6j82q0IOcol
EGvlrUL0WG/s85j+4AICqWB7Hc6A+G9ID56J1r+/8GDVIArV5EoHfG8nADtAqcP0
xsyOZ8IUCOF6iNNZN9QUIi8z+xOauvHR/24zl9rFcQmMIJykRvJLm+hcpobMtRcJ
lKdhsfT9A9kqKZWwSX16jBRNfh81gQVgMil40p0TkcTJExIeXj6eDhJEpE/tHY6q
+Z47ogxvBQhNZb99gQySciMOUfSsTXpgZcnckQmwefylcO6Ra5Jk6rz2MRoTjN+u
krrK9pChdrJJVF5xbVQmgmwMHR1KEnwT0DeceNvWzjXSIs9xybEVIdl78j4LrNPN
pn/SnnXgoaN3/y21kC08/mhkYy/dZUCPW+yWwWdZK/gUGJvJ6sTathS98LIxHfEL
XbDwElAkeAZ7QRcWaM/09byHa6f5hJWjr20yc7YW0NAFL8OmXZG7bppu0ca9xRof
XVw8fijbK9hcmlZd0HZthWHl6WWKv8yxeJMdngt8NeB++Bofn7Rw2m1vIuxGjwua
6uQXKYW90fGOI9AkmymMfFlW5qs6kiaYc7EyQ4d2lGpK5aDDNlmEiqBblvhDBfx8
Zx++fiLSnkgdqwuFXeJIKH4LJpcrzjG9CgvyWAvlWFF907jTx30efqgDrl52olMU
Z1kVK9Emnku2Kztm4pzmx1hL7rA9/o/uWKkBIL5gpNGdfqY0jzmMnxDsLTvwnuC2
Qbewxar8NiUR9YQq9+0RMdB84ElgcyexpJfvR7UgmNVqCB3xsMUPeD7bjZQyIzcI
2nudm7JHsAjyPVufQAKjguKv498xaOM3pC5RbLSPynae0Dpjoa2yo4lstFWoK3nM
tH7sCztRgPCFypGxmEDO0dpNexcMQJL5AvWl0nZfFKM5BuRH9H/CnFOaNcWRGz3g
ZMf17Js2EQmrpajBg6MWpsUnvn4qNoKenulk1kBQwXYIb2Onsm5zi7UHEbhJgG2D
SuooMyCRGQxC70WTKDJjIUTN/VFQZozxuiUx15LsbE681SXTZDHB2iDTC3igSsyG
PTrzTJYcOiq8iGA17eoBmcnG6z+g27G5juD+6XxWHCmGiLDSZUJKnyRppbJZrHGs
0/V9Ma7s/tfTK5R3bG1BXNn2U+yjpSgg7i8x40VN90TljI7TT5OQfnQTi1MwBkFn
YCOc88B8bPqKZo8g2lQYcd7CIy5dSYWTedMEG2aG8xQC5HKkcbNmv69hk1pkwQxo
CM0g/k2iCXF74l9XUOEW9p+yMxISKLWYX36eIX73+82CntTWQgIEZ6yaRW+N4ci3
i2YzD1gAiEABq/pCFvNYE31l7CzwGjvzQ/bIPuPgAkyN/P98GXGkoYsOO37v3QK8
DFrgUZlmhxs07KgKrfnw9F7URkiU0+L0tlpp3VqZh6brEewr4MdCrYe/UhdqQtsI
9gaA3VhyW2nDGOTD6TMzDPQ+vCGfFs+dScaq//aOhAMHBBBvXpxY9n+48VZpvxBW
uqUrLP5LRQojfhiBWO0apAIV3TlgrMeCa8HXl1a9g+4jKjtypcumVzI+IhATTdzR
gU7rNYCVXdNDhd0fM3yNzUwAppa3owbVF7hRsnp7rVeX7ocYnz2kRod55kuncdxj
GOMO477GZi/WKTYlkG8eW3ktxgpZH3RWjGyba8GyGwPcz9rcpTsoQ05m65kg9CUR
tIB9Aem7iwVDbt0qzdacayMppMzmCoTvZbSUPxx7O1Csv0xIUptExaY7WU3SlsJU
y1yWPAXQjoKQ3etm0s+LZTKdIoeGQQuFaOS6H9xdFInhVnkzpukSTN8/BXU+B6W5
7ySmeX3REjSlP7ubEOTFC3ZbIlSWatNGQno+oXAftbp6YIGETfQxpvpzDK0tyXZQ
siRumZcOm8zC+yAdnIL47C38pXiMj6kzII2URKZefHSUM6i3AVKLEPVervZ97ilV
gNMecOxdNbJKuV9kLqMvx67uXltIvc4YLaqvx4SMcdiqidZPmaAb0JRcUxcjYFhK
vJXa8TXQjlczS2C8mD/2jfVfl8TaE6KqJsxgn3hCGteImGrawmimxI92BHBNKuXH
UAb1DT7Jtkq7FvCOtPIrJDqTS9an2c71A6lU671+4nksBZzYBfDJoeOjbxoYBlub
x1ALB9EFxUqX5HSNc+4ESpojg8XwLqVxPqDSdpkCpuaqsa0VXcA3HlssbU85wm5J
D0UGThXnnQc/9w6w0g8pMtQq2U0/Ec1KwHQ088DXYNcKwJ5nhNgrHtJrmNYR+VpX
VADmgJ95zBGZuc3Z7gsCmRPvZwH7agf3Mg3A5zA0cFpBPagPzPdYuZAT/xtYcRII
KW6FRJwD5zaV7fQfeF8rChru7oXj/vWO/zs7XMjyh1UZC1aBlnVXXq6VRD28L1Bl
uEp9IbMpSB55csBuX4R43+Y2wxCDa9UXy6vlQPBee2p1fTKSClM0CSMbPqwQ/V5c
siXja7KQPD5AsDwpj40L2e99oFo1IZCGUqDA1GLpksGKo2q1h1xf60oIOI2E8kIp
uVSZV3Ho8HNxSJSrRHH7WgNUoIt4U2dWOhGk76F/FJtY0f8YEwZdiRrwMYVTwL/1
9JOmFPy/A8ihFbkx+819sOdsVoDFVhhuEiIAvI6Jr6vC0dwZO6hDi3ggCgZUoova
+Wm6B9B4AJCoskHY/gEZl6DDTOWTmVxUjYYx4I+P+WwBcYAQP5nAYhA65TIyMgD7
HKmzocN2c85CmlClUEWDLQmiTWAjFJdJNWhoPAdQ4pxLVKE8qiwYZXm4PfE2hlCi
zEKxvpJvHB6RXhn2GNEXLIm2tz91ocPL8Bp46xH+GGzKc/OtG7C78P6Havgd+s1H
mIzBlkgJjZ62ynO/izCQt8+/Nrzrw/2wWxwl3YbOUokk7tmDmv8tUAaV9zSnxUXt
ClM3PKuQUbQxbqbdaQwIh/f98FDPDQrQHh76S7SmUXZh2xQm6LmJXr9flV2e1lvs
1RKcvF9ISZmh+kaNSaCYzl+miqkGndmLKs8uB9jB1mXiDVXYvGdnnBW6/EuQ1BtP
wNLYJP4Hdga/IKbmGdTjYkAY4O2yRQf9B0DlpAAVxAdzXqCxM5dpdN5tytWA3EQo
nY/0mz2kRUzroLckRRIB9wCPNig0iocYgvhbBZaAolhGTmXF3QWZZZ6LbIv8FMKA
quAmkSq1Ij+uZv0rJrkJ+HLAdSUhLIQgGaToeZVPYy7zkQRYoWvYrW7t9rupg4ub
IvoX1pAu8i+LwsMJUAw8S9Vxud5PpBFlKie+L/d9eX/p2dLlGF6Tj7Ks7qpWgZdU
GJapfb9O6SP4MWlNnohwVfvhA/2m1JAGFn88Zm8wr8SX6y7UPJelv6yc96bJ+su9
9uA3qXgwYEaJtnWBOnJpUhqw3DXkXORX7TxyIbESw63paNRIROUstLumEXK+9P6u
FaEj0BwOmlnLoX/nIq2sxy/NnQGZYXKmGhQ8kMpMSDXgxtIgusWjR/wrbTyyUInl
1uKEXAc/PkdiYFzyNiAUFd/syUP70YEMqWfPRN0HZJeAGDqqF+VvBDxDH8D096E+
0oCvWzlwv0VPc1gMTc/eIxsiekCwlN664UbHDfkZccl53qyTvzO6jUPnMaCD4jBG
oUf+9KOOOz7csYEnaFQUskGu1k3xsesbrmFq+yPeZY03dpGU+wil2hfET5vf4Chv
dtGFs/uw3LHmTZCV8rD1IorbYEc+IjL1Ijm9vhtRii6k60K43LB1oXg3fwqi1Vbm
JM43cW0U3CVgB0FCFDFlb1l+jLT01pGnzY6XZay8Vy6Aec2NKeN0yz07sH6z3FAb
U0yE3wiBq3mwXVmTkuIbvFp/0zor6sxOWJpxPCNE5JrKRjcS2AO+gPzhET2glMjN
Qs7NqYKV25PlTWgVNnLZI9V+oWtgtxqaJLbgcaCksJhHELTySmfR4g5shBUVFGvQ
1Z+E2HL/KJIk8Bnj6t6TMIsSjisb7kfXbyLZNlnYKasaA18lu5OsZ5oBVlsuG07F
rAdVlLJ3mIsNJVrfEVQsNhSkbNkUouzNyIUqFoCxSLPU0qsoDx9YeMofQoU6+KG9
KrdvuVPrqobs54urJRs1AouwT7KEpB3YcqipAw9a8nkDJasL18mftdGH5KK1M7Oe
DNH1Wv8G60amjFb0c/tMKcGaL7a0oZ3teQf4d65582qgPvE4ylU10e1SRgOjuxva
64SoMHec2nnIDxABWYALlzsz+6UVoQs/uEnQjTX6tLlGOUjPb2ehjOTtNmVYr0al
ueSSwdh9D0QuS8FuQI1PX9jQcpLJ38YVSimaOIuCodfTg12nWUbUK1mif7Mq/l3C
6Lde+auHUjm/soULXLHimLNjePOOohbgs4X6reLKiZLATjriZFB6+DaSFMvl1468
wE9Oi71ErDYJUoW7Kn5FFDA9Lmvdh28EJmff5D1LxdgQmYkovX0KMw7sONu6zwE0
ifcvcQpDvgpRcA7IDWy14F+S21wqQI197iTGeG0yC/Km732BLpCrj+CB243JeOIu
5GuFYOOoAh7aWI8iIOnxS/RtT27OIUtpmmIHvEqIhuSlVQCUS6SRmJWgEzlReAQ+
hrdRwG2cmcQ84tKJlHnx7tb0fgb953twaw/AwaoedYlSlHlQl47s93iwjawSUM3o
1VrnmhA6tHTBBpiIPIcgzfXu2zxgXjs6apIfTr6RZaCgjdbekLnX1P0W3w6k1Qg8
MpDBaROF5gqhlvBvI9tnrk8E2TAW6l6Udznlvwlf4zXtf1iZpjy0HUfRCA/6yklp
T/sUmuUvENlQKoD3ZnhK4sM49awTsh9MfVxdvfq2PhuZfuDEOVL+eiNLklN4UKzV
Pe6AlfDFvkqE+VoS7QbjLKlBxsE1FX/xqmQaETC1lQChqLLiQkbXUu16cPKg2iQe
7yAeZC9IGRhWAwkuv+J6sgwFjoK2wI3EfkPbvj5hCsnW6tHTwPDMJaWRBmr93DpJ
AKFiQl3KklAESAXTR+aGmmJqSJbvEJiKo2pgGYGR5b6SOn0PnF+MaSQhS7F4Evqp
l1TQhPryTayE8OrfP6S2XGKDz4F5xDeJ4QnvnssjV5sT8XtYIPOKN20K4HCPMwLY
AyDhTXj01IkIi7nXurAaUlIF5seRkI0GTnVwL+P3Oz6V4Fly1DPok3b8QDMjfHfk
eugJ+x0E9xNCjwPe72SYZI5W9vYbPtJWTLcCcwXFGwo/BbuvAcNDlZ2uUpQ+58Ph
y1muE4yNS42AbZFbdYjVwrF+yKRFjaxRYNddFqDKqUvV+K5HL01B5ppwaw/7FOap
QQQfFkstdCIl5mzivOMZXigy9ToK1EPjP84e0CKIgnKVTKBUj2ncjNtYXFYqx0CX
ikkGLgh/j0Kwxqw8QUpGXgLk2nxj+DDcVej6ZIySrOlgWBaZKeXIbhQZ3lE1Zzv1
XBehHJiUd2KWNcbgpjfS9E6obqv3joEDgRQL146GDOUmmwJpsm7QBl6RKlkxVP6c
F/B7ecnNZ9o9X8A/980yrlP4CM9BxRSECjZCDhe8D6+DN3JIYRRDe4qZcDe6Yr9o
Gs60nQMPCrTqtLGVAOCl5d2pqx3Ujg3k2NBktBa1jdrTJW2N2owfSwDESKZxxeu7
9tT/4LjWNZPIf1LXIALftNSCnXo32YQHZ5JjR+fk6frepxtw58kNzUd+MPW+g6Kj
ZQcK+xmNDOkrFcBrsuw0ypgbyt+YoqOMjAVGrXejuEk=
`protect END_PROTECTED
