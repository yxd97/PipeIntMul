`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjoC9DBxAM1ZKSA4HXoVpTpyuoyOJrCbhvKONyisypPZU2eHby3ie1dGzF83SKy8
J5LrYIDbRTzYfaZEGV7ts3sII/UIIx8Rl/cMbpiGG1hABwY9/titb23ruk7j+K/5
EYtIIkK1IqkimmdyCwW+VZ/3a7vuKwZdFt7Km2InsnCGHPXvbZ0CjaeBAsVxTJIp
mXMAJitaYG9CXmOogaTBibRSjRRjljqtUIN/Nq+LVncupP18Ya5yzlxiNSRRHLND
hTuU1khORFE5Dc4pCDKYnEkIL4WsQzW/CIRm4YaAZ524Offm1B40U/kfF6hN5BNm
rz9KSy/9ES25CiCKrHMieShx0qRtxj3BNekFo9scK9FtlqNQSd1bpxnTyREgEjGR
kkHC2FOh5XG0asIjfx0LEAkUDZOM0QJV9e8qa2o2Dtw9D7CyCPITeKGcAg8ArxuJ
N8uD+5DZwLxwGWF0dV348ee7O9h5qeU/NIGs570/tIZV5CXI17xxbu2wnblHo/b8
q72DUhLDxVY1Nci+RS9+BtifF6cEfpzcmvTNcOaJtsrEJRedGw9RGDJFmXGPXwaj
9bLHnPjr42g3qZjhybHf2t4C603kU6HyJlxE6GO+jJyocMtiI5DTAqj+Ns0IzeAY
5ITDcq/kePpGx9ogzbI+7g==
`protect END_PROTECTED
