`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sKY/TG9Cg+HfVkg4VTlHhlF/jvlmMI49yQ6SfrXoUjiVD4/AUv3EwiSENBo+ELG5
SrNqKYzanoknR+hAECMwS5zixTB6e5fmu50Ca4C2Fn+y1so2NKcuj2VsEClRZeOX
zF2XUwRdQ4ixXcr8/ijDG0oypke9IlExWeOp2I/gU2rJCJqSTQ2zgO+LgLUIy11S
UzliJIbivsxJ6JGs4wBwHNWe6EwGMEs2XByQw5oV3LfLpvFLmI1AwfAOLMK5vmqf
5dKXTyjV9jqV47MteKWA6/ThLOAkUzh9WvBXjavrkHSv7sdvNyfrQIrseDqd+y+E
a4n3VlUcoInu/e73RZRwlUMp4h/m+GulywiVp6x3qkoIA6vei6OuXOl+PoHCUMQb
BPU7ic9JiqoYFtWbjiL69GW+0fntsuNGQIS5CAmoaLu/lI5mh2VbqlkAO9Eg2t6o
2csgwkAp+xm6E8OyL2pBh03sYJ5bED/yWGUK4WXLbX6L8reHikp+uSyZJoWryd1N
biP2heM4QWwmpOQdFK5wwKHdN68LX6YuXyqR5VN9e2FsGkSaPvmsaDajsgPtTnLF
WgP1HQgvfBGEVix1Pot8pG36lyfpa0yuwopKv015U87a8gwWixNKU7EDl0fBI7CC
ObLhHlsQeEyEmNe2BIOPBQ==
`protect END_PROTECTED
