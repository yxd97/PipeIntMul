`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Cu8gB7YrkgjYsBpQgIadXuSM2I+HnhRcdaFnqD6DZStytpmOJOmTAXs0vpjNOMO
6QMOUdWTTbv/XsKOKDLHnZyjByfnrye/zJww2LnAYXYNmjSW0Hid1c5kM6GX5+FW
r2NDc0rYLv8J6ty9q28oS22ptAguBuK1MSlkUrCRoYdLzl4W6zZwSLeQcTDIZ8cz
aTKf2OfXLcUj3J3Jm0Lp3sFmu2Axrq4ZAMLbMV0y1UH+dPXH9TNx/OQZRsSXWw1U
4EG6tiOVEbRiX4Yu5ajck0YG6w7Ksd2YTf7fycxxXmC2UqrViIo+rfVv+3NaV76r
YYcGH4H4T1hlT/rjXTCJUhxpoRts6SHtrtshKD0Sq4adq86+IuTkYcLWDItn44RI
EckYBl4oD6C9v3XvnJTVCz9iJwvn8cn9IGv3gYK9CTXuX7hWKRSAKmH7NhOvXECT
mUGy2+FGC+OaP6o3omtf6w12OzCvGHPKfcu19FOqjII=
`protect END_PROTECTED
