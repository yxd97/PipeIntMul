`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cta4smF/v6lEVMTKhlteqoc+ZcBRLzPB+aQozRk7UfiOaK1lvFvpIU1k3XJcVZ1U
nLb/adCBtmyoSyoheUnD+8yVdUWEHI3dAaCbsa5uWKoGO5tz+7Tu/PURg3XGW2hQ
6wbEi56J3ONdvv1PGb5KmS4SpHQV33AKtAqnyUXj56oZ3z6odby5g0XIcxCc2hqP
9mAv0ZUlv4HlZrcprBL69MktnsRCI9nT6BL+CZY1bNrjjRbHul7iQZznGsgJZFgA
zrTfpg0I3w+rU65Tv3WNZ8pVr0p8WZYZj+YIwPoHTqQrlSrGo13U+rKyLfaET4nd
`protect END_PROTECTED
