`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1kpDmEOg9Fy1ETk5seb0VKpIFSWFrqUvp2jrU7+nOB2oCADG16XWIMks51cAymo
9P6GIO0Ska2NUtVnxHBWntJI3KFBrv3E2720FSGsDkRm5GYfIn2EZaUIYwP/dKwy
EkOMESRKZnhEOux9JUmVwMqjYmVH7EwOFiIab3DRv7xQAC3n09U7wDRwrOWK4PkJ
kfceRgmwvZJC/fj/xyCdNA4Hj3TFhGwWvhgKbIUA9WROATgMP/t389u6Bvdkto6Z
aaAt3xgzswwE6XNQgUCz5w1Ly5QfG4EMgHeUikRgjUcrYXcHiFk3oX7n2hODvlzR
ad8PYpYeY/uo0LbtHgK3bj3zcT06R3zbTEQpg2agj9klK84RzckQa2+Q1fY6HI3E
xc7mH4DG+UdFV2sTkflnJuWSbxg5YyWIJygVkMaPJBYFCxfHzwLqFnz6ogJ+jsEr
T2BRhYbiKZ6CgE/lGXLFAnntAmIgLiP9I1i3a1gPRpU=
`protect END_PROTECTED
