`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pxlXEXAat0/4JY5KtSU7+6Jptc5xD35LkIZGw7PnyQXBzbnLWuMds/SPSCme95oW
OdkEo/V4CkP5H4YrQ2al4Lp/k7JMOrNn3hMycBaAXjDGG6xrfDC64D3OH0CMUlqN
t2sLBPgzX8l6fPngiDGa25lx5kgVHInFM34+HV7XdRvk2s+6SrzY0cKfal/bfBcu
f9Vs6wkUAHUBnrWkTQ5nVnM/YZbqW55TkehRW+hZN8S0APQVQexez+8pfs1d9l2B
TEpUY4a1l+mtczE6iNFlQvdxCVemC44O1KdWQvoWMDCTCP028vf2RfmYxwDQ/aJR
PHUfBIQOPu8dYq0pG3FObfb/ixC8Dp3VOzVSUgA1wZYalQns6gLFTLNJRVXWNCcq
70W7WEV0PHnLktvVn4h6L52FfcCgJDS7f91Nam88C4webue5jRmU9ayMeSV7qxr+
n3AHlHMbTRROt/RkxI/XUxY/u3lbblmGTjXQyeqTTaarpshSPhB3uE4Il2BCG/RC
njLp7wGpf9sov1SOElLepZmJp+hD//HggiKD/YCAvPsDbn9LRFLWWs+wm69jV3yZ
WDhqSqfcf60OhFTD4oxaX7i2bI1+f18knp8CNiXiwWfps+0NElChmHu1pXbVqi7i
BTYw0dFJDhRgFwafhhBFE1PNho8UjspkZ3SP1M47drlvU3Tr6LObGYpoRmWo8lGL
LICVYYme5JmhnVCg7m94Mv0XL2IJnCAuwc8eyfXBxOjwFH5SqFFpMAlY4j1fWrDT
YygyglSCecRAPM9KP7QnlvFPDAkRZxx3g/p0nOLc63QHgLrbrectS1sRY1IJdlYh
brkueQdgY4/OecajGI9p3Mt7+xQbTqpeN03DTw2pMYHsOHwCrAsNUyWQ0aoIQv/T
ntOKtUSkfvjBP6P/R4pzbbCBt5M0MGkoat8OmUwLAF9O6rywcCc0FEBYg243K5MD
ZUqc4/qkn7I0MeprAzdZ21w/Bc5Yg1lv8rd/CuGERibkjH9DQ1JKm4jbpMHp7gP/
i0NTNRCOCJ+XPDMyoOwsQSwCOfneK9aghkMdvKpEkvqaQPu7ILObNveodh6ZCHdt
zunvh25VqxMlE7fqK34qLXvPCxisojrQhDmrLorwXmUB7kfwxEV48MY11Huax6Lu
V/fWxVfCcF1v3Ty6Oi+PCAZs/UK9cbytmoiDf9LLjutDGgV2Y+UeZRu+3YvGTso/
1YhHTwpYsv5TiXI8RoMHuzMGLiZOb6R7oUjz0Bv9ATENb9/BEfOhoN1JhnPIgBev
9Aqy5pWCpoHqaUHtedPdBm33njD/MXx7kz0apf7gNk+Z0evza8plVfL+JB3uszet
wfS+JkluNmdeCjXbV3ZhNbPlnk8FENfICqQL/myCcwwmpYYukEjjUtVlchBu28kd
eXvpLjFPjwnCLYEQ70QYkNqpW/fKaRgpPBe6RxrYuGl9XX0++JMLQg+14a1th8x5
o/qdLMcJLrSOOXXnNd+MvW6QvzYxwByPSd/6KwnKmLQ9tiZZ9ED1EFPXQ/BqjjBB
ZEU8OAqsMSdQ83uzIU0FmWrVj3i19vvkVQqa0/48yeCynAhu20iCJK6qO3ROz/3e
87g01lOmv6G3brBo1fIQrfmnmiaHUP0vPZGwv0R42W7WgL5zH4994C4Jkmv1EqdD
pj98ow72aaz8uxzJxcrUB30ub47sCnY1zK0O4aNz3UyW0KDn5nm1Hz5oF/UYi70Z
t4b0/Ef26ClNQDTYN0OP+HDLM/GRcxoDM/iiaUgmVVXFfZ0SV1tRPd+btNlDZj1+
scWxxm00zmguycHOmX9+0VrcSCEA4J2BtR5KmCasJzly781sTAiB8MYnneBX4lKW
4bICdumbk9+FHcIvTQxEcbNPmJXOoaqeJsmeiWaTBpKq0bNtom2XRJuoeTONPXtr
h7fSuMevhif5BZE6GeEqqnK/wWKUVPsUO5tzbQkL1dEJTgb6SmSl2j2Q6zdOGUkU
kVCe8OfNyvHCZ7mDSsqJruSEwn1sBYSm+orOO7yiSCx4JtupKzPYCffpuMAIJan1
CeUTXTMEggBfiN5rnM+Rd1f7jApKhvBP0JZJJDSPBsW5rWQDAQrs6+Bdu16Z4+aA
HDbnBdbRu9Iyi+YqIHA9kVbC7sj7mvwB3l24IjTAhR9FfumTVfkqFhD59zIxudds
4uUB3oxTsVS4u7yp8PfiGNKqRHEPrCYgDfjAyJZTaLtH8H5mvYefh2WoyZRrYn1F
k48YUqOioZJIiFGN0CI7cmoz/BFVJpUn3EwVdjCUVc/rwQtQ6ABgt10trfCH1eEw
ha7W7iPjy/tdTgFHW/4Dsq0mYdiN9UPmjQWP4xQPhu/GgC6pXsiqfv4cZFUzPupB
omT2rouYofec51b+a/4oqmYJ0BE86OI/3dV0dUgrsWB1yRN7jA6DnsU1BKxGBQHS
lkf8D8kyGQMbZXmhHj5EU/g47RrnUK/WnvoMYDBLRYeGQY8GwF1VGBFaHEyfllKb
cZvkHBVwQxDqfS90Uqyj9+qT19+uJpEXXG+BAIlYVN1tT65XXKIjp5KVa9oXB76N
PsenR11p2v8RtspIO4SbYYeA4xBX8OHUrhqBktAwYw6w6gPT32OELDnzaiowfD2H
yOx4l1XI0yPfeomcqprAPUHJnFSq85hQ2PHqQBMM3g2VhoKWUS8zAUZCiQwOfUwb
amqz1jiLXx/nuB7P5yei7T93j+IvHv17YxiuqQICrZ/J6U+5SMXMctrvPdBg/LbO
sjOPiMJtA2VxO0rGVDgjaRueWeMGYoYe+rlRxb4cB97wKWw8Xb8E7gXdI1T8qOeC
PSXb02j1T8HnLnZwaZYcSgEpg2VHQCAFGpgJh7O8UAN3QWSg6wyXLwISFXWk2QGm
i9WV2dfXTozAwnjwHKAP4SBQ6vMwZGVsfK5zKeQ3bZlI4vn/NJpXwlRaAzvx5Ub4
asAw8DyQhbw7exzyJzoOiNTxVGf6HVUyaUNIlt2EfUJIJ+1gfZkE2QpxpKZGOcVq
Hbrb45WQMifihCtehiefep+ZbROGkqcR3Q4vrD8r9GfLjRYhvuSZhG0VTsnAUB/p
Gjk7qL8/89I/gErv18z6BCa1GKxPoofFhx+6rPeFRdPenlvJFoOp5E0NzIGs9qBM
OHgODHcYBFymuOTR0/KA8Dq5VgIveLZAtbt6oKfYCWkO9UmUXn/YsTLwwwWSgQ5W
RYGfryc8li83Oc4EzJTbTY9hKzCjAdq72gzZGLkCLEt+P1p7APFnuTIjntI8WYzM
kImIWYG5kKrzMZpLm2I9CjWsFMiCg3oZlj45vMi7hgXWANwxD94fACDphD7LpyUB
KW+Qssd5LKJwhnVd81XDDPLMtyjqTnNkF/WhGlM6/pQL8MpSAbFmZ/yHIxYZ8tqF
Dr0IiHSRp38Es6bO1Hp+JpcdUDV0HBD4j4EQ4k0owTFwLZDFsH2bC4thkMdIhmHC
LOb2hyyBa27eO9qKbT51Q/6iuCISAFJR5Xbz7ryF+MT9YkiQ48IVdOt/f4BWuthL
nPU1wseHTCdy06CHVaMaHJmhE6kZdYllkiQMTlrQXRucVE1gWSywOxUOQv9h73zR
CCOQvGMrEe+HQL1E7eE7zQ==
`protect END_PROTECTED
