`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/pt/1q0KLrz4strf+xtRUKVBQAZp5nfYHu/XP6E3qUCbcEzID11PzbMdGihVUiK0
NmC9H9qE/gGcnrvfhbFcvGx4qhA7CvbiTaUGopwiEYfebEmwcG/c7bWx/2yQoEl3
CukMXXe70497Froz27hTwXHzYyd/E3atUB4pEE9Pegv1qepJ2YXU2v//gHamjanP
HoMEXzXOgwSrMDp3qhkA6vivuTVEzJd+BgUYjtFuSCWIg5U9Wx/qt4MJryBzvH5K
kdYz+vmibogvsnEoc1mGHEhJ36S93vxYb8MayBdJ6ruBgACGUmBbWyjDv4jnrS/J
y/bblWWDw2dfF+kRLmh86cfNQa9NNq5aWf2xfBXzpG+BFu6mP9GzY7fhWvZQfUgO
Q9UZAmpXBBO7fl3PkVOcZCWTNEcy+Qi6FrV8pusA6jYKFnwPkXaXhpv7jx+62P31
7gmi1Wb+7nyUxY1dMxZ6OBozkhfme/obGKj9QXmMVEtXwKE/MYywZUpDTbaQRprc
`protect END_PROTECTED
