`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+2OKgU0kV5RIJ2fUb8iM9uv8N/k6TUq4Yc/g5qTAS1X3BUbfL1mgFX9h9+hU1n8
F/fYmEdoSSYPnXSOFC2oOxkicagbi+t6oVd20S9vrpJdikM6p8djuyroiS/ySJYp
U+h8YouHiHnB+nZGJdIhzsuTTdQZR1q8jh32eEbabOXawgHp+IxKMUyRulQnjdH1
HbnghwbwWU641t95yk2a44PWzQu9FTluMzmnG0jh5RDAyDfFywnechBEGvo9TUlX
WxeZCSMcnU72M8G4sdVrAwZ/WTO8M3Mm7v/7s+rHiJLNHXfXzw9FnGq/o+H3q2Dq
44j0tpxHsbDldAkKivNs2g==
`protect END_PROTECTED
