`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Ja85/EicQvG+jqha1xPCjV7jozNXe2tPjkKM8FJeTUA0BgBdi6V668dOJWN+gVj
wZBZEOHLb0/1NNWphjhuB7F/ewSq0tGNQ/ie0HnqFO3FeFYKeDpWKV3Iws8fYM1K
LNLbfXvesv8wxs/ZQ4CnRBgMsVWP7MFa/KEBUH5mfHYvCYUoMRyjpAhAUTUOWQOn
UhddF7KzrPp8ZE8OwArK6K+kQAnBVU21nrASo5v0ohQQGnikAeWFYi0mMTQRlMHi
ytT3Mg82KASgHE2HW/iM2hwHau02Mkp6YITJkYPB4rIWg26+87caDWVZ4qZfEJDc
3M5oItDTivQN/x3Pshjc0w==
`protect END_PROTECTED
