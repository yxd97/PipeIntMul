`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bevgJOuGPicSVAL6BIzkozkamg8oXRDMrT0Ao9oerxEJ+PqFa3jU/Cf2E0/9nrox
aMwI4GTPoBLQEfXwB25yM20ZTydF2LcKhdTUSiedebtrvAc+wesb5t9aVtwL7wD9
ovBMrMb4Vph2gjH3p04Cnvqa4JXa8utNKqkcta7R6peE6hY5rzipRX+fga9MtVDR
CLOp4cm+2H3GzTtyT/PPEOXsLtBke1uH82v8lpLjeZODvm9CV+gT8w5wyEmPXYhk
dBmWaQruywfR1lwQ3pWZWijaynuWlS2hc2lxdRyM+iv4fxxBL5SVz4hxPE56JW1n
1HOCqqcRloSujKCPBC4v14mdZF7EVKi1RvGAM5OeutwwDxMXMCs0W3w/nMwSJm4Z
CVOWWUoqymjIcnApUtWK86slQWChaOOr1UUOqgQJsjmIvJOFG1heKTkBSgMLic/Q
ZySBqlcu3/2yye9Zqv/JixckQogtgd/dfyo+bUII+DymLfm+oOoHgJ4H3ZOrv32W
WWmLWKbRbb8/a1OvrsftFOaSCXaZoJSzA0V7pQRhP6jRRNtL95m2ef26tbDFd3gG
NE4KTsG88d0lUaW3JaYyV/zqqBVWRQh5LpBOyqwUdop5IkQDJ+kF7MduDe2J0pFQ
NJ+9SqEdL+LBvZHwsaVzTGWyBs6vNmBpVZM/eRF18F8k3uF3Mnx9Ya2uLiIOd+4q
NOA3fK1pzythTCUYUQoxrkYbQCZVgmkiRYacHJl5jCz1wFll1oD/am3Y5vr6kHI7
hIR/O+26rz/cBQ4Bka/KD/ccAxfXwE2JH9ntz/yPd4toelbjiJyMrQH0zqs15P0g
45Pl/Y6JVYoeLKCDL0mQVKltM9oR8L8mB/qqQx0NO64xiUKEgVQ3VkLCpjDmc75h
UaQVwrwr1tz147dKq5MvicK4u3UU9CowxhwuLZLzjgFGNrYtpAjJ40hfCm7cZAut
`protect END_PROTECTED
