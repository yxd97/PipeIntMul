`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7L/dfUTQGku0p062vshLVPeQ5YUU6VjjwpulPP97YSCOtN4MIRc8JbS7q497eGsD
XzNnsDgDZiIF9CehlDbRoR57OxbXpKqS0iDTnjlHaykPorBL/GFpUhlnyF4a+cec
ypa/7wOgIzfRWXA7JZ8/K96zRo+3/ZLF6gwMk2DQoMU+cfsDT8sl7OySTQPd5d1x
7c3nbxoOPWYThradu9E3dJF1HWaaKEfrAgnMvcyptbX+jB8RQ8ZiU0ubEGTxY2ig
dAD4Oh8rbUbIrViqPU1lyX/77xxTCoMek4T2ceG8P7ZVR1qRMUrfUiVkmwILxuH9
Tm9Bvqr6GfUkh8UPKwPbPw==
`protect END_PROTECTED
