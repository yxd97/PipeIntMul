`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RO6JmWa+O2lDgHhSR0N7jBVcYEkDVMeMY3BfkxUGO3rT9bkw9K3ZZIpmw4xISO1A
wihZZg24h7USAn/OxRMvoY10W8vavjiJR6jBOXkK9NULYa7mQzp5guYmn2MTVTSJ
MvgM8yIMMMYPoLzXQhsVeY7YlqnoOnf38vWn6I+ef187kBMwVvrOAWzKeqlzDegC
kVdvYbGXxXXhs1UL0qsvXr3weD4gjwOjpF7M7/O2NXRjdWORionUsQ62burwOnkc
+pUvDeZej7lDK9/1qiytL22SOW+7kGX3+BPEEwaqzPqGTRUb1cUP7DZ43bNp2ZBB
H/Y/uLW4QKXTnhpSw5h5OWhkOF631pAJGi92tvuFIybxSPRRZLoBglS56tfCHFeR
C39g/1kNQ11tuKuCZth9JdDbrk6BEqeL4pFLdJVSpnXoRE+uVKlTk/JnJu+g71vq
C2OJFcHqnQ2RxsIBk3Oluu6ia0miRuh/myIkJ3rrXV2QR3oOv8tayawqJS/NCaWQ
`protect END_PROTECTED
