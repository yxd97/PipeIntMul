`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RtsZOeV+SL65ntEYOmth72hRs0tDyxXY1Rv9z9OAnq3ya3j61nhE3lGtK0kIZf84
m0mL0wDgpyuX/3YWIunMDGFJ8jlYo45vgMk/Glbq1OoUAMJ11fc8NemsQt7aTw20
PCnfZVJ2/cA2Dw8ACU7vSwa1f0zrIKQXH1Mh9VGYZs6pfYFqCEn/FW3DCoXaVnka
mIt+vySjoYJi4GZ2oQETWtrWupFgoLknl2H0oCd6gwv9OkbM1CuHqU9Pt105mnHH
71pGPo4zOMw2xtKSXO0VxwaPOgsaH2OZPBsb/BQbDeo0j29r/hEF3SDWAf0ZvZ4D
e7zzkCF1Blq0wH03Da6MJnVEzlMgyakZta0DRF9B4gAWZeGAOuWKoWOrfDFTWYmW
ecyOZUrMC+7HUxix/V0Qh6V3Hv6vDn9AC6i+5ioYbHojZs/ryj8sqXoNWp3RPS02
nLvxT+XhA0cVV1bw3lPy9mqWdUAWfvSBCawyXev6HhbGCVRHBWTp0ypLvJU4xPhl
Vn4c5mzPP0JgvzvHXnhtaYURC4t75LBGzljCQqiwX4E+d3iOvQzLaBw8NNraLdgK
BKwkX/cek0VSOZRT8xB9CX1szjRJQ/1wOOOYTx+Y9Zw//FVM4jxw51uZQWtVp9pA
cxbJTyZND5Ax5E1kabr2G3b3ksAscu5w9uTSHCFgg6i9qHKtHOLDFqOGgWrv/ua/
modyOX6VmLsIFSaomvUEid9q4+egs9uVy70QiTjzcqQH7KwYqY33I/JJMgNsy1Vb
Spf2teRg6JXkZof/GZ2fZdF1sThULzrg0S0KXhpVz7d+qSN9sGDJ5N4UPjLx4AaK
/p3KBj+416OD8gUkxQyB21Lj2EShkN4/zliM4m4cioHKTPZEF1OeNMMW+1UVei2l
w9t2vh695YK/O8YrNp6Qgydi2/1VfGYt8EtEXkpIRe6gs8GVjB1iF/lw2hapdvD8
7vTR8SHTIFIkCpcb0NUrEytU1rsZ1SroT96btwLWxjUjvc17Y8IUbqADUVbB0/Ys
jOmFqDcbgYvQ+I4dXkwpkkctUlFctfvIn5d0CJMyPUN7rsMfTNLLPYp5WrrC7rxp
ZYop+fpI/J391vsSRPWI98K/E9Z/s1quYsDTVEgSvJUpO6KhzB4BmNIH8B/a7phm
gQqsVSJYzHMt4R/Lpazp+imz+wc9/6sP+4ZIR0Llea2L3c0VtjpUZMc9NyWlq75n
751D/3kFd7oJB3uTfzqZF2KC2mBME/AwAvYi6LPxmI1oPWYNhjP1vFLlYx+iKTdg
MtzjgXnoyV/9cedh7rKJrkFXLauYz/8qzv/rbPNEb3bs99nYhWd0mhdgqrp830ZU
K4JvfIMuojPZnZM2wHE2Z8rjBEnNV84RPIzDwlN8Lq4bKr8Qyy7iiHp4f3uB4eah
86xGbexTrYNjwQnrfMuhqOm5wX2756CIMJeWdygKFWuA/HVnNe8xPGZtIMa4glfj
83o15ZIKrVYtwNCPxqiJuqdKvrm0Nh6sByBMIUczlmMIFeLSv3+/UyFeWllx/pct
iO2eMU/wXV1rhDJP9NpdlHZowHBzB5tPmSigl79rmzYL8vnP9O3v5c6nMlnF7jM4
R0/PBP8uAYH6ETGQPCOmt7ppsB6IOsMFG2z8KIyPMpHxzouOzmB31EvHfK9JBxs2
kBJvMgintBqeLHZW6EIYw1rFSQ4A28zyO6/d56p101ZS2V6OISHAv+9Dri6rzn6s
TOpfTh+JIl2n/YTSInVClWKB/5JinRopjePdMpVifQlnb0zJw1hYYdMdjJFd84XN
1WqJhAhxQjs2JZSDDQiK3s+JgMd+FK1m8lBMfxTRk8NBjBUnZGMlg8Ys4m9ySzAK
fbdqag0C8zgtFNJBUaGatqDfPK2BbC3KHxEpK4zO4sPRYsaT6/XqTbO/dTcr4C07
Uy3GKYctE/OhVUgPZ/mxd5uZ+lCF1tNM4rNt81s+6fDQ6LFSDCNMbTqcpnwTgpP9
pJQ8W+KQAiIyQhjO1kH20qEFuWBSwUNUUSJwDBn8XrcjaTCeZTW4XGyKp3hzwP5E
mW7+3zH536yDAHQoNJTuEQ==
`protect END_PROTECTED
