`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qpNZPV2tbXSjTwrGsJOpAtEs/4gfT+jrG+hb75655nrLHeewZhFZ/PsFToBQEXCE
OueHB8oCpPOYhpjprNwJE1fmwnoYg3UiZoEnqomhxSIkueJV4wBOZxYi8w4mMD52
fUo7C6f1VhKVn19yJ211sUiF5qbNf1qanrHCZ3l263jgwg4U3cZjaL/gvcTlS+rn
AxyXoXjmDmJHelcANMSkcuezbqhblLQPoV/z5z7Y8W4XVu/PQj5kvnbQLEaWQbJR
ikyHV5F3MtEGPfFs4XzZEkyLPJFkJgt5gTT9zlfIrLuEvsOj5JO6dBnCuSw9Y1LB
9A/9qTgydquBh2cqz3yoH1RYSWfi0ulOybYjccJzEXFy6kl0vB/MIW2/0IYhRA+5
cnw+huZ2kVEBsnh236+xM851PtmBi1MOPpDjz+VhSJKthw8BVKdWpBU/k5sb/kJT
aI/qtmpWLIyNdKxOyMLC7wD+KQKBJq6/qRvsJxY4W9xLHDa6VDbDaQHUdur1wRIR
`protect END_PROTECTED
