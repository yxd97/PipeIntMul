`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZXDDmCIWwgTYzA2A+BQiUqKy1E5Tio0XMg0iK/YC0/7mM6YijBZQslEUyLY/WN5
10mJgTaDyxhyLhpA/ZzqaN8yvwPaR+VXRuibInHFl2w5vewKwzo7VMScUjV3iqXa
mImFu9315PccnPGPkGgGYr4IMic0itp31tRVCyPUyFbD89hLvMrUbbqxsbKoU0B4
3YRBNHb3dQsciBt34MUUMge4Wf5vste/X0LtFrW/bs4K9Clr8q1nRy7h0bSQ2slo
RDaEPTKFK/gFV+JUfgGCwl87eRQ2vP2E5OdWr65OynT2oMz17mr58pTJ/rnRRSjG
r3bc0rXd3Z3PnKrJj44e8HU3ShWdIhmT+zG6R8kEB2qvh8ON+075y66w6DiV4FdG
p0edwpyDwZdgWNxheGyUNi7dyr5yZTbDPyVS8dxUoe1hycLIsR+2BlbGuYNCKxR7
1Pim62htZJk52mQy6hyga3W/5A57IiEk2pRfXkAHmVtLO/mrVjULivFleYSfdq6W
Dh3NpGRtYLnJmJ/rsiIi3bPaPdizCrEs9haypcaZH9/jaNeeSR41v7jBdjj45psO
KMPdSr+++fVj2rZ+KaJHnXWsD6SdLK7bVOPVu8Ee5bc3dMRkyA1qi/Y1i3uCIz/C
SffrvpT9xtSsseyBh4HnoFM/+jhRCbi9UNUXScXQkY0/CxPJzNhNjiRT9Qy+dNUO
WeZdyksPGYnoVb/CIOYna9170Cb89T/dbBwkxsa5Ns7n+3uHi7cG9FI8W4bJuW+/
w3EVyKSaDq7mAJGwrJadnXpjigFQFC9Bzaz5nt7cKBOc6HhEUMzAPy0EYJdkFEON
QgX9s/LZyfxCk5Ahp68N5ppO46NycVNzmLlh0I7skYculwisFHndS30+niqDnb9d
ek4Ds9kbhnRS8oeMZ9eSxw==
`protect END_PROTECTED
