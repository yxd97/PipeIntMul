`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhvfyoMTik4LXyTgBfhKqo9dUMeT9kDPYGsRm2Q00/Wd+iNyVlYROBgH+fjj0rSU
1hTqVgtZdgolQMGo6z6zw22q8HYlDkbl6lkV1S1+1dm3GuwoCDAjVbJaY+0HJu9t
PAdHU5L16/faLVS8anxTluH0UN43ZwEryavUqn5yTpesCDsX/mfG7xDNBmauKKTP
BSzd/h7q4MhUVaL47Tpl8jr4jQajyPG7es6cRqH1jGTst7zswy8XOXOIpEeKWHl7
TckMOcTTRgpI+a2wurBsK30oKSjEbdXkscWaRZyIWIJEwKMmVx7KzglqX0LtpadJ
F9WMctjc071IcOonxHb9AwdklEYsU71DcWbmnP6Ymq8eCdiauzGk9bzRJukD49gt
egKsfHbD9iY/yHXQbJCFCH46FyrS3o2WRo1NRHCKIFJvuCABRCtZZoVX9f1X0Mq/
7/PGlK6Ju7hzsQAjL5K69prNxwH7sl+QnZosrjreLf3R8ofAuVq9qlRInsy4FJSX
dTYxJ+92PaagyOb/9XXcP/PlN2PFATCTTES2zJIVfTYRmaZ2ZLAGx/E+aqWcNdsj
UPeQ1xCMVzIQHEEMOqmHkHSO5yH0A7La3h3tm476mFJpjOPQFNz9t0Ugl542IRlu
/IN//63egJ/fe6zODKmDxULLmF88o8Qj0rRy99nFKwkiWx6tbB+gV4ykN6qF99+X
tvo6BlUphybKxsU98Lx8CBFFQO/nMj+SncGhpoYDe/n2NieF7WW3SDpFONcd1SRP
5Mmxl2LQcPEWMmyWtSeBD2q072FgI6DY3hsAmFRS7KOZifGOQQB+7oLnYiYD+D9o
ZdqFgwVJC7mhkBQ178uyOW4J7QZ3RZGius+Vi/5niks=
`protect END_PROTECTED
