`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zYHA4ma+dSF+ekxXHkhllciYr8S0rQLgob1JGD0E/c4/lFz4p/P1o4UH4001dJ0r
MKiMrk2y/r+IYlJ/aPrJEeS6RVcqdfwB2T7Ucopme4t+H+Z4r21+uuss6f+rBUl+
LMDy2slcBNXfFjStoIySUBPux+r0gxXjzaANi9P1Q+Pc7HhSsqbAt2qITZ3mqlFT
8V/iX6gT6OFvCzNQPJhlcQESGZiqB4BxjCQh5ZlOwfJ/3SXWKRYnXwYdgZEwyPqx
K/02eWf1Kqxqnom/luTmRJ/6GuThv+aVlz0EBCdoWCkrnBvmNdc7omN7uKufAg6J
`protect END_PROTECTED
