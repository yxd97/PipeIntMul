`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MOm+RybUMOtM/okMHYaC4Xv7AfLlNX13y8IHUJDJeyYOa71C7JtZGKcxdZDGMcy6
DQJoJOiUuGtLmVknTQeY+K6c5NpMG19M907ERtKeMUgFcoYXX4yvpswT97YdGFFg
DDX/iOilj7KeRcaG3Y2rkNce8dRuEXTqTMhr1zwAfsoopz5pofCOdJNiVlFrXfRu
M1IknGx/LQ2zd+Wgx/tOVn8yXHZXRWDWKvEwfwq0uMBHXSR/GWtcOVdi7Rw2UH9l
/HWs46hvRuJVvb5et0HpK78ayJm8RK7Chp2drixNr5aultikwvYfy/PVi7NDloNi
itZQokoyHwm7tRNLGigep3PxZXEzvK6E/nBqUis57Tk=
`protect END_PROTECTED
