`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lNmDCnudm/I+R5K79AmD8wHfxVZnygCY88h+sPvTk4CKN1URJvfGKKtpYb/2ylW7
XzFqPQUJ5ORqApidT1dEsVY+yffqr42gS39OMczbnjkGSE4O98eubxrD2aBPWsKe
9gbAjv6DMHgJvgnhdVt+bgIKaq1dgNGCh5yIpiqW7fjxVsYEDx1yqy/FZ6a1aNIt
3m7gmT7sCdvI4GgcOsmVI4jY5PSa26YJdxdfukbzOQ3NGR0+vGOpin+mMl9W0yDE
D//01bj92/R64VhoKZJGc0xqTVlsywI2QRNHlR1agfolPGiOGdk6KR05XcPlQc+d
Y+ITy1dN9fK7k/vxImLdZSC7cxIXlZb/RpLImwmNRN77v3KjWxvsXLRpsXdGUU1x
2IzT4sO8ekDN2WbG/P+pJ3P+1cxevV16zaYp9oJJiMt77ud3QV2NmdU3Ne54lobu
N1/YmYmelKMMFbZYoXcj9nrYIvR+OJ3JTCjzuOh+1awHXQeo9iAbOT6cBDHh5nOo
T9NyIN9Cx+EHcLPNvj9OyCMBTdiG4VzXmUzfZ8df4hvw6f5cxj5cmWx8NYjweMSV
L8nbVaLEtJIsTZor/dXQtHwM7ebNMmOgObIf7v9yegSE2Mpxz+J7+O2ikopLCTBj
tGPcO74Stq/RBf4aBPP26A==
`protect END_PROTECTED
