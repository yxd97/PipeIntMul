`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e8PrOAcEiWEIIblkeuNHhdrAZKsbCdD0BctejCwK81BlVO3HmhebUzI0c2vTjkL7
fITFFsSXDCEDC5/rAKKudkOrO2UyF2u8anaQwmSneUlhyqpwMQlKfEZL2Iq+Rlha
BbzkNGLUXVyUr6rvyQYsP+to8KPy2LVvlKU6XT+JjJBhkBrJn5LDdpXdeKBBO98g
//BWhG6n/uAD5W0xeloUBDyPFHLOfwIs+3V1tYcrVbNUutaTkfU3dIZ5QbTD1DyE
zWHr0vgu10fDd4fhZ+dZoDvUmpnamBDrP101++GmkvFDluyITsjVLJekJpyJGQSW
EGw3sVP3ez8sc11BCDZkVUJvaeArEBxryG70Y4kSvvnj5dZd7WDO0fxgngmPlzC8
z9x/p/fMZfj16j5luaox8plJ9Eyr2Hp4Q5KjWgxJTB3S6VQmFhmlMKA73FxAih/P
LRAx+GZlJ7D34xVDh5kRu5Cnr9Lyk/MBp77rl/iEH7/ktqah9IjAeTRQX/73aeO/
nnOX8TJlBUwv2fwAbwTFydGqKoiKUmkqKg4pdDGuORuhIHQqcAkJQLeO2DdW/DQz
1l7cXWneovq6BeUy8usQSmlv850vcfcraWYHR1VxOCLgVRyj0JbDwbwAkaYKmgmt
PdfOl5nYANjPX9mbK2xvTyxB/PeHW/VZEKP1USXwQIZ1+mDZXER1sxRSebwcRFJ+
pz9yVg6Wk1ZZIu1WpV/9nKfZmf85lZTkqug0YI0ZRP7TEdGtsC2AJCfETk4IOhOu
mtVHFIxFzRBELhiJms8gonk7v6ZKAp0QMGFSa9JLSLt/kHwHrxJkjo2lU/27IhKB
gfs3pyBCaVcqKCXXZbcVTvsIzyi1fEDHVx4HjoNoiwRGuaLinoOc9tnYg0yPnq1v
mngdKdehwX/J9KWLYg4zWYMGCayxMD50D6V09I7L2wsNxPhQJ6k1x063BSnkxDEg
3Izft96saJHHwGrQUE+LwuoE4QiKQ6kuEZ/Fk8/N7air9vFUe4eg4vf1VwJw5KnD
SGHo8Icf23f9+0eOrF6P3fkJuDRWeY/VKaTzUioUsZa+7lrtZB1YlKT0MbLJC30e
`protect END_PROTECTED
