`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
va6rlZHK+jtS05mY+52XDAqEQaYTuNQIe8mQcs85XNJf4KmbieI7scjZME6xnLXn
fn0tdpu8HE0LHvDgBDs/ieLZOxV73dn2Mjb1kBZb+KV2PKJD+zfPrAPPEhNT4LE2
5gyDJvx2QIFiNWtDfAqHNhiQ3ClwbkWK2VpN3NTVCMtfRwFkVS7OP7bnGnNbq8gI
5PovFkw7d+OpJnqLFoTr/whpaVbobJ2tRnygvjQHom934ZybHkVBag4KGePh9yhO
ST3YSARsucjqxdubM2puEh/WO03oLvb7Zn6UJLO9wY73gy6MwccsKO/xQV8EKMVo
bmQc5PHqjpkqU6Y/FkczkNB929JTlK9OvfVwnTzzjfGG60SN0pXGU0WbDmPhY5r/
5bJfD95MY3OtoTy6FG+OoA/oZO/WRf9I04kI4kuNmX0/AiPiKsmkSySfns4w5Vua
+vcogv+mqBBjMoP8gM4O/mdzVgzfE3WTBEUhbT0md5UPfcUfwc9zV9ZoNJei0fVb
LvE0ztCvgh5Ej3iinNDZzn0R7MvKszJ3dDUZqaYMIyfa9UzW2bQXL2KHGyKRMtUt
puAatmAzpMgnj82bUwY8Vu0zyrntUkoLiJVoI1zrykAJj/bla23FfjoRSim+1Uew
xuqB4Vk3mjPjLgzsPqwWuaCbqNHhP+z2rrMRzZDjVkA2A1Kdnql6DKWXWPibRq13
zdtWfn0tWcNTLTzgD2yoTj8mGZo2RgFSJaUxaTp+HZCKe7DsLtUulMUICz0s9ioJ
12qWj7gcOiT7lXYplO8wBw==
`protect END_PROTECTED
