`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7nosTv1UkURckqlAS8cnYJ+gpKc87A+RIIehlxT5m9IfVjlGYWBnyy8qs6LVJtPA
Qi4SLDPy6+bEIc/7LD6v7kqHjp36ZriqlPDgDACsxHe7vkTPpbpazG4VqiynMEJb
LWX4gfU9gqLaNletRU3Dh2AbjaGAllQKdaYr47w6IVuVVLcKHLCBrgXgQEA0ijAk
Ei0OQ1jDewo5NAAdbCJrH+0/IdTDHOUDDbMSV5PDQsAsOG3Xd4Z1aiv4RnmIL47y
JeagrQjQ9CxbaFBNFPgPOace60Cv6oFZxQRScSv14YNUq4JSz4/R0n+5R1f09JQJ
`protect END_PROTECTED
