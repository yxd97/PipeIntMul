`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYU4MT2vYWOKXa/3aOucwmiQiQc34RC1iynkCX8202l+oH15VzMtEi571d9uDhrn
/PQ04k/Qazpd/DST3A3V50QTQ1ykQeUfrXZWf6H6asFzUNjFJU6X7nMCNgkc2o8X
95+e2OvKO0TehDMpT8x5tHzD763yBjadZkPdKGnWtd17Yx1/r2MMuqc0DDTDSldR
VoLgD/InNlSZcEWqPzCqgykblDCmL+jx136DUAZ80e+BHgMDtZ34op5WWIJlTDh/
PzRPGFQtMyJVhWScLF+8wXbTBeIeXth0ZpdddYsXt4CHz8gEqoVWh4EmOlCdG9ue
+6EXgF+fitt3MXHqoItaaJVp+XAp6ZDxO1ZgtLe1CVawu6MiLrSpemQ8UJm4wyDT
ZxgvdzsS8TDnXU0hveYsGZ6/6vTUH3tcvH3Gs+5CUAel0bJffpeLaa9KFjXjEsLy
A+cyuLVQL8lKEq9WB0zxuRkl2M8W2ohNW5Q2kxpvDhiC2cRBsIrkbmTH40l5aUTg
WRdjbPn195GcfvtCpbmY7AIMBY7BTVOI9jutVwA0+NuCuwAwvq1m89L7dg0Hm7Dg
0gNn2WXSP85XbTcAJ9OaO/+z97YSvnH+fuRBzh6CmgyzLnQazMC+ylXoejyi5IM0
MSC1W4onMwP6/3yEisPoHtNCT07ZjgNEiYt+G38g6E6TBkRdJ/kWi0kdzOAZQvke
snFXqvvGgjWpCjoCiBr4NuHOCDySwbKQNFaX2hTlro19li4JS9t0ZUhdX67/Sgyw
TBAq1D7qCYLpukVWM/d7Cye/7LRNVQBJOg0EnL1bQ1KdmIbezVYl04s7R/A4EzTx
+y1BYwRUtABuvYlR8o+/ggrPzU0sCLEEljZ4hcxz9gzqBFu6LFoMr1jWU1tkT1PW
1bu5Gcmo17I3RYLnMNtZr0kJWBNYHMZO3mbVkRQypMGlZjbXdA78Va297IKig5dB
Tj+xs2sHT/FitcczIpiyW+1uqN7UHH8ekhC8ee5CEkhQc2aU6rjXD2H606ym/vM5
ThOKXGpUocy2n4pGmV6NuJ2ae+1/VmRk1HgnrbjleaSZG4KGp3R0J9q74U81Ubqt
oQ1Yik0GT19P2oZfa/bjCQQQAz4ooVD8i8g8KGLYmM43l2/lDX4UZD6gtSXNsC2C
6QvLd+OubkshWvR7hzisaM673ZyfJR5TUPmxRTLdqtrUyvsLt6TbpbIT3gsY/eJw
eq0bpT4Zowm8E3WX6dD4eCcfnXnvrMNGDhC1JjAC33X3KSSBWn65H9jjbnN7tRDy
c0PuG2NjQ+jYkDQELBLlIJQf67vnFvyDsbSbLWMo3iYBdHVTF2hJIr6hSUO/bkpO
6N2s0xnwdAh9QLOLn/8vBLxx3nqxkFypD12W+WKO5d3UcyIx32yDR+hvJbemvXDr
Jm81tpFgqFfL5B7SXnL5J1ud5t9V6Y0KzPTJHkutzKM6gamlMTpsldzc6b0CMPm+
daeiUb1W/hugX8JPCzrNiYeN2bgwUvEHMCH6sGG/WkSQRmFkqdFp5q7EMnUPIj7r
yp8Nuit+HHI8nTyXZKykFGdiXBSiKzUpO/fcyxEkJ13kO2cJOnDqAvPgW0uWG0Ep
61+QgQLjsF0SWaOQrKMnsR7yaZF9cu/HHBOHtoLz1Ib92c6P4AmRBd6C+L8zexiq
sVE2PLIYzKd/5Gwa3VptgrHyUnMaCEu1YSeC4U62xPDFG5TN6w/zptDATxaEicUB
`protect END_PROTECTED
