`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vj1SP/Xd8KAYi/o0UlGW+HuB6cB6wjW2mSB0BskuR+MVbR2gxhPxFhq9JS7DOa6X
JoKEncn4rQtjIOFhq0VKTyMJgVBlYBrWvgJOlQtZiCIPbdjEET0IUeLerRwp0b9a
F6WtNnGLkDDMXw2eeBIS/WDXltub5F1N0U16kU7ZeWNc/Jbw+tA1RFH+gDsa8Q+R
DXXVb1pXoQ2egwR94FB89iaktNg+Rrn7LaZ3o1Ij9UmiVcpx/30blQ9PsePlq7v7
y1hNMpExnKphUduIIOlooByn3SRMzjsYJ1rKIgnpsYGupiM7bWUFTIdL1XURAIj3
w7NASBgdJfHUg++BPvztsVxbHFpvQO7f6JJPCcrdo/TlwY0dXsz1yNLmt/h+7CNQ
+pX+Xnd291pOh4a9ITyHV2G/qJKHi1mqwT3iHD3BbfRzmZY91Zj3vzivT0Ak/1kI
`protect END_PROTECTED
