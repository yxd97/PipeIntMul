`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84pjK2KSpgUYeqi675Ck2G1Kb9LRLOxyohaIBx6uWtq9KfkKXI9uqZNsE4YKlAiw
jbbcX6Lefr2xFmPrNH7+VNMoWBVSEV1xCf4tJrtwnDHwHZcRKzO+qKQHx1E4r5RB
YRTFZeziTA3U1xLTIVyNqoBbKo+O8ypqinWnZtSbsTDjyL7nJv7RKc+wRYJeZiR8
9wgZkRvZM1cFDV66NAFlOmVO6ffuYxTGJeBs1t3eFRhLaGmVv6yXTEMEOTyXu2Oe
ZHWkvVYRgIkHCJXL1UJFX2FDRvabKtq/XXManek3BJki4H8m8S7LIuGv6MHn+Vcw
BjAksLkrUTpTTPKeyEX8utW4NR0T3Ox7irnsIs5zUkgOMk0z+34dEmzv7sgCXvdY
/CendKcpEkGN3oJcaFLwfmWLAa+XKBh2gV7tFdgjbuSQ+6rQKBvWmVR4isrnO51U
e6am6XSjhEhRFbU58F0CZWmiD/5+s9NtBUpPUeSdPGDtAQ8yffJxYTMw6bPhEpc8
l+ewMhIit5S0T5iAdibEnN5lrqj2CtCaFn86Rns4fUjWz3qeOlKvHY/vqmylW8dT
JAdfoggnJDW+3EvBFIdtzbyy36/LGOPNDvi+UZ1bNKltha9CsdKUjqBFdYeEyBIB
yuRVUwWEI6cuewrRHzqTAg==
`protect END_PROTECTED
