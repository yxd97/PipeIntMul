`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rRbni+FZ5TLpvGyYpE/rLaNV2PhGndL46QQgL9VvScBEeuExU7EqhO2hiaSXC3US
ofB5p/vbbSu+ypWjvltj8AbL1eidaCdvzI6ILt2/FgR20gJyilYDOf4pFnzMeApA
Lpkw92bvPWyq9TcYDqD+g2sMZQSJPOQC2NoyuGvMfIVb0Ro0TcmtHxIg3ycUtIUb
QG1Nv0Y9BrGwKI9SycK21u/+FFRwVXCpYou8Ora63/FAr6Mq27e7sBr+JyKAlQYc
LDo2gq4QO3u626XfRQY9NrleXONAHwZcy1N6TbPEF9CcmcfGvpWoX+c72j7hqZd5
W07r3+5xDICEmu6RwxyAyrDEShA7aAztNZ9rXYkz+pQJI6arTi1d5+JuPvnXXErG
9TvtdW3+NVUiNWzxvusga95VCDO1mRJ0Izc4Kad51mgeeMRetK5bUxJw1uKUyQHo
xMEOcSM6FhL99IVLxry7F7fDeqm5+whvGDixpIHmQP1MjTUctwVmrsMgQNXBK+11
YuFkpaAQNBjjhYf8Kxe6nzTj4a1H35uI00MvJjx6j0Zk1vWwpyZNUR3bl/9mKKWb
PcMGa3/IxyNKMw60mOlwksdGKlK2y5chzN2vQLZhNrznzKozznkBAIabr3rjbhJS
6RbjJqeX9x+mPwakqS2bI2Lj8AIS7Qxi9JtuiwA790bbotfgaa6oAhTmiaXMVQHp
zwwQuwxxDc5fdn3nDUU6hzs9HtUuk9WRVu8Ebxk9PkTRi128R5gFElw2acy7ebIB
MCRF9mWscOSQnrfECDrHiUpu5t3W3B3U00BZefL2VnjL3PQiyxS9VIWu8jVe0sff
A4k7YYEBfl2p3OtGE2HvZU70jhj4PRf07HPUpomXwoA78/3n/cg/k9KJ6ej0YVjQ
6Ufdt6aIRkNs/SCq1wit8In+25hQ3OQ5lsZFH+JfEIFQsUFD31DF45cuKIqSLPUn
FIvj58Yo4srII3AyK+myVjTG6nsVKQcSsnddJrfLJfz6mh3kBODsrN1s0EXqLv5+
XERngSUaj/okixJ4sulQ+Kvd9UvFQTtDGpmi8PPIMWKagJgubCyzxHTCaHoq85Lh
G8fFMlfcDJeFVzmE0aG5V7cOumRGXT2uxEnQMNn7eSe/hU2XGcGf8g3t3PkEaN0v
UkTxMW28o6sZvoY6yjhTo98gXZ5cKlqQaixrhKjkRIUBJZW3nP2YfPtJWv+T2qrk
QexWhoYbIf6npwRqcNxkkS7F4KYUlC4Grdu7SqOfOh2dKPS5XliDIrAwbMQHMgr0
zPFyBwGu5K7J9wlO1eJLofFoL5JT2bwg4b8RVmN7FMP08X4h9Xg5oh2Vy7dUWbTM
9MK076JxCNKoqfpT77RLJO06jLVnj/qKusQgI4rFz3vjNd+GcB3Np+RBVnyIOhcW
Pc3F76jhyW7zs8BrvkGvA/jpEER8hEnWXlVwaXGlHODjtKa/tzeseimqJXbVK3Zd
n21Xumq3XXa7mbO2lvIow5QoejFpMGAqlQ4oOZatZarFJD8HY/7v+c1iTjIrx7JN
icwoy1D2z8wE3aiaZ75BYU40V0f+9y4KCAlPiL2mu/JQi67fCRWGBMDOqJ1po2DE
sSKt3mf2mvyFF0CKHx2w1WlV3vroucZkpLLGZrW0W7ZUD6SlvEFnI/z1i5f7vHv/
tQinaMNOUlPU6uVlH6bvMMAXE35uF3IwnL80JsqrUx2vkiULYlFLDApcNBHBKEiI
/vNh0YUtWamEqgP+vfUE+QC2M59hxq6/rMy0KeK2R8TvbLzSgrgPohFSSMm3lYQN
rK3NevX5o4UAQSJxXamiNdM6lA3PygVffBYG/b95TTs1bCmY962pmsQlef2VcmBf
xPKAxe0rYBKxNAwNRPudcSuCbK+wV63M2fbkhMU8JyHFCLZzOm3RLjhke1FJ1ZRU
3lVMVojDMrEZiISMhCcdFhfzU3nFK693MJyFhXxAoltPH/YXx0tMEyWTCjBurUm3
0fhEM+WtBENsvG6TqKmTR+KL3+xAxPiu+GdCd+EA8IGwewP7IAP2WJqlvawrroew
h6Ozb8m1yjrZJ6eLA5z0xqrPa1gQocLi7oekXg/juiS+rAZ4bpq6+M3jaa66ItEh
bfe6RkO/ugjas70GK+P4p4J3uP2d58E1BMHuX92CRQKHS+iFvYd+0n9lzVU3HFgn
XnTfUvllufR4OQvlW2OL/A==
`protect END_PROTECTED
