`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGhKB2AniVu1xLGCagAGCe9+AF/XNdlOrH1M2R6WUrhHXVq8fJx4s7orEH8wPUaC
F3RAWm59LnMkW+ZUGT5XmnObP5fdDgqz+TTnbvwq1wdmLyudqhXuNzzc2/HijrUJ
IUGeou904D4tKrdCF4ciUlO16R0xnq3TJTYs0go7Pfsl5dWXfz/HZr/AhZCJl3TD
Kpy6Cxn5zls9//hJOhqmsJfZBZNJh9TGaW+4FzjIBA4ja7ZxpWoM2GktUcDhPNCe
ef0u458Lr2OWh0mWqTI2E8KmVA8FG4HUq7B0vU+c6eFfc6y3Nt7eWnoRPTq9JeS5
Aycx4Lf1kDykvFQ2LcxXCNGxZhxuq8f3JJ0l+PVR3CLZswUOwS+Xj2f55QLR2KyP
FVOF4UgDrb6a9UFJei73298hb/xpPKKBHsJCr1NzNQbu3KCPURFZIyJWh9/DA2nM
cwEZofEgJklH3Eb4gYYYwtKTF5Xh3xjM2UvO/4y69WMq4V+Pu8UQWwgMWUk4E2cc
wFB8G326DDjSNVdsyNtHGZDUzsveHWvRNAAf1IMp5ETaT06g2RUUIcg8J6hR5/SH
XYQfSU7R3hmUnGf/XLQJ0c+jHtukImQzoZTC4gXoR3NAoDqOtCxu/dqjpUC9vRTL
VXwQ3AVgQlOh9C1bDJqwQQ==
`protect END_PROTECTED
