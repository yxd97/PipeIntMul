`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YJ/I4TZ7nlLbSchlndnyPW1T48rKJobqMnx/4LYB4q1qp8D96IUUnJb/X7LDveXL
5nd5SzqD2CGmbPf3wweZJRZRD2gZAuPaTzGuEHU7+zrN340coE8GgrP/J/aGXBod
pkZTLiN6daVS0ZbBBXuToujoRGOz4SgyMDozuanLwoQ0B1/ElkTTrRHq3MPqcVpU
pZGZpj1z0kGhfQWmW8WQOKAkxSqIfZp38yRm5kQXGjv9XTMEqvAnctnbR14JJ3mc
FlusaB5ipmI7SUBY8RM8KcYn5AZKKdPmE6mq8Fnednkk6/TLboWMMgGoA2ZIkq/T
u+UruEC8zTXxhVtRQePAl9LgBtruLeSV+1FM4gMR6RZcsoxpWr+7gsWy22fFaYtP
jEWWk61KLUBjgHgMe1QxW0Pu/m/xwJxvC8pC/DCrPmrhNT196jyqH5BkSrl4Q1K5
z3WPqq032XtkmqpDV50b+f06C5TnZFnPl4pgw2auWR4W0ekPu/dKVVKHefW3KR78
`protect END_PROTECTED
