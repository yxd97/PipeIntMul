`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8+57Xvph4PV67wrAjufBu+9Wj3Z4AYNrjHHrlf62G3PKsO9qqLYJNiFoxJEm9r3
KrvUUh7OcDerfJjoIPyBdtykX89LZ9hs/z1uvoyy4GoFC/nqmn8b+VHucEVZ6CoE
ldaZ8iYLEJE7ajXvZ+hXfISvTWsWXurrKlcLbpHUegI8qwC8zLKk9ci0ljAUSSyL
hnWzS2J82JQzj9s399l+id1aEzWTrYLDOLJwd/tkbPcL0Lz0cCp/sQ5hHIc5tpXe
jPpaaKr39e54kWxRCJZsAcrU+3Wk/L31MeuuVg9LH5zMEbzl/X61oIOuF4Z6F34S
IpzK049wh34mj5NzZsYXO6v70V4yJ1a0ZJtdkH8zwCwAQiHV5i3+CH6hNLIZ6nT3
ZprHImaIWcwGjmCm4CMU7IE8Tjkiv7cT6dQNx7epdcbW9Y+yv5eHEBcUzs+Zfmhr
qDnxO2ExcoOl8Ge2eN7pI/FoBpNvckpOm36pMnbj3qcf8997Kn8gyrRDLvTcKweg
hKeUcr0xpVHdSzWYvCmGGGE+oLiNls1v1czWWiRWIvQi9E9ek0646ZJXwCdF29Gr
EYO+D/WQt4HYfk1T73w7AuwCLT17U0Osa5wx1q5xmytSrPXiJOrqnwC4t/yC7Aia
YTDX2j+SAW/QPVLkm1TnR9sgNT0ZGDOw1H9CpucWfyzdIzvrWfR6Pnt3LKX/74UG
MiWmIbFTQmvQG0qiF1xPLvS9wAnox9bI5ibsskQuO/OArVtV8RpyUcaxRdppE5yH
K6vqIOz/K0muRarDxIDvmdi2eTF09nzFX8CoZ5InVqg6+q86JRpMMgGTnVC1LsIn
jeC4bnXvs8hiSlYQhqkgTwfQtWevRcLWMUSsam3oIplgaV2WKjBz4haLVKLel0DM
r6gn/jxHtf4+dCG43IkmFZWZy7qy7Bicl6sK+f//6yTrHaW2HVwMRA86Tc3ZqaaE
OwzRzBX9KEH+rqYMo5JtUrug+Ia3oVkTAmyAWJAHQIU=
`protect END_PROTECTED
