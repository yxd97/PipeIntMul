`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaMgjPgEck/+Uyk6DiT/VkB52VQhR5rS5EfK/uimPXvFcb2OxDGbD3NWRcf+iBG7
lX0FVIFlpQqfx/AL2RYXU85/oYNAAUjMM/F4/mN5+dBtLSNRDA/Yfuvjrb+XB4T9
zLTyQuWVQ2UU4JPW4jV1lhf04u39+g0KV1V3cEQvV4jV0vVKkdkpiW+GbVqtudUH
W7svUN3BnbJVcArJp3ACuvj7zvJ/KhglZQe65tkfzPtoyU1/4Y4ubuNwDh43ZPOI
gGLxtTT0qeIN+zbVWZJYtaiBYo0mVqcmqKLETsL2scRR3ckDeGxDlpYD5bGa65fH
In+ocyyccHbkxCDaPyMxlQ==
`protect END_PROTECTED
