`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzDKIETWQiCnkVa2L4EnDme6vZbK0JDxYo11fWN1iT5I9xEzCfJOIGVcQpUmUNiF
ICUCNkda1w6Z9mjbKvyfN3QxlePPitMdROwVZgoyR3me9nvB8NNvvMnpo8y7ztcR
D1zJKVb2nEPTdloB+JRtiWAL0GNpZN5bJDNgHwYsuuOw/dG3ubgi9bHNkBki3JXi
+sqYcwuGvt7Kj8fTgkJyza6PCWLGZ6Fct8W/ZInwiFQHtiSiupuBttVMBVwW8WYt
WssH3vHcWI7uxDS+nIIF44sWIiYXnTSn5U0KI+zfjsI/bsf3UZ84fMw06NjpXkBH
2mbYiqMeQwh0usY9dd6Fnw==
`protect END_PROTECTED
