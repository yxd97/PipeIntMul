`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zGXZ8QtSc4I4b9loW9fMJnXDPHk9tTT9q2Kchwv+vKtHsKzmIIh/GViK+nrqqvAo
uMm4zgJGrzw8EU73xvsm9Wg9vtLiGo0L42bsyyHA1A8GOme+1+h3Zd18vkvKO2Lw
9+4M1NlhIz91Y9p3hgB6aQv3oC4Y7vxNQ3i2nJAefYFS6Ow1zR2ddt5bbp7C6q72
Uxhc0LmFET4I7bv6cQ0Ir37o05QcumItf3FmQHwIc5hODIXjm+7sraW/imlHh/uh
l6SUOfYgupw+kQxOQqPfQ69is/zB/CKid+NLdG6BdYsZCB1YyzN2guzYuvu/1obK
pE5sTBcFBR0ho602rNt0KUN9msSJQnYYuAoy3sWbbGlLdibHMXN/xD5sqfclSfRP
liSnM0kXT5HZvbmCWX64vTd38WbrfGexc3x+gwf6dBwooIOELnqYg2fur0Dxqwk7
f0sJ75wJZknJSsQAkrenJd+8Z3a3FQRNCbXUgkHWUG3jjG+lhiMMxKi9uuovU6YZ
/JE4GBxJSnd9LD51hBUkO2KfLcBV077xRzNwk2evrP60VnRI5dY7eaFKCnw32jP7
or35VRGVOfrZe6SP9BOM6FY1QJdShRQILZgjjNO8RSo=
`protect END_PROTECTED
