`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qZcy5sjkHa3hlHlG/3E2AVRkDNiCra3CVHnJKuc7zCe82i70fAYf9pZN/SiQmn8C
9hg5+F13gybZu42fquMdNB9cPrgX4YZOqW1dX//i4eNJklfGOEWHHSn7x+7p7PCl
FbjxHeozPHPb1E+TUos56cewaDckB6EbP54MieOCiricwT9SiKupEiLQTqnFura4
eqqlI/cRut7Nceqvd2i5FRBWZ6JuEaVobp4sNZ7ATUHKHrwkhEaNOhaN5hnQaCwh
bMJxXH3G/8oJKoAbM2zg7ljsK3KBD+ztje/qsxO2/LaoYubv2Yj6XMqhjonFHNXn
mBN7Uk5E0MltiZa+xVNMgyGktbXeZ3sEOIKqn9AQZbL1yGu11L3+nHLVUdzxthO0
yRtTl6fhsvYXZnhn97qLGtHb/lfjPKT/PV020z0n7GJ4ZSLMc0ChC16EVFf/eGrM
4FRksQ1l+edzx2tRkNYFmzZUmQG3JJQi8WNV3I5VsWXLWEp0VZ0iJuTEp02HqgYX
Zzz+u3/hPRCg3Ez1QWTfgk8UCKkzM5YEHg6Et/XEBD4iVboIVzcGx7v+Ji1kJUlm
L9F6wrkqUHfZBN7Po3Js5r1yKlrK1P2WQAl67Wm17mh5+uLm1Fpr8MKZa8fiMU3+
EPm+UqLsvXMxfI66un9t9I1XV0E1HKxJk7LkKD027JowX/Y3OK55QWrccWQYoGC4
X4fTUVLT9xFEs7UzbZO2FS1PYs5p9dLakKeWDnR+JFK0OSwSOPvwxAdQFtCwKlre
TwsED57ek/px4225cRHIw4TcSAzFNJSAFDhVkD/dEO5Z4bpyGeRW8U7mh+e+fIE6
Aqfjl1ob8WpXIZSQVlRpx+TV03kaUo+jdSkAL1pM/YWQoZAADBsCB5CbDIZxAQ/o
sFxMgI1waemTHi11VjSiQS1qpJDjmfl/47fjxI18CThLIcfpFA8pR4hWDiLClcnt
SBWSHPf2OdXdV9BG7EZ8Y/JdfenZYDrSnZHGDbModXsct+J6V4/i8InygkQ9jNon
e2/rCdtCUTnuKqum9Ws+JuTDqrFCVGIacYWwxSNSqsV57NENqmt8I+6xvE/2uYob
b1C9LhX7tyFozaQKfzjjE42ggnNXOL9DRu+kaPkN2mvevM4r9DtWPwMY6dMqnF0T
kZ11bXcAVcUs+KUri5QbB4v9Je0vA4ITUrhat6egXURUY5BUonYDrgapU3WksY7K
pL134nzu7NDB4LbSgqRCm7u/DDLGJJw+bF8ShcTXPIRJBrQVpqCtVk8R6kfQvXzi
Qmu29vzLN7g7KNDpfAqd2oSKYfeWJ6gZVsCLMLG39jIasHMCvrQxVyU8VKuqxvif
88vbAM9cU6GA5iY8sCs37dux9a/E5tLWZVNZVNDFobr807PXxWIMcdyVKX99OFyj
6oZxMvR9Un6NUYQ6lhr2g8rwSXuoZA5XK/SCtytTDoj8VBPQSYuymebVi6IF8OAp
TSTRyN4HPrNwo1HJxQVLKa83gNXFUMwRQoR5nkbESFqtbfHtKiOXLGZ7OtQkno/K
df+tKqbib4cggoWx+g4JqLqkUGuahkW94u4KQr/Q9KGYq51G4e/m/3kTiatfu4R0
7HqS1U8hfb95na+Zo+cA1Jc0w0WMiGL3dlSkB7BC9Yxk5p4fiBk51YfchUnMCaBP
Sj3+FSUEWB4iHPPRBDr87M3N+2L9rRPvDBbjPSbMN31z70uaxP4CO7d1/Md+4HsM
Mn+ayUKWtIqVY3BtqT/6iPNerWBpO4vJlVvnwUohTsqRkwWaaFTcIiEMzizLAC/k
99pO9Zebz/jSiCVQTm4axw7z/bzzDC4fiODURhQ3Z6XzrOoU8E6VvPdSTgzNHmms
qb9CMVmgagjQu1382McmVNUC23xb2fBptUCZsYFRixbZ5LMn7Ge3f185p5LLkyPN
HAKG6k6J6NXJ2Vedlm/Oavq9su//kE7lGPvfWuHS/A+ZV6KoHN4/SLh9IKdmdgmb
zdoLTooIUYxqMYoteGMdmu7aqUHnuAq5Lx0zTJ001pZLmmhbC1pGVNcbSdzLFD2c
BbYSld/lCIz6NlHQ3e+CeA==
`protect END_PROTECTED
