`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AunbdN2cWj9IPLiccBVzISGSqA7UJx1uxjaciE8pxL6U6RgP2xJQDeHUbLupUjmH
Rz31kShPm9UsL1/q7t0mJYaQFeQJUAUoDrlFDSQqkB9kUNhTiApveNi5DY2CT+lf
3Yc6eSH6tBi2cTB5r3ldp6DvzYI4++YlplUxcSfBPL6kWgh2yviIZE9MCKO5gM+t
tlRKcJbqRyGGaZfQXW9LJNUgBFVANdQoIkwjoLi2B7b2vek7ZahVe8N7KftAZ2rI
vWyRmmBRulD/gtgrSmzg4nPskgkA08JQbKqVvLcU6Jk1ZQlyeAU25pbPA4vZxV1B
eduzuhTWsM0Zx0996/pxeZBypN9mNW5IhfJTtacWrBU8Cya+Rfg/+POP4ofXfoF6
TqVVD98wzIfxv/qfZYpqtuagaMsPkfcQyvCyl64drAuksb4uHdYGJTpt/mLvYYFn
AqBMQBR+r6cmRdKbctGyPMKnuwOfqZlgbLI9pt6C0rJUNRrTGMUGg5NQFV9yuVOl
BCJY6tc8MccV2IzT+FdRlYu8r7LoJT52Cb+8bUHlzRpa4zyC2I8kgCcbUPDDu8Fh
Gw3yFLWRcgwv0tgaK9kJKmqfDtMad5aXVMTx9RP0ymP58QWTHAqWyKVkMPyg0Rme
DfFNwAE2dQgxyb884Oq29QtjS+h+25O5GbHjVqnWmC9wSA8RSV3uxm4VlNHoJKX3
jOZ/LFZx57e5fMMiXYtwBcLZWTGOFTU/ktL7rC2TsuZRSK9lIo06934PYUuxCgJK
NqNjeS7QUUDVCUHhEGtMXoepYWFX+zdbb+iSIZaTfBQgQ0byJgH9CprmmajFKjC9
Kfca8QH3vUX7fjo0nlGcMeBYe7Yh9zjngfyXw64ZagL6JzzVEazM8384ZdbgO3Vs
cvS5IzV45ICVMH+/VX4v0nn870epGuIZpgCLKimXPeF1Ah4nY672SUC2MZcVAFXH
XTvM7n8YpRn99+P5hIFrnqkOJEthBYPCTqyfS0byCJ5HfvGyxEz81uBaZT1VG+8A
H0Mb/gq9CBq0aARiSPbt1pAYboe0RMTAv1TsBCcpwugtUTOXWt+nezYpNbTGkZ4i
WMeX6TfrVTDp6tdMk/bGTKF9SPJ4CWUBooHUkLUiU4WJ9JI5vJaKTByZqQCqRyOn
SHf8piSP29sHzSJx0l1NiWXDzqPyP37+cZmByzy9AkO2KUvgNK3emVNZHgUWfYKM
pxNXJ/eq8sAYqrxTYTv0M8FNnL+aL+JuQqSppH2z2gd8PzD1gTnoynCfcYE/Um85
T3/xvepLZtYJFjuH8pbowg+wFwIxcwgqByUqfQkYvvIMkj3NKpX04KG9mNKDoExA
MCq1nbO8DMw2Pt865MvIOyU+sUlosQx/gKaH53UI+9oC4SLyO7SfDOsXWC4A4xyE
HMxXpIJFfflCD9ChAnkApocTn2pqdv2l6jkQw6ovhhcb1r5COibyqSR5NKEpQBo9
YCawbzXyA06zm3PUG0k7EsH1X1/y65gjrREg5vzy4RwjnN4rHNErbDyF3R3KeTt1
eqhfc4mR2XZfVT1WCmkE9R7m+ZjSTPu2CpuiH10gQzXaoudXbfenHRPjOr5kyceG
VHZswHCoP+XbluOyfQcrPeC5cArn6M77nuFZfuXD4dbU9Idw5uSZYoyIrhE410eq
rp1bt5DedGRK3IiCdSmJC6poOVDwjLmTa5fiNqTMOPUftgm8WCdy/cc9R03NS3aZ
i8OuE6LZNlaqQAllfIhKsiQP6SN2lpdhC4Irj7fqmSUswzTSCo/PHg0zQNWkZcSp
WJ6Y+dAuIIMXLYferPcaovxdjZurbSOgqoGwvZrfYK32RDdH7tfbTXLwN2C55Y65
AVpTObMYFHQxqy4657JTRBmpyCzeSBhRWAd2Py3Q2AyIP6fbigM5uOziuz8Mk7am
fqah7NzCXZ+GGHeXOZAxPOWHDCdLQaB1xu8vwVOn2+wPqilzPZ/LQwtqBYSqQqKP
seacf7+fyGH2+It+dyR0kxZNPD/f+j4m9YvX0RTqEi8vfI3rWo7WJjSvv2YkJVbl
PDJHYyMBYUGhXBFyasJDlfYF8MBEFv3qnIzCJfCswDcQEnB5zcWRHKJQ1uu3RN3c
p+qXIM5dMVW4x0sMuHWvmUiRWvx02J5poaSyzqxsbmQApuvvuYnjMqXri2KGy/ob
dWauGlpqJq54Z5OHxLzDP5X2lPi2Iu4y8hz7iV2DRxbTsAyCCaSZtAnbtN4bMmBP
xwIT8JYikXBdO+XrXos8DW5qqCVJz05kURP9WynqCWqCjVlfu9tKRuqzmrxkaEOZ
w4oBg4fzG90+mK4imHaOqy2mqMMPzg2EAR0sBIq1q43lrHMlOLRI8rpoFw4lN88t
x2atHuK6aPWIzOIxIvAaIY+FiMrIE8ZuYNiL0ypNsiHoilvBBqyoCXWQ8dcuQnrz
kFI/QEpfcflo2YCANHy9s00oenRUzezhlvRjPbtyQ+8ESdr02IQjXQmFKItJ8fWg
4oNxGJ0HAA3+j63tPTVz9Le47+YSxKQ8IgJppQFI/oBBGswceBhUpsSkCsGOQUzY
Hz/JJl8zXZ910wWjOB9+26xIg4iBR4wa1HQWEsDRorWHR8b+ki8inK6Q8qDNG2g9
7kHnccF72mlQ7yUZsvfF8vL3Gya98G0Lqz2C9K4AusOlEoQ+DGIQsUP2dC0dLbLI
cQehOcn/KOBW/5i5gbcxLimcxOwJ7W5Bf1bGVNx73hSnQs3VFyrzbIZ1jwBwcr+Q
HbcAkcrbZNHgvs/3HbqBiDYNYngp8kFP4GB+k2UuUu6hxXIZRFNHfZy0zlK8wsXH
4wgm13mke5lLM7oNlMJM3ClcjIOLx6SlmdIKUTEFOzE=
`protect END_PROTECTED
