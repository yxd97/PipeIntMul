`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDN3i+Ka/qL/azuWZFhoRzMtC8WB43ZcQNTYI/nawu369RdVNtGTuc0QaPT+8To2
EWpM9fp9+Ed+oH9ngoWy2KHzidcimcZE/9VXIgohM2zVql2a7ep7HHxlDo+UvcKc
pqc37rLPhvsKUOU2lr3jWlpIToDcE0rOfsvOo/gmcIQZlB9cDFR4KurFbpLEuDFp
iFVW7uk3FjIXQNJUvGIQH++Me/Gbb/DITkxW1Jm9gPlElDpbwo+CNYDe9odIXGJN
mnq/deFQcCGLBKMT/7SA6f5y+TDNXLPM4QAagCtWcdVcTURXMIwn5GFF3jgNWb7L
a2QaTeWsiZc4tHbCb/Zw22fe8/4BRVAChZh9A/p19rgsG5AvUdRwrxbSnui751nZ
48ZTsEgQnz3dtd9ei92hc9ILhilpc9o0/bxWFwgLwuFDjwu8czQtG29T+yqor+th
BYc6dos5vQI5rtJHLcRisHHhW+ehNr6ksPk48bUJ/cuwJkSFcWoOrA3vMG22XUIa
L5/3B89GMQ/zGdMpnKBIe9LLPAQBqqn67UINQk0Y90vSqoP+btpMJIs0Ggf4oQho
KwIKBRLfTqmMOL/JG2NzyA==
`protect END_PROTECTED
