`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DsGkGQtA4xtPNN5kcEXdaphoHkQniuDkoP7Vzng9tGntsvNUjQRXJqqKQZiAn3a
FDIvZFV3O8PYsl/JAQ+l1AbyampFsqycJ5JUcD4t/HIjPxCH1HPZjAqBD8qwyj3y
2WXRTw3DHT9zg4ZgprxIOaO6NVo/wc+0Wls1TWa6cX2YrrnBtZxQIc5MiOXrVt0P
K/FMRauCqq4k+uiheB7DSQprxnMx6x/lHqkFmsfj6mI6Erwkn/qxruF4yepPRq9X
et22jv/7xiUKppn6dBioDc/k3D65kUdCpmOfKggKwrLFqUK+lZXXB4YU/yTeQfd7
ct5Usdp8yzAclIaPhqetNeFoQrVtsAx4LE33gjdNDrG8AYiSp3ORVEYTH9uckIPt
Zy0+9DsNu+TP/wVqF7BMPmCKxIyIwX+r4t9F02t3+43mfuCZWOoELlbxo6NKnGxh
`protect END_PROTECTED
