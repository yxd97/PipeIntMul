`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cegZiuAR/xTYe8ofwql+rUmBZ80bqzvIi7egfF52K0MmBfvTgdpTzxLl0YQiMsm5
l58O8ZGO5cLTPpRk9bdymlBPLXOvZGmg8ojJ5w2GX2Nb8sjrXOIrcGdDMAyT7/MQ
fCQox8MIIsQWzVpiiP0LKuL1vPY5SfUBLZXIeCfZYrPYmA1sgqPoRoJ9LE7EHSgz
NcBwNjQhCHOXDarU3A2kdPN1wxNsL9o4v8SUIUeMI7TN9VTi7DUyXpwKSWUlz9za
HA4lWtBvoxm9jxUHMCn2GbbY/ZcGbByyLfv+qG/MhpzDaVeoz/WDqp6bbBYtN0g6
YZDPHhFvHymCgvo21lpTrvgc1SeOi8hKYGjtxV85ZMgfTwUzQmKjZh3icYgMh7cc
qPHJxqfiw9j2kCOlAoGn2QKvERRoiMmLa4OVChyaqxANGMUASJYkhlywezuLNuML
41zK7DNQSVmH68G0jwwKwD4NX8IacrZIKBdLtQmsTa3YvcdbHrOKXNopap63EVs2
seuD69+ecUG8SBVY/ecqyWp+kcg1l/sQYHO2e7vnf5RmSJrlpU4IdBl5kJ0dz/9i
QZl21p34FzOuikKhtYjXNkl5dNqV6Z71HE6djU1dGtLUji+HLFYw6V9ScQyDwQfM
FvWqKmmCq1qRhOJaCjX0WnTS/UeOWASkAylEa6rzF/nxxa1/Hn+LsaL8uFcu08Sz
mMt2NbH1fFyPRAOBha3UEbbP2RdHbGeaxrvbw008q4I=
`protect END_PROTECTED
