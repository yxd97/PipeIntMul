`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mf74LuY6+l1m6csLSSslgK28XC9U9DRjmqTw5dVgciMrDTNAvkdtNRP8UGcpDOnE
hYN16/ecZ+1nysx+FxnqKjNCKIzykABjcriPLqHZA5edJ+5sEBmRGsXECgARt1EF
YnC8Qo61k/RA0xThkt2lG5QmKO9FoqT4rxMU9qILWhW0/QtK0kQNY4PabjK2Upf/
H4SSfGXtO8ZL1rMx2bTj8cvplGL8h/sbEd88YeLW5MtuXatLWuIK38fpwnWNmOkV
nhGFeJyhEoqmVyvRAr3eFKcqxjL6Q9WmQdpwvTUlYhflx6s18ek8JfL52uh7Aqh+
XnQDpRlvuHg6Ac0rHEuY3oTELGBEYOLGJHIKSW3yUJX7KR5xJh/HAhvDop6cXvH5
UMvqK0mYSBm081t3evtyH0kfj1/98nbLLFeBlbSyHY9XFi7S6bKoaUOySpexN/Ec
YGyWjLdz5u+0LqjSQZDBYE+sExhYAXTzA02nLPSuckkY3TcWXTG9yq+wdpGI5zDN
`protect END_PROTECTED
