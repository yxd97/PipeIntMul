`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GzWKv5xgXcRT+6HutrP2l4+3AKIUt2ucQSmp13S6c9cScmyCyIBmn1Mmna/BXUS5
eVR9jhFtTWlMkDgm5GHlzR1v2bR9nltcCW3mqOUE8MbLxa9bY/S2rr9ikyxPTa0m
y1yGZZN7bOn1+tMXhmhHNHQTlOm61+KUG2MFXr4BsefBN+XQHvI3pgr2jWZI+Sx4
hbKcV10KFeWxIGmYnmDM3QVaclt7OkJuEb5Pna7V4IP/rvWtWKCKzC7/osarT1zk
DDPKJQOkqxoFWORsBZZJGOOj634uONYhebsHv7LoHlEuOxMLxIQDNR/KL/13Ue2l
GyB7fz8PPrBOncVREoxyhmj+FH4vvB2tQk4Jfb9pfWABPp2lDwWLWjwU4eQaP7I6
STvY7pFsc9LMXmkspJ+QXaID0+aa1W+Wd/6t2CMc3sJkL3R0JypGNL1gK0uMsY/Q
uZsWdbtubIvxfMMgKeD9IpHVXSw+CXiM9PQzvBoLlVT8NMceOqbnNhCxTYM3o7BE
6IZ4lnq7GIRBLG2ltac7J6JDju2V5TjZjp9YTK0XpFENLzLpXYy/qD16us00orqD
0PDb0bGB8jE0Ddq5LIxRZOEa5v5T5J5CR7CC8UWnBQzqcj6Nd6H3P85DP/Pfqpkg
+rACirEDtww0lSW3KR3wFI6Q85GbA8YFFyFl0qPZG8Q8b6LEZc+fKG1zTVYbi0qs
rlrHsGdJd3/Ct/t6z3gb8WZ4v3LPTykoKrgSLVjFiT92QKFGyiw5b2+lWx8jOYm7
+ZP8jIi5W1sQz22rtkopQA==
`protect END_PROTECTED
