`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QpqR9V6h8WkNMLAd7hLR5oDrnRG6FFMVaRwQaa82VB4QtY5FhzJjtYxmgeffk6ZO
22CIZY+n+mGdoN580XYG9VmQvpWBrNtZ7DqMVlOWro8eOrSg8kTtsvOLesQdTtCg
H55mg5EmvRsOQZ2TeI2fDl4qFfIoN1cLb7ANn3yCmGgFPhuAStHAusfje+1U0Jze
ZVSunqYIUcFP2QyCG+6fFQgWkI5/7fGP6Nnd6akXOSMcHEQKH94LdbEbg6n1NEOQ
FTj/+BMStHpLBAGCkFtdf5/CP/frj2SfkZ/xaTcecnJ8QYqp6U2N/QvNW0EpFYpZ
oreFeB4H/8TBOqYCtROhzgx5dIWx4lNll1Fm5LNdzXmBsaYFFCRIJ1TWcn8BNCEy
kCzEWyFYNRId2LRpLF3MJiiQmw53wsWlaCq3DwKknkVj5LKrq9gI7ZoGnXWP5t5W
091re/Qpjp/fHQ0AIfjw5L9PA3czZyki+iY83MYTTIP4hBStVh81HXwXulw9zTzP
nAbeNqe0d2OQ2I1pUc56MGGUz1z2RTr35UsP2skLkUbiEbLuvKFsiyV2DO93/9J3
QzJTGr7bckjRn3QtyGKLYMwPyJltTYzTnxPhr6FoqldGciciBQELef3WhEXmp0He
7VDF00BIjZXaxkzHw8DZXDOT70VREu8u4G5h/q2/oCDyYTdxGmnToKGl+LmO64ly
+2PR8Tg0RrdKZGluiWytKfdAtJsP1rilhPAqMweFJTep5ClcJ3jLGPTDKAWWV70G
orOuuf3CgCQMvUyt53mB1xpZQnbYWQkp01U4GO0GYmITux7Mlwp/GGrr6KZOtJiP
CpAIzlnF+DxUf6ETI6OMyyGRaczOxK3nRnIlhBRlyUncezFu8wB8ZCsvXyKTEDVE
xXqZWS9ooalGLA9QINyYVU6DRg9FfYstN3RdXiDNXoISEWyhH/4+rv5UNRv6UCGt
BKndcg7AQ53xDg5WqScNSwW5uYey25/ryg09MW8LuTWiDQsIUpkPMmf6V2u+3dj7
0//BJIXvxVildjPYPZggPU1kT40Y89WMpx7zMrlw3onP6f+hcsuphliR86+LwFrB
X2MqfjNMM6BXlFM9316YouA40+cEjPhBxRw6BO8SQSqGptH4eDtJki4khRkTdNwu
72aPYShZWu+Wkssuy0gMSxMQPtI97XbrUfo0hcO4TeaR6r9fFz7EmFyqHSQ+Kp8n
0QWfh4hYyFlghBH4n1JXL5lT2VqceSaWZaADNmPZLIDn8KVjvDu5w3JHLHT41IHt
3UQcN7gvKpbp9t5k/dS2dhYjrEwyHIeDyJN3VSI8V2gy/FoauxGV9E06oxNT/Vmt
GEPC7YtNsqqypUbVOm6nbA7igCby6lcno/d0EW8p4QNFKXeLEkr5FqkSrlZuJdn3
`protect END_PROTECTED
