`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xH7UzVIjsvGJ2AtB7u/wDs84b3ISZ3wGYoyN0z6PdshZ4JiOuQPGmVFdbUy3cIBw
GAYqNetz31b/ylawEef0T/JbNSUkQR4q3JZmkwISAFjxIRvxVpxHa936n6QWGggi
Tk5jEgaemmUStwlxCfbjOFxEPO8/dyTawnsmCp52AF24UYEKZdncWJgFEt7Thq9S
jGSWzgsTQKkW4Vt8Dki6tuXD8Qgp1OPsbOr5pQuwWZ0Nj40nfKrpM18JsCYGzJ6G
vhIZ6nL3ennD3rzbHCjUp4v2vQD5QpRw/EquOdaKsfbgMtJZL1BbMOlitM9ZpGo0
c38AeJku0miydv4KBghF7Z8d+d5rHXkx5xiEEmfwOcwlWemE5A01VjDBZ6VLE0+H
ywBvTX023rOAS3IeVJ6FXw==
`protect END_PROTECTED
