`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Tu9tav2hjE+rR7DBQ6xuv0CSbxwo2OBGu+L8BQLb6dV4/nDVHagG5SkScqrk9Qw
InYUvZ+pboQ7iXy5cCoyoXWx3+4R+tvrZP6h5utpYPuP4p9MNp8o1DkV5vN0Uc0E
E5Z5JK9NpWnWPOVRJgFJ8Oe10T2x5d4PzluRgeU7xi0J+pHu4rEvM3vAEEAkv1CW
HfOAlyw9knQ85xzWqaJGBrAo47k3eWZ9SPaFVAqtn7/g7h9xG+A2WpEMsf0VIyc1
WVySwNgaLcwWvWzL8BJAYuiiIxcyyk9q+UCEyIeN03F5UbDYusou/K0xaoCcd6pG
bt8yihzsZei9K31pGJYfkg/okJmG4Q+UDqITb9CImuJUoOhBvU26gtfVoHTn6TR4
TMm9YN+egnUeWfj+4VeWe0fa+c2Xdi25VQu9cOkBoxMeSz/zv/CCuQXD/PupBemU
syRw/LMzYkVoRcYjx/WkEQ==
`protect END_PROTECTED
