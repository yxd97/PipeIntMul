`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejX4LRSvN2AazCAx8TZR7b1asV+Me6CKfKK+RYCpnXDxZCb20te8bBbpRh+EOzQ2
VJOPE1+KAYOAFFCOWDEKrI5hbUUcAtG1V1GzBVkLL1Zi1n/KL141njO4T4k/VqDU
NQIdK85H5fusbr8xzAI/R6JxKCb+nfPA7WhPmdC9+p1MmNVrhrCKDnqhmijuZxmP
YvrcvtAXRYFvCvDgj06LQqKFY/JLMOh8lUqpmz1GXwjL9360tuTSZ4fu0NS14nIm
XipwqNl7MKJWWda9ueGDGBwKOLw1uO4Nb1ZWm+ocUoO8EKJxcjaU4DPcNBDMnrU0
8kho5WBFhr8yAg442QuMdj69ZioSTjAtJ8GfqLvtzMI202BTQRMlFpt0Ys9kRGml
CApKuqKGPtw6u0o+LxwufvCXdZvx6F7nQVs/2FebfnC40juayYL2abHweomQ0YRX
/8ScMFQHpdW7vqSWT6DzfDIyp7FNeC3btUyyLCdrxmNGZJnHgrN50isZDKPyGHOw
ZoW0SsNkRUTDNYt4Djpefd5g2sByNT5hSekfG4F8sT8XolOauJ+k1TfsTlw6GrR5
3CdA3IGnrlHG5bKCgI8FILwm86aUuSIU1vmK2pp49rbu53KULGP/fipRI/hDgx5s
5NWaKQdgSgml4e3Xfg72TrfGb6B/z62zwX9DhG02JDKiM/xGCEY1JGszFVFZxpld
sDGqb+bIq0dEE1IsC0OUFG09JGJzEBHY0amAB3ww7bHwLdc3DVg5E3hfe4V+56Xd
y26Wkqk3+qtJTkpUZweDH15gVwaObhN0AEBep78n3Z3fXp/Ee3pkTSGbBY4dew3a
f41WleuZ8jG7xc9/8yGLiQ==
`protect END_PROTECTED
