`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sX9gU5AnteiYyzTYPbmgCP9LaXoq4cF5H3kP0cGRXyHHArG/c+DSw30GegLIjf3h
OojfRmMLYRqfd+fcDQSH+hiFG9uCsq+Y7Gpg+MaE+U3aNdyIgoH4uhYuB9SjZuwx
X7Vr5tUpEJWY40wqU2t7BbdraNdkMPjvXzysw6L/fNpwB9BYz83lgvAUDH3VfSkH
55NIOD/HnEfDml/fK0UEgpr9IpDA7mfc8Hz9WYOioBI9x+sFGic73IXxoTvQGXet
C8jgj4s0DZKIEN4PXDni7EVbgNJTyUzvXEqCa5PmczahJHVIZhADoAUeatbGZbRX
QhPkazP5q87EUEm/q/XQ4KKJaLonUiRO+0UTWcYHVTlbOYbaypfES3ZvyboAXbFP
relw8WBaa4OH32iusy4EVOImr9EhujOQKAPhUOgskzg3LA2LX+CH1BVDk/PaVd7N
Gp7ZbOq2VGVRohifgw68NsdAakqDqmHvRhUhrzBagfnjN7195PKjV0pGHNn50fmY
nuD6/ybdsWdLl3ftI0dExwqqkQjR99+1cKsVOsMNIeA8msNa1gYwUUBT2cHm6cjK
88wJlWM8xJtYZ5wx3nDWdljZz26QyJmnP28ISjK5BoecToMqeEbmqIzN/B5URSZ3
AivxMFfrArqKUIP+QLHfweZRTGlFTXgC1EN3MC5iN6MF2gw4fNTN83WvFoQ5KGlU
g27XbXkXNgLu63xoRIJlpi/NcSyl+4Wra76xedSB0oGNQ+a1XRiOyrNL6np/ZFnv
Hz4DYazELCUuL1hjrHwoS84TINaCd/LwQXuApjDQHQV3Ca04rFPE6NxORxKqWLWT
ZZbJBsqui62fkRTGCXnLITL55Tf6+75VNYzmXbncgt3LGYG2AnTrfsxaq2+8WP5R
69FBedJfwaIAH8okp87P9mDsOzGJL0U/5brBuWyKoxXwM69fZKeaZiH/bFhecFaI
DgK51WE8nkvoZ32bTfv8Kk1IYkD2H/ssWYSdzBwYALcnUtcdKB2o3XroUQGv9Rxz
s+hTUH1hTlJNzUSnNqtLHfKYpoTb7jbBPoK566sOX22HfXxgp2wyFOBMcHnSCFAC
cSZN/u4qsM5iK5N+sBSUn4dD135S9aY+WfsyOKwiEoixiAkt8HdsNaaBpNIN9iZE
9klc9c8dKL8C81Wr+8XwHZ69322uVey2G4o37K0I4Jrsv3le0awJVOWFROs4iBwy
dhDWde+Xm+OunaA1Eo+p6LFuO/TnrzB7jac+X29MFB3Jy1OjQH2yCbzNfYazL1dG
j208HnQLEZE5PHGTWUCszGwoHIoSed4vY2Ivy0XumYxqO8Tt9Oa/ukkA+ck4U65N
2UjSJJf1MVP8VtkuFgQ5KXdOqamDOarT0pkUtFzAN79EZv1xQTksgMgg544GFwJt
E79U227M4ALikvkoacUEjaHEojP0K4W3WQ7CK2LsuSE=
`protect END_PROTECTED
