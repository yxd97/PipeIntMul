`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZyJ5DJKTSWSJvSsdJIhIc+AuajmFb9rMzEkaOkbZME4X2k75ZMF/ncTt97pROqF/
/d54AbUPIi6kqAsWVO9EOVU1Lk4VIO8iT8T5oBgTEVoTzV/1ljKe6B9hlfY3gMJB
sWzNG3xD2mbZTwOMwWS70nIWLwn1ei/Fi9ehsLRdc1bTWvJHKpoaYW7bSDwb7NJe
GfGh0f/qyZgBvNrO972Z6EGiJNawjmg2tn1WgUlwp4OcqEWp2nmCdfV9MkgY8Ct1
p48vmfwOAe+gJxktw0MgILwqO+u6wH0rSCPLgP3DNjRTgc0lEMVEeFq/uDdnJbyI
be9ZP3ym2XV+wVI5B53kfA==
`protect END_PROTECTED
