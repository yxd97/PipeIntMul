`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AKDJCMDtE7gKlDaYDJO+CziBBsWH5Ww6NmPeOCcUczlsTW+vwUSVlnv2jE2BW0aV
2n4qtNugYD1ICxj+Gx/pqn9iyjlVDsUeSxGGez0mCkwX6XS1Xs5bOxxcdg1tdvFb
5v8K6YWvpZaVQhM/tki+GL2AxOD4syYeBpGf1Leyv6b+9lDKjENWvW/wN6VOrZhQ
uf9A+aM4k8Dvim+DwebOwezq2Z1saJkP5p++nMUajPhxp69zIrUy78dmI52eysKX
0C5IKc0wR1KcZX+3hgudyd1cH9YFQKz7s1ZqqVdtHxXOrDl8CLKf3twukFof00eU
hLn14XqfXLHyoRNV0ytYMyntBptVevbwBnAo/kSczhEEXDBHX74U3K65RJlKDAlT
jWr/2uQ2CNzlBPCaZtN5wpstPlMGljk6sQSsYCK/BBu5ChRM+c5CkOzvwrWlNR64
LYARR8xpLeQCX++1hKkTArqZCuH4E6oYn69okzn99JVCf2KKRhF/4u+J3Pv5bTPd
9skLLLmgx5ORSV5hdaBblyP7355EisnAEhefFiELFuHYqqZYpMBbz1ToGgbOMSye
p9QlYz0MsqKbJ0HlKoOHRLcP9QsbYT7/ReM4m89KEEan7y7WLBs8opyuBjDo3F5m
VOntrNCcO1/eU/1pgYRQS65IcRPj/dRBz2lXRF0mecCe9b0lLQPyIYb53fg+F1RK
wfkaZk5jnPRrcVJzqHiDbQNbtqn6/3W5JXZ/N9C69uAGdPipRrj4Rph8PkF6aTgp
KdUa2I7NhNg4bAGdivrbGVoKMIDuNH5+Tcdk37olfNZmbtVEhFch5FP/dfy4+B7C
BRVUfVDle8Dmc7Az30H4lybcoOPX7HVu3y76GNbdEQngwpZbfGpRCnLCaWnqHkN1
3gxOLpcMz9scNimqNENcQNC75Exnxh48OmvRV0KL5JHBSn61kxJqiJ8RNKhqLzLx
hyjF7rX3iOPEdZl8NLgbqkOFQIyrZ02zvnZAyZCifULvQp/WjPJTFrK18KAFebV+
`protect END_PROTECTED
