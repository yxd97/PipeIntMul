`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9PfiCbsPEit9Ifd0QY/n9P+pexQrPHechTOs92gTBBTNTTikJdasW8XQNtB294op
2e6Hki8QqusJik3HfBtwgPOwrM6Gad3rM1frPHTMLKb9iEkEQkb2kVu8yZuMFnJ5
QTseGDjtxCtQohQa2W5V54OXh7tGIZ+z5xcIhj2QCbDfyerhWT6egJItBAMtxCp4
tpKK5iFTGFNHhZ+b+/fTPzD+PLcWFAn8mfLIAwvPsL/uadz2J53T+/m6AieRtHkP
7KLgwuZiq7CxqwPbgF+PMqfq7Q6XBNadf4mHbt/OpnM=
`protect END_PROTECTED
