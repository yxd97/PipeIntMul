`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qedH6tXvS2uvJEkUiRU6QucFdPifh17A13qcrBpBjw5Kg+SmwClw8P2NW2Jm/m0n
AeeY/QFK7neYQx6WE7PvK4dr7pFu3UOenylCOd6VOK6klAJR4Q5al0slUDFwTd/Y
ek6xhJew2vaJaJ5bsFlx67RE2NohRIrWYAabgtRXJ0XuZYYFUK9+hZ00Y7lO786Y
dIY6EElinRuHCl3efrzlNslXwKgiZ9p8YHtd0iJjd3yEBR+1b3HUpsHwWuXxus+f
w99ABabYspAkvGS2Sb4VlEF5TiYOiSg3GocAObYsXgM=
`protect END_PROTECTED
