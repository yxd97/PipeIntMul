`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x0dtMlR3K/raAPmNVhJss20u5voIn1KQIWB+Ec1ZipOoFH8QK0DiupD/zwbIGclb
Pr0F3yPmV6xBwH7Idslu+JE0auEhdSZWnX6qvASjAAEuw7u2gP6a/kOZ5pBZ6uJU
8BEmNG8BfV8Sd/EVWBx0c+S3CbOzD17ccYjHsXkKUaMz+07MGULB/FUvQKrO6sO3
JTg5EhobAJDXKwTdJYbBtkYdC4gYkvQvOdRuLVqC0vqP+SaXIlNxvdCfn7of28/r
HSadbMkfO9BmvdQAjh93HqBX/bKSLr34oB85zHlaF0XQUbNUXfhEzsmmHoF0ceqt
XbLEWlzMMRVTkVShr9juNXoQm9nwcmfclf23TIuJ2zOde4M2HNBH+dIwy7O6faEp
8P98+D+DW4D5WHlOaDvTM1SNX8fwWF3a52YjBH33S895S0gIqybjTvWW4oXlB/8C
+J8lduCDinTZR0yZNJed5Skm0QbJiXNlkolCjpNO1yZ4Un5hVVkGOIWOGKHfOE3b
oX2XM/+hzKydfaSKmfX/zttmGDtT7ombEbeMRgeysbOF8rDY386F+BdR0ixzOBAn
jQQ1zhTd7Oi413xy0ItC0P3AY/xky7PQEqVdcaWmQgBKKj9FpqVR8DCgtOBobNAM
4vzLGsiy7Tb49ATN6Y4EhihdWwvL9stXLH9HjCZBFyj22TDWkGgw+FDw3QTgkTkC
mbeOwa42Feoer32WfN+ATTYFXxYw9DiKm25pXlfQ5QNTYb6YFm6J2xgl+AzjYgwv
F8jibYSTT+Xadr2mNxmg1g94Kd9fWi7GtS9S6morMb+WgIShom/Z64cjAKUp9uaY
Bqnd1yh5g0Wkai7OoUj8hJXgXY7Ax+/jCfTx6N0jHE4CBerhnudVeYc77P0ZJpIl
hcAPpL9r2FeP9ermUuPZPEE01ill9C4Lf4m3u6zcYhXyVb4W0J7StKrmyyirvLuR
DjVV2Nq/MHI1/TOqUNepTOnWvvwbz+Ji+QPoMyvVeQQ/mElhB3XpPeLxMUE7WZg+
rKwUgOLTquYfQadG+JQQCWDF+/KsnJPK87BQGPB+3NmnbQ/i4HGw/riKG6+epVrn
vAm95EbNSDkzKHi6JEvX0sYVIwiNf0Fi+Vtzp3OPQoWbYSBz7PYE3hpcIm1IEIHC
H3BKVIbsX19HBJhVhwgJGPtBdecxuwd7oUTHbb0yjCQaUjygsEfb4ijOAWlzsap8
xDDZQKXZ9cK6feMGI1c6DsMeYnCAkv2Vo3IMWDem6RdOvf385QMU8/Cy73LWoS8N
4prThZRF007/nHbKFqhRGH08zzUnQpP+ph66wJq6nnszwftnYjIkIZEmPWXBac9I
vrlYCw4bRaxE63u1L93rpuQH395K4m3MZlju01eT82kZ8ifN96xa/NC+vXMzSUpp
dvxuqrNhH3WqQ6jfhmtP+cLIldfxCCNoDZBXLrqANGVpVzAmT54c8gd0pZ17lVaw
Bo6Lbn9t3iwJww/W/I+HeIMf81eU7uD2SSURZ9RXXH7GfNKfSlbvZYrT3QZZqE55
1pJCGR/90yF0+AwSiE/GhSUrXswDwP02zlzRq5Y9MLdbat9aFPYdcONlxj1uO6QY
ZPc/yk+s64PN+NZKTjXWaVLkF/8qQmMSmg17uv6QHxAYsPM1g5fqJl4UHbFGOwjE
8j2aBdl6Nry+utHFKjUJozBP9d313C+axU6n9A7SNp25lK5j7jxxQSfl0ho1WF4A
EmhaPo9/YtEJaLLk62uxlNu/EM75c10J3IpUqZxOtKQu5opnSu9zZ0DkFNzkmmrs
nRhDDb6xh+9seEUlayAEur85slBx+pxpS5DA/ccQr+buwpxh7mCRT9FuYvCejCxz
htCxWVHzaTsSKbNKwSubV78FFNSFb1YrvSrvV3mge3IHZq57P/rUQKucweiVAo82
ou+kC8ub5odmWIRXLVxeEeUpqXDZXWARTh0Hj9sRs05zjs4rLeR6Nk0DuoS+HaAr
qCNUV17dzovHDDTWL7tX+WGATZZQHrFSfTFI6j7mSesLDanbKBqFebynYQ2uFqYu
3zYd2UMAJy1ifFSlmDd2akv9vMGISqthOl3Q1l9Mor4ACYPnu++Elm2AXtBqCZ9p
/kJXgb4H2r2R/GrjUeMe4HiPIUJer3IpE9BNsE1fuZKwgnLDDHWJIHugdgyFORIr
f3bKpAoseBAX8R/SQ1Ab4HcNfuqiNOGHQGMG5pkdu+IoNdtOknjsc7Nfh+1iCaHG
zfYLo8MqzPjnHyQobHh1ewV4GBeAPuDfDcSdONy0QJ3MU3y0+JmF0p7ytT8pZe9O
kWVuMi49gKW3X8g4w+27OqQ3ZilVkr6XLitWyhL4ddcS9kuzneEUzLA//FOIBi6s
9sL3m60Efoof87cccjCKTVI7Pa1AuBNBoMbX2PlqE0Zv0fspPRd0JwXaE71f9bxR
ZZx6/Dx5f7TDiWjG/QhzxpedLEqFO2aRrXB+3+I9wCdWFvhu7QhKO+mp+39rPxRr
gM2J5DfK3SukwNiMCcjbVd5XcMQjPaqiTV2AYozWo7hLnLtVATb63ko1zjOcnkWl
H6qhOome2WLMefLvh1yItRSLZKWVf3UziiSCHAlO2DeLWbEU2zrlbNQbKYhHRthi
7ZrGQedXeNc/75UAzz9m8q1CKICkLU5Is4mxtM9LlfrS3r1L3YbvXZMCcRUo3k+7
aC8N/+9sYRCxEi5u2Eo7ZgHybuwCqp431WgiID9skLK0aS2twS/XdlymxZE/8iXA
tEckqCDZa/RZxmtJ4NfnBlwohF9yfO/ntYH+pObrtND7kPATqgYEcl7aLmyA8OTC
LpGma0SS6bqVcfz4rOzHRdg79TJGdTqr5MhAXc46HePgXTOyUwsO60RfgwtYaWKR
8kYtGDqh3h0iEDHdruD3axwN91g0hhmBngoubIL87obKBsdw6uoyfAds4mA1rnv2
KndBb7Xoi0QlUji40lcenNndidQeD9T2dAJhtdIr+rD8RQoMXWD0mrE9bLF6kPTm
f3MAYcOyMpQEfS8T7C4modmnaGpr1QHUpM8PqoeZun8SY2GwfaCpb45UCtNySNZV
PkRDp1Sckp9Ta21/MkETNVAEvNQSjsPBJhO/2Epv5HixIFpaDG43QWypRqUC3n5S
cbi6rDy3ZCd9+9eiWJ/SmvT3QHZyLdljsvkIJ3WVJJEWea5EzNmlJIF4QgHrr0V4
M74zYHYIuZKDudiYdScSd2nvs9DmMbW9zB8jKq4k+Q5fSuC2UEKxx70dsjVNqkme
UoqCU+vLx2+D1BmsOKMwJ1cA28DbzMkO2ourLmyt13mPXloKHlRRmN3yiFcA0eow
uwYWeJrCsp23NpCaYz2lrJr/IVJ/fctSVRpf2aRGUas+3SPSZ7wHO3VYCK5EXvwj
64rUb4e/Bh8rNJbniBxxj1YDDqHxOQqdWooKRIlZocr5uf+pTOMvvHxGyeQJJc+c
H8V60wrjbFowkzdYDjN0yDIz53fj44TdjLx2cyM+22ofsPsp5LnviC113XzAqG0C
5Zzz7h82ZyzO/gDj1X9rPk2Adj/qksRrJ9RMZvmsJKKuJb+65DpTd7B6yGZfFLuU
qU3cYbWSCu3PkxhBMHykC1Ee5iCc923T9vlqLUM9RB+lMiK8ER/Hat1DD+TWhwYW
TH521NUhV3omr0YmpKatAlAgHDc/g0XY30ljJD/FfOzj96SnR2KJV3zG6R8BLGFb
V5w6y6uQge+1c1XITU45MytJxwuRt50vtu46EB5gVGSK4qpwXa4ctIemFkEe6xhX
gQGEvamnXFg85OKaev7WTA==
`protect END_PROTECTED
