`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRb+zIOxHtOt1cJ5/c4QMCAhp1SK2fHCMV9jLsn9YsoQP+Zb6X5BaIlXPfzuNT5P
6s4UpfuRswK+9WxSThM8ov58X8WCiiDgt2ddFsSakh7XgoGd6Vw4Pb84Dov0wZnG
xPOFVyKEQ7uI1xAyfS7Af4mjmontJ0XB71eLlxs6LfJZ8chBNURWilvdm05Z2ei2
5KR1KvUrwwVsrg+YWGoKbrs6ir8lmKAKCWOdml7CXvCXBe4Vl41eRvZqC/P2FKWt
CYUYNyMw1Qh/Dg48dwYgNIu/oVrqK8trXhbyoH5lyU7U07v7eVe+DQ1528OBmxDO
4whiC1rsnURbt+mv+3sgPYWNY2KXP/Uq1rEpMdXvkzEYpaCo/5W3ZPrU2dk41noS
c6BL/kSfnN5d+v5XnPyfq729Cl8Mi5+bkIdTwFsDcURsqM1OPvjFx/wJWPYlbuFU
VEh1kyLCT9cysRPky0E7Be6zNiLGK1SIDKtKjWor0ijPwohAiTWJHJmo4AFwa8y6
`protect END_PROTECTED
