`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J6Wc3Xga1oFQKYRsgI2OzSmTjiIdEFcN9C4pVir83uSYdnKXHKKZ+1KXd+Akw4Kd
qi6bgpe6Ei4m4ACrOXgswqfwrz6TuSn4lUFYA/Hl1Fpkl39efDv5cGL6xqHELdME
E2FrWUaYnjDF79jIOtys48tsa1c/v7gQn5dfScRM3OcKhI9wYH7fEZtRWx0JAgxZ
gc2Sddo5NI1eWggfc3Oii9m6Fru+PIVKqG8WKwib1H3V8xRv5HjEVjc/G1TlSZPq
X5RrQ7I8DFBM49cI53Ds+mgH8L/RoXWTWqRJT5G4V+DLVInTHJxv7arqND6ec1Vr
`protect END_PROTECTED
