`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8K+XXCM9vATYNA8zGq12KVSx6yLPSs4uL5uIoBeN/A80yjmE7igQz7UzToxN/Ic5
bdwb2uIe3+pv8+3sDP0w+LtqbWUJq4crBqHYhsN8hsaSCPxRmr5ZR3TPNSPJPTm/
EY3mfnsigVoqY5f6iNu0fge6pxP0UO/V5KZIrvpScsdnCKRUkK7ic42bnV0ocg7k
x8Hf3VJgOya7OOlw+BrnOmabWMpZKVXsNxrI013GKqb3OQLa4HzRA7EM5JF2jU6I
Pb5Fpr4L146okD7vfkHe/KK7+0JcZ4Clsv7RR+VZK9ga14QALJbq7XxmF1HPlE/o
qbVM0zEazb0iijmOzNkjwFR4oYijDZFNy59d9+SCSd/8ie/MZUbUn16QnDDGHY0x
`protect END_PROTECTED
