`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
faxJJ8KSPK/qX5an5bviVIhbt6BCi99uW3B2J6uj2DKzzalD0chDwtc23zfsfBLz
/whrIsTaoyJAkXRKj0ZQvvHlBEl+hQCCl1T9n/Isgykf/kLPaqxvY4f4UDyiDcUu
1YAi0Y/M5gZMbeJy7c1xOPY73r0Uk5It9shgBV2lzeWfPymNdnSn4MrhCtTJ4b6U
gLTLyf0Y9em7TMPqAjuCwrPpgAb8AiCmnU20Vtq3S9BHvYcBbibchaCPbt3aVZnT
dOE0DUpiGxhA6TgI2uYPzA==
`protect END_PROTECTED
