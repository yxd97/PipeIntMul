`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EaKi3g5HttzxRkh1XMEkmGbaW2nMpxFKj+idrB6HHXLXT+7kkiPXqnzqfUQpg3PQ
Ks8JDBoaH+I7q+7nP9S9LkUjFUVkNeaoP3555/J7RKyxqlWuSwMVYAirsAACtM81
nStO+yykXLbqg+2nmaEyhNh84JhSfoJlTgmvLgHWqtTGV2djlQU25ssNLazhm79w
TPCcwnL9M9eTNCmbX6iwNz/MjBpxTioY1b1ECm3XBSEYr0j1rcx2hx3lTzCGDz43
hFr1UYJxdk73JTc9iEA610KQ/jdI5QmAdg/BYe+W5G4Xl8+Kb0dIJI1yRS8wAKsn
B3x9ZXmqNbITnZUKOO+wNLeJB0y46qXhKj9OQCWmoEcZk1rR0o5ddn05w6bDfpOt
judF5dSRR2d2HXN+tmeVG8gGlxhePm3N4Mm9/QjeP51QV09WWmFTOqJ4ILZ2rWzX
X+A8MrvITJFoAINOejGxZUCUDqvtgFKePUVQfredPinfo9A35yKVDPtZMHkQns9f
PLjeGt0XqOC5PhvdHLkSvA==
`protect END_PROTECTED
