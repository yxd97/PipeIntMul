`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmuFYAMmu8W38YK4kk7Gs7UxvDAUBuXW04nLZYpPRI3FkQi6aMdyUse6SEQE51QS
N2Hy1m2d40sJacjLy8YrPYwNyUWxWVCr4V08LB287j1jIFN7jJaKzVHhCMaKNuEj
PmOC63Yuhdmp3E71vigzcsCQ8hr3HGFHbLNYvkUZaT4Kpes0VvZ6ftUMyz4hd2Jq
0KgmjJyS3WT42uXnknnPUfxZaaEMY9rhzLdcS7UFRwZmyzDFiIDRHcQRbBhjShs/
`protect END_PROTECTED
