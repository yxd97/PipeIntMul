`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fUxNrcsnxnDUkQQ2tUfkKMElnFhDhH1VAxNEU3Tzjk8JbNlQPH3s7EVDSfjIg7hv
Tbl4PggEr8S0PPA5Tk1VaJGhVPr6v862s3jJ0Qi9Nz8DEN38kUis301AagS8bUBx
iEDtkk1K7GZB/uX2hLQxlgpEts9Kz/ED/XUwNucVXhCxddzMHmNbAeU1JbXv0qjY
GI+Bu6NAfR4prv74FUvAhiLhDP9zssq+/aaLKWS/NhD20GPnWFbF7GkOUplFwVo7
x6pLuRIW9sfMJ8D3d6k1O3a1L/8cFKbQIc2dRSCjUAxnUc2G8kula+SYEuPfwRwh
2qysIe6mdAtKEOquMjhLk8mUmSnsZMrDl37kTK7WLhfKfl3QduJGqvQyixQ7/SDY
s/9XasoIRSQU2wlqyZ/qEZI5u6acB2tFCF/diWEknCAuckVLe8UCcW5dIguZQGhf
8D+6rfLlQ8ORJSrgenXOpIhDGaKn6bpez8MT78c/qGF3b4yjGp+pvy+JdwNHnFbH
n4yxiAdNisVMgtYf+s2D8RTfhRMsUtoLmNIZDfQp+LZHuMCurBAyDNZz4w4gafuE
mh+JRQnhJbT+nXAKdnJbMFBytc1tF9Mv79Mq9Te30R1G0++a0dtt30+pf9pf1oa0
yFcyme6bh6SmBUWKBBP0FYRvDsMQtOCLPMlv/g7K/C4jro+iq5Gin4Y97cjHBz1E
7jG4RnT6o0gu66eYa6wbZ4e002FvRuL9YeG06IfpwqklGRhNB1M3Z6EziXcQBk8T
eMLuAfti/Gb16f7N2VGM7A9ZnBwiHSMxRrlD31KZPGgUED0wMzGeefUbM1copBHr
6QDpYTN0x6Rkz6bIOPPdzbAjQwJ9zoTC4TYDl7RNoONG6iCrv0MEGrwrJJolPH9u
jLpEcMLUTc4dLNyeoLw4NKhB2KS/RsiuyO9UrsFeC/KMvCP3eogkMliZ+2ShBMNV
8YrKf2CijAmyRDhTzD8F1DhZHRLsmqkeeVr+NmVRcov8IOuS7ugGtgwl83Xx2oiV
uoEg//SQucnCDpeE63sP7HmA/joHD8zPIYl+dfYAQruPStCR4D9zE/qYLEcK9iK9
jhmOboVLf41iZ4yQa0OfCkERHrUSLAmGKqomNSUv6yL5k2xqQ5rl+pQ7VOn9YR7Y
sJ7PGKqBzrIF1pWuMzEWoTe0O+nK2mHOtdmcVoTcBW5XM9lxXGrgOb3XCZ8sN4dg
DSSZlcJPgaQNsZJlrEKaZHRJ/8M9b0ehs6unEgb6VSTzqtKZceAzhTG+QmV+2LFi
JYm/D7ZTtfrq16aduxq3vzcCRlryKtp0XfGSSH14YOeshaTxuW/hUilwXdSETBjl
wBpNRyetgSEWRJjw2kKl/uQOpnzvjOQU+hq15RxTEbU5RYPVHUXtygzltmGYOpcV
6l/rlAr5n4LkOllIkpVk2SST+v0EdTGhXoCJ95BBEVSipZYCmkFwJe5HiLyj2Wod
WluFsOXJ5+GNosQZNIVIWJTq2bNE8HUTpBNPwuV0nrNF3Jb1JxfrYsk7k38R9+JP
VECi7oLPQfThKfiC82ytU8ijK6Ull8m/jvSxFSCLhTHJRyJmFBmPvuoT3Jx6hKvb
5NNXCjLKoVSZd4W+PWz+yJxFMlvc1kalY4lWgnRkQ0dVYG0Q7SFcsqAs3DwMOAaP
A1fIHn3pxFbdhnCg8391vVor/Kvk0o/WHJC2VuizGzqsXQx82zp+oZNRED041qoD
9DCf0uLTK/qh0UFDWFZW8wQpF2CGwMqhR5++V4qrHDlIMNehO8fbWwWhp7w7J+A5
slZw4BDkjtL7BxoEknUy4GvCVaWL8fxMRJwToW3RtsbsunlPdaXZF95WwD2HrK65
iTJsbm4VwutE/TgyPZOfVQVniLzPSbxUXn3a/c21aUKy/z9HlZDceicVJ0C79M0p
4ml64Iih3NXjCgxHVwdRrw4kT4JJJn6sXoBK6Nvj1dUaKTyXnA22thmInop0PCFa
WJ4+jR36NUvtyjtlSSFtWDWxgTLaO+ujGyRXdx7yQiai+sgWClcRfbVQxKAibB8V
h2hMxguqDUQOeaPNJIl3z4nzb4M97V2T82WsgxKJYv21oLxA94fyZpVoSC5a74x5
NzqxCdQoRcKLCUnsYGVtaOimQUZVb1u8lWAbO7xBCGFmSZk0/wtH9CeqRpowX9XT
tJ9OhbYqkCJIFUgkldabiRvI4r7fhe1tcRRdgpQFZbMAiO6bpHkNn6Eh/B3ypbVO
egt1NNXVexzI85UzY44Sep9UIPZ8oEjU5mEPL4qPP9OLR9i/Xk2GJG5Glr0psTuk
mTjCGNcqaDEJ3eA9EYMFLxmFMUPs9vwszG+fVCrnx4isx3+9Jn5eZ+jL9LN2eE41
ok77GZ2eExnbrrsyKDwquD7pToPsP4FycEfZx5mSCw1tRe90GWlKN87UKFhACsJL
pzYudwzQSKa6OhJQDA7+r0loXZLhZMvuBvs62YIuLzCYbnX3693wovvKN5qnVTbj
WPmnIcESYIc9rFbtA/ft+pu+aac3kwzSh1b4qBchVAh4b5MhTRqYKEGpo3ATh+xK
aeJ8dObBXPjOvjm5iGmwzruQmapi5eD+ggYqzFTYHdkvQNkVJ1fCJwPwWk+Tfjc4
rT+VPnhTZ3+f5jDU+IEQd14XXEAy0kaDpjp/do7NDpi/P0ujIi0bxtk6F7PVRTNn
f1afvgndHWOdR02FxtlgbkrE27o9EhiI6Zyh6xERaiDm9vWJuJ+5wbDxoopy5q6T
xj9NC/Jqnc39ySB2h6FROTHCSZMzHjJz5RFV+hijreATyn//pnVH9JBVPURxrHBH
RnrLzbn5u0D4RTVfD1vRK5MSB98Zew+P4YFRUwISJRy7VR/nZmX/GyGs46lDatJ7
+lkzuerQxF1+sXHSEjpX8bBtozH6fnU/QQMzXOSc+TA0kdmY7d4G/aifjyYWjUcC
f/IZ67lr8nyKVbIDKwiVkJoaHvxzyDBTfzAmfg5Ntnkd2YJ1JayCscLc7By4SF3j
beGhD9JuETi0VOo0vVx0+iO3ZTzleMDvmbDB3BYtYUUnhpyhoj+0svY7cs3WbcEq
SPK/QvsX3zp80drSSuNHoUKDQnegZdZk/x4qZCLWLIgNmVTHgBzHMS/mNrL9UgR+
jzFEV0ZgPeJrZ669WQaVUGz97zu2dCIspSCGpOW6i3cN/BrXlhg2Xs/ZCq197n7M
7WJetTyJpOG88cQpY7WOk9SSBNHIZ1i60Ct6psF6Mk3fPRG7mrLtTeDJGAi7KGmx
GPfSt81ihyk+6AzPlWQ4yB0EAvQRqBInAWDt0zEcJfzBPzNjksY5MUWKjqS4M5Ux
iLPxePGEk0WVzfvRAkOKKhJUhx30PBWm/L0Px3Lyzm8F7bsuSHmrfH7/2ki/rPvw
Zz3XiVVMqv0hWzvEt4/tdQisGqGPqOaXRDo5cueyEK4AZ+A4SbLVcU/RVCfy1n0D
OUDVRmRITIrwJXEd+f8cmaaAyZEMy7K2vQMet3DhRHsYnbyEKYUyEXlJyRq8nupw
6JAiyCI4VM2BMNCHErQ3VZqfpyRv4UmU8AJoTcQV5hqRuJNrUAK38ezv5i1IbhdP
zUTSswiKCEYC5Dqj+eQlTGOFdmVcMFUlpZ774vkWVG+7AIMI1mf5ICFsYTT8TK3v
tBwVjMUXxIC8Hb8huuoWkgKTm5kojKU1MbdKsuRIWU62eTM/BdkEyQa3lLxBnX+s
p9FJdWgb5kPlSfnVOE5OcvqnAKekLZQPRAwN0jtw6cHKd3uGfAhjbwc1cKkmmLKU
RTyzICQSp3U5GExVzPomscU+X+hfFX7JlzxkwcCaEparQyxB65A9AHjJoHF8VXOZ
mbAk+WhcwHODPybUlPAsUsKWHEg9tyNNJmZmrCAIGDqTsPfjTQCjCfFlZr2GjvWy
oDzChVOdWph9sm/KmyGBFBwL66qVVHHRvWcViORnhUM/SM3QY1islT1Vp9XNIejd
5zMNilUJDiSfE/3Y2dRA4CSJ/VNeuP+hwgHdb0BOMwTz4IWtNHTswbhpsTECMP/M
tfc9gK3AWCTzSVj70WUGWD/HVMryF/4hblToUZunduPCmevL7PaD493vgJEpVxja
PYJS5b75i9dKQnGe0tR2KrcjL5MA7+KU+2qRQFyjZvYcSYV73zOBD3+H//+D4E13
1gkmI5LV9yQ9U8Ph+6ighgPlj3CmxaSnDncc7OaX7JJ7b2WiXUph/CFsQGSANR1v
jasuoKJYTPnjUARVOj26a2dNKiG31JtrJAzzldbKmem6sI4q0jfr8DHeOKT700BJ
MGWcRQzJxISjYWFptyum/lMDQmYt/kbzQKo66mh2fyYhaoCs2TJoxUqUExDsQQzD
4zizumbvWVuxtKqp4foYpaQTmrJjjFs/VfGcS3PSwaQwDhSEnayEaeD+4ExrLZAq
/VtAnzYKkTmGJ23TSdWGozqc/XQ0VMf0LXEzIqrl5S7ed6/l9nF7x9SrBU0EKiQu
IRY14zVp+FLj8UQe/qu6ECRnxsrgDrjlAczgV1MIQOx91677z+8xuio4qHoEMiTz
oNXsFFD/L6/NHwLvP8CUrG2q503WUaEjWzlQTi+GjTEReUBh5CMhABwFuFHik0l3
w5X0GkegJ4KSHgwC0d7suz55S8Ev6IiilFFL+pJ9WpjpM2DKkbNwGZsd3qSQmo1N
8HT5RudZGhImbghhx8bg/B1evzNScNrrELtX0IyTuEfsHyTy/+ydrBGwkK7ssoFl
TbjdaVVIk5AyAwSu9l/COjp/w5JW19s3QybroNtQZKAI0a8HMoo9KW+YqbirAUX6
aAquOnViKYiZoWB3tdEPvFbVBYRJtItG15q0+GuB2JhapwJqPQJLVDxf0OAm+FcH
Z9kyCnlA/O0wpOfu0WBdUWAAvEjyDvla8/WnpjEXrAWk/TFCAd6EvI9G4svxGBky
xi+sA/HsMVqua4PWQWgjAfg3e1qqK4OaSJY7TOKwaNeuOV5PZXv7jCtWhTGRnWjf
R50R/ZDiZJMSVFoMP7Ivktl9GK3+bEvRGMQgsdkbwBu8wMjYC/J68XlJ3tNg4xRP
GOVegzNO5zvcuzfj5MlaSrfP/xu4fiZoCsHqVfQAt2APkktGV8BESwVSZMfmH/yg
w9uDbjn19JMRhHt2jeR4kqPP3FM4f89LHYamdGjxpYYCGVDd4NzAcmes5H/DA/2d
NCydT1fz8fb1LYxRfZOhRPv3VZmf+D5g/+Gbmsds6OLf4uBieheAosJjHSJcAKoy
SqjOcJrxYgiU0sob2ALPgMQprUnSaHrhup9uV68MDFBLSO0VNiyhrEnL2pCn6Cm9
f+V/tZwfpgfeIRGH3uK4vJlFgAomGpyKi4mNGhk1uzrN9djoNplvuqJMEULc4auc
YBsANjYjeOnCZAL9guFFD9zpS5DdElnjyWSMOOcj8//TZJYyrTx+5WeREZ14uIct
2zNl+60rNkcGiEBG9zHqXBgINbCCDgarRvWzcKm49oeK1vKPdGgnp92Q2+d3xj7q
80DJ0wu8s5AevQyN2YvU2pwQZ1g0oLRW7toTCiSEplou5dMg4HsyvepXWDnsDm6H
RcE5JjA0SwadulWxacosV3CziwTTjmW8GqEtq81Y8Pxp1Jnp79HpLsvrU2uoIGhM
PY8VilzeeYswSmg9uBXeklKg6nSJPb5o3TKKFfP+sfSROj0Dd0TBvtDslb3M8I27
9+Z5VwXLb8M3FI+X7yzLcnN5Sq8bmD8P1qvBTALX123WW/udDAx1vg16qsC0FvYW
XEQ5iwSXZz28O1WQGQ3YjcaSq1liOlbgYDyeEMcLxF3hIYGixtK8sW0m0bxciqZX
wRbK6Cr7WXmuw8CynLN1mP74A62uz/YwboWZyQKhx+PaOwDmYTY5N4gWyc5ndXy4
s8wVXes0W2Ces/vYdRjfB7C3oM3kpFZxy82ms331f1ZIt3OzMm45DZWmza+/Ag/t
iOBonUiK6zFl4ER9PTTPF88K0hrqGgQbRxa5rz9LiBnAh6vYzQh7uuKFx59uziTd
tpRJew1y0EJd8zYz3sRpgmXXMxcH7lvpgcByasjqpvFUPX1BmR2RxwbI3NI+xHyc
/qi6tHVtFPKIbGU5I2czjHHfWNqRadXZYFiufGZuTNtg7d4gcwOLqy9XOwhWBUDP
mR8tUSCTqddCc0fM588vgjseVnLYr2vMN0XS3LsqXwwrYRSVgHbCvZidI/qqnBIT
QeUzN+EE/uhAk5iTOUEMObBIQLoqc+nbtyXEGdxl1ZhuVn+eyPZG4N3akV9sF+J/
cVdiHScRQSarYvL2TADHIUJb1m2rrt9j431aEtaFCjBsl58rgiMkbIl59aivbUI/
cLN8MCKhPlCLTGoMGgXeoIqghlDQJmr6BukGwoPNT74z0hqJp8LS7GrTBGBQa2nc
lwuncdpo/i2Sgmf0UpiK5loWV68FgrQf0tYWd3N76CE+COkHf/dhArrWesL4VA/F
WS8TzVmQjIu1Yj9PHtn57PxRdWsh0mcMy0TavpSb4Z032vE7AQfH7dgmF3PaXEXF
nBOWdrjPMnITPlyovKuAJrskZ/oJpYoHd1unOlnwZHh+9oaRZZ2ua7LiVZN6tRRd
aG/cdkEGkb/Lt89AK2HEwuO/i7hMo13hM8bX7Zn2Pz+PUMvu5lgh4YxqNSjmOBog
eP47njTNfwBsgyrgVp0M5H+5Y7hwZxisYwEEeeqUbUhNJ5gKWA4hfaEKSgfqLZEw
y1Rv4hEws7QY5ZTlP4Pek1muDNLxOMiKHAY8elBJlO/cxzvnCG3BFpf5bdh3pSWR
0gj7aXk6akCHGvy5PUib2aTj2xNtjw1lGXqbLSO1hay2Dfyckn1k4c/6jrYJlFpN
yGfR2Ez8aIqpWE54Ui5sEucBjxRIRQi4z6Ma2R+8CxhR0ultO9GjMXKsqpTWhQig
Fde1K+Okra94vUoZq0WSoEnnb58QNy6u+YYKMNR0drl38PGqZi+LxcYWk6jfen7l
mF+H/U8jrIf5u9G6TICVMvlIv8LM0HS7sfUicbQIlRm1uxN6xeEEPAOs2Z4jz+OD
lHACHsDio6JPkZQMGUPsvYk9fE8ECTH8n4puLytwwMrKewf14Xw01pS5eIk3NBl/
pYD0iIZOSdqtwZRDv3/cEQsyJsclL07yp8SCDRXREw4Fu+AuAk5WnNSWQuVxiJC8
nPUqogzcivQvTGVlE/XcvD3sP/7cKUnU4ano7pbwOU8ZSGC+yNiZFCCFmwOjUtLA
RbTvdOwMPW0wsokbV3c1XiXjCdHqDftZYlKEpJdfh3DSMwKkajdC20IwmvDRkkNN
t/RHAOQ3LzOYTOKYOKK8WiZz4UFlJQu/9ZaNWVQKv/H8cQ23WUE4Art60rSdyD7c
xBC5eotjDxdJApx2HoR06KDhgsKFjJ2qT9HYBx5JhDCbu/vowDqXo2hkltJ2XBO+
SGBkfLwvR4nLHNjNmU2vRQ9KzkKt60JXJhRn5/z5k5UjUAz41SJ/KKLAAOaK5dR7
RMwLjU+3Mr82DSjRx4RpuLhdLfGnjrjfVAne6+3MHUFzeFuc64H9Dxh5yM1TqC8h
bHDodIDoA1HDZVf78JK8j5NUA6oxOngR0OyVdbVMlZVAlDsYXAFrU69JExeOEw9p
ETou3LAPJRYMc7TYLcA4ntEO2dDDskF7MjxXDUfTW45bpCubRaTEzZxUg+r5ol9y
uJzCTNYZMmTVVgIWTC33Zmka8AqwOaDJrr8I2QoARvKIMNYYTMVZzSroLm7K3tdp
LzDW9rNnmF8CUzd+8Dwc3j7viucs0fy+Q6x99WaiSpYTijysaIg9/bLzuZYqavj1
Fa06AOvAa532Op5Tb6uIp/z2R4T00Ris41MqSltP2288P0wcmGRGnsO/sac8Bcx1
iRzMYuWIe4LRA9/1KNWtMoA4Z1NA/zULvDKxM2nSD44DUtngWiUBHmDbRu6gnvZD
2XENs3wasVWg9/+Qj3P5aHQ0aQkjC1jMv5Pp0EHc/AR5yPry9GHe5TspziTJ7urU
C120A14LCCkerRANL5yg3QZTviZob28zRUTtuRsIuozpkNss/jUWjZlCgvlmDWie
RfHof7ojGOAbtGD1Dzp0fyVUMWx/ofSKwS5XCTPZsxDD+9+g3n1aYHlNem5TRVe3
PJ5csx9mcVeqJtagiFbaa0Vo/kzKMWR3G5qVUCX5Wsp3xvUCmEictdueqe633Y1i
7bxT6CKlou2IoBWIeuanAZXnrrDkYNc0XTwDf8Kox2sok2+hkd3dAgPikIDWmaIb
nGzAwdj+J4KJfyiCPd762BTzYrSNEZKr8S64/VCaSRqKdyCwmlSlj31b/6i6tfag
hez93S9L9magM6y+KSMEH4BZTrK2/nIlo64SPc4ELuqdSkDP0Z5DWI+aE8esmfnS
GatKkP11/aHWNjilcVyReyG5rYWeLHYU/N85ueXmY2Nz3d4JgIE9RCZUB03lOmRM
YvPQWInjgjJNuF6+2t3SOrv8Cx6QPqcKc/5a9CEPhWL86AOHgNjZKsEy7rsKH8dU
0oxBpPKTbI2eBeTiW3quZByEw+Oe1z3LfrsM7erObo9sAvbPLaHHLeyVh0m7X53q
YT6EurHm16Rvg1dlgmMxDjg3nhoQNCaDO+bPx+ASRdCt07UtCGPWIUYSFp01xsDL
9+B2HkUebALlW+qUrXwX3ppN1xFtbUD28wTGmTs1Wefl6kMKMB51mF9DgjA0W0Cz
hu9lmNL5Typ18IulGmUMp5bzJuyGKX14Vrq3xF7TizvHlsMpgIFJD5hc34kQwvPj
RKrVor92nGbzjr4qr8f4Bv/K5TniHv6fl6hmFno5FYugTGVh1Hnv9D1jx1H/xE68
4vwpdk0ZZM4+BW0g9MEUNxt34o11cHNBwDZdOiuCK4aOAcSYIFuOlHrgm1wDLdrq
E3Saa7mqttJZipKMrSB7ak5iVTNgOGFVDqWd6a4SUCDNHuIHFzLdXeRyRtJSS+Cg
+710ylu2nWddu5XXm6b1RVN+c9eb5IECYtxnrpqEhGaiZVhgHD6d8UEJYdQT41Yo
eNcuIvi1/2pH9oJymv6NwwUqgmtXNM1U6Vq9MygWNAlUuVIMKjNLa9nmGImg3Aa1
9aLWpqABU4GhvenviNk5K0YepzUFSg1fGyV/cQNu9V7Dlb/UnzBn7Lkx26NgtDdX
psZdngdWld5qrVI9HZffKd7yqZGoopM5tYZcHZaycbKJjI8a5b+j6HveExkAoeFE
Li/SRSq1vB+eVj7mMb8ELi0kR0Gt6n7jDotF3hu+Y3lHiRSxHSdHwY87S/2Cr86P
HizibuNfqKRVgpDfR92Ukk897iCjKgBva4HXG4I6ng+rnPkwjHXFJdy6uk0k9iXU
M3iO8SKZtZqZzh1D0TzJ1STAKGeGui6f9CHztSmH/iYyxItUwHXS2c+jbAzgUtX0
dA+/WSfounayx3XNCeJA/TBOmdwuXUmdtpWl6Wn8FZARtHSXxddivkr8WB12vm1b
vLTz9wy2yrYoGlKbFacfyJTyEcB8/xwKjOnvGKsiaJ8gBkJ8wDUxvj3vrommkQb3
qd8bpPEcr+m9BeHOHAK53mwJ7x5mzAewnuEqqZ5+ympaFvky9gRb57X02ZgqYAUM
hTbTdPzQE5sh3kXgCWzr8BBoSRVpNYCFm2AE1E9jsizcyTrGOE+wmvo34IS2d2M5
setbeqMShcUnbmYWzdq2mR6R7uK41Mw8UonsmIZHuK94NmLzsD1oyBUW6BVawU5N
hDAfRO3wnb1ihw6OCFCQLXp9HLJvDTWu1x3TLQhHJO14iFepiAPwVJxqwu3I6lzE
cxQ5zFvIPOj1D0YXzNvFFO8TYgaKWvNBIaKxNNtBV2rBQ8RJe/PqRjV458CWRs1g
7xF+3NnAx8uzjnWv3Ds+19t+z1BHzn87ZuHuY7ooIbA2RnsInhkmisYHKx8SNPXs
T2ODCNB0FanA/v1obNTsGcFi0W/IL8M7tjrn8Pxs5EmOFSm6EEa77cF85vB8VSn9
pRLE/jZM5mk6ogdpRYQCD01cghTqhZeEoKJ7mMW+rYffl6kgSGUjrxX/KYoORmio
Fe5DxkK4ssYVOVjo3zJ2ILIZ9KnrZg/ncopB0POfEmFOhaCs0qY29iJRB4i3lL60
cQUL0UKvZ2YFTMzy1fgwqFOkOobthD2xWW5uMsV5aKE8IWPfbE/w+FvWaZirgbNI
nCU6rP/5zK6+CyiU8N6pivZkIUwPrLNTWZuzsWdQ4kNErz3c7ws0o3NFtKahhwyh
Tp+hEGasaCX6WR9DUH+kcWPrrjxoHQsuyUgsWVeSfy9fAOtemS3tJR02p/MMvJ6D
M6T+RJLWtieYr9+16AvVRVUXxwWxUqwLGp+kpoegCNNm6zFxv3PdNtsCTKbHTl3Y
y6KMn/rf4E/sddviP7SMFhehGiKbfAbv514pDdcybSab4kHwEON2VXzQ2tBwv9eu
m2ryw0zAWMoA2ISPJ11vwcHncx5kc/Q1hsld+gzQma3MpEQqWQ0gF+yceIUYSd7F
6Ba/vN2WApFOkJV87edLiAi7t28sjj/60VITkBD8Uf/1mFGRQ/LREYgZFxyK0jQA
6VTXrOEsQi1fdvFBDx9oL/i88x9dDpRzK/oOWn42Lcwcvyq53/CCHs+1pgA2+9OE
cj2pqdUAtnNF1RXFzv/9ilNfB/luM3BQtE4/MNBaZWgCEMOb/a+IBa2X3TjZE2Sp
1PCY8akF/SAwaCfJAFhxr7V4kpScTcsC0Oq+saIgmDdqQGB15hAoaLOVzNVNVt6y
/Qq3YecY5V5IL9/hoC328Ao1Ym08MZYl+uXcoXbsNKchm2ysPoQv2OrjDVSzdSXo
f9/ylDMu23O5wRnh6Tqyb7WN9S9k3UkKYpyg3eTMPABf6qwHD51ZH7IEXjsOongp
Nwccy46k3MvNjiVgR1oLwsssX7JfFFey/2/wpCUj0DGsi7uakumDkVU1dPk538ip
1PDAn3c3Rk5k0EtdLy+oux91u2UWiDMXepw7oXDgQrm9E+Co08RVqqO3kQTd3hp4
zaXcN+Ecma0RarhVeSjVfRN7snjxTHxLRjEZ24PORRQuWeVHZjX/bthMuEsptswQ
fQN1DNanVmkEL1UG+KcpEXg3NhxVdwom92FUuEXV6IcC6RT3ae8BCJ6+o5uyQqE3
t8IjtPYBqRMCVbKHN5kk8R1Dcqkan9gNChGzDUDL0IAUlMNT7cHh0cGdxjNgk635
9l5IaYeMc9OoPbQzqSXDl/SwcdIDfR5ubVh4cs2VrwI7oHUyd6uoJuWOiUTkI2vB
vjeXAlyJc30yEkTgXYngFDn5XjUVVIfmI1C5Cy9fuJIL/y2CJicGnj9DcUCY8joT
Tu5SddaITFOnBQKAjrFEsjDUAB1y4d/wDXwqJAeYu9rAX4FOm9L97y/J0IdG24uH
77MMdqNQ6vUFouNysDLPptuehntnWGI/qaFl2/BH71R4W8hFC86h9hpX4E1t7AE7
38FFY9nUIQduu2Gn7NYaFjmSGTvCRqQ8uWsV35rkTFU3DUUCqXTDS9PEwZiokzYJ
`protect END_PROTECTED
