`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMZYDXtlQTp2Zu8YufBbhNpWRlk/2jkmROy0FziUG+LKbhe1gMKTR4sYlBktIgxS
ghIsRCmCScFkznl6ulINIGXT+InR9JxNbEPRrPYhrSl6S/fABUGYh59OmUjmnevD
GdPfV62MHB/AOAAYL1CLnyu/LuuHitfEjItIIz2fR2f/PkPBHhubFohdPHyrhtNT
yq9A75gYQqa2Wl8DBDz5Z9WFjS693osgcUVczt9x+2jksAHKVYJTlfV9s6yQAPDv
eim5bZw7TCkj9lzPi2/8iDsHhzWIhghdKS4ZUgxq+iHKbsU3EdsfObO/HBqQVU8T
5fk3C49UGEpwEx78bidAmXGEOJHFALgrSTRRFlWiKtux/BjZPNAIZUAvN5ftgJDf
mYvwBhm2HNGwfT2GGQpmTvhONfHoYVDsg9spwJHfSwVds7GPx5PJ1RSLyQY1O6Ih
`protect END_PROTECTED
