`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T1voLQZP+PCIlierX6DMqvCU/I5LaQbSm0V3qODOoPv4jRGvSR8PaEGBYjnSmgZr
UfPebaQaG00YKRG0FIyV98xHajUWLTXCn/Qa2oOHu1BVl4f6KZSxlN2sPvdDu/NH
Suksf8VLfJ4UksMckqZl4fY7TuM+8fGJwVABuNUgGogDt66gJ4L2OJmq15XVYecl
wL3indwJZ97+HFl3ZuiIqDOGXHPe/eGfS7hqTHMQbZR+RQjJ2j60F4q9qgNJgX4l
DmUSsi4Ea8D4OI0QB86wd1/1rAEPt3hgHqG9RNkpIQuOhYmtsuR7kM3dfUnkxfdj
uRVLpPoLP2eBCRoiXZp8gmqSa92ntbOJLILNmsSLVa+oIRkBchrhZW6R9SLN57Ds
xlQa8EvK6B3CNWeO8Iquz2b824A4O6UgsKdsCkrx6xcdJk6uuTObJIen3125PGiw
UO9mX3T3h0H0pue2bGLmfXIVLxqsfOVAtOOMs//BY1kJa8sKaRHeDgRM1zSv313Z
qeU0qQ4E9wW2EO+ZmkV8aXQMYqnAQDrW0X8nah3qmlVPrSl8PRXZOsHA3JZ0EyVO
coHwY1vnyMiZ12igmR6hKTvTzKy2w6+IRM9ET0P6QORZm2xQXHJ5vKh6ponaD5VT
XR09CUA16dtCU2SIE+U09A==
`protect END_PROTECTED
