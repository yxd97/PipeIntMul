`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUgSM8U9iuNoTCHdTmFwRO/SR0XgUEsmDg2mv0JDnPyNTOi17KOA3PbJ2f1y407V
mf2AsFFj3ONZLzupwvJOBO4Luz6Ff4eVMmzVjSOhmftaDXHt9hh8zlZuh++/Xrv+
D9y61G+eqP+eh7vp7UZzzABBTM6+QCDICO0v5Ib+ccyQs394ssvFRkONLe9VmJGZ
lEPif0Kb/i853P+HoOqqLZbdP5lyUFeaTN7raInNnFU70XfMEdMpzP8hXsg9SIs6
Y3xUkiO4fEEA66inVTowcfvMXc1O4FOKXEOojVFSwMgfSbcP9u6EwrUghNUkCipA
ITzM1TYdK/NMhELwx0mwwXXCp/Z4KeiK0rfYlKlYdwsWgb6qMRQd451wr6YivfRV
cSZXooRsVHn44tFXLyjCdAduzwsXijXi6jd9CYtIzyQTyUJpV/hufr7h542VfKvt
IiJmhf45Q7vBllReeHDYij3N+nwDwntTx/FWIhK4iMpgdzhmenSLmCsCfgyHlWEr
/I+/xsfSTyEC45/ApfuAa1DRl0jQEseXCEqa6AbPUIL4tfAzRqJpmz5lWjP4wRhv
KiCNYHBAhJJwKwJSZKcPdtIXDU5ytEI/nBWuTvKBKQKPQr1C8DXI/v8O8vN60Wns
cP0VuopCrqHpuCb7apo1tFG00/hPz+PZkc3qIinbLxC3T2uYzdI3h+dIccaAV3ZI
ry+Rj7stHNeDIMIdhW+gk5uWDLQ2n1DQ9+q4PgAb8u/9ngfRuPNxdRpno4o7O+8w
OM/eVfNh/N13DrEJx9PF/53KNAkrtKMRBU1fuTKorKEMQDo7KCg9gdCCBPmI7SED
w/NXPHJajYjLXvhzRG22S4m4hprXMbyilCEUmEkctvQcMsXnDE2AkRf8dcEGIDo+
IL5Qh5wE9cs0yzWlQFYfiZDVrqkuF/CM9/1xnXj2XIKBiFhEIq2nbpB/0GzH1gjb
o3fdFEsVXX7f684qGfGF++8exVzJ4giODJTjL2Vn/PUmzPVQc4J2uEpdchZLrN7Q
qsF11pUXdU5PQTHzlGqVM+zMYTHlnP9n2w/NJ75C/9owXROZ21WkkifDv1HTNejJ
NLNpkh3R8CE2iWAoikfJ16Oje/YbDuzzp4Aalyv5cQLIUhCPIIG3qTwg0qTjSuL9
NS4zk2nd5A/EuNalKOb6wmY8tKl6WPANnWXdnirbLDE7mMW0+cu1In6hwe2kkeQ/
g+kR1SeN2dhP7KPazQV5YnIaER5yP58Tm/7V94cP7hnB0Pv8AX9ohELgenUZBs3b
9nSv7KJsIm+krupeqUZetrjILJhTK/H1hA/XSGsD1xaDTbKnoN1K4CZAgRgVo79E
u2efkhH5zWRRnXNdY0b2VPldw5VP6KIEL7RSctmRK9S/beKyFOXlBgzkaj5AZjVC
Zfe2p0gby1vp39hM3Dk8wWVSl5IMvGbD1NvkeTJOLCFCiH7N/nfyMfzdT8Zur1V/
LzDqcrVsY2S06fb42SVWE8xKQE6lUlp7YaHgeTVbOyzelBdqwIWpvTQHXgf0ODqN
ZeVPzE+egsGKidYGiwWztAHicCc2pkWuterUtGJz0Tw3CCXiWsGs06gPn/11MJW6
GwLmNO93V8zcTR0SiPQWIy+tQuOchoAK0S4MRK0AXciQLZ2FsCnye3zFVwEfO4Oi
ZEfz68ubigGn2SkHOAAPQY/orXSNlmemez0Up8R3+VxBHYC2HzLHyfXNHDtodcB0
Co/3JQwV4/B6cm8tkLqz5+ZV8WsYPkJ0m5lWC/VfGJd3gwBSjZtTk8wLsX6fh2fF
MSaBloatr134PvQitYTlpRo5wJTPyB8NXhdGKQcIFTa2ewYxUB1qq28Bue/dHS7z
ZzDYrvEALRxNqrxBj9nIliGkd8EObkxcnTJ7OGm9P5I69tXVWrZS54dqD6d+bl0M
P88P60K1LIy1ElqcGnK6teONtLOcgIyCExSw2X6Kx65j7MrottqhM3BYlEw8KMYP
ZQsnjP0+kd6DSk/Zgbtic6sIa3esHpxxGYZm+NPCMt2mWhPhEJnP+kqr1lThwkTy
hi3mtlglo5mYY9OZabLbQQI5aqoxTZ35Y4p2WxYUlSkhPl4VF6D7NmblUB2rhuwc
t+hPSsbuRpfMIG/UwcKEA9mPVhEKsX3GbsdVZyPOFG824aFv1wrN3f78hbnGDcVe
xoZW0BaYIW9r17fpZjI1FwME1XHhrO7J+OgwcACTOSU+OZJDoL6yYpihzGVlNjIJ
chWxxrApCg+R11SMl4QsAL2sYa18dpDU1F8vWWBpIVQeCBDZnbnrvzNIpfPbyWwa
hTevOmSeMxfosCCwixHXzGGuM65KubbfVptmhgyQ8JaVCiqNjimVz2e53LyzXTKy
hOnaFwFFP7nSC1abgXmIEyVlya4QmnVXOG1cNg6ncSLdzbtC6egeJMT/XWhk9Z0h
wpG0n7eM9c7+DA8YKPjktfT6sbjZPi/X4MUJe7K/q9F4ysPCRkbxPFMV9C1yLDRv
LYA+sbMWdHq17LTW/56pZVLL3W2Uf25BLdIkN2+I0OIQDE1IYL6YHHYztJymlhkV
QX652RG4lC6zOdLYNV5SNCzWkSmsBFqVvmd8bbrmY2nx+kISJTQTevTz2IVwAx9/
63SeAD6EUP7MZb6Oepn8eP0htc3bxgp8t23xkobnXkXsd6bkAwo/SNQutP5T1T6P
EsB77xeB+eZQlb1G9NBMZzoFXx1qR15r8rmPE4rZzht6sgvJ0ckKNWjVyQgD2KxB
1lFUyQFw61Q43Sb1zHzt1hIim8MCz6TcpL5VMIe8zpm49buK5FTdWNAWUnD8qmqq
NKTTS0I6q85OsFZdN74t49/ET0WMrxbeGc1GQ2xbygQqPLBoWNO2SmdbpFFLlX6n
2WV74vAGE6z3E6cB+b5Qjz0v2Q9oG0Ht9zac+yZFnZs9dBDy3BBK+6AK/iQCo+zT
0Us5GNliw14Ow/H5yzPlWK2wLZUi3BxGr+Tss1yMey8xHrw6S+1AnBF5qtqyDQzd
OvYOLpl24dRV+d2BO6fsQJVPMvZ/5OIBKAs0PvMMEkq+53H4LsyWiR+68UztQ1ay
2pIIa+5KMVD7E/+48MZ8ShUlydgIUle3sRyeoGnd6EKQ4XN8HHRjz/EiVbOgCAbX
W3m0q/2PSMz0rOOj8Up/y1FinCxFtZHjh6DT1kDYvjvl3U9nu7ox6Ztz0Y6s8gp1
546eKot6In9+tXpOckSwUHAg25zNjCj2N8Z9c9Ieiw2B1FtxS8XCO0+ZFjTc74lB
AtD64fSwNOvuKXQkLhvcUeK7UdoRde5nzpMEFBmhICaVHZVhXE2XwFyKQ45Qu54S
D/b5ee5TnOxCV/pd2mnHbiYkSBJ2u4hnA4QfwDnjfNIZxUiAEfC2j/hiJXu+N/Ia
7f9B46OUjVySgvfeMKznj2JrQ8Wvx/Hn0dXRFwamMa74HDpzoEsOH6knDu4SxnZL
mj/0rlDY0q2ZAh8hyw8FGRZNfNWiq5Vitn/GMSUkj60Bg8bsY9pgmGi5eowCK0i/
CkoInyxyuICG51jvhJj5mSFDzIlEkU6oxzpljpIIPkim9HZfRjYauuoU6kXXjagM
fGPsP/sjyymC8ZL4xp9SgyEgcFHr5Nj9WG0bRyIMZKLZx1vm3zxXwxiBo1lQOg92
`protect END_PROTECTED
