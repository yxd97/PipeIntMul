`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YtLOw2WuLBLGwpHVZ02++TKbmCgy7j4I5dSaCUoJkXWtXObjJUf/M5VJNorHc8ti
/2Py+W6j/wWsvGg2j400y99HBtmo3ZAOvSvLrXVY6OhlZ1Pz3Sh6ErCiSguZJuSA
yiXEPe4DbjgyOti6SLDHNesikM96qiH380lOQHMbO7JOVQELCCB5vrGxr6bnPgr0
RHLmzNmlQHL0c7fOmuPbvcwx68IR3PqTn9xFFYLs2gyoOIv225ZFFHfPQQrQvNhq
qMH0J6B/JGuR5e75bvMPfRvdNh6ppFd+4ttUhLGafPQPZNeP6iFhDjUrVNhOvs+2
MKDhE9JKAME65S/ivB7FsA==
`protect END_PROTECTED
