`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zOmCk8nkX6DSRtCvlFlQzn5200uixIt5gbgz5f2bdu+SOCJA6U6YcWFoTIjjsUjq
Z1y0aCuQ5XiAez0Mj4tYyXaUid10re5BF7OkWmUo5TPML463QQxy0SI5EhlXe/TP
4pBnhDJnuzpx/ohCL8Fy5a5tP7WkFKS9KmVLIALKVYgGzw1mG70kPrdC/pU/jpOk
SGVb0yRQbVkA+6hVA5XXqNDvVpxvahymXZpgnDvi689NqAtKyuk3Mq+FuSlWWo7S
h4pY7oGI8VbFCbYxH4aCeF42ra4Sgok6uBiaRZploETy6pMXee/B8ICoPedF1wM2
E8Sp7wpAjMP7CM2tviKDXm9khavkfjFaOdOC4EppItuom8MzgQOv6aScSfcczj9d
NVdVTf1ks/0Gv5zldwG9nqdJlSFJrRvMt+5Iv6XuN0oXEQtuCepe48yH04dj6WOJ
iToc8n3qWC3d4x9WpiTE1pdist88m7oq9xRYze769XPmPu90rclFJTSTvNnf7Qpd
f3roZRmFEy8VCQ3WvyJQDOswcJXJA8319k7h2DXpxSew/qKdAn/2pShTYPr152sh
+Mz34WuKABXW1fuAIigDFDRXhjpvwRQUp3DXcCTNlDkNQgVJOhPgztrrq2pScpp+
CsC/ptB7GZ9LACUK4n8fNW//8pe9kbm23zFSem6avTZJTpuo0JMQpMkt62FB6vzz
iSBVmt2BDtUfbt7opUg4M9+278wgMILqcrw3hSo/9oApf+/PZo0fMjP6FYR3h6B9
s4Y15U2jMPCmND97QCqryw==
`protect END_PROTECTED
