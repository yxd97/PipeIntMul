`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CszxKK0N/jpv8Y4huM5XV5iwn4RNtDiVhlZi1GSTXCFkVa+7AVwVmOMqCc6tXiUW
F+H8KI7v7RUbkOfo7uEAwSWRFiPvJUstKthq2rCHgW2s9oU4AoPv3Gz65Rv8gp2h
HRV1k5ZJWJ4LNh/e7YFMI4rHa6Gn8TWEhPSslFwN/wWDSFe86aEyJU8OjlTjI4ul
Babxv7OFrfLOKVF4heLJoquxZ0byEnbOQ9/SmWCFcDuLMR73vhqo2QyT5wNyzRcy
d8jLW7mLDQ8ItRDlcrrOCoZ/XAJAxxoBhgE/w+MGTYyJawKxxnlE+gfbfwitiNGH
ClX0aw5ZITsMQAnKD4RgwQkp02EJ7s83MjU/G7HfZ00QBdlV7sacx4/4aB3GOFlU
776hnPgrugb8FIUbMW/mp0RkL3jdGXCP5elm8Y/2HtK2Qx4JOPPgm6bpYEiwNC3a
V028PNEAnDvexDlwnWaopJG6zRR2NJBcDvTCNOVDygPR6C3H006yHGJ+jrQd855z
2oSZtng6guY2iUVOIXaJ1hhDJtSwWoPLrlTbyreKr7eX1XuL7gFufamgkdPg969R
+rl4B+9gb6rRPNWiFjsRCLF4NPvRIu0NRs8zY1jRd8GBoCA3jzA3i+6wNw27kces
vUbo1cl8KXnqvLHr09FX3dYaTiTcfPx1jxOmP8soTx3QqVBszRqqQxTTOC7LhA1A
44/Eol1CPp5PCSF/6nmwJDZuVoF12WGQLjtj+6oTnbY=
`protect END_PROTECTED
