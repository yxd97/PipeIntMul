`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A53M2N6uvQd7A5DVi8vrnHfRimnaI2uiabk3W6Vip0OGnQPgPjBmy5826IJwHQNr
uOz7FQ9Kk9Ri0npiWZ9WEuPXj31UCRP/Ypu+nO7Hvs2/SuPku0ym8XoOv9AjWobX
20lwOE8bmVeA+I/ByhgiLVbPNJiP5zm3Cp+3adxZIpjSOMDAUc68qYqK2f2LeA5T
WtLx+O5sY8CLMgMbqHYjH4xIj3Q3G/hKlWz7XwfVmXwbeV1711STxFDYAckXLz0V
+MjyBnQFvptNOzL/dfGWDvn3oZC04gmqp/dhlpGD+8gDGLwwaCX7Uh0MtfUMHRrR
eVxPIxoWTT3sLkaNrGvN6t1U5U0I9jmCiGcYDk/0HEL4O/SMvP0P/coya6GHYa6Q
Gd3XX/LD+LpK9oNHyzMnWYVswkE1yY0iOZcR3Xub1NEIBBf/P66quqZTT8ym+nK/
AMgXc7ku7CQCIJcznhYejpzPW7ifGLmTtc9SjUX5vx8OEtR1ZIDbtaorWs96Xzg9
w1wYwGmc1RWfo71ElypsVZ+UzcEbJzFDv4IgxblDKXUrYY5lRsUyDxGOyVEeAD+0
`protect END_PROTECTED
