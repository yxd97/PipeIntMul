`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/VJAO9WG60uZJnoa2rY9ZsAW45NjpSmQ2tGvdWVC4YPvK5+gN4F6zhD789RvNzD/
Gjdd+OGRGCyl4B7inxvlEwlqn+bUWExi+C8JmYAZ9WYpuR9M7xDBBB80KlzFjG9k
3IP+aQnbLTw+YbDNNygU82Rm5raEIb7f7uFxsAvtHLTr9kqiHtiAMBRUjdRI70Tx
pLVkQsQPAfOALI9ay/3gbgpEcTYu+2dsPGlp+6N6OlMv3ya03xJQkfga7a8CCCEu
MrESQiQKTr1t1vImqsQwFjp5pz87ZhDVAvsWRsMSXZhUfKzTLfu9jJijU6zwjcUV
9wmZPaUdH/YQmhacATAOvA==
`protect END_PROTECTED
