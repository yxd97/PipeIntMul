`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RtV8DAoNak2e7FDYv1kK+7MiPO0o5+kixs7Cchwe6G2cxmzUgQhrq2FwgrxJONcy
TbDHEksxn6O46TMkFSdvLXIk6DvltBbE2DUbzSoCEkfr/RsMN9UANvXwtHPoD3Jx
qNdt4r5jcKsfdHsAe4FeVEHEDxOTe5Gk/0omSBTwBCMa7lzWkwm5elolUi0eQhQI
i+J1pNaiSw3xzqOR/05xP9FpiPlmbbD7PS0vdSYulG4C5ubOvK9K7AJ7JhLFGFV5
HCpxNxaeqOYIXLhtwzhKdMpMnvmsgEUqiavs6cBjuwIrsuaX62Ow/WzrUcC+W+zx
4lPxDDmVyOnYvwXOW3z35yk+QEpcQeL0eOZi/d1Zwe4FWy2vHPLdlZ8CnBzGlDJ6
YLudM/6s0z9B2qDFRMP3u8JFYz+e+GthAxpmX3s0od6tauIwM+qgZ9+uTtxnaXuD
WVbiaUVawwFVba9juTnMl2sGeCYQ9eMhKHC1rFdEuzc=
`protect END_PROTECTED
