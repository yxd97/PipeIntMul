`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ogl+6jpZX9zDdAlDY6ZiWQHD1fKqpTrdDte5jg5wN4phoYzQZHANcmKdsqm1Pbsd
me8bZnln3ksoWf9f/tX74JCLDEKTYpBycdjQOHE6lR9ppPsBQYzVcBV0W883such
aMSqFQSB6Ua7F0vMSFDe59GVVJIoxFeL8+sehX6Aoge/LqHZSMhqcKo1yo9wta8g
CqclnoYSj/k0SgENHyVqZ2aKa1PM81X3EwLRZQsmTAfzklrruqUrEKRILc4jxSWa
Mkq/5DcvLvN9ZGHKaPXddlAy1k56hudhDBjCclPMwteG7lv0bLzL5DU9mGgn3Zqg
qyA7zOxaO9j0m2SzkRRuLuTFGLkqtUtzEsSFyyDIrmdv9ig+h2Q/QXntHAKU6YfJ
I04S61eTbKdyJ/yky/k/MDSGbFsKtHLxwGBQgI/dMVbcIVwh18VSBXlgcSpTqmXN
g4bPS0IKA9Oy+tEBDXBTpI1NBOZZ/KKS5C5wGWw/p6zmDEBmUjyQuE5NmeKldlk0
5Gh9n6n6qU4RSs9RaiqgPBJqji3+xIWhvcSVo61G7XR0+cnKmbPjqYcQENZq4CC5
QvTAhSHCqFS1/5Cap+VnwYxjOivgjVHVFqD8kb3SH9ISJseAlXh9RguE3nII4Hcb
XyExMPboTyif/VR4L7Au0MYD7uQVOI1hZ49yLP27daM8j0gsRiDLjmy6Nh7xB9r8
k4VFxyXmyzrRVrQBOmUff7s7C/WDn1TEX9zEHVz4uzyH+YVFN8fNLuNkBeoK/IiO
NRqqc5wsRbLP83wI3vGtJHwGdWOhfv9AWhxTGcBoGRScZosz2JPtP4nk0co3OHNb
tKg/4M1q1pwSjkuK+znb41IMpmo53Yq/BxJax/X//cwo6Sn2y4AE0GSQbxdGLXww
7uW3K6dm1fK0BWKYf+IqIg==
`protect END_PROTECTED
