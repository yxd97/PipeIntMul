`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LO1cTj9+TSUGJoKjjUlTiFz46ZnQ4vyJYDXQFVKXnfx/Rz/UmOSJN2TXc/GE9PH5
A+B8/xOPbspM+IxcxkXQgoL/8sB0j2WYlmgRAlKybRmm8RkfHO5vMZaog4ce6WZ+
STr30RP2nye9V3ZXsxyZRXtlIAISuKje5faqcwU00FytXnvea1hSIVeHZ7bz/dnj
Ga5dJWQCwTR2sFf79RsSUXQWiUEUAegE/rT1XGUyGsMZ6uCusHhD0pIV3b9fa/o7
m0+AjiJZJFehjpWG2SgVs4sPmsDMaL3eDsyMPvUz09YnvZZqyM9fQVLs4k/VBfN0
IAHZP6DXiCyq7sHOyOFOwvimrYHqIM/2pcvbinni+5Q=
`protect END_PROTECTED
