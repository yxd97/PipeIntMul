`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4NR0YRLsL5I5vqjZ79HUP8AfaVhWRs3zwV7KLz0p+sxOvMS4EyKup3YJXx5GdksQ
g4vzEUVJsPShdbjUKhVxjInwEKVbZ2D40DLNxfYYQ92YEPMnMiXiDkdy4ELewHcc
CxhU9bB1XmtKTahUnqWMot0RIWKxfSN3XoMZIoChRYbriUtNhkf8vUFsX+wPBFDd
9rpq0VEvFZThGExyN4g0XyJSxFxB7wlF8h2cTua/W8NmcbIkVg2PVCAzuwqGFjJ5
wFmYP4CRe8jv4fFHXO8c56JkQVWqbySGB/9kWgnssX0re5lwAJpJgRDvmipJcmGo
nbygFlnE7T9JbFUJYHj3qjtUvSYaQZ4LQIVGoQOk2aG4BCvslskWca59JqGS5QuC
MewAR6xf5VAb9X4imT8ZxFA76wAwDZ29Zc8rtci89uoyN8B9M6C3Ky804jp9UXwv
ByrAS3g848YLFlQI+U6nCRnK/IjXc8sOQGaHQupqqt30SuAvH3UndBDSAHJF6G+b
5FBrdRxYvrq0nL7HK+VVbGEaZ/Wld2LJk1z/0qlSwuZbNRNLYE+L/bI1N5bOhMca
R4/mJKHR2/rIDqDJRYQFWIAcDhI2g8J3Q8pFZlew7942U4ZjuWN3qaRM+TSgHlvt
1aHBTIsjq+8auByeT7rnmg==
`protect END_PROTECTED
