`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41P5aIwjav+BoMBxLCR9W6iJmrq1Qgv2UBJnweUvNaMhhl7gywKFPDU9k5/+u6QM
WAKD96YkU9SXtmir8xet9T6DLPrKjJBmt8LZ9l//Iu0PbBbzC5lp1Qhz6fKV77yB
4iP3WBeVWjgRYkKm7it3fwgsNH8gZJ3Wk0M5BOH/lBW4jcCx6WflDkEyp/2QOHYP
MIfrFWIzAvcT8LP92LxiGuSWnUmGL4AhNmQBXU/7T1XGpDcR2AzOc87EI+8vcQ+e
Swt9nZrgAalwFW32lXrF9SXuZdu4+rgsH0urfR3oJ7lGZaqAN5rkwHe8N7P8wjYK
pQpaEKlx5feV1dI8MwKTXjS7aiFwHgfvhmwgGNqRB2imKVAz9VhBnS4OKMY0T2x1
d5PJ1nfB75xI7Suz3cazmApyKPRx7F+mu6QBoSZgbpCzI6nzy0vzj2tztoTZrQdy
XClleL4EmL13UBVUpciUCYVsceTff5EfnyvtRxnqE4QV3D4XxP84C9eGP2yFe31r
`protect END_PROTECTED
