`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5lpMfFPuKb4FFqkFYjN+F33k9aehnpcPT7Sgq6FKNyPTSgoLFfGgyCJMOvhvp8L0
O0inStFoYeAqffaTj6zYUyw/22BFzHJr+KDwve05dL/O8yPBvjnbdA1m/AcuKdRg
qxzvbrym3R1pO47+QWnQvaNh3ChSf6iUQxG5EOzNENxGNqts8j1gsge5xi5Y089C
LiS4swkYIOqL+KinJdznN7GQ7MjBWsSN1l9bJ6+M6e90B1C9DHeC4PgP7rhQr38n
U6qnYy1/vHEUpzXy0d5FDF3B6KIY3lWNJdJyMEX9GJtesbqSPOsF+6EUA/4ZKWRO
N8Kao9+6h/0dh2P0eobD9/ptS3UiwBhQVeGXLEnggnptVn2FwRQKSuLE28bEzB93
7RdML9SdJIKZIhAD0EpNbjEZgQ5YXmvh1ahz5LKWJ4a2xO7guNVmgxgYsX+h0cUC
f912yvtHpjLjFjZQAC3Td/IwZOlJH/fii5duDhCycV46EC6BijwZb/QYv+r7FCT/
StG1gYYdWvZQE2h0DMTGFKzh6vntm0XePizRIQwxKLBpfPXKd0eL0sZUuEPMDtWL
2G8x5BLly7gxGe8b+nIPAeisndfVUxyL5dxon0pFP9NEbDAxzIoW27Hke5vpO4AU
raUakCjX7x8yvEVbGbTFrJxtxWwCBCHltCWhM9XK1B7n5sCAhdI9UJnkZHJk790a
H98BH+fVCQ8tE5R2P8pHahxsao94XWlFEKCqm/GQC0k=
`protect END_PROTECTED
