`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZxeWIrDmeI5BGHtY6Sm2rZSak8La2TWs91dGVmBFUMlZuGCEg/Rcydsre26BQmB
+Sk3tQBVHwh/ftbV7ojoKxrySksEFpk3gdcuq3IloZI4H3vwyS2mcyHg+a1mU+IT
QG+tYDceld76OPiG7z476XBEhREAwQdU3Yiue+dbWtzbpYB71GtwJQr2EqyWFj4T
SaJdrFPX2U9LIdQ4KTlDFzV9zEdNVDDvEkv7xOwSeS5wrum3dkNeGmkSZfhZF2KN
9aCTf5aJgHN2CyZXrg2/veOuowp0hoVns9q6dFD0WbiSK4Uvzg91jyLFKldjvlZW
Ve4nBHy1DgS2Mi8uPW/Nw1C9pAMltc1QlvB6BHCcHLG6rTZIDr133LxbA+Ftsr5/
tOYxjAITognjT4aLVUELmDuMj5g2XuA/2J9tLgYCESiSNMEvPfsKWdCxltTcg39K
2zG+SyL/wR3tcbG7XX1ucZwpmr2CjVoONMC2mKvdusfLDAOdNd+YaN52fwfhrqEY
l2ss8OATnzktWK6vRwmvjaboCvTn2u0wUbpy+lQSxMx5QdVjGNxUCnaIEb4HMMVG
HFzmOx52dCU8yTPJa/YEYFAlGU5OO0PQAE/RNXn3dFVj7EvAKMiiPRDjMAqj6tYu
D26rvlUPDBgXq9d7HUqoRa4XROJRjKR+dlCgRDcyNW5l9qAjhoX+ZnlmI7OuVURg
4isIYPk6pHlVx5Keyy2UNK/xJf0WAxlPcycPtEjyaL/769ncK1p51eLVv7K/Dp5Q
M9xKqRpiZr+QH3g9QvkyLbU4+e6GDRlI+/X68hBEJZ/qNHdlBvqGYOk+FUT58hm+
IwtjKOJGwpoTIKdXBqh97W4rKGvstMCDNjK34rInye30jfQtTffCc46l93ADNR1/
9E18mqy4/SXia80LCQXjDYmdEWpRm8HI2TVpEN+Thm0BwE4w/JmcTTeKi1FR7H5f
TNc7eNcVtQXlfhPA8iwvmdUAwkjYCUizyi3sRRxs9OBI01T6nLn8sVuZUfAACrF5
a0O3exJXLXwnhjo3Rzx1dA3tsX3urCcvwvtzKWOey+QeiCGH7RacBl/4u7UFRJho
lIpTRWvceVcVLahOq1K65aoypByAlxMR7xhhHERSqtY1kBuB6kR+VjjDTiaxL+hp
cGhF3uWHRbsn6RJTpdD6yPGh2MhvuC/B1ohL9pZ3Sj9kIGF422XVBQxiHrpzvvIT
odCXWL5ltjCtP/HiKTb2nSjwtT/6OmrBMlt2IO5pI1JsuDV7xA5FUQBZndJQq1A3
7LZhuOhMT+R89tTc/ou+OhLmUg34bu85yYup2FpbITrNnLQnABoiOEE6JKMN7YSc
ytkSKULqsAUypUE4UwREMsnmrZr0ahP7vAaxhTVayIDrfMjiDHi/zykGUQ0usKyO
3JGIAs3UWUafqBP88qTnC/ZXTY5CYMSxW4xfK9vtzhQ2iKcvbxYCndanq78iW0Lm
ekuldsefOLtsFkJwQF+q3z/bk1iRqPN+iq7ihnP6RuIyqRK39+O0hq3iVbUCCoj2
2dn8MJPvAyRhGFL3xmsKvpOsX1ZTBCKA8fTZVde9yrQi/D8uxdoWnvqU5GcJshll
n0wMmY5PQfBKIygvOm2W6NnkCSgAJkxjhDWqHOd1ijHzU4uKlBYGt5UkLY00SaUu
t9mRdXFsx6DzO7shgoR1j6P6Pw8NjrjKRc53cN4iLAklEzuaiDDX5QtNlye/hxcs
OjRcxCmPSzcrZK1i6Apm0+dWMiGzM/uIDqkdILSSiDB97hgF5y91RfnS9rn1DeiY
Y6NkQkn6idnuxxdFJ/Rt5syDjl3maynMIXolBc+g7ns8CG3/FCZVLlWnMqkJQ2Lc
X+D+Vph+8Mj91wEo0PgHRKiNMV588L57qgZkAIgdVcRKDDryr/W6BZPwETs3MGr6
2zFBToP+z9x5F61SIrnnH8xeTU7w2jFdDUVUQVY9OXnMjo0fCLeYTLoOHkjB8GaE
iV44g+boXD8dJNahzb3zFJXECDCVWnjWF+kqzNP0s+OfCCzQLDHxxB2sBlKjZtIm
VXuzcYlOmDqaDe/TU08GwarH8AMb/CJlUtd2mvTbUwx82LlEapvi70NRcGNSFNFX
1vNe/tfuY1gG+uH2zWvxu4tUvdDBmnSKQpRjhCsyHhv+YSdrR7MrxVWuLf4l16MB
iSVQYBPbfzGDn27dsbC18eerEDocG1Z0s0tljsBadAWaaI+v0MS29nd8LHxG49fX
iA9m9Y+DurqoL5+z166NdBzya0UIIVees0ghyd5Cnq+aYPgT28bYKTAQYds49JiF
m6SqTOdBQFk03InyO3sR9Ko0P39siGOHLTMSnoEtYM3M1CZO/T/kMC7d609p03dl
ScHNXngKocauYouJQZpuVMzg5cdwGdZjtqRR3ihfUu8yLJOfnmOr29hr8GFqwblO
XYCshBzb9C6rUJw4edjinmWYYGruC1NpvSxczxMZVJvNpuF+LPwxQydNTTNOyMm0
evGQiXlzkCI+zI6td9ssmCpf5BP4xNvkZh89LxQGyHs=
`protect END_PROTECTED
