`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ta5kEqnqVaFAi1drc5BKZwyCN/NrNCloiUjAYTHojU0EEr0UwXbeRq38kVMy0xJD
Er8l/Fka0PcV/VG2CfKRt/wmP6AWY+Bk6DL2SgOLfSaGmS2RchXuZleinMH8Wthu
stSTmQaNoXWy6Zy9wYKmpCXqCZWdqZziOwzzMO6AMbYkQhL7sl5h2Uarpko/rND9
PglfbjmFPsm0GJKuaYZRtJZQL1ioxIHCBN2z8P5RBsKyt8dzCMmsXiBXSusuG7WG
+vGzoLXnEhNwashGS00rb0QXb7P1FqwrKDiXujpLHOs3R8SPKEqAs2gAvRiks1E/
mdzzP2AsaCg0+DSptI7ltgdWtKwnzYNzYxNnhQug42P9h2qC6xY7bq9gesReOVoG
zWX+/vvTXWaKekIcOCPpfv1SRVWpiGXPRkDc3wmnTHFZ+9yhJQKb9UKxyyb7/hyO
GzcIg35HSVrfeI+qiWe5KlymufGtBuXv3fgwmH7jajZ0hQtM7f+bXcqmr0ikPKp1
55n85azeBP1P78tuAnh2YK4lApLsa9AQWcotzXpvjFBXXzkELoUOOO5pYBg84rtk
k3fUp2AQ5MZ4Xzd+ph37jvFnrELE2rus59yHUrHvNDZgWOcgOn1aklPLsKKod+4N
TVZPaOzpRu+uHIrQni2fdxCLcd3S5QzD+PkXGlYhaHDFzoom1xpU3B2+7YImN7t3
tsvVvGMEW06UQyG9VG+mvg1avBA3dDh77QT6pLQEEC8qKq9uyG4QRejRBzN/LsUF
bQ3PbdS1f9pPfNfCYoKNJ0hsRVIkCokW2bHps/j4+gFpRZun/t5/Q4HoSDHaB74D
mUTI2fSkVGiXoZ+ZLGK9LgMbItpQ86X7uyT43KRWpc5HsTb1Dz13nlvVBoqXTIEt
jzGhR4JsaUpdfQJMXGxM6svyVcvzRbI5e/4VwWRUVb5qwc4D8dopDOqtVe5E0GrO
Mbo4xkLsN/3hTmax7AtGi8xlvWc58pXsQ3b0Ye7b+OlqCjqVCV/l7bir8qWc2ivM
j0Dq8jRLswaW+nNfYXlDfYp/nCIypreUs8PmXh16D/U=
`protect END_PROTECTED
