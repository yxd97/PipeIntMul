`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hs8Roo3GMCJ4re3x3rvt1Ig/qETI+WxO2aYPvlMGpl/rCMsHloby/YO4uUi/auZu
earzCVZ2yWCKGv9p75Jo97wTagckxEUZj3A/mFmvRtIA8XaGB6ocExEJXX7o7kg4
l3CqbAc2MA7DqdqQ+GgBt0Ax2TYA9PTjQlQqPg4EhlRiGrEWFe3RM9e5rKba9ZDo
ogIWEYKWOBxc0krRE2GDqwb1IlgAfGqIzxzIHPbXOPvh/UPl6Fbjn7kpM6+8dxm/
gIb2HiRaDxpCbepSZETcKh/Jedc/NgcUjIWl0+fnL2yp9c6D5qkKy7F1zXvh13m+
Bq/lh/aaH0F5wrKY/MpmlXEgSZ4d2eETc0pBQ+R3qoGBYvwffNpmYpUcjaQAYDdh
W+YOrnh3giarBLrEF/jiHIVr6T+STpt4LDFfYzLRsl0Nl6OrgCZN0DhuUtlO9EeJ
BI/Xq4hHqngQUpxhQkLaOnit1v72ZaduvVxGtdb8KlWKryBLsCXat5V7cTcaQs/+
+Nwn6bna+NDrcK8NRguh5VsLqyYA8QFTHYKqqNRZ+lPRV9G4m5K/lmEFhk44mY73
2Dxa7wZOsfE/Cn10FmwBTaroBdwpX+z1cLveRmeMDN/0ylZX177+CVyNPWJjPws/
`protect END_PROTECTED
