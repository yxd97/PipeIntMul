`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjJv7rr60aUwpSR6XsoSaYZEm4p2Hmf5Huof1LDFw1qyQlVA8dN4K3MwZ0vreBeq
bATeskbpqFwHKA5Qkzx3MDoJ/zoQ7yHh7yCIvdrjDtJfD+mBFQ2R2pC/FGKjN5lk
S3o75Nznu4bIUcVAp5nRSiDS87FeLUhPGUHZyTH72awc8PoF2bkMxt9Zf8PgdZWG
JFcwq/gXm4DrkWqVnFwkRaqHfd9BAI9iQCp0uNPercDghL39Oe4XHhE2OpmNX/O7
T2max60bzTVd3bXpmsdkuEJQrMEaPPvOOWTrJlOigJXPRq8Mg+uUajAHAOoijHwi
mAzlxxuoAji5fXyyjcXGaqSRmPME3c1PF39U/OPL0qUWYHeO190eQbsLQouC2F5D
SvmaHwRI3dPcnfY4mE5YA0pu11STmUfX+1QKwHAtHQ2wLCujI5rneuEnzL4CIVrs
GA7E2X848qrWxt+8jbwJCsnOHEmnRDSaBBcaYz81EiDJbnusUSxybj5tbD7FDYQQ
3uykHGZxcPPDdw4fVdg1cH+KIusNy+PAPGR5qNPyzYXX23sY3Wqe0tzen2/xBmXO
6t3KX+jEnHwFQ09Ki75urA6hCTvRIcXgZvsH/mUfg+xZ4LYFgJiP88kokd53g2ra
SpaBtpc1RSJWO8Rv6uJl3RxicIpBxMBiHSMVjuaL1c6rU+KFQJyaUa1czGCQJWjp
HvRH5h8SFWUHqymjF3TwZcIHjIcoj9ZyMMnLYSj1sYW1KvsqgReMmwhmUb/+Rvv6
Jg8UfT0ZMw5eU+jpu84Tzq+Vy6fAzsOfSMnVC2Heg+DnA16Vhs9W0aqxqxziXGwY
hPr3QPOSCA+PO30+q0PS3hiEU5+hlwokqndOcWjknrjKLKg9+QrVsp+AchFDtxpj
l2M7Wn6d7H2C/7mFwqquR9mJ3TYfXDce0GOUiSP8Erj1avES5mQkSlFuHmQx1qUz
MYALm87cJ+fCpS6XStw+07acvh0ZJHhYKt3q+gCX3VZgMjS0seO/B7FcYqKTJNra
40sLPVew5rSZGn9wWsJ2sy7Zv68oSCz/xxu1JuoNarJ1MwTCAo2XN0E/7t2GnQiT
u4uISGDGqQZnrcNugSRcSA==
`protect END_PROTECTED
