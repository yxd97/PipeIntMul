`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jH8DpxzOOz+Yk8gcoe8BZGuqysPlJSWBmNG5UnfPVL+1IRC7UIXHRm+pClzrPHAN
mlkHFMIykJS8CswsDchPbE1p7fhw2eLd+yrbrqb+HKJ4zGpPC42KETi7bEHKAxNq
zPDqZztITyQzUiOn20HWS9RsbrDFXMwodoNSsvi+x7u+mY6kJE8DzjXbgLhwzx9e
xJSv2JsiJtaOdQrjfoahJ5b4RQYkxnetJtXluAm0iKSDwKtHoEb5tl81Ll17C9AM
t6fMGckqmI3Qh4PA4sNbybnftB+zGDP3YoM0zOPGL4DZ/WQThqPcw5to+t6PMq2v
`protect END_PROTECTED
