`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3V6iYV1i8Tp+4q7VaQCWdxiV83N0ifmnKGlI7xNPi/FQJnnDBPmbc98qWcGnJOuU
AX68WOElt/zhQfenfeKOPhPbHSHwKGK6sCLSvdDeX4Z8MUW3La8KZvDP6aokBFTV
DJYfYK3mErHPuBCrbTYOAI1Sm9RAxj07sb7fzQXQ4vRXZcGm8eDQgsrrm4DfCZOX
CdO+ewhhDdH6v6DsGfRRKe2npVszKSSDZ1+r41Enuy1gjA33Mt/CfkdWEMaHVa+W
Oe726x7ClqfuYADsjndUPXEev7a4p8Ci4g3iwin5tqmSeDBeBh1/OfmLD03mDiYb
oIydEGwdDlkfSpXyNP2Nkk6MdY1WRma/3SQ6k7bThEso6uPw3mrEwJ6fMb+monAG
lj8ytk85PQnhD6ac7mm938omcH4dgnioq9P+f3Bao/WMZif0mtsPsPvT8hgdJTDE
yHn1AVVqxMqk/lKj5XeMtxuJM7RZmKz7fu8gtwnoKani2W04oimPB8lq14qLBC0F
nndmOCKdFsMp6VRYjeE36UTKlg6/YGOL5nFukXgZxHW+7FlE85Kjw/BJso81budk
rp6dBsU/ehS4Y/FyjhgAE9QqvmzgFNs/lpbgE/x8TLn4c+/3jNH/QgbrOtqGl35E
HZGHej4EkCcH3B0f5pCEN4q+NlML6aza9VTcxJcxd5g8WJID0dj/64uaS2pHKG1E
KlAj0vn8QyCc38mIIQLqzKCPLd/zEzo/Pz4Ssk2wnLR3ooWqa6elXqK+bJPmyNnQ
fMzAnnG9+JkMVLp803CO4POXMJcAx8i0abyFqlprJX1FFDK55cETSBFVM1opbl9t
6j+CGURJnU16UUV3TVn9D5cDRLVOQxznSgo7hztG5UcXNPdgkkRzTJgJq0xhkGOD
rQLlFunURvHHMhg1OFGIu+0X50vUBwyfFVxZpfIp9V8VtWpPo3nm2qQ9kscWrytf
zC9dLuqb+k63QT8SORD/Bb+7tIoSaX2oiu/4rVy/OWEituYaREIoF8gj135fOinr
qo5Q2HTAfqb8irr8LdWuR4nQlsszKbfen0JaUsCZHlxqpQn3mFIi4HYv7pwbELwi
8HUJpwQKcPX8QVCTaMl1mNrdHcNJqQv75s4WcRyM+6t1iu2C5zRnG9Vv4Q7ko5Gj
pBlfg6Bqg4AG2Y9pYoxZtzAbzrmxlSdNkOhj3NzPMXuut2hcmbGxnhbFx9Zls2dL
yD0cAWB56PHl9BJJE3psnsvSF39a8KGXWlcuUwtoJsg=
`protect END_PROTECTED
