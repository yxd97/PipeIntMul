`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0QvfjF3wbUGV3KVdFP4jqY3sRBmRrZWvH9yH9lKC6oD3jHTlEIezNG0SPHeh6C64
F98FYufnHa+4AkcpqCYw4B+WX6naUtSrHDhg47qOTuGbrsBPXeqBl6UMCE+TQbUL
S96yiJPXKIyLpSOE0c2OMfbHw+MTZif+QFQAKUcCdqZD3w4UG5f3ZbiBh9+90GD8
9F3jT/fsjxg//HC9POwIG7Q6SGlufxGRXXQ4UQ09kDKLlEh1zwxqxRYIsX2OOqt/
nIPgwWz7qwPtmKxXlNdiD6SmYf45AWdBX1FzWe0Qvw1d48OHSlplSyw25PdLNhsL
H2yxCgSNwGMOvY2WwUfYEoS+78ksUQniJb3Y7rLlm+pLflXQNDFjSmiP9lAcLFs/
WY8vtUX5yLm9O6zatIom+e1ImzSqgNIUbrEaqEZEn9Hb8NWLfAuleAK/kpDbrj4x
46obW7GZHxOcQow4evarhsiR4lppJuMtRlVBcLgzteQ=
`protect END_PROTECTED
