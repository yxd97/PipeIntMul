`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZekrXiGD2YMccey8RmQP1Ue5oEzZ2l8xRKnyos/Ub1d49CLGkdUYfxAm3FoZwtLP
Cn1aKxHZtK2OYGL0nk30P3ioQUW10OBgYn9FkzP9giw2ksr8RjYilmyDWBam/edn
1Zgucpf8Fyw7hjW8PeKyngnKFqOlNzKduTGfbtTCRFBM+VObMH7CIxyuUWtpqIQZ
Q+o9S2wAAfEjres88cssuNTPb1ChV/aziD+ak89k5eUij+KLJC+iSg/CR2tZSA0F
n4yrW7zf9Xke6iTOpZ8IwwTLGoLKUt2zS2AWCDQuO8pIctMbA6f14wq60eYlyaTd
X3gAuDd+4UBX0bDRXNfohuGetINZCHpqG8qRRSoTKADtbuWajF+7Zou5imxyAjZk
SUepGDunOUag6Es75JvwtRFJqd9ohnJgVlC77kpfI944ahHxV9lVGQCEYjfqWStZ
UgLZp/j8IHvYRy+I6wvWagoQrTD6VP36Le50S7Whj15kBG3FkXJkP5pIHIwjGO/p
9cLuBmiQk3U1LXlLWuRctTBvAzUq/ifS8vBSsbaRe2+X4VA2eyuQ7qiGPzcjD0ec
k/VO0CxwWh5qhg0l7sNCDMBODNlNiLkVqrLvQ3B+pWnDcXO9lVZp3AEJTDFoTDOM
3FotaooYUtDTu6daW8ASGhTaGoO+U2ycuX5uKhOb87dK9nG4Jb9yYjUXiSIx44Xz
+UhOazyy/23qKenkBHCP+TE0EOBiBPgg8HK1CjtDDofM4gJO3R7p3mAVTTUvdD9y
DtSvNksX24gsKDLWsIgv9rMppbnGIaRtMmcNL6fDZYFBR+DqZl2/H4HG3F4xpPfX
OV7Vaq4O45Gg+X9SRrTlKh803jqJZRSo/LdS8PZb46xLSFdtwFS70V4gRnrU/YPA
cx3xGLXHKdv/8lNVQd/bX9vQwL3qrprzGBTPmfR+UCG6DDMWttsAFrCWzwVkIT3y
O/3DKTNg2rKaExHWC9vy/tCsP/RCvd8Hw2PEBalSBbbN8x0/yaFACDJ7lYuMXjsw
AFVe1x3/GVqQ6+c2JmuJciL2utFgbO4TJwZdMP98rHZjpBsilQa6R/ksgTPksgU5
55TVPfUzCH49+goPmsQMGg4wScwJuHj2+Uk7fccvFD6bvbaNTfumo+oINc8UHEHf
zh2dCEPAVviEv3r2bkVl9RILzcn4eD+plLxzQ5MBKuxqq8kpVUg/jGuNQguHz0HO
FkvSUFyox/xmgtZymPBPuhjVla3s4dazTfTFm46MGN5LMj2cfHi0XJ4KwgqOJe7L
ScWLydsqT1SJ/t1GGUXQ0CYsjDIiDsLGbGzE6CUm0MlyIghMvgwsakJVydDxoqfC
5ZChVXnSGWZD4yIc0FruP+AUc3lakOqx9nXkLEbb2tuXf+2WbozpXVA5Q2oCSQ9n
vwdlErowo6FczvNfITjumXPkgSvaNkx8cCjto9x/r8pygcVyhKADxeILfNUU9rhd
HkVao9PIq0xTQvyiJZpxxU5mIZbT2e+FuFi1hZmy4skv8L1KZRM4LxVF+5aYzY2J
e5YBZawMpIhpNrIpO5qiBmJPbtbOWf8Dps0hyuwSIleISDOOs012nCoptK4mgcy8
CWId5Z2ZDlQfrb6G1LZokpBJndIIcCBR6gfS9GBcBkLLZQEyRZiZXPpBFkhkny6E
kU9XFBd17MlxSJILg6EjZTEvLoH3/+eooeqqUjesi8Em8+X7pajLz+5jzETDxbW/
E9QfN/unJ9EAxv7XzeWi3NHtTWtFLH46fZrI/En1yoSpI+4eJY+Are02+8qW58kt
SDPA94n2/gnM5cKH8pxWByTNUMMwKeeFXu9f3WtWVuqRiG2XrllmFnyBUjrVMt4x
dPQ9M1eA7ys9BpNhNVBHlTWKIZaES1vq5bFc8ngrxDQMo9JxR5/11V3YLsJOXxTZ
S7Kzgumhy/gTaM//9f9rgyBEuP9ytJvkkuIYQTbQNAoLpB1mhBgCeK5mTTnY159U
Xvz8T0XLXXfzne3DEYMrFoz3PH0NoWraI+SX4z9zKzr7vRLFVsBpdkuGZTrZj2Np
LeaenFFlrkm4nIv72oMNETdF/3sJcQb/HEJIhURI1+6MeH9tYfYr164wyBSj0pdo
wg0HAbW0hMvXeAmtpajW/i6MIQ5Uj/E540aWl8jDMAGRQmvDHHBoFkagXBYWJysE
Ehm9/WelDV7I2Bh8pFFpBKUPMfjE4uRKDl3oYWq/UAOkaU+SOCQJLcp+0LY8Zlsz
TFp9EQH3i6nj9KS6qcTqV+duOQYceIRbzgxr4LEhD+Q9t6KDaRJmb/fTKl6Wm+kA
PnNkEoFEaWdaPMNRWgukJ8ajLMTjV/WEXyVoj2MW8LthVaA0MZ/dUfM00pk8UE9T
q23iTiz8i+oYn8s7JaZMzNYITKQLi1dwpVzJqzhUIUI2lgKJf3aVBbkT7xt8MomA
/7aJO1XDNtZL3Emu1ho+HLdl31hLOc5jT/b1rQzJl3b5xKCppO2Kz1ZWX38y07un
AZTP6gedNz5dFn/Gy5D8SGu8Muj14lvozPr2Xgfpr8UDCXU2jTBh+DaatgD1WeH5
zvIuBY+R3bpxbI7xrsxhJxSoJR5KOPHDtIYE8nTCRZTbTjAA0rJyeIbfzXmcWt/9
UqfJPxMiAexiZgenyLwoxw8KpCvpAweB54Ou0s4k8DOEbb5m8aCj81OhqK91SVoP
1rC/STxgEbWveEOk2d2KaC1mqWrV/yOU+ParChJIMFTBac6VazDyuCXJXvdkiwJZ
hkHqjkEPdPHsbC2TqTyisCZf3QE/U3MZwrx0gC6yH2QJIxdhJzfvwrlX6SFFKSDH
TWRDbYESXqI0lhx+jZFA+ZSph+fyNg+YLQm7MlaH32Eu/WNrbdUYkSvm64FB/9OT
lfVDA9tpq27Sk/9uzU+zsl05XjzBpGOGOtmiq/zg+UWtK5KXsi/3klh7K4UrTCm8
1pPNHGXjJu0LGiSd4HsCXilFjDsSWfewwSY4gzXKLYraflj883PfihPcUWV2fmdG
m8I9cOcYj+xE9b9dpQnD6rpzASePMULFpG7pU8C4LKFHZF9BmVLl6R8NwrYdCIRa
lbR3uKJWK7zFJqjWWQuj+wvN6F+B6OcVSe6GSh+ZKuev3twi9Eky0Oz6SRVzM75V
k6At3+OlRA7fKiWCEPg46qiSUGadleYXQAVO+bjZEtK4QVZpT6XyEwLJ/96kUzj7
jXkvLuDebMk2r09MDTOz6+IuGv4kFk3pdvaJm4wy7mzAZhxRIL+eFZZgCMKIhyDI
e6lMJ/ZU3W4D2iV8UuB7TwRBC1lU38y0GjQnWsJPb4RpLVuS1TFv5+wqW0PhjcbA
9Wmrwu4SLFDEpOXOBESuJkm17ppPzk8xdj6BPY+eULAfJtWwP5aAAiXdUSlsJR9z
BXF3ZKkOhmwG/CHydlVE0NC5YY65fub8+VNnMltXmuMPgCkgehNFdonv5v8awePB
J/HmY2uwiRK8xvB9QWU8HIHq3X3oi6I/ZHwSPl9uLNtn3zo2ac/T6q31+evqvn7b
j28k7TrAen9hkMG+vFKpyNRdA2pL6Bq/r3jeq042ynqEPZqLQqZFGBD9A0WmLhBu
nqjA+BC9MlHoyyyQgTfLHQtSLKdWZ3mTOXrnlljM5s2Oiys/R3llXAcGdgdzSzfH
NQebd7OW8JjsXB7XazHqYlFNMKTNiCpbR7OxfeuBBH2c20FLgqEVMZJdx24rVbse
ZyuuI3ZfvN8WIEFdklmV1y6bHh7SSBnuXobf/Nfg745reRWoBByDXocQQnrXQrI6
pBy0XlzCk+a8xXce0g1FF0Y4uSiRXhhq2RuBOpWGqoChxKIMxGDlDgiu9clpnH7y
xlW9fxDaHo/UHJbg3reP8r1LwShjkXNPbIOGAldXBDRkTAB6Ec0n3oOZuS+yTXkk
VP/bNrl7sbGlr0Ua6pywfJVa2CLo35th6ho/6cPjXsHyuixebfk5C9q3GBVpmA3M
yAel/BGxfpEMKsiomj5tCI4Qfo1pqgaQIs55FIf4wcxz0BnT2w9s8Uh0Rxu9QD2O
YP5UJpX2ivwdFGasVmqgbhonFOYYJazj/vTPOEzZrGiCCzb1nVY3NbC4pU7LwgLC
m9h7TgA3Fpw322WmQx/tl+iU6rdHzqMGHwZKaxCgnHraNU56De3LIOhMDpllx4Z5
hZujqI0TixW66JaB+sAmLsOelXx8RGgoQsrJvatTZNLHVc5/yTsTPt1YNu2znbLo
xHlORaGL69vYhv8+rGfSWuC3VIRiEIgrlx9qMSf8doarm2GCDcuH9DPCxcqaYJ3w
gCY0Kp1DQtZIwllZjYtsOPIy/Og8WoSnJN/xGs013xzv7ZSUYG/SbuByz2WeKtDU
vCBF6vi+6lXi0pAlCiVwBBRj2F4mrfmMii9TgMBmyQdToMMrxWoW6CkkP4iA5xBw
ZQ0Y0knPqXkFIpatJHfvClhi/85ClwC3L0Ltxn4KdA9N4f7M1ORnQYDowDyroTtO
8eyNmgro9Gf9i3vhfEz9zEpTwVHibaRgpAdAE1H45Ky6fm5bmPhkMW5jZ4E212+K
SlgGg2pcMVn5PNf8yJZqsE5KtJ94N6LpTj9Hg0lkacQbRtl3GrZDnY7ADWmeZG97
YdNim2u6cpSpWyhxpm0Uh6TlgCQAzwyTr26zNI51HT9kg6/FWPOhwKUnBXy3oEmB
XoW5GuVsGPRuiIJ4ptRiLy0dKHh6Lga81zI6bg07mRbSsOhOxRyVHJJ3QBcnUf5M
sC2eEw3LdjIS6Wi5E/jahSSnNKxkYFIKNkvVP+LgZvIzTZ4aLUbiIiYRgxiWOTtE
LBEo2qIadC/zJQMXLEsScDfqLwZCwmjPd2KgKztBEu4m5TQjeueNxrYK9xpwsr4s
yW42lZlpORu3Ddu78W7K62UpewbLlsJ+nguzbkVA4MfJH2KSc4P+OdeGSNL4LM+9
nzIienly5fQCAOvWck5FwUc1XuLgEJUZOQllIDbpbPOMEwBdqyfxp8gU7EjDbVsV
Itr748uCYUfr6o9nKCQyTBSjBb2tnSD0fEJMDFvCcZK/Jyq/xY+V2pQS6Obuqsbv
kTGM64k7bNd9oYTz/sse/1Vj8vRtiFjoQaRPn+BALkzeiMkon9RxeKEitbfFlpi+
XfYnEb/PhtYNuMFLFjQxyPEVprTmJG0pCUaNdxa4M+NpAoa7ekKxt+wrNtITt+jx
uqckQtnufBZPZFcsrDSKE01yysHZ6UcxBPelXjUaM13K8jLrp3lCOUx7pIQnPk3w
SGKK5w+XMbSrLWwVU8BoXxlgntTVRnUhNsvhTmNurX0Kq8R/Xp3Ravmhv3LXSeQ0
3kttVu86KY0iTNlz8iGz143yRj4jRAQUgS2Xoe+G9xMOKaolFK6GOdOPxBCWXsF+
7vcAmE4gyYZi8XsGIKERmC562TStdouNRx/uu+hOgGjoMBL77XS1qOY89YJDEg5s
DKSzuTyIaC1bOPeUwxF2qgb/HwZZC5Y4EPE55EMr5z8q8RsuJDT1XRnswK8dK2Fj
LU3whI0Tdu4HZ2ZJVVh1xTAcKZI6L5oZtD9kovF+Wwiz6J8TE7MEB00GXi6dK+1j
tkwi7fquvR7g7kooBjZBc3/HOqVJTNXIY//vmgoWhOqbRZymE12Hg79WlC8BP6XB
a8XrC0d3Lw6LtfBmTE4Sr07B86yPrhgz5h5eGJQYnbS6FcKNE39a24CS8p4xubOc
Yy3nk4whoh8C2gy/e6OgadDQ3ZiX3/BA7PzVL9NOK1pxAw6/h+YP2tkLkvLtiGsx
VRpILE8bWP+FUeeV8318LyFIefMSruiaA0Dt6aJFccItofZ4gHC0iY3dJtNnwA9B
fTZAa0N+xnmtRwDskjs2oB3PV6EX6NT5rMfHeN7HDreQA9GMoxarjd6sjOIOtAUm
mrycpx1ZxSqayT3ZJthrVtjW0YkAyzvTyHaMtSqZeMtFLY+j7jgZsfyDPjowjJNk
knOYd0Q7k3L1nMfApuJ5gAlqN32CXsNAAZ+4b0Pp6Fme3KvWZFv+LCeLRajJFgsn
7LYs/ZSqVwEiOUqccAO4M7iXp+8xRLtKLmCfaEl8j/LVExGuDLaN1/U8BJHX8Ckl
uPLlKRjcvekcsk3ziEHjXAF1A5kmdEw4auOpTeu9WNa7EyHjS58iCXYko9kCS+EA
4Jn5lZxSnBwkj9wS5wK/Jf4EgFf8jZdE7QepsTWwleJAvfuYcmObSUBYEnzgBjgu
Jw93RfW8aPyw40pD1e24YWXgpBknBUeKktRyVgI5XfNz2ZqTer6lu5AR1XbUvPqF
hcer1qYZwFo98EJVcoVhzOeLPa2Zbzxbyg6mBvun8q9lToWnWeuxTyjoaFY+odsh
9odKRQfATq0ex6vHrMgHGZgmjeIEVMAwNodTx8MPbmJg8uHxgEQib2Y4SscoIn76
XDrsvs7lHkHY0aWiA4oBZm2pD8jxz143Hct20gzY9L/jaW+ZYH884Vl00n5skxY0
dm3ZhKWoMZYXS5WuliBS/IUmDfa36fS6vWUfmJ+Z2MkPaILWlhh1UhJmYfl03JXw
cubVOeRaDP3GWcIyha2q1HtJdkXcIzD6U25DWnnTkJxWWfX7KVcLcvuuhiTklDP9
NF7wrWplRHjSO5a7pDi9yyoJ6wMd1mt9+AfDKHpb/2BtQJcHhmBmFZOBCqLwycdC
xXpKiW2VypxojP6hFtl+oR8QwLVh9HCtqqJrd2VeZcffo1VmFXI+dZ9LLTf58pZq
oLft6AkKTj2Ls5twzrJoZu+iQ20mXJSexdJwppFbUdH7Y16tw8K08XrR33aY+dNy
+k4Gvm0LubaZN+dYV2jl/yTCRU0xnb4O87GddsmYl0Aa/orZVz0Egci/+eh1FS8j
ipaAmBe3P21ZxL5NFMfk1a/RxCLOPZV0poirnVCjwx+z1w5g3bfQEA8x+k3vpdif
`protect END_PROTECTED
