`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMdgzUR7hIajo59z/lmsXVId3MfdhHo3ACoEMieBH8RXxgdMllRfYmbBhVyH8lhI
EZ0QOErH9y0E/+480IDuSEBmG/uT7+pKD3nHIi7q6Rb7zBJiTZupP8/98ToYuLQc
5xC1g32V/n5OuPQT2mqIjvMUUMZ4CEmDzkFm9BFdVDaEgWyp2QP0ThcrDEz7mcZo
+rUlj6o2afAh1r1qwxbGXfYspE/F8CMweAmQspQqVgMR2n0wT/4C2ERykEcFiCDE
tXM1G4Gby6DQb4iGRR7lnA==
`protect END_PROTECTED
