`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rROt4m/gwv3eT2p34F800mzv9MwCXRWDYifaC6qfOHrfh0pU8pj8EMha2ofER76w
BP2rD6H1dZZWrDfN9SrPzBj1m7XVpFjDQmuds2JEBNKJFjD+azgqHotV1aGVNgZl
ympgY54VrgVcwlrrlJhlZr/2Y7Zt2Mo27NgT3Wk7R48JYL6hiN7Uv3mY77sY8dM7
AtpjBmfq7iHsGLSWCzpG7du/GMVm7ujGUTXyg3TeSxFM80elUb1vqvVq1UgbHzYu
sevdBAnQ3OAwCibWuIgVf6tBfa4eO6pVwcxSnrSkc/gI4SKvTePo59deH/dEg8D8
B7S8r2/HLvo7ypCUARo5f+BpDcJoYEh/HTh5sspgXESaiDYSvEyl/NlFi6VxxNMu
DYu+JxCdm0xv6J2hD5aRqiMwkHyLzfZ0bKHHf0AgxAR55wGOn3eGGOq0bW22dNVN
`protect END_PROTECTED
