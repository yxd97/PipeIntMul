`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6q2k5Wk/O52J5fztpHhED5/w7vW1R2+bCAqDmXw+hvCYcUxqNGckYxShxghRzc6U
bnjNBhn+CTPhFut3cWwZcbGVzinPzaoR+QMWhAlRbocEERYRoM1TbTzPyfWjoccc
5zaQxMouewIFjLrth5z4k4TLDTiAgWPYit5roA+ZCX1OGmSHR8mmK9pv0lp/TPxU
hUYzit/akG0S0Fw0Eoz1DGTOjVpB6hP15e3pHm2Puu2MVKJbONaILo/0ZGM+bOdL
mgrvd3BlyIH3zEqqEwF36Q/Si9USrtHcbd+Iw/+nc3jPdWgn5ECW2YjRz74U+Tg8
eeOcaAoLcPe1TlLNHwG7fPkaRs6R7QKAvS5xqjo9sXF7FWzjFi2YzttmGkckSqNJ
C/t/OUknQYBczBQl/x3EFcwLmpBheAYGobM1xGL6yAKkHtYVaa3fNFwvoSQdf9qd
7iC5KkA194k7FT6oCpL4XNueYwWrKM4a0GUaZvGyZcIbSjD2Nu1Ht04GFoafOxKq
EhcrsKO7wq0kh1+Ls9WWRjEUJsU0TVR+7HjwE3juLHjIdo4qUVIgakKMEqY5dWrt
qniukFCQuYp5M5P24EQfJA==
`protect END_PROTECTED
