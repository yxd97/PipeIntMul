`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/kviY+G9o8KPIdTykYkj4EYzAx2XbwEl3hJrV5WWkEkxP7IKaZVOiJmWzIUrS6xj
uJnzP7JXVOsZ6KM8xiVCpk4SNkCLN5TRAtApa6iyFBjT78F4M2ALfW/3LnenxU4a
mDJUkjaD8sxz99wG18uKoeDwwhWAw+bWQaoiQLIJPUVSHE7EcBL/axifUIAy2oW8
iX/4kr5YJKJLomDE8eTeS06RnHT3ouorM27qhWkmG6IlivYNoHACCR9DHdfXhNhP
oywV7S2jup2QagXrpz+u0DRfaAGdYZK7jiKss0Jh9q5mLMUb7c7lijSlQJzYIIti
fInfldcqn/YL0+r+EHRgfA==
`protect END_PROTECTED
