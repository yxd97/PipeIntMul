`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zSkK1vPZadHBFfP6Qu15SgbV92BolN7kbz7cARneo7aLezzAxw0oSHXJf4Gmsza
qRtTHgpYv5OdsKvEXHDxrVvFAMSKgdZLzJeiLXVKbK15wQN/+vvoQc0nYPieLjyB
c9kkjBRK4DL4mnXd1z/H1tZlv92qgsMjSgIpO401PVDqGrkNxy37l78sh4XCMBJH
1tHt84TfcJETb/uisCaJkFi7dB54T+48RefYw0RhEz+ONiJOZOl2IPVtgoKKiWA4
Xwmu7MM+OaP7Gh2xcMdmn9RnsqlJHWWeKTfh6mkyU+kSEkxEjYBLrVuo+NQ6uFnp
S/X1pdSxpKQesqbVw4Ll/FalTpCgyWbcREAxjmoptRf1UUKzquD/bp+eYcm8mtea
2Y7eyJVWTjcSmEg9SzqjpEkyY64geGu+4f89lwUrJ6TkHvW3Z+YYAwH2nmxshNuf
VSA+26aCqckO5S61/Op4FJTINOhh0ZnEPNjxO9iWhR3TxHkReUXV6p00ujSWnNGJ
qxyOsLip18d0WMMpr16s9SWEZOe0CL+wZh9fFzrCQA0720GK6HohM1dGTTRlZRbL
hlpBE+fxVUrGUkYODbbSqUoDh0iKd4yJjQuA2J1iM31mwsUfUUDE1YqBhulHYwZ7
DXjj8OjXFxhq3YT+15wG3pNkr2XaltMnJaNpDIvSfHXRNG2+KQf98LUWD7J0b48M
FRL/na/HObnLVH7NYtwA2LYdQbuf+n0tmNOzdSxrurmNNIdnVMH2eaoYndXnnqaA
vJ5JCpWqLcxg3wQZSd8NY8LPZKIhfuj2UbvYVB72sxA=
`protect END_PROTECTED
