`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Fk/flbSTIN4F/pMLZby1CIeeILz/TfQ1S5BZbUrMzoaBScgZcGxe2U6iCNAJajR
ZbDO74md8THOCDMqEJRcD3ZyId4SIvkBrqMXQg/oj76FfDPL1AIbg95JLEwsP2eF
wHoERZr7EwzlQ/N5w3Tl3DLCQ2LunSaYrQk6JsKleDxRMILSZcy3FNhem28wtpFS
AWSLkLdy9y9zV1vg50YzBkebdj1zPPalmk2EKeCTYarVstFnpPUUpezjiMr2O1mR
xVuckF+KSLznX1SXyQz+rQ==
`protect END_PROTECTED
