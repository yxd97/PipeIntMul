`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
erf6/sF1d/1qgtHf3US0FiFRO9hjd7Aij3wdJYvPk6mYkmyc5YHFax2b0lKUDceI
CGoYAUwDYg2+hc9tNoXu6tEVG/hQ0Alyjb/+bvbgCuy48kGT9Ysem/Q6sGvY83hj
Q5anAJ0sMm5ZWaAZ75OaVJ228zuooJpOWQPJe8lHsiyKX0aMh6vJp9z8lVAOzRZx
Z5Uag4ePZ1Q/YDCPORsZyyz+qy1yXOKB00Ev9A0MPAijGM/IsrNyeUx5ixCujs71
cANADqd+n+MWWe+TiHAiDJ1TqSzirlf61T4da2Yz5fAEoOyZWCTDB0fHMrCfUkTL
IvRi1RrICNSCgit8mlIfetFdepGBjGY3fM9L5jK0GsihG6ir8KVeTKkR4ESrkJ0J
TP/7npztXXtk6cDwF+JZuJp9l+PeBIjQDjCv/pxZYpCHL1apun1oV9yYyAiASq3G
dhEcUkmWc31tZEhb+4OoObF1B0bCx7VtP6ViCnd5zR8=
`protect END_PROTECTED
