`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
msS6ufvI5XCs50AR0FDH4yjBERzyyotvKLwDHLWi3mmAowvjzQp/TEuNZTj3HN1j
TxVsDASUAF6nW53BfcK/qYP3qbyIYDM0TJ+3OIzLaFTxqlV0hWL5X4MzdmvtTEz+
h3MCo7qqjWzf3ttBWy3YCDz/r/wjEx1DXtm6eJIVnFqtFbeAoAcHRSxI7iDOqRt/
JqivVNgRL/hrIeHKe35NGcETYyjojxMwujVQPRS5fqJWM+U2hwyPZudQFvvJpLGL
9jHu6cpkwvSVeuj8N1L4Pg==
`protect END_PROTECTED
