`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QuFTVHDVPPnqau9cN0KvbCNJwSm4Bz/eVFgsqCL8THVm0tDA+wuisRRcx7YdYeC6
xXPxhC0rlaAZM/KG26vO1I29JFn2d7Nv1aYjR0AcR41bclfPTNhqp5GzL+EZDPEy
pMPOjBUp+l7NYwp1NyC2YdLs6ZqU/f8UlSq6tBp0FltGlaGAwH5KE+xlpyMhzMRL
itMSVkW+4SIgw44K2k5iSMn+A7LJNEedUDfVAA/3xvWUkD7Net7qn96ark7C1enA
ZufomgCys4t4Ey/kGi6Ly2+9gPNSDojZ91d2bLPC/IgGsv5bha840IBQ8sWhgU69
UW2yAywaAZV+v63KEtAZw3I8nyeHt4B4il19P064cLUGSEK+BwUqfskM2W96rCLX
GTwg7ymjv3NPkUoHPCGk/D6vj9beAoEOwqv2Wl+W8UTnNmATCiebY0CCrjrwk1gp
b/9gsoalEj2QiJopC1ju7/QCjbJB/Eg0o7RzhpU0xNNDGfE/5NSNaOFqBFpCyx0W
ccJJGNH1DS7w8Xww7HKIaBM0kRJvO8s7xmsi7UVq0EEjVAAxumsS9Bmmf2Klp4H7
JGOkntdb3dCXU4EDCp314YfeKDEtSTWHUx7EL1tVna0+rnn71e6/umbe62e8l8kw
tflmAyjMCd82vZIDl5tK+g==
`protect END_PROTECTED
