`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HPWkBTbfmhwfO6d5bs8TeAvqboFYSaGjzlvUK4bVWTGqlodFLnCSEuF9zJUj4ejJ
3VlP0T0yNk295ShTKihaGaZWGF3x+BT3xfbtzUpzOiUO+kjJpopHc7LXGzn0vT9S
9KWvHyb5Vxwcm0Gq00p4HXfFvVUI/lZjQ4y4aODOBFLUV7gS7LHAwrPWFCUboT99
90EYJ0AlFH2jUFeCqbhb6HOebVSIdKepbanbJMEYbBMgmsblKa8Yu7rbQgx3Ij5B
OtTxhnah9O9WKqgskRL4HfScXjanMx/HOppEcqeE2K0uqTabt3EMNngb9s2D4D77
rT8CFIhJrTgdHm78PgflSl/XmUFc6Fx2NxFnCUm4qzI=
`protect END_PROTECTED
