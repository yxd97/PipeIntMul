`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cf7+LggivjdPVpPqfhC1uSCeVluMeCHVG5YCgJZyaMlrWKlV2t7v7oY/IP2vb/R2
CEqWBCj8YW8vhD2wU5gkJlHM1XJ50swvAS4S/2UpR/oLjw9KuARDBgWObGVHMQGJ
IiXWW0WxR/UIR/yFdaIEgvs357LW/5co07543mX3TKdo4rNzhCFjeb+k5BGg9uC+
nThN0ypCBhj1B1ShYeoF2zSHY05cy2w0GBS9nfiRZbua3TBDFm6H+ennzfcAWJgo
Ro/AykM55W6eztXQpNDqme+HpQ8AcouPpZBrS7And5yIZqTk16m9jG4MsnhCVgW5
dDUDFadIYPpsJ/Plt1+mvkPWm3aJ84kvfNrX7XJuDMF1NTKwEbfPT3IwdR0j/7jh
Kn24GxXTbONUnxheak4VEzDzycVNqLrRW9G2srjGFR6W/1k0dLpAL08EykHRfcAi
rgLM5MUbUEaQvcibix/Z4PnhwiLd/7/+7h2wa5NAFyktkN8I6aJojvbPGmcI+KOz
`protect END_PROTECTED
