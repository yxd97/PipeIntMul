`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MR+a+qrTE8tvIvBSK24TdDavKF3q2X/Pwk2J3ONPn5NrrCnQMpd2iZnHc7A8DMz9
q7xZ1Qm6Zya3HWHURUejwvzw7y8pUE1DCDSgZuJEItXIsKRVa3yPMEdJu4lV8D0A
jQ39hRaFHOHmHkfUzmq4WCQt5GiQTc6izfDR1If1NI8kJdYYCMYPaAdwzJrkQHwy
hd/yaYcSBYKVDLEWb5yzU9/PwZss+ZnppwwpyoqWorXGnIGYCmHdmVzm97CFTKQU
x5boSofpKrcyzxt8lRcxlwuh8S8J8wn/PbvPFdd7kcEOiNeQiUeqmTZ6iPgx3fG7
xZn9vXgIr1tB816qzWDq4XcEwH5jC0NDenuqgF9v894YcI15tPShw3x7TzUgjn6l
wRRKQcmEz48AWX28UQ3HLWOwFBz+mieYL0OAh+iQSD4=
`protect END_PROTECTED
