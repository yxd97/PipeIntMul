`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0LYkjxy/o9ZgE27j3gVGJ7OO/z+YzXomfQCmqTWyfpcVq6oLhOu12MgnMHthGk3J
x4GkJl1cpha9xMCO1s33y16djdCHico2Rf0V0At7OFzUXD7bNqYo5WhrtCjKQOb7
dEdB1iT7PktHMv4YD1nZEZ89bpTm1/YE6qLqm3JDV80LaGbP0Novr0i5fa3ID0Uw
q50VGQ45vuLTQw8L8LakOA==
`protect END_PROTECTED
