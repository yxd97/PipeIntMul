`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMF86zufQ5zp1EGsZTB/7xFpM6Y0fJUUfS8jAYZE1pksFkUSuZGuy1UrOJuG5CmK
f5ERHN+E/puC1EsN35Ji9vNDwKUW7aLJlpyFARjqENJ55cUAIEOerRbTM9vBrH+J
31id5cUtGKZdaf6tP4xwloEfhdHqFgwmG5mau+UaK6dfBVHViuIniIeBJgCzN5KL
4DBfW4yYmcNcyPQPTu2G+BrwwjGMiTYivDKBJQZoiwNhgAjYi5aoWk9JRbRwSJk9
qRlv5ProuDH6aq0o/RXl0W3PjANZkRoUBaeAmiIFyJHXbzOatGZFDXr/KEzH3/QJ
ViOo63D0AWfYNXBOOxAdq3hdY5EWjec9n8CuVNgkvxMxyxT9VAS5sTb0tX9MKsea
WxsNv57F5rl4SQueukT0nOQW7kKk0bLCknp851Drl1OOFTbsjRy/qX4j2FQ6inw7
TL/Qdld6TCqL0OaBdj4D/mDXy8+YIB7xSCGSlQ7kMWqQVKn6KQjuagHP7F7DmXTk
c935C9EQXRWnia5Lna0LeqA4dBN9owDERLXR3Oli3nngyr13CU0kKFzVFo43AUM9
jqc+8NVb8Nb1zKeXpcoWFNRl54LqcgwgoDh17ODd/sdK88e07b34N3p9jKYhQaOg
DZyCop734v+6GnGAJvaQqX3F2KNgFvxa585jBLM9dZmY3wT96yw57ezuRxWNUPPW
l0iwia/Rp12GsFmtiRBQBA==
`protect END_PROTECTED
