`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s5tg7l+5FnTX9W6vKWMNNz11olL95TG5Rx26aQKHh8YWz0De+zBBU3bacVl+G5ap
hRWuviG1wWJPXMWvnazRhZ/TSGTYyNUSkWD88Gw0haWw6FCERHLljUoxYYFaOJXc
9jw89hjUWxW99vsh9BtKxs+7PSjD6H3hJLxPIy339+X/5w1CgcOGZg0LKOgefV5M
v5c/PYG+gY6RlqM7zRm9N3jpMsyB3YbT2pJeOHTsjbWdNQqnJWRktidz4hX9ByVH
Xb3P8LswW3mfs8EFqHIiFiWd9aVV0cozjkYkP0lXGvn5JBSNbiX6C2WmYgV90b1b
AMXFcGbTtnkY6B36MrRVJg2+74gjon2mluwaam9a+rMDLt0aIuZQbhVY6+lDuRyT
QqpcV/CTWXFoyUOsrfCxZ+AOdkszHlUgXERyLez8/oBJOBMRMlxMbMQxzLmFbLl1
jIcj9T6JZzUM6MDAbTqTcjMMs56nhs8Qk5tHvcUl4E69TuDPKQAGPsByA9g8W47S
3RzyZU7w8kzgp5NMwYDIg7zOwEYGdxRnSC2p75CT7aHNau9G48D1AM0hb71mrZYx
5hBEzFYbvFdgxJig06gfso2w1DuMcoLLUbSyLcDgBHYHOUNXDYA8/51YT+OczhNf
gD9u1mOC9kh81675ocZmlnAUVgWz/KVm9wFjlmaY7evZcsuHo0vW7NrAYndch0XD
KzUicOT0Ix1xNmdzSLoEHVRzvFBykeVuP5Bktmz3DF0=
`protect END_PROTECTED
