`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbbSpYLpVnr4hwXu6SiLqFcpg1lo3IQzwvwB5rPujh1NDIMoDep++xZ0trm0lFIr
G4D5ktlWX8+tm/t5PIY5VZ8mpka89aoz8RrAwt3DK2yLC9g88Qk2vlMyuWi4iQK5
bR746c/CTExmPTd1gn6zNeVocUXHlfbkxWn1pczMLUgc6ufqpiPUJ5ZY5zjsMOTj
bvoX+jqA8AbThs41+WIb2IOJe6F2oTsvSnVtrOsCopcZPvqbRfhgZqul7mJARbw1
PtR6YsN+PC9OcfHliTVBXP0R77v9kOknM2Wx0h5EhgJxmmQKPKzDlxVlko1d3vIa
`protect END_PROTECTED
