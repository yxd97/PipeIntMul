`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KosTMnwcN63jPrtkfCGccLoTGj//8YIA5yCByDZawuPPwPB3P/dUPQdH1ehMmCC5
JQdnq2+gnyuModjjNT2MR8I7R6kJpffUyvPdnamYWkBoXmrg/AudOewM4iHyipcH
LbGHOvptIr5N1dJ8DHMwlNorqWT3lxgVS/B27mMmg2ym+lxDWLDNIR3ac2y3TdQ8
+/o5SxscJtb/24p6CLgSEVxGVH8Sv/4yEOEtKvPg4+FQNaUI81Or6FPUWcg3vPbk
msfNIYM/hY5jurioFErzrHbq8vYEhCkz0ZQf3lZ/FQWfZsYmEEyKRnUf3aEr1idN
Ki3SqB2Erhs+jntPgOV/tl6AXrRNTp5qlq7oXVoEho2RtDVjH6g3I5dhrlCZkZzd
g+Tav3sth4QNpp1KWZNCFurfdtC8D2pTU7lJ8XEk11TB9/brb7w32Ez800RgX2Cq
VMFKLHAHw4LS0WX/O2QeYFP7mRN1+lG8GQceqGHQiGLrWaZzRmXJzbXM7nQrR8Ae
iioBa2dMrXFzO417kThHamUlJ9Cv9ZiRmO8T1AXt4VlGCxIn3c9ZMc1+RCHv5/pF
eaz4154b97fFKyg0Xqyi9Q==
`protect END_PROTECTED
