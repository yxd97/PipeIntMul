`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TmikmsjRJ1S653B+eWHUBLEnjSDVJtX+kNXhckdJq3hqvFLh5BjT3judVLZMjww9
s0wt9fiS7qvBbXJchzWujWb7PmodFq7EMI8BYYbCJl0LgSSNRcYhiRugAXG0eAPD
dlLSyLhnlm1+2+7cMIi+QF8gV8ouqjbRrN5iwZkCAQRoCrJItNdYg3Uv7+YUoKbD
JoYOczYazAhnTRVFU0ge+sCiMWdZ0eHYmwwsMpDh+r8raS4TKbQBij5VjtiuQSF8
gerkpRHRBsQycoVRL58bpnuTdoMZCHVPUbgO0Ii3A8uUy4ijsFzhYQZQrNySzOmE
MrWbEIOZ2UQug393zQHYmeuHnJuDk/X9772+j54cvLfAXZImthshvXQyzaEgggFk
VYsmIknPJZE6WzT7WuNu5MUXY0QvCZ/S9N9zpM84vvZN8/ob2g9OCoZhXXfTqORK
AIEdrn5UYyvCRGQOdG4p4IyR93hzQx7Hqq1m2TM/N46V/LgA9d1ipplMzI+3oW0a
EztJMzv/pQj0iRSE3WDk6eE2aiHetvDqlambYn5PhCnguPUjDZlfeLq/0fv1ysGX
`protect END_PROTECTED
