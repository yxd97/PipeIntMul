`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jemJdkXom30SbE0+lDmXMCz71MRkmJwtM9rpqUmkLG4qMvtCXVmjcHdQjOghEMVu
Cq5FKR30FWKNDYwnBUnME1Ihfi02ClStLELZ2lqVDtX/Qgn6JAZTkiZyNk16P/kT
dWkAlOBRLiOMotukZis9waxXNPSfFtHJZTEcVNK7SA6I8McJAwUNEdJcjecZ770w
WZqkkAC7QZ1habooaP7/IABLMCYZkHHsjY+3rc1H5nRqG6+g47gX+rq5ejYQFPIW
M6EsGr4rzFtlHzza4Ov9YdehiYCNSvYCWA0fSnkOXYkZ5ZznQA2peO5CJxpv5dgf
Ybr0f981uaSkv3r5dC4zdL9iglEnxujZut31bM/v/q6Q92mias9GG8Owr+rkVXQ3
fj/L5zcvv//b4unDoyA7DgPOFs7FT0d3iKgzb951dZHYhxw12yXPIrKqJsvMaa6R
8dSlwp+LrLSrIsYAPFAaL86wfC4u9ZyKuIxkMEm8Ow74InkSrlT3m/os/liiF1Yo
yjAOIk70zYskbUo1DK0aQf3KSHlQV4ABWjlDnkqAykuJ4Y23U8Q0I7wLEhSQNReP
qxvg0/f2jW21YwhNwGQtJAbc7/W4Emyb0BzKsovSLl312FulG7C4ciGGKiZzMMmO
QCB7rSPnMDXdVoymQVW/C9bPLvoCfzjdLXic1M01p/8kLCWwg5gPpxgMqCsJOgOp
H6DbjzCB4n2UN5GQbFJWyVjev+8qSvqap2FzYayJM0u8YvwJ4IPOwjO0/2vDdsFk
GPZqMdLtVtutunF8ROQYmjMWYQHrrwfz+ldeFQJSojRY7gtqRIBiHQ9076zSnGvj
GR/c1muaUNEsJfzv7mZktKWLonpcU6JeznjJFKI/qzaw8Tt2q35pzEob0LDOFQI1
qj39PUxqbTy7IBtCkzAZPSMemXRJXBROGciExrIjvIJVw90MXE4PesO6A11lQvP2
xt+hT5ZYx9ff8dU9biy3q/DFSkr62ogt+fsKEIt7baSXC2Aqe6xMPwdOKTKrBH/q
hWUGqiAiYJoKm7jaKOw4iIaEm/mJqoxj1JnzdoEl5oEhqQVyWttR62OiKOdPuLi+
ERhbO86BebBDub7hEMntUwYPCO3a+17HC71gJzRzt14tWsz2San1CEjifIrp6dmS
xPumlyO84Qijl7jEFCZaWwoisSqI9jc0WLAUTJYKqggCTT7DuNJKQzm4oFqiSsvE
Qi1rlT0bBsGrHTmDnxUKncmqIp+EbuTBAUuSlGsiVaGIP01vHhgktF3jRkkLlKV/
ORrNTlw6TpeEztVi62LOGvx4ni9NmGMqsIjpyJ3cFxIicSrORS/7J2a2GKfwKxXO
x12GeRYo5rS2XNjZ/3mJIxTHcm0LOGKkO2hvoPqxuCUsTkJ0T6K2NwtsMwB0WIF1
5hfIL0Ql6mEszCxsxYs1v+fsLy2NPZV5QVbzSgsOpsgUhBuhIHKYBO2BjnB58N+h
ZJFDUWEcBpLEB92MNTqUqtTAmDbX1Lp2fKz5QB9v1LZQ3adcFegZyAs1PUgDF7cW
GlEa6ehi2TW7pUn0X6Mys1EP94eGYG1xLK6UVdZ82yM49WimTtmyAzbkaaXQyuWC
fX6PyQaBokraL90WC2vu8hNS8OCi4cgCqkzd6JXIjmTp0GWdhduNmw+iUFHbWQcl
QQn6Co/6Cf4oEyOjRTZUvPS5et8d8O5E9+aR4WELF+RiAcwqxNUk4eSmvfKjxE9F
MSENHULQmrt6wAudcZgawyq6fBhk75Xe4VIpKbong+phQ+tqyfpThMAeBGIEiKbb
YlivYIg7W8cndEK0+chxxYS78ZDC0/Ng9KMCbfYpsp93PajH1P/69gpZTSsydFIn
QoH3hLDIxfQKsN1oE8tjuGeW/ExP8qI2JpjjJCkoZLfyB9ruqilJT8GXHON5CWcx
8TZFzvdxPgId0v+E72X8+nNTyi0AiGDIFkR4mnlt2WeJ4YGEM1HReaLvOUsjmETH
nsoCkfO1S0E9TN+QyMV17ftBZu2WMdWSMJQtDQMFcesb9JFbHqjuRlFUOI36teCB
vZYiHNoybzS74qMl7vW2a2b4s9RwErI+l5ZwXYr8tg9bjo2lbGy1UGLIWqNl5IKq
8WC6kqVr1qwOGzwa/ESJF/E6keHVr6hkm533cQ1GrInNBIBzItBWOlXDcq7Hb4sP
UyU3v6xk5xtJRkuOxRBWztYT1j4zHW/XzbaGIIKH+J7my+brD0CKF1X2Nca3WTM0
rmeIrJAk+Lu+IGzHsM/bTcoZoFldi00adO/sgJ3kM1FQrYHEdJQLAb8Fk4BnqYP8
mfRsGplCtGnF76lblLJht9OKEtbTs28R6vRI4xt/DA9TkODLS4Tb7kPcmJay//fs
zJ/qTICk4/HhNAdOCrPOeNVY/cF5IkMfy+6SJA+OrARCyeWbiLL6K5AzaTpvw+nY
4585ykVoOCX09O5xZVWwQZH7LYC1HUUz3HmrLAvcpj+jDtd9YFQ/VAkCNHWrs30m
a16QX3SOWTHH8De2rmhEbu8++5i+e4OmUAAGB++myj2dniK7649MqMw9rSDNzU0t
sNXn2THyL57L6bF6lbLLYyAovQPf1R71Ol/CNZurDlbLOSOZCWfoTRpmkNoF4KN8
0xl1DcUOo76ol6hORZ8TfadUF8pvqWtIzBO3zDdZmH1em+PYrbxegyuEXOqyG6wT
NXpUkNvnQioGOhCuceZY9MQhwdZauGPEK6vo2WBsIqbmRPbxH/YKxpL3xV5JxKEK
G2z7rFoo6evZQg3KCxKr2jPm8j33sdb2DNgFL3zWIxut23L4Q/eWCvfmJe/AZg3w
cPHWHHaDQ+2L101X08IQTfHFxewM8MEMKxy9KP9OtDD8SSzRJzg8OWsmHtJQ5vAR
suiWjTmm/MRH3SgjogUel91RRS3Zirz9ZfO/TtFbJ71/soTwwSJlIeZcrjCpaVGS
iikDeJPV9yAWEMoK1fcwIlRZ9NhJuE6o9BX2q8qETNnBK7T4xAJH6rB9zGk3n1Uh
k75xI9lD/VuDOIREUt5523xNI+UDCnCPs6j66nhzBTEc359Syl5HL5AuzENbYVWb
wbUqrGhnpzeSuz39M8Hm2hLw3oBIBZaOS+ujZcri2Uj8ieIP9m9k21ugjFtNYHyf
usyHV6gzdcNSkIY3+6Yuwd6Pi1Pw/59XxfCLF4y198QsnT971a3QiM8uRSLk/bQi
hGOrCBctzisiIeNR3R2iI6XgbKzoK7F62TJm6abphmjrYABqmvkkkxyx6GyBVFgj
oYP72IGp1ib0l2PvZjS6wN55poc8WjhaUMfb36Ni+tlWg/T5/o+fVLBPyCu+bpOY
qyDjs7OJChQm3XmlbQaNqq8jy/dmWfJ8q+kKXHi9y1k6PXQfTIU2q3mHo4TQEDD7
/BTI+JxmejhbjQfp0JzjnveXzNUY2lut20YjKFFpydJqe+5SxHZscoLFBJaJcPxv
BbaCxeHZDO4KLM5kzupHcTeKrDMuacnRITscaanX9nTcsO+fFTmomTWeonMs9pcC
Jt1Oy0NxrMGLEe4mPEzCGEDjOQohSd9H5OHNkcNWSdah3KboFLOHZ2pP43c+9FAp
2XNeWNPmwNb4j5opMtELdkWpH3NOd5sOVgDRAk9SFLFkr42wDr41N6ITU7dotVYb
QOsxI4ooPLQolBOzR6YVy/6JPJMVAX0k78QME73bJjSdnzAeaOrhJ+xhZnI4me49
sUhbetzbqUqtRHRsif1EnYI+rnaHQkk0UZ7oP6+1+m1skJFvQu8mRUiMEa+CxQzr
uBU2C5a6bPN3auI4V4fKI8NoIZ4s743IH6LsSLUP2W5ATDOfhy1Z/TeKbfMTsORy
+M1UJxGBw1rePqAc4U+b6nkPwK8qHxXtHcx05+AkLc+WKfuXSBtnevEaOHzRGXar
kdTyO9T1ugW+72ZMFqeh7iyN4934KSSutyLKIXfhLzuQqZ7JoANw/LNKH02YsAQI
18IwzC8Dbb7FH2RBmdLwQUvwE4rVqv4xKva9sBAfhfy/WBr2/JtayHQtEvcj06RT
4reBa+6smjZWzGBaCB+F+MjHMnnb/rZfI7rDn7239QQXafS9CHdlsg10rAmUAjiW
jIwIiOtr2xJzyojGw95z2fsfY4Uzce5bjqHrK9iJOC0y6TYS277yETWeu4aEjqyp
qqOhE9oxmNfGXmlgspdjR3mW3yoe+igjqHG0je83TxdzVqGrg5s0QCmT9Ni2EN5l
dUaz3zW4aHG9VAqH77Uwnqjp44doLguI7pyfN+86OV3p4txfFhH2YKc8z+9QINyO
h+yKl/nUs+seZIVhtotzfA7inoNAb/bXngRpRZesxLUTVCEWbYSlBrk/wBzzBGpM
nbwMA55ciX9xDw2bdeetMvW3Dwo2STGZn11gLU5x6nIYOCsbwqJ1v3CNCVKuYNj2
QT//7BGo3XkEXzm0Qi2HO32R85yzNBqBHtXhYnUWeZSiwad8AOVmLzgRKl1ZKjHf
K+N9n3XoEyTaSWF/mF9fiQ==
`protect END_PROTECTED
