`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g34vsRXqxFLqL/9aVpp3J4l77cZbxG/IFvowhkzedQjjYezpT9VNzerlKE2DUkre
oq0jESqlMrZYZBUyJTudW9sPwQp1NjKcgtMdaa3t+XoPs9pQZztppz3hycCUYsjO
6nVJK/vLqdT/D2GD1bL7QvvqIk/h8zZMYDtiYr65C1VtmbHfUvReNCMkRrtwDInp
f6p4QmOo2DY7TaCee+pQ4ihmDVFtfLs13eY63c9iG0eu1wY6woXFepNwuQQNjEC5
nycLdg2I5nEeV5R3Lna+E+/bkf2RhjA4h2ISyqLSTUe/OYbfWPOxVVTmPG5NNK7Y
TW9OH5v4iwXMPOhpldAFOQBrsS5cIU2egdBG6FP9Xiv6xFwrqdcCO/z37MDF7BsS
ZmDKJ1pnXEXdPpV/y8En46QI2Ebugrm1JcBhKQ+AgeEXVQchqh+nfxhODCO+EDeL
LDvHvCi4oBQJpgwOdaXoFRoF23y9WonbwAGfnZNr9oWFM5GP+lzyp5Awo12iPUXw
TDH0Li7pfF+sB3/ShVNmDdWsgyH2eLB5SEATgfQx7n9SSKtKiLJo61wC1e3S4Y+/
nkFWFb5C41QmcALeVXLfof7KBXuo1QDs2tTLIZmLcEfxUiAhVmCvarSIq/6Dag2T
c/chaV4DkoaYIEykAUR2z5cPmYtTjeCXu808EZIZeCfmGYDxytBNxfChiQMD8It5
FkuBEKZH8gRdAIxBQHHhViY1+gRj8wErY7sj4py+83/AHCkzm6eTarb9ukD60hzz
FRQh8WpVPFUqACB+sbrkWPlS9DeXzzvlWSzfXDFoMOWWNZpm+RIkdzYL58AXm9xf
mXeowq2IOoLAQJL3kHQWP3EG1zy6AEnsvF7dmKpM/3o543vSzC+bYu1P3LK3PWFl
x+mjfB6H2/YO82vBBRR5BF6KhLL6CPk8epSv6A3AZm/GGjVxFulGUQxK5EaJlT0v
sya7CLYpelxnd+iL6MHUlawPJtWqCpo6rUtGF0nPP6UIeU+eZr6saem9dXMNUzq0
FlX+CqqbzhXea7rR7J6lMGtn2JldDLP8tmbeU+qCsb0Kc6s7y+K6zC7iQ0W8Cabx
Bo1370T4xXnEt4c6PzjifdPgkhQ3WcsYAc79Y6446DP/OjTEUvJlmPiHjpnKcIwM
QzdZZ2o0OnutoRRh2vAwiOB/CYfY6NBKa0SRvnnPW2C7jwCTjYifx81GeOQdQJcD
ioZZih7Zx/tWI8y6ltnVJ8mj+yZHy+tEUFw90Omo/cPHbS3BMuAKZ4Cv7dCRKW8h
qy3xyUoCWZMsrwktw7bj/dJ3Lk3gsinNTM9985yN3dEQoQfSmmqeBIUxJMocjZZI
Fe9+04fjOsITyk+XH3SwkOeeWvbUwlcmRGKA61S70rOjUAK9WIjjkMQt3xUdWBvV
cpZz5LMuLiAdi80i8tO1xFmHuDxpWdsbsrrBV4Kg+kXFAys0EN2rLRzFOYIZMUbs
VITyvdgMhR6nYOCEFlQv9MdLU/GcrTJmswwYR6+K45lGD4Mlzk3fScjSIHGupyva
8l5+Zz+UQWTGoit5jMHGLG5lSw50r+rPLH61w5xV7NHPLSKHJ2vO1rDgCzhY/UCa
iLc5vKvu1owYM3MCia0b2wOKceCSBD1kjlZqOIUT3yAoJdfa8CDG74BWYLGLTu/J
emdtXe0qWfiFs3sg/jr0cwqPU6kavS53vVvGG5KW3qbpfGEjoyUpK+FnzysdYebX
Q343fGjuw/XEaXb/bS2sghEZoL5xl9TextIG9kfF2WC+2ZVwF5+tUvVPd/1JDxJf
YvLPeJbrpjliQiinAnJgoW/SX2CvZqAxFIVmEupVxlIxGDRYJbjwAn4DAoOyj9TT
EzDAVmYjYqhjYgEUjDZAFv/gIrxNZvo0T7s/AfFLbAOAinMoQufr8R3o9XOHjeoo
2z5GDQk5kCMk0jG/59aA+cPTQCXX0eQNSwucFfdl2bybKZ78DJI6sILwXqXut4LT
0i/kbCaGcQ4sQu4J7PCRr9wle+VRHBuGMmsyhmj1wavYFmSawkap56sfHybqwb49
Jit7+wgeQrcOtSzz5tU9bLxYOe0jdXrV2XcDP1ta9luuQB7SXtI1EQpeV7BvQ5gu
8BFHjNHy+ePOPlDh4hUMfRa5U82EEwVc6g5c9vaIU7kDLY+XSRgQ7vT9t4ry4GGn
A1oI0V8G9kA21O+NeJYm6s7vVUOjBJMgFqn/iPDJw9bvv1Q1fQ7ZksRaT7FZuIn6
IEQDw64D4WB2m9q1Xnlws+3rgjBbCBJotbzQmQGlh0zmvMLcK/pM9ABC/+74IZHk
NKP7sSRyrlljS4598eYetKCsa0XdhXsNVTUo3mnj4D28xJE1CHLSgmcCgOVBIQlp
RI80GqeKm5CYUbafKCMqPvl4Lyz5NEWn+XuymFa2mj0/1gPkv5oaTnxBqpnyg+iL
SII0eZWXjRviD5AST+Ih3XSkOljeY1Le8zR0wlwaFrpD0Zq1gatsnY183MT+RVOR
a/ExDqxXs/Rzv4uFJ6NPz6iWgIJetJLyd4TCfMssAF3N02r5AZuhm8kZMCp6lRqu
In20dOuawl7IWnGsBxSuio0Pqi6TtWmxo4btFPuCFL2AtIyO3H6S0WtzGjlzOMCZ
3os2m2v7Zdk9vmZVw1bl3sxaFXnbi4vxW7mJMvRbK7cDqQbU8EOW7ASZ+1CmIVQF
7Uenp2eKqOOhqaexpKGYbRuRrD5rFtqv1yri48vetylgzmc6A2agQ3OltSE2huLk
dM6efRAuU2gD33jUPdG/ONPnrlVnM+YJsITe/OvdUTAH4y/IRqcFdT0PNqiihMUv
lKkR13y/L13sgVmRCsE0ez3uWrC9eV0P2Kh0rSAtYCenQDlodg9g+PtPSnDSN3Ov
aePkw50LLqn+3OnllNWFvEPr6gYe+WdHbAoJ6xPjgZxn4OU1aNm4SFATmQPbwa60
zMjgJbg6khNRJU7rmwk/W08CMr771hp06O2FmnEjQFw29kWW9KPoP3XKDfyIQR4U
DWGHmBUAPi6JcAghM1P9bS894FpnXCPfIbgnHx2gaLdEgwI1ay5YbARBc8Bg7Ngv
N+LaZYv77rk2WxcRqWZAvLm2wHJ22/FtojTdH6i0XFYsIv5OO7/jL+9Hz+LiUvJx
mI5pN1wa0cMXEuBrV5GomJNg4HmiWnK5w1y55Kr9G9Quye5Uc4YG9oMkeTB9E/gi
tnhOJZULplUDczf/dF2S6cM4V4NgDZb8WGehnqJk9VP1WjQfh+Or0t7Jqf84Ukjn
bRcWJPCWxrkzMIsQ+V6xImDc2mFE8zXg7gxmG1bP+dtru/RZ9luK0ctan6+7cVd1
9KQh9rXUmzVPmNdajKv9Qg10oRMfa4bwKR3iOyzaPzhenLIJ9dZdVi+gDw5apsI5
R1jQLWu0uSh9i5Vv2OLy1j+ZokvkHrEMn7vNjqyqxq6LtBirUWh7gpfxY879kEsv
W9Ho36EbYO8uve1a8mF1t2f1JL2swixI9/6fkzV882bWVCKYikMhM5cpJ17nZXXa
yTZrsTpR4lM0AupmdGCT9I8NxmJ022B5xfOxJJqE+/spjAEZmVpwKjyV8XKdWTQn
B79diIKSL5GXpOVpvSY/9aZQs1l+RMa/3dt590iENwyfLtd7+l90cjc+k7d8cGmL
QSObSCFp+QL78o8XUVFsNmpV6EJFMsur5fdZQrEWYJ8ZyUKtmmoZiZMlrvdxbbU9
FEJ7YkSkwBNiUC2MlHRtGjsGHTUm9jghEFmDBDnBdKqgeJdWMRYIZSR5CoqQYYmZ
tdkNxYtR/PQSsg2rpPcF2BRRni9K0gNq94MRsD8VoueVzz7w2nbs3t0TpM73kpfT
0Bm3HjYHlGaftKfdawxSPxkuv3S5amxBNk81Dr0/xCkboj5qgqO2686ZKQgTBolA
OA6CX6UYSqEju1PgSAR4MB80ckuxqyCdVrR9mMiDhqn8MOrQA8WcWlwwmuQg9o9a
dw9uPg7tDpWdb5H8Y8E/S88IZMZ/xvCNnVjNdnXmNAnWbixbQYl0z9EvWVhrF1rI
iR1unyfTtilc9P+p8IU+U5skIHOAgthwcjLJJMlgzZr7nhKM46M+gMSOMya0HQVm
CyRl+d09m4s+pjVxya8ow8n5AzhnO1N2qaEMaKXcNVJi0Fk0NHkILQAxwgkgFqV9
ddxszeC0GHJzrYa+geZPwd+kReHtDb9oehONAItob9GxtFWMf+LqOU97GdzQcx/t
WJ5mcAGzXhgzOI141HEu15Yp/0OJHnwfWOWzBfDswB9ZxDHJzj/RvQ88S+L322oM
jReXp89AVMlPMESEcRiVDyH47owHLRmHYgpnh3Vt/6MA50c6g5FO9alIVVzkq30S
lLarkyr8P8s46Ead1F7AhveQgaZVcwvkTysITD2YAqNfn4lP5NgC3XlaF4aj8vSI
qaFpJBP6pVDCFVWU7bIa3/gm92DzdWxjdbUN7kdkY/Z3EhjbScnB5ydgtNDoGrt2
DUgIg/AwVCMJKfTxzzh5FCmjnJjjEq5rgxw5mbgf5XlKK2FblW1r/GCV+qJBlmSQ
OpXVKRulodLoQDlzbM1xU10TLaRmT7UpRtw4yS4qwOLvauVj88D2VM20iDa018xw
qgQhJt0qJveOnTXKv6rmawQ/WhofbChfz26KKy8slmO8a8AEUB3YvbmrCDRHJGH5
86c/cKSuGbON9WoMv6HxDWhnHO7io/QaLWYCrE1U41CQNoy7di36bq+LRP4BsXQ7
R0BfOWbFhAvNpS9SJXrCjOSfnh9A0Sc3CD19KbSCTFYfJWy6qU7ewiYq8PZOwRT2
owsKLV1Ke1bwAULyI2uWfAVa6z+k7NY0fdK4c+YB9caeTpXrlNY1lY5yoGsUfIgN
INm/i5XVlOCvD2qNpmxR3fk6zutzeS6iwV3o9Clbg96/+1zejBeD/snBdAZBpkiI
aRn95Mm1Rtn2V4WUC5kLdCh139phtHPD+UrFntZ8CzjgtppYP18o9IBKd0A2nfHt
Vk70cs0dbcYQgfq6ZGu1EqWaUhlF0ILFfTGYGej6tWdn4ZeNSN8ECTeJ8aTlKdI/
fdW6PKW6lJXFV0AwKBPHa6t05Af3Ady6Z+8RHkioQ6SQR/5BinCIWZ0/iFr+zSpw
U20m1nqm/a/XoNbvh6rlPRZ6433Ud84J4fJdy1Jgrgc5/+Chyg4toblCwhdvrQvG
jIpWLEGOrznmmlJcDZREftB2fOwyTykqWiC3FM+fzxECxKXEE6Z9Er8NZV91cIzf
Ncu5FYgaWQM1WXGJk08zUhyrR7VVws+5/HbdP3xwvjjxBB4u7IbGi/NlhjooJnHM
LxwL8RffQ9MXq+4cpBQehVa7Wta87JiQChToqzzkcRL3gV+qr/o9N2HGeX8qlndY
eP8lhT9Qky0mQ1VZGsByQBEyyWJBROOv+AuoxxFAMG8XY5JlLjVwJvLzf0b8V4Mr
uyAal/C9RLwP+KF/G3JofhcytnVCraEtES6cHkJ8kiItNopdm01cciu/SPzDU4/N
Je6wUa4vaeu9qghiqdmI+CeKSxC8xhXy1XjYJyuTL9mPfIQ9yFLVZ0ZFja9zkrzr
aDprNL2/Cid6qT63Wt4LcQp2vMFs50z8mM6r0qD2IpcWhxkwHIiXKpd8cJo8XXLn
D7dJQDd6DPF174HH8T8Q/PcfbSrSs+4AI2shzJ9Eah6uYyaTmF4GX+AyzvCn1cPa
PweCLQ4SJif66W0cE4voBJFazIeSUHjPlYnbPR8f2Awaj3xhEGaI+VQVoyzI5EEw
8CMkO8cJqq8aXLyHk3glaWPxbqZvEMHyfa+NgIDqu0yVLA2wC27aVaOMocb5o8oZ
dpKU2kFg5nfxKN3r1nSGlnoIVajBTL/WeeMm5H6xQlYo0iYfBMwauQeInNHvtuhn
2kYcqOxOQpg0JOEQ6XuNM/KsR5l8aZUeIPItBRuJmtOdbfFt/JVzZ4Zi9koi0afT
RcLL76IPfGR4ffETU4Aseooabp5aMJ1xyLJvkQSs7M3nbcsEgMs6ZiD+EzCy9E9J
6FT5Am+7ukYeI1aZSMAEwTn/Mwbu6C0Qq9GMsLMioLRB3hpx1RoyuxYL/m/r93y1
UCGPhuF7RJaBn/m+OSA6upKnEjHcUYba3AutuScHNLd5tyrpH69QTjwLPtlUyT9V
vqvCMmMKEDhPhyzp3dzZPExHNK2nkkFsTzgkuapYJBDUJN5Q/hiNkSKWYMMpmqfV
6FTSSgY9ViUBK2TrEmG6KyCuoxsLeBeugytOWYVJydsAJQTD9tvdMGhWl6eoEk4v
xINWDjUHDG7HcnvS9CIbavntikrGTSxqCz2wMXg99sd67pokv6BXtB0E5IKTwEiG
mWtcZK0ZVr6UnSoxR5BKFemfq9YZqTH+Dmzo66nBbmz4eo/3YrOZ6ipbKPR85fJ2
Pf18GcygK/OzE3T9KI/c/hVhEAJ8q8hmNgtwOU3/ARLHRZbAKjKUfTy4vLJOkLk9
ztDOxHnD5VjFbjtV4LT/tzlrnfGy/Ut2HvT//YBtj8GoTOn/3QrVlge23GyDEAyE
fi+CMYZvuzUSP7QGUHSPN/M6tfYn3NodneWv1ymllYC2g/l3qoNT4GQmla0sByae
ZA4br6XDR1U36M/QZiKVnXkEj8mItgOmvHEz8IQpCiKroGpfZAx9y0ez6QEXZxNT
HOXVZzgE7bi0ngFKeo9r/mBOWS2Ey0ehP0WzrQC0Q2qhADYktF4Ms81V6eCd7J1A
KiEJFgfBzKnMlp0BG2VTA6n03ujWW+m4iZ5sQpIDLU/4J7KUy8DD22VxSIUjsdTc
OinH2jX7XBmjibSokceS9OTRKOKuImGTwqGvrtIgk8YA4NJlMIoFQFODLjjYV/vz
RKVxanLV68BJaBxJ8sf6b6I0/ShLqrOZ5z+HN23+xtOCdzgDTK+JRP/VBcbqv8tw
/OjeHSqcTGe3dsqx8L7T4VZCh/URxK7wj83sCRNPNzNqk58i4qBVpyr382d2CVd+
TIMe8vang96U7rWe8T5RJqHZVWqni6/qq6OJdixqvq+LJ+u3IPbYCKP8ou3sn7dP
Er2jBSfWza73pd0I0Xxsw7qcEuyDOEeqrd3wv64MxT1cbkGEZt30DqYd9u+RGv0Y
xYsp7tAr1TJggmLEfRNWtxYP4gq9GalqSbijYRidCmiP7JOrYRzdgnxshSOH+3u9
2a/ZP9CBGpZuZs8Vo3UCaCdC1yGbG07pGgNDG/x521Se2hRQvoBVy3yPUMZxDM+f
3zDoUqIeyrwtYbvETGDhXuDTzmLASf65dkZ0soAKkuY+0x9zAno7ZRkqnac89RHM
nH+tu7q9tK+QSwDnq+qczXQECyKcaYt/z5x7L9xLXPZLOZxJljsaYV7qbDlYDMC0
XAYuhiuVQn4WRibybLzTUqUMc1AM2ZJIivH6pdWe74mJQ0ckoXnDxWazd7/odUWQ
jLsDjXRS9RsM7HYKNZrtDbtSyRwlUZTzlbMMotzJ0FLKs+chHr4NnNHAOleH4a5u
endqnslSdaxAJe1vuMFcS8Pta/XsQMiwmuVVAL8B1ZBjWd5mzh1eIMmwV5Sj5cjp
z30paRHJ8OKB4CzH6LNGugvtgIpWrbmZwThU9qM36mzDVG0nSJF8FrYkyN7Hd1aq
rtUYBxI5hYx288wVSdhbFguNo6BEcR/7VauOK9iqn/nkhfZ7VeybSqmNqK5RDmRz
FOnT3mkom92/l7425Rjj92LKVz1XpkpJ+Ty7u3Ht/ZqzwR3ble7p6+GKf8nkW1ks
A1/C4wlJKafoy4gbUFK9VX6u3K90Ll+2ifCVe/afrteAA/0szMpk4/aTVyCjcYMo
O1dm2NcExxiSHH2JEedyZneZ0kyG1JoT+tZW4B6CJziwk1TNQ9RPXBBh7ITBVujN
eebMbmkyEBWjMA7ytSooctES9H5ned4sGpZuV12wNzZtsOuqrXZTXnOulX2x478J
Au+6NGDsxX/ENnZbwC5cWh6I1NzhsvpoINVqgEIIr3AADCY72pwPwUzJLJqxkAfR
KRgVKE/D0Kimxq/6pqdTOcqXYGYB72Xx0CooknMWcc1SlsyKhGYjtnigGH/9+ddz
eMigTofIiKQyD8/E7eLO9q8t9v6nhK3LzMSPgDecAj3EOb8oeDd4BuwYIfxstb/w
1CK6ni/W+Jz9EYEWWJ52403MIuiBaCMSs1hnVf7q42VQh8K/IFIAUlPGpQWq+EWN
KBlPhWb1HNs6eUN03nJA9lzJJxVSyGOTYBJN3OwM1oy6xEU/URcfAmwKzQ4vBV98
rHrcShUgTphv3VNVVdVgG/BSNfSJ9MOewocbKfYIxGeAcNavyJTBroyVpjC39wqG
8rg8cdCi7ucRWpeWRnl09v4dgvFCO86twSFkqjbRIZMn9bbsBPhA/broAthEjZPd
toot7dnjzBQZA60ugfUJAwCAv2ywtVCb4Wrb7mtQrYasJVEMNKlyfT9HsJrbDu2M
CHeFvHeXVXGmeCL1hgNbgcKxkWMO15llR9wZLVaGRe9/GHfXFj3D/zt5llNiPQJ3
BNfp+I+jmNnbkfVhvhjwM3j4xdOsAkiDPuJRZTIhYPsCH2xlEzKgXwsC/17CX/27
/03K3ptAYKvwUd3HU42/o+9eKKdNS9OEda1LMaS8eCE5VDOPK1rtTkUkfnXiiuSD
A+7sgJh7JBwy8B4pqJ7xRs+xHmSh8Mh21s1anm44CwykX38fnvh4kISmih0ey3hm
ZCGGU9YN6sbjuqmj3WFrSvlWU9ugTFezcBgV1pGPA3Eb5X2kHJKuZ9ozm8zMcZVT
sw5prloRfaNfVEeA8cqmXHY88w0gC0KqSdwzIwUC9Pi/+RuE3ymtoTX9x6mweb/P
wLjE8X97T1hnYO5ZSyOva5eTTfnCRqybfyrr0opeZ3ynBHRAF0dqLewCwlhZ10qg
gsI2YmDZC/Lxw3xIi0l6E520vpFwxbueTWUebF47ro3cu3Oetqw5DmxCeMZnIl/o
kR8ZHoV7gyqmqYPdAj1JuU/B2lPNYL5sXUbR4JB/00yCm+AWIrnu9LOJ3ldV6Bsv
BQdsbEAq14c8uoaHG4yP/S1Heo/b2Er1wfZyYc9F2VkFnDSVsvED5MFjG7yd3mvK
p7fwB696g3GdeYoidlW9XzStn/qdRqMHvgGmN0xhXgOAf3J5bveFogfmXdy7ltnB
pxr8+Gew1LR5ydZyIcFk4o1Q10if0IXk0U0mojdnVk/MYaoIjmGYCcWpWNMMSElJ
E8dZizwggE1kR++lL6ltgdnSYpbmTT8qvV2EqCICJBM81rEjJffXR6qTHKQMYQ4U
cWa/PPh6kzAxY46zmbX5dEUmDaD+/820DuOzN98lg35kg2r3OFyf6CppZyydU6oU
736YF8OtIuzO/bVEV1bbyCwMnK225PbJDh+i2U/pu5vpw3Eg78yj1aUru0sNDkwx
AWp3bBC+hZQjmjsj/dP4FxiFIt6XTRbFBSYqnRpimMdC2xMWa9wkhNTNZ1DSqQcZ
zeSoRCN/2EGMPafUNKxsrjsTZq7pwYyaMAF2HtKq8csEpyVw8Zg9T5A1FPCVtpj3
I0brc+J8UnjuxckO8kQG2+aUVvt2Urj+19H5H13XQuPrS3Vk4hUD6xLE7NjnAL7p
xUuesd1CU1u8AWbrMK+b2mSOFc+AZSJhO1U0jRYcX29QSz+bueBGOnyDnkYI7AuK
gZRvsrPPvvWvyk9koCM0ND8U3QsDealuPn5sGJ5InDvXDktx9DjBevaBy3D8Ruil
3RPJsyJFyKBiXDp6DveJmAlUjmDYrQ0CxqZZ/ylNBDvwOr41PSLgZIGWsbxCp4d+
sNf79wJadnLDKBGqfg5fe4FizB5Qh/+BCcQhcZwJYFJloOPZjSonAOuQ4rftHc11
nuCjqLxarHPSRLPl4v1aFdj3QbArZHRJoNOs7Jxh82n7oBvomq42kd1UuxbLpPuT
r4fKN3/+0rVaB9599Br1MysxzmJWWAqnd0Fa1+FaCqB9y2zu5HD6ahxk8mn8CSbm
3NXDWaw+w0bgelZBE2CiflT2+0vjXBFISYqV/pFcDnJXPzThnOvZ2RiKzBCkg+ht
78tZCFhXynjTMYCjIeZYK6fP4nkfHfwYO3Ce9dUMYVodN5pVnhVo1v1XrSq26gZB
85Sa/E+BehKpvxokMmx6GHfFkupXBLqtfXcp2WB71IWIjubONxSoiblkcWifo6uz
pHpHHpzqV6avT3kZ0ktwc2p9HTUZx62Vot8OiAmnSpz6KglMhUTOjW9OuMTh/7zm
I5729mq2gnYIpjqqo0gLy9BSzvO8h4VsES7AmVwscn4CpvTy93ptgiFmTdwlg7i0
ysAlwnmaGMKqv7/FnrDDIW9RUUnSe8NZJqOW03Utc0em1QfAGv1G96soSqSjeVFn
LgEZTOxgege3dJ7l2DstEs/dtWbbMJP64F0KNoeRn5AGoDovMdMfUeOrgxwAr2DX
VT7vBV4RfbrvFeBntGOP4VhqJlqfjSznrea7A2+I0tzeo4/gc4oe3Tc9nuQjG61B
VWC+ipxhlqdJdMxTrhaTVlcbXln6buoEm820LurQJv5r2fWKwqaZfUU33YlW+0sW
DeJp4DLDq4KFf+qF5LZv0UoL+n0BKyTDnazGOAjK1QFxOi2mWohnMSK9+zIg/IJV
BSoUfAyh6YhfKSOMdsaa+t02ErmfevbfYUP0S642d1CN0WG4reskAvYuC4Aaw4sJ
bV6XqUEFluPbCKB/WWylXpzC8N3rsDWWjo3dXk+UZBCHqYsX/4CJ8T6sTpQOaqRQ
euyxErv4AKUAm5gGDS47KLrE2u6w7zfdqYlWYS2gPuTylAcdOYQDAXssAmdualbC
M7VYBP8GmVDcQebmpIrCkOQZqwQYth/gO0BHRzjifMK467GKXYylXc5JjGHyHOTP
FkyrM1lzbf4Vmedt2Yvphjsb8cJ8TbCmtSh+umxn/s1e9KE9JzgIq2zhoZfBySaC
+QvEOQ3nhczzi4q/99Vmj6bxsVMO5d8qmXzQ9TYNTas7ppK9oSRv9XK4QLnkeb79
JitetaHHYBVStQDdIdnnQj9NEQihOl7t0abYTzuoDwMBkm3BYudjcgJ08cNQO5KD
u3oH3m6xp3h20+/hZBGzDoAMUDU/cUGDLFN9tZWx3AZUTJCavDtCSHeaDpR7Phuv
N15mTf1BrAJ45WRMiPD2ixX29bEzDAyfFf+LzXNCMh1dz+OF4ikazcMoKxmN8ree
ty+Ag2zLNXgB6pX9mQqjeYRjGK/6/kK+bAhBP6RZELsrEPC0+HB1m/7yN5nKbvsI
9A80liULSYevMr0fccXDbhavuUl9jqiJsIedkWKVU2uYyYg9Jn2uzMXyXiZhgrhp
yu2vXPAF4AV+uE/V56jz9Ej4GJQZ4D72iGa16Wdj3+NSxQ5NTBRp6N3v2GK1lSgM
gpbY2g/7lt9hLyi2Q4qiv52oSJd5UkfsX9tBJyCV8kt4hPYi5iEGYrmNwHvFsC3U
kgvhrYvJ9ZIEkdC81vj32UzLxrk81InhQ461lU5AM2QB9wzGcj8oOl9KA2UKQQHk
U+1iZmtktQR2N7jYB0CjlILDtUqeJRonqAdMkL1AwDZ13PnZe+8NoGJ2BR8iJ6Ug
cc4mwVwNh7U1sUj8ZV+PJZn7MEtfvIRJ9G6Rrj2KXWJ1S0UU/v5ZmZYWQ7r8F6nT
pm8pTSmxLAMNndn+v090zJ0ScipPomoR6yeJLT+4EEOPGoGe/HkemwIl8c3U9Nkx
P6VitG2W3BYkDr7gPS6YDSsElVdhGNZRatd50NOH8oBKaiCjkMt/Bqe9s9Fr70K3
vKW41OxAfRlWmZV6I1/PPvWgvz+6kkkf/M8ShC6HZBWpI2J4eV9tCX4Lbmb5SbAi
oLf+iEx5QTagCa8PNTZZW7Ta+4SmB/nH6a3Ra+rpV3tAUyIx5v0EVNXqDttMF2HF
7WWFKaqaEqVbbfmWjzw+FDcq+7/ZKiJmFOUprynWXtgCJ/GmCMzyQXmJ/TPx9bwm
45pQesSwcpJkr8aZh4nr7vzRhtAUIRgTY7D7AYQI7oJlGZSJfWp0wPNHz2zx0tVM
QMPvoDNvH0VI+ezcrGlD9MqQSYBg8NCaVPnHAKv5vv0nUZ4OFWPoADspLqgxbFqu
VpKW6eFziHk83g0pUivbfXw2ZeGc3PetFLA8KIpNB8Az4dZ5TruOrLn+LA5+ik3j
o9HfVUZzLqVaes+ii1gTeWNcTH8xHZuQXoC7WZaX7Nu0zffs33bFDQiGmA/tRtUR
gxPgeE8lEGZvifIf+zi6KirtZNrjd84rtVFgBWp3jfrsYL3NdGn730x3W6q6bpEc
HUo66hJTlrcjg9g83pHoWtRL5yi9GUK5G7XgKYwFr6NfleTd4lJqEFxaMgf3hQPE
rw3YOZtQ6s6K+KVxkMTzcoQgTgbl6H125AAQLEhHmPgFnnidoUlsvsZVNavn9NnN
nHmn8Jsuc7/oD9fO1oZIiXbOeCVqX0iVFbPcIN9qzaJFZctRXJ8SUqolwQfmaxAB
ogAjzN8DJlFB7mG1ijtNtqEF1IKlM9ntvoYNwOSyZxgqXjoh5Su28ywFz2mi8sG/
n9C+JZDMjEqWzULEqsiSqddvnNf13/1DUrEWPLua2l9y+xzb0OPcRWBvhpL5FYg9
ipMYe7v664dBTe2bq3/1qmMrzj8aOOAL9R2c6y0uYSutSNVOE05rvFcRXRZWHvEl
Zfn8yEsN+dO+jVPeOgbNA9PoMEc1UO5cdYj4fAwpLM7YCghQFCN27cVdTzICcvRZ
DyDK8wj4+SUW3v4mDQps56neBipQoTXXZTxqndVDfzyekdbDxQmNTA+1yfS6HvKJ
tRbO2slAoxKNJaAwGR/XeooM66a3PW+Lejums801eWC4/Zyu9/wuGA3keprOhQaU
uzaPOxLgSTmgy+3bTGm0cSE46WGzA5YqRuXRKRZO8xL5QpD6NhyR5EGy00+Ds6OO
XFhgXMwm2tRozpgH+QNJR3neUAUrPjjlCeix8X8DqizOfh2VzjM6yHo5vkshmGB/
+0w+CwOKWRHrtpDB9hPECmp90BtKgIQj9HH7z/L1LJ1Rxumdvdr5iyo1k4LaYN9E
CnYyMQg07KkKexR7Zw8gCExttM+Mkrm6VRIAk7spyPU+mmaFkkn4Z5iG+MxIOIM3
LWmawVXZ7/QClMpF5Lw1iGB+tq7/17yABcawxCn2WTE3UlTlp7+jQvOtelZBsdnE
PEFkTGAsoaNgHXSR8kcBFyPC9pBmTZKzwNVHxVLGFbAobbuVHBGMPqg2EUAtI7II
V9Nc3Au49fj/TPEIUUBfXbEmg/i+Cwu97KcW61WBHeUz00o08c9Mi8zvtkBonz4u
I9W1gNy1jP/PrN472owngnDZE2FGv4yl5S5CgygyuKIdboyFM9Fs0j/0JCQ/Tnf/
AWP0VHE827aD1jbRY6oJ+UW6DO7XXmsLBzwIyFQ7O3aXUZxF6Q49I9hXCxact2D/
MS/LOMRZ8PxMTJ78G/dglNenzkLZD6xr2v3WphGl/HbTWHDBboyhfEvluis615U+
u7oia4FQPgj3cpPPiMbIEUNvuU7R/aTERFg0bqnjROd4iFNn+bFJ7j0LU0TIWipv
VGM2f7sR4jJvdx9X9dpBS7/4qCHtJiiEyd/Tq/L4U9BntuSLQA6GGUk12rW7XXqO
NyK5AEWgTeNsNxPYr5BuHGAsBveeID79Amr4Xph6Lb03Pv9NkjU4aCt3VTMyyyAk
t2fUW/vsRKAWsZFmldbnNjBZh0uUp+9fJCHDJjdjbHAcpHPjpUqU+iwhygapvQVx
JnDj100egdW9uA6Jcs2YYqfXFw2YzDNaEBhtM7QGKvLd0Z8d6XALt1jmLjBRUrfD
rMRuwKNxI4voyIn6NHlwsoJ2OOWKyrK9vyag6kXTfqIcsGZFxZr+HkQrwac15bnG
FwYGbctdhGwlb/5IIwWiQegIwf8i0GMihCAFYgcbk5AiHUT6vnjI8swlWvudFPo0
jDjQRPBBnrWfERg0xdOQwFhUY1lgJaFK3grgPdZlniVlvQLv1OtesJdWJxtfLend
OU3qtFxUgHROAJBVqV9hbwTBy1S2LVA08rV/NLMJNdCUpdW2J89bmM5x+xuahU1I
e+fb5D8tlKCk6bc/sowPH0/YFrPt+QowQwFg5zGsW9AgI7Qb6kXi424ckpPSBatW
bsddeHM9fxN9SH1lVh8J0b4e4tfK/urFCMaPPD2qg1Qx5k+Yj8xHgoPEuKsoVEPT
+vL5c4sYyyjWw+Lj7LCHadDGzyEYY/7Pw1URf8BpSb1T5KCexvRwvaSUV8o3Xi4j
c2Bk2ohF4J6CDUGiXscb7SDAXA7HUe0LbdE8ZMytQctQGM/Dv3CM4hb49Y7oqaQ9
tq6ncEc204fz8pg0UmNH5yQ1jr0mcMSgbmJsVpC4pA0Y3cj+fxWQElc+eIH6R4le
tqg3TRijCNNWTKiJatHi8J+J0sVrUT/DjYRKi+Sp8Tjj9+iy8AxgHwh0y9AappJ+
h6Q0e8onJuF8xb/R4j6I8SmWcvEU+gQ3ZN4IrkmDcoMtacFls0hpvJWrUJ/dRz7N
0L+lScYVKvbe0ANJ6uzht5kglh2gyFuIEPHkReQCI6WTfLJ/gn05QeICr51Mv8KN
ZiEmUzfRvkjqoSiMFIkz+3pWIJ61hb/2A34aaGYzYG73dgxDOxdw+OqBI/k0g+Ie
PgXul0/kCdu1vxoM2YpTpde1tUMjkZZy4rK0zdwXh6rMLvU8lGgp9S/sAReiON3b
r1YmKSypU8+yXyiSv7peFwXVs4qGJtu0JTwM+n1Y4fA8O6Ff/8dP5JHh60e8bpq+
It8B2ugWRwLCZquNhSCxR2gnOTC2bvTXsT0WGDhB8OWLExCv+0vJjI7v0+ExA+NB
uOZ9Vr8DVzclAqH+aFJjd2TugCeIpKR/FVHjtz/sXqZftesQTVKHFn6nWfEVXtVc
zLX4h6TV/zO/4iItClkC+30SlPbx5GqWIKiwjdzjReDOj5zXoJkU3ou2cPwOcXjv
guEruyXcZRmrstbGYfbGYTg7EYhpxgyQPBVTD/oOVHhnwyHHRvsRDrq5ilPGgCxy
iDYoqi2JD/Toq2sLx+fVjAubwQ+kimt0TpUmzjOOy//aMS/et0k7dv0tyIvhfSUW
FLoa8y2RoRZCLOWnnkTPPpWybLSRkPM0jjDhE2nyBnnrcYoQvJ7YKrYYr6Ui19f4
r0M0WkxVb52Jxv54Kh755oescx9+fuhiQsPm4AAxFn1YxRPYi28ZmctrHmfUxpXm
/8HVEBwYeuRKIARY7C82oxPn2sd7UIdZkxsR7pDCkEuG9O8ECys9J051EVIo4tnt
tNo+VlIUP8SRORDYiLmJsXuOmOl+JBHyUPvbSjZbCXaOMpX28JvQoe5rIkuBetNK
KdrNjms1Ew/TiW9ejtAWIOAgO+LETvVTH5Y2cxTmKbIqvXpQbipMpmZSu3cOOMKa
2mvR2a/oEJ4EsfT0FtqQcIQPXA4rTdrk28MHU0TwQuC/Etn985cUgsuKlZWF1DE2
y8i36UMApLSGWjwJxoFtMFz+LjGhFmKmltwW0lvT62111C6cCqOFs/5AM0mErgW1
t6dvvRWLKj/+3hzUG6UTInEi6kMw8GD9qSNJK8DT95bD7exBdgv3HukGYII/A6VR
WKREcMx1+CPqAqGi12bSzHr2iVY7NPiUwoBO+S5v7vMp6PsUHVdgIQf5IBhRjDxV
f5g3myBaIwbAoVPad4uvUQBj3jkCKi/LmVz5g+8iRiQg4A3RNWzyYGxH8jMum8hN
kTJdraVg2/d+pFpAOiL5Il4E9GKd+X3DzkAQffp16HDJkbOFAguSafeMDgnYSH2F
ejEfDPXFDllyhVTSDWP1mYv9L7aP0jlKZGIJbZXzdpeK7vRfGT6+hIR7w2FMBT+b
JlAPHsc6FHTn0Zx5kyfIrukeGnTGTMLwYGxqW0+Bv/yfZRwV7kzv0xS/MdWsGNZR
24tqRmmzwAoSrcgmPe+SyQwmUN6xHZuPgS4/We5X7mLztOZymemNEeSt7ayhLzGJ
+MU7DhKt/hA3GS6iejdk7hSMznYmZSGkbcr8mH55xJchcMtAWlMGPUEPexPaBwTg
bJFY6xEb2VEzGrjmwfLZqawoQsEWxScND9dD4cYmAMvgtZH4FWUlprYsFMe9OQp7
F0pHysmCXqMC+9YD4eGh5coKFH1usL7NkheOxLEJYnrOyCEKfuPQ6bYJbdsPt0AX
dLQ+FChRFs/m3KLBfi4Ym6zb5Bo7a8Ly0w7sMaVJIPbnGD/wt1JEMWJB/VYzkSL2
/MzigmDXFL63wOJF+jlfzWGNtGiqf+RMKGGeg7MrYIYLjXwLy1RpOKUS7+KbrjBH
aDJhkLxR8qHnJ8BOoSYsmHtCmxu4UUQfltms9VIVOKVY4G3H59zbf7Rkx4823BiR
zCTjGBV6W5y7UwJsyBgCtI/YhpV+614dlmNG1QAUF+ZByGi/omtOcbyO7SvNvocM
PDnfTPZENXqDOH5bmQ9wbUnUvivjZlm1yJzh1K+jz3XqK+i03fxJktqd91zxH4Ae
p/Q8WqnsbShLMXWKnBbfd4R+dDpX8JGJqQCLbZAb+cqnGhk3xu7jqxoIRz1R78LW
CnVb5ergb7xZe2uo7jah4r27Me0r62LWcqBz3AWdV2JVdcHZagutOURCw3ISt2EG
f1dtZytPsE26ZU6g3+1HPZc8iU98pUdFBcz+Sn30EgJHYd8uJC4m7iO4Qi/llnwu
16q+4+lGWQ4A9HrFuU62uuTMIO4wW5oEW3OYtAgUTG2eLNSWM1bv4sMDuN61pfyc
VblL6PwmNPU+KTBj3AKPhga9WtLOCQBhHbCB04xzXKpBh8S5aSEq1eJn+r+MZ04o
BjKiW9bEKdiOwKt26thXjT+JLhZSxjrgRteguNfTWYIkj6YNRuacg6grkKqpq+Di
A3tq/Xo5OUoCSdYIOSM9HfzjF9t/mxLMFozKbPpwz8UaKZl7ca3Ud6CQcznMvSM6
0SEmqFE6F9h21KVaRbMQrqDzFBOMRMXJ0mpCvM5T7l29sGW2+HwXXpXyFaU4gh3k
2qngI7D+t3RwUm6AxG+e5oy0YghhF5Y+x2JZGHSnfmuy3qbTw1ETXZvt9vQvtP+k
EXO9nLKdxpa9pnr3ptshbnskRFxVu1mF8gbU4pr8eNtkDGdvG3q8MGPWf9DZtChy
paTE9x0z+f8GDFWQvN2bIAARmmdJoT7+xdz3ln/44AfAVNlxGrktqyFJDHvnIxQC
LJBULAE8keDrX9Fc5lytIdSKZafloidQWXbWWev/wzd4SuBHx+6ODEhSVlgvgffP
7kWPtxNsM0OkeK7EWy3ZEKuJpBnogJVuVecBkolHebucojBmyxQTJ8xAbPsdS6Bd
qkSuz2+TYs6I8WYJ/9OOMV3p6TvRpMtyk3s6ZrdaZwyfbR2FIvxxxjKvmseJ1ACC
vL946ahcAHA5Wq/AhZXRmacNMOEfgZ28r0NZ+9jKX5bmHV0aJJgBjuwCKd+inQB3
NKUV+nbRWGRVlzYHRiZyBGtCakP7Jrx6KlKnaJLlivBoWS+nNa8mpoXRqOVJUy/K
fBtq20Q3Ld7+Qc6yV1RJ78JTC62YAKkb8TnR0qYq6XraascIrRHtWWWAQAW2Yr6A
U0RVMz+ILn62F6bSPM0jwDCQGxMKBF06DmSll0jsojStqiNdgBOmr6quCgBh0LN4
1JftEpJgzEBK3PIx11BFMCd8gfA0yIERIm+q+VXGaJBYaMGApzrmPg9ZnfwHUa1z
HaEGc7kcQnT7/YEChk2cHjnRRh/cE9WtFSByU2uCmHYMjdviGWeKhbR0oejvmcg/
s4D2ldYalJhjmgZmKk7ALojaXf7sfKaBvTdnQUvmqNciEiApwEmJcs31xA6krHnT
KdCZCTqNhWDlRORZMnXv13zJlbICgJFCTqtl0ZnPFUsbOZ6e5nb8xt+faLC/c0V9
ll/t3fJ5cw64GXssKlgV7PUnmmYH5fWPz4o1OTh5i4yPOMlD1RyqIE/5ofNangOp
l9PM8GCmmPrsPVKaeTKEdXj5/ViPmQM45rJcYqXXaz19hz2yecYvnxBg+vpaE5wp
NmC3Tob3UmyNAmSZiUssjUSPhb9OQI1Ww3Q7EP3DOtWnHUwYQFk4HFAfbsQEUaWT
DYHlg3tGfdb3hsmXn2NhomQwg3JHxOuyuSQqTQiCFTRxB5jmYHB0XlSepn9pIm45
MsUXXvDB8UL2t0sHNo+cgbrfxkKu1E9QNb0f6IdXLJPi4OxnAyEYcL0nzKUDw+0X
CLDcHmnXjfyCpPRzCkK1BJ6rZBftHdyL1s17CgCpP2pBQKmWzXHnyDVmWQYe+/9z
EyItxrJgRRsltx7eoeWIBP/N2SBI2tZorts/equdKM6HRc6A+syoXRta21vgNxLF
7fGizOmeMokSGjhwkCH9KFXK4RHONme9bl5o9OulemR64GB9BVPJxrt0MyHQcfYg
EHe3mMJOdO2oSHX59A1XEVmZ5J4gM7puMW+s1hALyl55NRnL2UQPcZreOZX2E5wi
8H1TFUjFc7RTHY3DuFox7bnGq8/2LKYSvnaGJtvNEXnHz5+F9+rUWIyoUlejEg3c
4IpEsz6JFKKeoSDXFXwBmA==
`protect END_PROTECTED
