`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sk5VsBqOzsEkb6yYvPOYUm/KYnwMSaPK4nYOVWeNstnx6hgNnZU9qbro8WHZ3wtW
hecPu0cuVfYOE4hkhuAwKR104DNZJcVkp8+syxJ8Qkc7FXHeYEk4KZAzsQJP0u0M
9Q99/5ZC4le785KV+Wb/2HEwXyUObXcSVH+/JiwnsFd1dTilhOakpWTbdVt8xzCh
AmQTW3qX6C2vL5I0jmLFdn7Bat7VJFyP+U636lry+e8x2qppjU/VZt78TDMQSPZe
6gRfDmGoQxSOVOUng0TOlumrJ31AR4pnfBFWcOixdBIk1mZF/k285oRSIClh2R2S
jZ7RUjjdDbzwNcjj31O31ZTqgl7piFEFDF6Ox5RbY+tF3o/w6rLTXwCNtwt6FqAC
EeLiuNNphL5HyBSQEJPm8m8lj2M4g/sZWm3sdxgKxa0ILR0St/+mODVvUAMhUoPw
HdCJxJjdJMuL1w+X0c4aIBRSsdap+FhYTpJXNujb3w/Ud+x76b91q0OPd+0w2kBH
xFoJO3lGNcTpvQv7DHHgTU+glFyl/1hRx0cPYMvNfev2zo5SSlgN5OD00mm2EOu2
`protect END_PROTECTED
