`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JLitLlWWIGOH7deZe5jF5OHpcpIuRYt0f0S3/PuotMAb6KFxRPavApftoOI/QcC
UsXvYKYjLHGV/8n5DQUHaCYR13TD5u0iYvaGfaNdbkrA3972PlS+hCQMfFDArTuf
6c9ubSMRR2i7x6/dSy+sqfW7eQHDKdugE61wP9SSI/phece/yF/ZUM2vmdgYrxrs
kKKs0rjwp212p5jwXuimaIHgaLnAoa6Ee1oVxW5pz38tiqmJ8fX1ZELbMhPYnWji
VvynMQBK83FyUQsjVAb95k1UvuH190PKTDhJDse14HqQGQLZnbKDeg3AmeieZODl
NV7tmOJzUsCA2pmA48Y5Ur7ZVNPwfwIMIBiuLDvHz+TjQXgjgEdImmR90wjlCKi3
`protect END_PROTECTED
