`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euTDeXd/ZEDPsAAVsg91dqkyhhQN2DTlanVO6p1WQJzo8i/NBsTN3TbigCI5b3lt
ffft7uWdXgYLyks+68AUubVBy+XAg346UGo+u0zxrlZ013ruJhfRkQnSWZFaViSV
dga2WIDGUOWGfuEf+39fuRtYIRrlp/OL0EXUQ8zn2fVvU8SDG2TJMG3vYg6ex2ih
SELWQPqoie66wTaXA9oF9GN/FTnLhX3FDG2furMyVZ6ODHom6x0tqHORe3ZI79cw
DNxugJYVejq6lVhBSwt1qDDA+AXtASSEnBw4xs5HuyOyKMtwuq8fOgqEapl0mToo
y5OKwmFFxWQ78Ah3Lgd4kRLIr0eHBYJ0FwD5HdmZn/bK+vM0JnLWiGgOymxIUQSt
vr48iipPnxaLrd+ojQavFzdHPkwbsnSugy/XB5iz8M86738385vX0UNJC6LQHS4E
SayTT3YUFiH08izZw/httZ/KcpG6rzjDtuZ6k0Mpi8uWd7DBk8/yzmF0nEQCDtXJ
+3k1Dn+Ntx+J8S40zrQF3iSq2TpHNOyqj5hilgltAEte71a5Awy6jnbp4Eu20IqX
v1HpAM5TW8jySxNSLjzFrFtBdiaYrfS3x2jDQK1h+rVQSZ0om6WBUysTDABMyB7d
OWO90ghGXLqf5R109otb+Ns/paAiqwEso0dI89UBerT6XD1JX0RH50GD9gIMFuZd
qydGpRORG3TM/akd2YiUrEXPDg0jP1Bik/qnepvcwAy4RB1asE13LSTQRrCg/hga
WPouERPpij6SevMiHB3e8RsUK9NmAj1/eSE0Q/7cUS+3gaYX0wTT0zGL6Cp3VsRa
vr/d/ddh/t05DhBS3mtoh0WABBzXBSP29OTfRP0KkdptEbc2hO+TExW7qCLCqgd0
8RVhBxQiEo6gTvM2lg6PlyhWHJYWfwACWyexgzuHvIV9v1AcpY6+HBk8tsf47x5j
afN/ztQWNT2VbVifAQyT+dBJgbWE349FHv8/FegUAJBHWzad3kztYkIQVpMalhLo
cA4qZAkezw25wm+o8YU4OP1CCuX1uHfaCLW9eDhq4LNbki/5MIJScrJvPYAgQvjy
7JpwmgckfCSgwn05rJ3Iukm6xissd57u56FVbTF/TAMmoM7qaTBmk24LIoBr9kAD
MECHmAsWODtjEZsZMmc8bWsCo08ijTz1Y0Rgtwmdo13O0+2QGc4eY0bRusdOH5pt
2QoEL02p1Ohqx4Wlunj6Pe3EZV0a0/gz6EWZvtFsk4gKPdyONSAv68TlFkuIF6zF
YLOWkEtq6FcLKAlipDRSXzZT0qv0uK3DEuXzAS3NkqFbXYeI6JBa5c33n3VFOkux
5YGkaO6KY3pG9FUxplKCvYPYEO06B18Tl4C2nSL3Klt3ehKEwm816tYy+hxsTCND
gtIbOzTS7QqTOQagJgdhNL6LbwYiMJ23DYZPDTqNs+zuni/mcWzeoncSHkFw4+4U
oL/+sg89ksOtT+qsnMdPCedO1OtY//Q/iHBCAFmOBlVfMplZriVQhIhYm4K56qLB
u+wECloKUv78Lg/bohh5x5svxAXaiRp4T7iYcbbZevtxeYxkuZhs84WKzBVXWHj+
QA7Q616R8VFkOhazZ9Oe14vtUH7vIG3fIqpv69MSrSYCMRdQIgYxXbYLMHd6tZnQ
AB/QiXJoINAjeqj8BHS5DNXMIoUNTYvAB1zswJ17nEdtsAOT9tzO7rKagde/uCgo
V4LYripddAmLI+iVJruvpXuJ0LgaS+/XI7C0iIeXHb3PUt4gzi3+mdFnM6LG2+St
vMESnroJDjeOBmeDpOVqDNiY2nhwcBSc/HHlt/sRbHhG2T45ch0yTk18UJPAbjg5
XGW7QpFFa68tKwtud92JT7Jf5LAQbex72R49dHGd1SlyUfTk5Jv1U/OTZeeTd9vp
s8g7YA3Mc97+ObbTPpnOcWZ9pu0DOY2YEriziXhKUKe9I0J9OC6PFovIoCcZ3l9U
4TVVfYOJmKvxtoizsWYFTg5KOFPTlrnJ6wXOo2tt3q0bwg5foAkgK4GV/2Dw5vE1
qhLymshlovEO+TIkTEjITYsTDENrg98fmzQUU90HhKqER9DOK8E/nt1o0B3DZvzO
7CCaKjk6eEH2QS70mYsuLBOSeXfyLlC2KQQR7NSpgL30p1sb6ut+F3rUmDkvak/K
biKQPJcqKq1HcRRslgEEzbxYfcYy5BVI+hKMJKE4+HyS+u7fnCnvr7zXVmoeWMIl
2xxO6PrfuIrfSqk0ObFtfWW8MfWAN14xBlLe7Q/bo9xRlQpoPcnmQ2HJ8XBSx8uP
cxXDlIRTE9++wRd8ahgLXsxcy3cjP6ILPQLSjgWaOxknDLLk0AhylMeKZ8mwhEO3
d7ugafhO9ApgLnrhcAL5UFzf0Q6hscYsfXmzfrSdAECoYXcapAyLOA3gn4FfG3k8
RkbvvMWICDKKz8LLWrfvfqmw0GqzE5/TSuFaexCVe8l7+GVkaQb2Gbke/pKIaYC6
WGhKGfTOqObpLt0Z2wWvcFWetotynaS760c+yNZP1Y8H2Hjxni5cHxHdmandq85C
v8cg9GZ78//O/VDrJB09r12jOA3BIOzAmTbiJDpshWw6o7bzfP/MidSPXC4cQIPh
wNENwbSqnCcd357SkNvkNIaY8GFAdfdXAMW1eI69vvR8fNJp1unnPeVSmsaQvzz7
EJKMr0NG9UiBoqe+XNjTXTVy2Y8uI26kqA6TN33Bi6Q3im280CN/QT3ICZ7w3aa9
8eMFBZtY3dBAy+8fItO4s67n/S4vYBS7MYLb5SLVV9+KKJCLWXTbpUWZCOGYbxcN
lSKmKuV9XJlfSyzf2/bW6g==
`protect END_PROTECTED
