`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ip/XBooF+meGyYYyVqg/WNyi8E2Ip3DvkMaJZTa7OllyLvshQDVp+yA81eTHMgAF
Rr7uKC27C/u0QumiQSzpo/7qC8KIO3u+GvNrxwtGHlRyeiGPuDYnPvGliYaOIssW
64HQ70hzY3Mmy7O1Zkr0o5l+7R/47QVVREvcy+3xPGihrbVOWUh3j1dRlne7felY
Ou7t5AWwbMXDMtkTS1GgA44BuiYHr3rU+nJNjjZ1j3wNXWLLWJ7PAqjTpCxZbxRA
rZSw/jmmW0RmRx0bbHwQWAN3qKQLp7tsBgiT+OQGodQUHaCNcTT4PbHjlzlYg0oz
TC3fSV4ZMaTf8XQF04WV/XkxBx4dFYH3xELVtifzbxqphIZx5mdWhhq9njPF5Saj
`protect END_PROTECTED
