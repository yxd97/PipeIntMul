`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y61GacWAudNEw1GT6yxl9hjCyWu915nUwH6n7teqiTIVh/GR816M0LYkeosNsEam
lu5h6q/lFlHpXFVq4zvW84s8LFwzjJKDOHl+6qha6IowD/uyApiHDhBxSo51XwsV
rhuf4r+3EH8+axRPUNUcFdwpoYBhDyOMc1phSHkU6fawz3cOlt8wi/Kyay7wABcY
h+ib4w6Uji+h4YyvRcMCcE8DVCHQ9l6LgFh//+eFdbWsKLhRC3OplNnfZwZUAjSg
ykl5MljTMnvHIB2oyY1X/4i0pvwqgtTPxAQvBSOY4RngnGKRZd83A/MQF/WU2EGj
YFMR7bbxKWAz3ugfc5qMnWFEa/+ki9APlNPAVKtLsUW99HC59EvZ5FIP4eRBwqhw
hIlBbRRQhgfVEaPKGCmfY3q8HxSPGo1jWd8aAXFLMnKivB6f34vwPEOdyU3ADg/M
/AxqbS69cIL3YgnjjE+bAAzU42DA2tEIVHTGUScvrAdHnsa/biIicwcNur9A9Y9X
0OXHmqg/64w5ismV8rWKhS/Cz+Jsi7QWjmC8f8ZdMip0iZ0rn+VnXF+8KQi8EPTu
sRZQpajldAYTHC55eaIt/uID6Lqw5h7wov/VlfoI1mTXUEyl9LYg96ZNnfRlHqEE
MT7Th6cTSZ7rX6/9dDSTnTiCdIjMI0Kv/rf371HoHiDp1aNUWqJNQ7LoKtFxU0kO
2Dl74h+Ry0DyrI2XsduCKndQgUpg2iY4Worpgnnix5bYzIn7ztmTAi+/w1K//l0n
sMGEfI9o2Q512kAhnNSV6SqXDYfb8uC/0yPxyqKDNXUZ2P5YDWs9OtwLtgiBWyfS
jlNZ641B1Iz8Z9aZrFSYKg+VTUK3TfmiDMrqzK3ofVpw/oiPo/ME1yG2G7chuLOo
8zeokjXHIF6/2OsRLnAYbt5xeqXZCmmEYn3l7go9PhLR5XIynDhgDwXIjSnav2Uu
oMLktFS4wRCHnR8exZXaasxGMOxCdJIYK4Xq8OceS1adtv4QzAgjDzY5YT/GOIDW
NPBlOd9L9YVUIXqz9c5be5T0I3SCNY8cZmfl2mLiOw3c3E/7VeJl51DRTk2filAy
OZh51jbWRzMaKKVoHdpE7g==
`protect END_PROTECTED
