`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7s37oSKG7L4tDU4bJs7KqoXc/AxFyMN83lF1ZEOj3ySos5oH1YK3qDaG7fMUzFvV
Bql/P9R+FwFFC+c+pfTk523BqFSlKc6I5qcdCAReAfoadmBcyGYFxQ/W38f7w0Z2
5ZTji7IG28NWckRwpYGb+zOFgVDNN2dRZWsteQ06jgYucYnEsrTNC1jJfRR95ygS
WAMnhPRnNwxyGUOHBYqgAZ3Vo8eeqciIAAz5Bbk8zj4uoIbvzdr9Fi5fgl8XxazY
vTlKpjmZ/TWVzCnlf19ldBqE/mA9jD0zZN2OcPdyhrEGe9Y5gxfsPbNIwgg04Uu1
+O8EFfOxz7oH8XT5NaQBIeE577sT4B2IzGLsVfEVwombGnPDg5GdIWFLI+jjlHII
CZVuT34OWbiXm8cStlsnDHNM98FEm6h4DgsuYa83CszhaqqlabAXlDKQNuj8IA+2
7DPX1uAK61/bVRBBkpUWX/BEluOjIUMZMboVi5Qp4mkqvDSF+0GawJY1KtX8cIUi
aCzkXcoikb3PNhz87N22olnWn3kAh1OntdWfE0c3cj0ZKcQl1Q7ctumn3Lvjganq
+VX31FfYv/ew/SpkiJ+Y5kCPpNxlRUZwsA+Ay9C+ehKZcJXB0CkrViB6Zu1D0N0x
UV24FO42LWY0sg/FDsQZ+LIG8fchskVXnIy2xRQWg2mhFwp21lr10kBMc2dLdzvZ
V6Rv75/37iSnLVjF06s6tRPs7HYfkRm1zY6st6dihRSoG6o8ch+bz3MZ71co5DtS
UhBXk6Ekl24B9hp5I8Ex2PvXLeqQwOTfBIQN+B6oqiIIDZJNUMngeCL3HuNdnSvT
8D73bMgqDwdOr7An7bUZ5TC0kITzVIok3CL7dZ7Ryq3Hn9qsi2lKjRNNuizy8LFk
`protect END_PROTECTED
