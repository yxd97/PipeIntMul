`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PvFE6XMg8Fl3jogDxf4D57a6N1QOer+umKHTIWuNLi9xWLelje7ZRX9vti4OYZnS
cOWGl7MWu6BatFFFGI2kOFC0q6nHu6m+SSmxar2iDWkwT1DswlGHT6LcSA2MpYZL
zUiFh3sfG59atgSce/3xGosZpvYD6FKAQUzEKBBn86NgzaAOYhbYa/++RNC5Fz6g
SNIzFiTnf7P1nYjWknbnBWznByDRrUyg+aoyRxSFpAGPRzVlra2YkJRtUBtf0fsV
cpbkXC2tF56v/FCUTVSSGXFag11xriCccUs3IE7JDxjBqIwKApZOXuCdjTLkaweP
CNsQV+8ATVJHasvo17zmHDCszt6ogcMO0PpqMQnxRzN5nbIIHsFaUoQvcSKgQUZi
wihhmBd2kUfML75wFszMEAXEXD9g6rueGKpIvn1BdOdUcOTQT2TDYzOugfZTYrjU
EMlqy5mbC4vdv+5jQPcP7n4tclXX0N6RBznvIh42x1LKmmKEoUeO8AskRq3GrJ0n
+hVNYGOqG5s5ntEG9MVhtoKNPuxklUPdp2v+wR1Z953RCl0EaPfi/GwRi9h8u63m
F3ap/0cdGSxxla+YGuZi/AmQvtZ8OrF2dxdC31tJi/vy6lJOs+CpRJdDwdc1QPHZ
rRETP4FzLRTUQnq6j52IXwFLD2Tz3l2Gy+Ni34gpWEMO5HZlZZfBNuC4txJpd1wY
MgRAEaVSw4ynRSljq4Am1OKTTIOFn24XqEO3J//A2HIkkUU7kG8jY6cKvYbDjbr/
IWRwlNKcTQ9aMO7iwmrrQ1iwKuG18nvVF9n2HV9rKuO2Q32Dp7IyJ3mKj/jFrYY6
JsalxsWAcZ8vG5q/sxZiWIbzaH44+ut7rqumuPosi757cpM365ygADdwS9B9UXoa
KhUYsBRR1q3NcHUl6olHmsw3yikRO0db7Q+y2ue7i2pmUHWOL3iWh65zkpGMwudG
dPSsZOvQgX7Tlm3Q2HpECLVE42IvY7MkI83DVj0TFq6R+Lzfd3vI1vMERVfcVSoX
oqm1Sm9/eDN2KtIDPfDOnHy7Wd+eOmsF6sH7+Zte39P6AlYwvNb1u+E3CnvK2280
YhEE8M3IoiEyG1XAAkrXhbt+T6BJuWZWQL6JGdrPpnVQ9kZ3rMW5cgGHBGK+Iz72
dAr2qNH1WshQeXOs4+ueISGzAc0I1fFsWarJXhUTEMV5yTXL4ilcOwtO3Cqx/4dq
R6WPLbv0AF80fIfZNoSMvypFWLW6tOfjxkRGoVRjzjUvvSntpVp3zph8lomAiRzR
OpZO2bdfphLy1s+pwe09V7nCukhAxEDpyx2GChCAPJGDDovvhWI/JV4xhsrttry2
l/oyfNkQmLNf5VMfw4FxapemHoERx2YwCJdPPNTckHXiVHqyWAYkfeJlLJLronnB
NoZF3trHOJXXTHgTJSf402eUjg/L43gZf4IGB8Ttku3SvDvhB0iUZTWIkg8e/xbB
9pcN22D3MzhCGSnALx/fan8rgS33GHVBXXUJNCIVR5uhKTWMX49SVX+1DmbsUeXw
XSjMxorDe6qaV0EEBq+vfG9gKrURaUgcuVQGsiwz06FHSoBP9O6FNcaq8S3HZJ0s
YIPeq7HbVFFv5AAqJJqCVMcAeYk966vTpSd8LkhnrtmJMmUU3n2ObePfEZyMDPqs
7GRqM9260nwxnC759KLonbWmiDJr6FkPGrdHy29sfrOwfetT4rQlwznGUZNdwi9i
LQZovBgY751Qe+wylMPhmPZemoDqlMjGTZw/11QORro+LrnrPZhJrBYnU2DQTnFc
p7lu2VeS++sItDZp2LruOaMFJM58o8FsMUxZkWX92I+UbPSyvXS5VgEhDh5daMjq
P5pyJrLP/u1YHmoGh//gbJBoBseqRF0hgY01yaa0+Odq690vooV8lZyPnktZBKJ/
RhM3iqZZMOEaZDcj6WPrROcKBMHhMT3mRc6vJjnA7wsu5rXRdx9drdV74ufzFDJ8
3sMnHc0KVLy9VSlqaPgoLDpRvsSfOzWoKj1dMooN+Q3n3xWJKOfTsREX1quku4dX
NU1aEPNShA0DpH3rZbNFWi3G69Hi717dm6GrpHQF/0bosOA8TdUBgRfwqA/MHjsD
zhujjPUJyUYYm8JxQytZN+tPqenapzDXsVqnv0qXy5lJsrtCcbVNjz8XwpX7AVOt
nHHNvYQl0f6beDNB6dV+RPK4KvD24b4VeXwBtDR4DcuAnj4P09i+OQOWh1D1IXnt
+McHxPXkur2Ln7GZ8MyMTwAbJZz0UYM/JqLo1P4+q676rlMsOaUEOE3XN+LamByY
J3OO8MVTEAPl7HqhmDASJKUTIRtf675sjXD6WXu9NAza4awutgwnNTHjX+Sojyj+
MLpiiR2yrmGa1fbb0d2aRfXxrDjz2UDYjDkIhYGmQtVNfOlio0eCItrlJ4F3biii
xl3rd3HUntZ1WegD1JoNiVB4o8TV1SUFClpiTyJ0eT+wKR4MR6E+RPWXwCFqFYnc
dCIJJp2opC1z+qdniRGPsSfMvtg/zeZbjYz1H0YbucqRNDRTkGC/17n/LRh7uHuD
yYpPLhPTryGL3LWQyY7Mjy6zUQsSpJHnYvWtjtS5MnclieqZKy9L5OaxoCJqZp1A
CuTdYHVDeepH/9/f3h1DuOfHRoocwvGgSNcCXD5RRCxw6Gd3csyBFUHKY/wWLU6a
Qq4E80wJR2dp5F+vVEv4E0kHxXzC/5Vz36hudRk/sgRHDE+seMdH9q7kJkVsB30i
7lhfxAhp8X4vjInFNYwYdn6J/l4ZpwiEjRrnRa37GlsCud6Q/Qfi7os2xTatOyby
//tzeR1BIwDjpY3UzMe0YZ4ua16j/xgZqIot3+/HzJTdZ52DerUXjq9op0LxRWG2
Yfcq7ZYa1EaHMG638ubc1M8vNIxVTFZVwtranB5LGCoOCAMZ36KpzAkMM2aKPt+M
yJ1R9lDyL5wY3XZaBrbI+z/iVqgd0dIzfEAioYOFBoHPRs7RvFNXEWRZYURpTwkm
kCR5JXHxXChv0kW/q0XmQ+wlKhlmXiz6/DRuQ0J1LKA=
`protect END_PROTECTED
