`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jf09NoKlFzU7Iardq3wxppLI2yoq5d90tU5i2k7A/2howXoy02KWBqI98/btp7r5
CBWdH6u+Em3RpgiL5nvnYmQDN+ZHHZQov8FoLPN0VzRkkafa/9mMLGQ9oPLDWEiF
Bo6xsY/ZC8T1GgOE+qWDu2Nr9T8o9T5o+Ah67bcPUJdiuA35A9Y2W+uWiC5j+Ou8
ZK50VETK+apUBFu/Dp8VIZ/nYiXeHz9LDziOloN+tUC5fxl8/AaWlzK6ikh7WKFu
7fj2hgAaSfJYGOdu73qhJJ9u7NYVhETOScBR/9679FY=
`protect END_PROTECTED
