`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vVQAuXCqZZ7dmCdIhOpxjqZWngt4g4Ng/2SKiduIb+Tq/hrG/b2luiyMFmpykmCc
C+/7yfdb7ykMWyrZO0be+gxYQ0OqeMwFhmdtpfAujg6lvX+fGfqBQqts8WA5yyiW
KxNCPDwn9sgzMTuxN7Sb4kdbPDTsY7Yp/j3lJcn8oO1vCCVh11VWM2UcQT7ZeCVj
MPMibZUtUEJS8AIYjfV2yL2/OJWaro34ZTUi96f0A9Q+HRais1NTrIokhGwdmLOC
0HW/XLOerUkQynjba81X6Q4igQF6JakmELZ2ppUYharZfE7CcrdNm6ka2p+yaOwM
oDD/qz8nfOSGCOWWlreU9fzotzxBNrRfvSmpP9lA5F9MjkP0AltKRfFgtvODMNqw
W8bgeIbCjiE2GUDwZd226g==
`protect END_PROTECTED
