`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLNgU3b0atd6yASfF+Fy2d9xsegt/oXr0iNYu1+WHswMYPzyGxYnmoA1UCGhjrna
Qu7KsFPpBbTLOpFxmhPk6Il2l3FQD78p+iXIctkNWyFcqqtKccz+ncdIn0q0MC8e
aqQWJQlMu6uvEBh/8YKc2nepNk65Hogo6fRpgyiGS8R4oirsedFYhAB2s/RZVnOw
1FlbVNSm0tUZVwEp2/LMMQtUNSVdWeCbwu7zXE7mweGwnEIgN/18e+ZgQmCENGkQ
wG4d8d740496Pbk9a+vihc6rOxe8NvyUozqww+yl7FjNEVRpGyikGVbH2s6qW7nw
rTHuptrVrh0bQQ6IuOxFsBcsNUD0mV/EjD2y1k6RSm1enYUF+yqlH6/qOyyEwomZ
O+NEL0XliVFnrk1a+fNeU0i3gm5MSb93ZKgpQBvk//1AJ7BkP3C3TsyMtYvo7RvR
rjLsPHnsTEfAR42H9PxmyoFFoFzPdl6skG3GWDya12ibFaNYNUkwQ0YRKaApIbC4
RQwfYqwoYKKY1AICiYKachcxQS2RcUj28Y1tQYEkzax8H+GVEv0Z48HkCqPiHoxR
VALKmyze1gJ4SZNliB8BJ4JbRSi2hGXE9NZ5AFc4fIBWLscpYaPJRkVQQjcr8tBE
xhiEuekh55VHvp0fyLijSEVRSFzEL7BjDo+w+BBh6vpZmKCVB8N1lbYiazPX7v2W
nBoan6P6egJmbB7W9/jIV3f+hA5xRTvx34h6QQEHAdz8OTJgEhAN6l0tawHGFuEW
UzZ8EY8KgZPy739CFk5yur8CeU6o/Hk6s6uTTOCjDabFMimjl/imfQPG/4bXf0NL
aD/l4KmyLzpBpOiej34yyw==
`protect END_PROTECTED
