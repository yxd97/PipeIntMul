`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1v/XqYrBoBynG7B+JvMilNbz8yv3B9uyLmUTzAUJqm5SngzYQG3WcRNlZ/M+kFhT
JC/DPx2ZdEpyee3dbb84cY35l/g3S7okWpuzp2IDB5xQGXVsqdYIv/rCEqlX406T
tlR+tOa63BQwixymOQjYzQyu8qh73b9YRm6LpMKuYSWC+MA45YPk/JKxJVXsvyr9
ym8bnrgP/QCxpsZp2f8TPN1+BSO+QQ2SccaUtXPSuX5sRQo2kef+7mKKM+kwu82E
rA8fkogfWtSQS7satBqirzIjvldOKervRdaiEMjJVlZVGWqa8ycKlDO4NjcVGwFB
Xic+S0V349W7sHM1qbsffkssxwd+4ypfQ8UB2fbWZs72HXUOFADUEDIiHlLav5NL
KUwhPNke+H3InPv1XEm+wyuPQK1b3Va/jzQPNSQ796H217VgE6eUge7SbXhfZO5K
bnbuIXOdWKt9XHQAG1Q5Ux2ZVEXOuNoaVxUOrmMeDi1taZKeKFohMLJjVJPSnG/z
h4ZVpz5HiJ0f8ThKUEJXAne52eNt810tfkTBUtpXh23CXwcxIJe+LS9EhPSO6UCx
X2Tyd+oay2+JIX3T+7jkr3Snxl3glcsCrVv1xMjOS0fIHq+pt3o+zQa/3tz0pBnV
/N+4bx0XFt1ayxwbEObZ7AgaVIZCBKGEiWaWaZUZgsm0F7iKA05DpS6OfmCHLezf
fSgKH35AnKyNpuCyvAz21rWHKgEE/LPdHdd0POyBF8HVqupLrYGozTb97kYohb2v
59uthSEjOWCUDGXEF1Uls2kXrv8cXFtsTrQXl886tXmGpoB+AdtanI6uDLf/EOAI
DzrzR20fydR3y3zp0M5ldZCMvCcTrINxWVVOM/wizRY72po6djNbNwXUnGrHbDu1
1fppNQqJgd+CvIj9OYr4xpyBLAGu3Axx+Y+vl6VSONVyD+F4mRuiJkC1EUL8oDvb
UGcmXytK/E0XLUa0gWIBZaNhpfI6k9/nbhhMJuFNUhTnO43IAd+GIomhaX8i2sgu
9LmsirGfB3FUHS39nUo4LrTjO3Bs9HNm3sqjxjMIUFR/2vrNDi2Mk0YyymvjX7kV
5XJz58wb4g7aygQeo4smpfyUYMulk9s6JFfqDJNZU6bPDBql+GikDRH7THryeWBp
/RDM59A7jwu8ilGz4VdtrVOcRPoQ4PmCnBfp0K6XPbnDyL3XrPpqP0uSUb2wnEvA
SPOswObCQcIAMtC+4wF5JaunvmMHe9+sXeKpjrADJcrQs6suoFfhonFWqKGKZYcP
luEG825pl7SZFso15WSptHawMg62qN+GM+2UxJBne8ouTM6MA0QfqNat6EJ7gYO5
oU34bO624t0ngcSKOrjw9PJ5jIR70H5KcmPGw7d3nFjjQrVhTngrgGj0DqrNoGh2
BUWiQ29VbJyxc7T8O7bJZOT9FL3hn6WOIKvwgFNWV+dDDpj+vY81PAfvg6EVufCU
PgPqScrimsU7fqq0YpcP7UfiP/qa49NvSPCy6tAXhNJM8HET1BoLhkzrlgkSipfK
AC70KFP2SE1RsDaz1+hojcYRc9oQgz5zxyaeZGkLe78KKn/38H7eUMh4nqimTgTn
FnVu9iTLMMcWawSCnNVac6RVpdz0s/NpbhzReYruH66Rkgbmfgzl4KK4spVKb41k
y7la0ktz7xn0y8G49z+uusTFAtdgdy14TYvUXfk2o+UgJyRskcfvLPDGvsjSHpcI
SxXzhC0N92mVAT1vu1w1jSDJyg3vgMi2ffjDa4LEUQB5kIjygXeDI2XefZcVf7uT
o3fiumAZSem2DKpYEQQv88u+1IlcVk7UCvn+PStLWilw29ccaiCLx35uCbGLp7ZW
yzpseHw+aoHKmrSjwyIUdvVIzIhDTL/hdEUMxh8aJqnx4otaI4haSzhfgnD/iy7w
HxZr4ZpAQfqN2hKpbKXAEQl6pN9ngnBRUckeX7iTIjcaqPL17dJ0pLL4YwbciBnt
+SYgx8lX7QP9jcL5p18iaD7HKqO9vF4Yws+qzwYiv+eacoyUkDZr0N37R3OClCAl
tFCj/hHmlO+L5Nkfr9o8AiYUPFbdYZ+/gnPljJC5l/DTVOf9enJrz5ByIFQ+1QPN
bKsbwcqp2xVxzzTBC8K/yiESyeLT8nCsEDkCPH8nHPgd/H76GvgrRJ1xphK+DCZS
jw42ZcucQ6e6Jwg59CjL2mwWQkV+ZUWgWbe/wBe4hhNH/dRN3rJUoVzYe+dY4HMM
rsiOlEV7KpH4db3o53bQf/OtXLRk7Fn36BIvIUZdy+YhMJKBqZ+mds1ABTH4yTO9
3Y/cRqteg2fM4VwtpdUbgyTbo0/50UYIEBBZX67AdprOwtVx8SthasbtTI5wYKkz
0m5vaPmAbqH5KK6lU3g2U6bSRyPGs02Am6JQs75lOpK2Ch8WzYMSVw44lW9OS/h/
7BMvNNfkVdT1a0OYh0Lv8UzzqA8fiL+qCPtos/NkPsmC9ektPX7KiIMa8jAJ+oUq
1TUm/OjX7Ht7kdD9YfQ/IdVm/UpzvrJYN+w0YByZs1P9UlALZk0ThAG8idmRSZvv
h5vuTexJPtoWjJaTx7vLOczemWs/aDdWgnqvN1LWOp6UitwZ0Fu8vuhIN1oeBNuA
KXLhECew8knQ2xgeZ8GMtVDWldeuP1IymlgboCJdrNAg9sH0WO1JIAzQ9cmUYldA
T9kolk8I0blV6Y8olVwhUPhUDS/tgeXVet+xDWMj1ccKumxo0ICyYyfjDY9Rth9S
27sLFc+qD7xcaFPanwC46Os2xWymvOmZ31qPPfa8uxqA/fv6m4Pm8ewvCmKeN02F
47c2TyhBJPNWzxV9XSv+JaCV/xhe3nQKqK/8Y2zmag7eHB91kamqwyMJHcrVBk69
44hp/eYvsTFXBYr+FENIaIXRQOUEP3bsCQb0eWJsd7JS2UCDP9fls1CkfZVxtaD1
mTY/7sw/aFbfNAZG6cAq5hsywtekveTl0h2y5IAyjSr3sDLJTmfeAUhLEI0XQNf1
4uiynkRniP9NjBZG/S5UTlqkEWd9KxpNydlEw01NTnIvkdZ4/hsolF/5GGzyzoWt
rKbExkt3idLnPHKEEfifyZYXIeRxT2A1bLAoEqRY5WzTDH7kVwhE/8m/e7pkJXys
jErH9yMBBhK11mDxAzeaOw==
`protect END_PROTECTED
