`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Te/lENQyGyMwbf25W7VeM1aWeG5ces92nHhV8jkwLfFZTY8NXFQHdHsETcxGv1LW
JfZP+Mdys7pvEk8BMWtsxE+uEVQE1UF2xy+PlfCWvEi9IQbnQbtCainKXLyiFADK
UUE3zf0Nva83WNOa96fJ3JzqztM/+EFBeg1BRlozVHKIPy/0+3pOWls7nyMowL3p
2h1m4Vm/BmEKTCoEJT499ToCG/JamiHaebmqfaaH+e6bnpAGo/D8w7xgl106Wqce
Ay630/Y2f1PnYInh5lHAJRUrZAYYUX89cI3H8vYKXAOSGbQovHyggA+vWgEYtKQQ
i+NUoB10+MQAu1snc+R8uvm9p86ZPb6uHXFBTbh42iYcjhqhiHlyRQv5n5/Qdzhv
g4jBIFebQzjzuI+ZOwDP0r2JP9XTMRvygtS0nFUGS9R191a2WsXSNCODYizqoUYK
a7rAtZzV2aNNfltP/NL/jW7mDAAFl66DE37NOc9hIJstHMJMVSHdHlclCGY7TU3H
/pM155AkMqbOTfksfh3r+SaV6/xF8MHicl7zNFGENjH8MrqCt9yCHnEOxxd8v3HJ
TwyThtpjQmqSsoUBXxGU23SKfuVCUKh61uwEqn02GivkDgbpey7gYeo4P/19W6cv
3qvPVOgAQwK1q6CkOYc1ouRFP+RUKo2fYVSRn3owFySL41QkMsMnwKfY2vfhLJwe
4K2gaa4xVv4vMdITt98FZEpPR5SyPU/24ODs54AFm9KzrJQmm+kxzMH2bf4cI7/N
/NdR/NPxmF2KyeEZNny01OTckYF4FB2POYC4yEBZnOROO5KQm/Siq0Igt7CNf01j
RuKm5FMoA5GKuWwEp8EMsyudGs2lNF3D7aXIb5K+VNnNFJOWSZxdHz2vhuaBu07t
8xmIkZFnaPTBytne7LijR/ChaWVQ+hhpM9zPESmcX7QGNB0lAq1PCTMATLbvyqkY
qeRljQLBVllS3dGz9k8qCouCH0i6mbLLdIm3m1wOSLRWjhPFarL/XFfe9A/n7zw8
PCHgz1f6ljCDOxKIgDEUuMO8BrjZFDINTJ071Mj8e+lsc0cqbuaeXsi3RI7beYVs
mqB7Ob/Mn5S5M8G00xjL7sQ1lJPoRHoQnVLpYh917UPaXzWPPxyyOsXOgdzbmM/j
aQTrmbIjIrT1D675NX0GZjfYXsMgpgyWo+ZLnvGHdsalMUOKRcEn9Na2wSloRK4h
MZiIBDi+GWz4ly65CX1uzeEEdf8zXdYQ6R8ldQt9bHrCjyFQaJ/BO+AC/KnESKVL
aWPG6ltFWbGfq3MApVZ3orY033tPXAPLSdBVxh4No74Aa5rkr/IyxdHKqx7ioHnS
RFxRqyaH6JAz+KN3zsFpZJ80xGr5YtN5Y4HeaTPbZRezJPyMqwPG2KpECTH3uggx
3zy2t5WhUBQ+PJAj5uNam1DVimAY5kbwu9WRs18A5+iLZSFLpLc/WpaG2Pj+0/z2
JVbpWB0s7q2J6dIyOAlTBBZp4kHIn0xSk9q+6ivMIVJfjirVjNWJIS0RoRwWfehI
UEya35Ai83EFJKEL+YstYK3CKP5ALor0dZW/6Lg9Pe6O/fKSVvICHDZRDNFtgw4l
dPinUEObqhJ9MSCmzvqR2fUdGxEFYzQolgDmtem1akSDHPY3qlrPa1Urq2LpLbbC
E2FSmWCbUngE/tFKjDIXpWOyvZyxvjv6gk3eTPuA+DOseOw8GoNsUSX9xXMUpj88
9GXWI8LJRtB8AzFvehxxiDRaXo3jDFM2LlN2LzwMXgxWvf2cBNnlxBUin4lNX9mD
bq6/tHxfm3tlnmbYvZXEKPv1DeSpihAXwWDoHgOpV8Reauu9ysaCsmKdRBhYNivu
WXxqLJdv+OA5ET24XKelgn8Des+nfqqnhF+FfelQ7VrLANT6IqqWrzgBCFJTsi/b
5qij6PUyJAfZztywSyeeRgnlCkhTKIXatOf2MNWZqb3nSHMsaUb+EIiiBzlknJTu
rM+4d8CnGK/1GxHPZPwjVGoC1gWubfEMksPNhI28At0lhFdv4anI2YCvTqGuXRWx
DKc0bnoYnexL+GH2Yl08xDnUxRKCyM8dqjUspcTn1BQQu6rrr9FaZ6+D8e1yeP/P
o1rFNo/VX+xXISk3sr9HwqpR/3vYRwjYBCC+6BLsM/iWlRgxwFm8Veqi/RYdjwga
ovQqeZWxZ2hTDGRcXjzuPi3uS/+EwPDCUhZDe1u4zSNGqBrJYGX2JdsUjTtRRx/D
mRabVuofz4zpMdsG9PSnxdtW/NSkg1Dw0xHVqbOuQNOTRZ8+LcIymv0DoTOGh7zj
j4UtWXuWmsUvkPmBIBoY4THzvVRcrU+xUjVEzemJ1lBPlxXIucjXLPmYVzdZqRcp
loALY/7pZ5vJOZTl5cJjlY1r+3u46j5UJY+WwFaGZoF5O6wagLA7pRrNtsA2Vm8f
ppzrBrnWShsYP50SV9WSIH0+f+BEFDGDZ+kbFDSzTUtnvLESp3ApLgWZBTrPGPfT
uCPN85GqLeoGEbvTzcGftz7V72fYHKF5BlGZ5G5AEwOROJcW47ridvijOzEMArn0
H/+JRA9AExnIxUtbxkreffV66u0K4sGGBUfTGkko8z4rRlpZDzvAjrkKj49rEDYk
A75JGLf7EGIlx/S/KhCpymLLIBDEJNpHCw5ETugx3Ec//RcexIsDXebG5WkVo7Yt
I1KayyFtxV5Uaks0a+MAPg34dt1E2aURDoFFVecsoJCMPsJmRNd6ZBqCGhvh3ADf
fPXTUxmSyrD75hyRBKnSRs6UjijnFE2Hg4y4ad0mqm6/Oz0LgnVKoo3L9ymkkNTG
Nm1Zsy/I0RHUK8DS4njtpy6F4Mw6IEJe9kgVWpIjtyH9eE9jAgjf0H8R4tcd4EEg
uLFcJ/LEWEXLEbHZEkuRibetTK1duWsdpZEbymMq/o8by1FmIkqsTOBAJWzvscbT
q4cNeE90XxSYcsHLgZcrRY/ns8tBtEFCyZWfSgm65c2jRliwoOJYQ2z7odRkZDMW
70mBssD61Fw+sOCjgQ7hUjQ3yfYFTvwLqx2ZbTznXpLoOzrflZGsh09/IJR3Q455
/gGhA8VtEKZlIZBSfc5C9OYUpculW3SoNgoMsWSb2tg6LvlRcdDkZ/qxN6VyMiZH
oxDBrLMtFTOktG6GPGGH2vGLnYp3EoEDaFOVFGd/g1ggITPeZNTGhqyYYG6n4MPc
WtNDNQKYYymY9nqaaYS4jDU+lBEAhgJM/m7Cm5B6yTWU/9bTrvqC2sGY7wsaTuvv
DDo87/Hzk7kNsPnmY/XxE+wvwonLuzCN4XvwXJGEWDjpUpgl4ny39IsOnPgFw6Ws
Xh2men6gQPmWzwrF4+s2ZuMzBrvmMKQA3zUU3kyIKOobndl7tgMKHQ/6sGAExqsL
ZIoDTSeHEiVTHkmyB++/C1DimB5lt8hbFXZMHrqMy2uzam3dZTj/KD48tryc5ixK
GxohHZnhCLA2iE6HxsmbxszSvLvbxx32A03aM2c680/rMPUD9/VkU4PFo/cZrxKO
yf4UkI59YSfp3Tjdgrgs1wOy5XVixTBuAczCAe0T82jB+jZ9fbaw/dm5Rf3KN4oN
r94mC75UYyVNuuWMF4OWK4vUWLPRSVBGONONDPsgjSsvGfd7k9QJ1/Tiv4HABnzQ
SFhDqTJccX5CN/Iwaiqfe8bPud3puYWIwBSOnVSiO5vNA0D0Ue1ydp2G+kY/8r6q
fdGX7b3x1jUFqwydOiXC9sgvPkPSbp6Ao9SRdNdpW9gcWV/HisPrKpWIdTlFSkg3
9bXuZZAO6XN22DDhxdm6WKL4w8QrGbt2zmLAyXZOJQMEDjnLHdy6jJUuiwT2h6cF
ce0+N2XNyVFZsyVTo+ZlHPQDiEKYWOh76Tx4NmA/Kq9lqfAXV+uWuDnKKM2mvcb3
U2+KXVPfQweYWw3Gc1Jqu2QjUyVZWcgbwpw37F1t7f64RSLT29Nt+4knjb3Qp3yt
jrOmKuM5l5uXs0+69DiIw7VsgF74GzvvEd0RsT04mAYN5Xm/m7MYp0xV1nyJd/3W
j9ZtmWegvM3PwtkMyPtskdPWqpHU9RTnPRnuzKy2GwqlMMEBP5SqiklwePw8xH3f
qwlJVTrl/StqqIWjKgCIPmY9t0YWfivbsOZXAJQ4YOgKZOeWJ4KuY9gNtBkoS9Up
aygdWcb4Teg/XgMv3HR3centCdaM5bQ2gJ5iUINHMMTtc/fWgk71phDq/OIj5OGU
r6MXWr754OcV+svbcCSytgiBHZpohGwY8AJbWnrRe0vOHxoEhRbYogTR7uBywlnF
9uuZ1h+BQsB24G0UHQW3qx9CeKRUOpqP+rNrZqkWJkMHOENsUWwZuz7hnvvTOUIu
3MyYd/ypPbEGJY1Lek3EZ3ftl0RrrWu9YYNTXz7mYagSKY/b0IjDVpztHO0hboZ8
u3LA7XLroEn+FtMYd5FJlVZiAUPYKlNHr8iD+PfoPGUZb60wRosRvmyG/hS/8MMV
WqhTfGrn5MK5NeOFNX8yp3a6LLPRcK8/nGdZIc8R+ayav0hbPHRqF/J6IZG7yii9
rlfoVE1nhmzYcb33yMfB/hJ17AfBufUHr0/n+xG7YgTcrvSZcMiYY/mCn2WmSXMs
HQzDrE5ZwYLluZGmsDCN1kPeahwD04mJZvN00IhY/RCL/rFvD7Ord/GbAPDoHQ+7
Vw8Csz+ru71XmnlExKGRCUVwPYKlgqcrBiHDfTRnhVqBpE11ndJe6rkDbn3qzuIH
/Q1e3wIqKU+ArQ2YjG1aegAqLC2A5D1GG+KCdpobCwCdVLQhZGJkcqI1DVDO78p0
4liV09vzT+37gKGlrWUcPByiA8iUkdo1uip/+8ub2qwf3vj3olM02tz7VXLHQxTq
uCSzSjOuqUQoDmwnSIjjqc4ugZWYgWbgQ0XNpXvZG++fzn7jqHVGOcePHAbydCV5
o5/gnEf583vEtYXK0NHhjRdtLi5qwZpQnL0tRrab1je+pjMAVJ0qcgEQrUKNtgdX
LNpRicTU5DyHP7TdyD7aVbCD6MDzrPlCWni3FdGIQs4tdcrtMmj28PUocBIUuaxx
qP3HrNSUHsDR9L/rWm+Rv0Wmu2CxI2SKgl6L6kfpChSkwlYmdexJFmABZYKHXJS9
J02aWOK38VQzr6IeWIJqhh3Er7yfYlr/x2cTkGl8DHIqDbw0OAnEMRwDAhR0dpxg
SPXdOT2HNzrsaAcjlGrAOWgTNTmio5w/6+ifUq+phnKq9qnGDH8AKbnSv2nXbN/h
GneWgJ4ccFgk6bCMNjGjoCGR0AM0Cfe3P97aqbAn76tOzRDhOCAjK7A4LCUsr78B
uJVvKkowxPOIiO+pyom6uKs5e2dChzs9JYLRxhWCZbf0NuIe9siagdeQpcx2hLJe
zj9Evp7HxVxnFdcZEuaHv23ANFV2hoUdk1cmZ1xF9Gyja7xRMWdrUgozxe3K6Bzo
27DM9XmiBqIFxi3oDayAiUw8JT8ERN0RJKXO4l4m0uT05eBL57z4ZkcX1HPVV12l
WyTCw/0AFd7BMf9y5ricXJb7K+jeurYcU03x42uy17D1lIDy8IDFZuxGaiD+tK8K
l5icr9e2f7VLAFru837tJHzt9BSzHhKUfa8oWiL9QEe7z4viaGyb2GhQbADGQwzF
3GpRtW6rXNSHoT7RdGZ2BaF/tpOOh7TAHCpEY7vAP1RbDwQrd6pZPjRjcLMQtwlG
L3HEOdPyS+10mtPk0lJQILflyarw2lIelC7dMOiK19+NGR8jndTCPOPuzm6ChwCO
GhRxYtXF4JvZBxYOn39fLUgwmFaEqfsjITQABKNONCDynns3GrjjrNcAd0fghS9b
8YuNzmAEfnCcH8G65J7mA/QoglxLePbhZ/DyqPFba/g0ch4e2p9p1+dBeLNIA54n
ISvPASNXpA07gCaxGMYCziMGzyVnw29M3M/+fxuwf9doB8FWVf7uXIJe+JeQXVE6
gDcu4GCi9T+X8T1seOsAJKgp0ClYGgHfg5HyV6VZkAvw181GsXhm1zKhOE2xHorh
gxLzlrKv7TFV0PgPd2YRmjQziw0/aiCtduawM+Ab2nKf1icivNeBdZeHgkjJaZks
0PFs81pbse3w71clJJgU/PDorJARb3gYKKRe9Ls+gpqUzmk0j3t+Dgfjqa+WWARD
Vvzuvmq9Ym6seyCJOq7znWVKSI4daGvSozwS1YgwRLn09eXPAOEqhCMJBz/KkYhN
xUiv/E7DO46JTYB7eY+R3nUjUJVOmTbodgL9JAX069E7E/wI4B5V+IaYIfldpovC
i7ySPRtoUAouXwvvZKtzyKqBoxzEwZxJDV0gDky8qG4ew5/7LmYmbsammGHFyFlp
fsdfFZtX0udgmVS3CTSJJ0zg/hWAEdpv+araxq7HiYtZKymkoSNJ9N/UgHIvJ8tp
as5V4dNgWJY4gxKJftqoEwo/9CKYngtzZlLvBguVRmgOU6YtObN/u77p+m1trvPW
kOaytZuA9g31S5N4kYEeHx/UZs3B/X+J3gsHHesAbUEShSUcDjd5+xpW76Mn6oBt
t5xuEGIZH3+Gx8WFU3oNEMmqjUogJcjXXN+Lj00bbyRr4rWnhz6n/4q3qxTgc9lH
r6Eoz+XjJxJ7YznjIRNkltlVLA8iU/udvluDFsTJ1G7kW2ta/MbIUckOuc7j3lAa
KDd3DyHd+GVtBWzwpb8FcmKRgMGwuHi0vdariuzsRUCI8WAr03+nsmb0vBTiiB1w
uiIIOwsDtYZhDzNadQScHDT/OmOD+pqufbrKFwMTN0GO8XSpG5kfzgO7lIc5LctK
daGEL0+FlbpuxO21GAlFxCFDfU7xBpQ40Yx1CXgPQRnBSjA/U4Mqh3e7FTrd1HSi
Qv9OqCbJd7m4df4u1kQ/jYMz0wFVfydzfWNqU7c7CEsguuba/bcQuhLvarV0P9e1
C/BbqEuh+OAaF2UOw8y26CX0mg/n0wGTVcqFB4kpMzf8G0I5pTi2kwnZVK6pOFPv
UYHrp9i7+1H2K+T4/ns/660gy9w81AFePCsNAqUsSjRkJSvQwnt4KTRN7BByXWQS
ExbK3Bm+9VFBvn6SSbt4YN5bz+WMhfW20OlunNykvQjtOvSWyd73tqKG6JddQmyc
/z6eacsl1iGa7pCN4Rto7i7oaJUVcGJgAani+H7q3Mf4ep7kjbCJsIOKUpSV5y0i
tP5ppsH4Pemp6fdNpKXRJG411eb0V0lrgx3ArESaLYfQ2jNUPb0V6qPENF7Xf0cV
d5yRPIXjkCEVTgDACtQcXSHOpLux9yDb6U8kkR2ktfF8kJKoSYq71cxLTWBq8t8b
xPW2/uTQxckdvzvehaOMFYyOmwkXsyIHWj0ooKBkXvmrlED/vTrpsiMsvdMtqVMB
37YgX6jrXjMK7pNNsTXPqM4rdRABfu7yh3ZzKhE/+Z4IlCWteh3MGBksAXySy5uZ
TZyk49W2FMV3R2qjjo7RHSuRJ8ilEOXDZUUpKNbRMQvSOu89WvmbZBTiD9f0NhJy
6OpfVpcFWk+So8c/F213cdhDi4sjnNnSTkg8px2xzZTGQWqr8GeNvFRgOVzoI/26
bWvTXj+/RFPeVebc3PyFp31tEjcA8SkDHv/fLYB6+03THABFXuLBULxwSGojZYxI
4ulJHueFaA7eTVbNh7V2hCgYRSsbEHoqsuek6/XhSZjO3sXd6QLBcnzdmxqHsZrw
QfkO0WOfOw5jeszEQ+OWdCOrfxS7GGBk8fCT254VOGy1z8tdffJdDuRgLG3hrump
0Z5uGlz5heCbnnXeeA9mfn/pD6YID16Rx0dvB7jDB+0Kvx2CvDPg3h3sG5kE+H2h
ZNClmLY/9stxLK18HxpCGeqjsjQOUuE2aRddfuuUIrnAUIMhFPSOHijlevVsUZIB
xq7RtiUDwbOwA/W8i6PLwTUepLh18cCoSO2o2AM8qGyAL+LB/sQoQzH4pZi5UWdk
lanIGZ+I68DMi2qm/QMKMIjSwfObYsy7DiGOiqlzgBV4UKv/78iOZYt6eBOz4Htc
DMhyCCFUukFcU26vI4pjUleGh+CG3WDeOfCU7110bTGUbK38xJVvctCLGCcC59lq
xIWv0AgJILJ9yos8Dd3Jl73Iba0WX1zq6N95fg+CfxhUulP6VdjYSSwHHF0CsJFd
pLUDCagA2WkEpln88AGvEuRwzxPgNtidwFa4CebiSIwzCgB4R4WvVfRfCSbsbdgX
AryysCVVe4fVYSvPD8/H0LBHIXzlmdt5U1v+0O3xQk09seUkJDshu69CVhpVGf5+
WNW7Fqq38PW2/BfOyxl/zDKlc1aaYIOYOfENtXxDooDalPdn5oDDR1Iebq8cjHs/
zUYLaTjDAIyBaYL8jRsk8oFi4Xot0AjomoOpaoEbTzmojh7Z1V99W0fFRMk+MUQB
l1hFkAKHLilA7RuqEx/gjOAZu0Bz1xkzK/f63f+eOyx/AUNruX5FFg8m7hNWQhu6
ak3gMcWlhg1u8OT+WBPzcuqa+pLaUfKu51nQk5/H9jLUxWbUKpQJVEPdwg3JcEDy
m++CY/aNLMLcsF3hzMgt9j3OYMXeXxwQhr0VIHkWNWdozBnZ6mZniTpjOOvn5R9S
gvgJBn/YxWZwpq+YSYWGnYIR87LprUEZErsEeEvMwb3UKb+x1ZKPvOJPouHBGGdK
kPWbbBNzq0ou509I/2V9Gfcw/SOc0B/pSDbxgfutc0leSdC2TqgC+JlM38LIh1tx
tMJ2Jhr15gxruTLDkRrGWIeeDVuKv6EF2QmEahAMBcBAAWOK4nn2gWP4PMHK16b2
VzqrXT+MJjnD0SyBDOTmftgOj3d62HIQJNYZD13kcdzsBN6GrBatE2laqGuktZzy
rHgBCv+Q+GJK3h+IZocsaU9kGjbdYSqifEbI7/ObohwccghuevscnR7oiGKA3ezI
2JxIWNRDPU0I/lOmktTwf8P+NIo0Vq9Mgvl8a9Un4MoA9eIA7d6xaCuVIpgqF/+x
FlPdQu6cnkDmDPtFhI/UycW9o5rrfW5DptrLJMUfi1PPopgZVK4cJqmXnQjrWp6e
1YOkl/dFwSOM1VSCA/s0xxHZfyHZJlhUMmrGVMX1Y4+5anPNG12rEpLSdFsUfjyA
YzqaFx0mH0xuXLhydvH0ozLwl8xtnDz+xpJlMxdYEMxjwEu9bD56bW+Q6QKMnQnY
ltF1HtS1vDvjkkRrj9tuKk5uuu5pIhspPtAKbIY1RYK9Wp5aQXgX1TLEf3hBULlN
9sdrPDVc4yMLnE/vW5Cj/BD60bqti2qAopZDl47R2uJcwtoNG+6+3yQFbyk+WIJz
a5NL3cQZXKBVCPW7fhT5EuE8pOM8RpRswZQRxy/JKYhZrooINwJJz/40eFbSusnJ
zyCCbND00T6oRdcoISTL3fvxT75Mg0pCbAo7KrLgjGNfmEwFcHg8eATm6awnVpeP
oe8eBuGDbr8uIM30ZIvqgKabyp1xuLHNoCU7nrEVTD+XFqm0m4vK6XCeiGn8EXAc
+KIOCm0bxjveBcyPosFmfWW8XyyhgCUPDS7CVk2KuqENu3ZSPhP5aoCXWerPhqZ+
bobLish1Y+VHw5A4aql6H1qwZ+f2qCaCl0VylkrAqJcvz+f1JlD2CnK/cLu49FPS
rnS3Wx+FeIxJZMC9KyIcQoJXgBrXTOjWFyzkOxG7Cg6fTUgBIaJDNpsZYp1sqfin
v6x+DYRWKlnNAGusyPwltiL1EnEU8wcO9aY3cBCPEDPMsF41P6VGC4AVB+JCa7vK
XPfAXeR1ZXokpzkB7WgLWbsVxY6CsQDG8GdJTjhqTdhcTCNgO+nKTE/x4M5iVd58
1aX5TXrcYC42PzYVc4oP/vaMijLzVUDWDgH9S8WMldgArGptZFd/S2xFLrsgZFFf
/R91iUNFVexRrBcalcNT4YpH3BcNiHuiart4iYwAoiUTGb/IL2uMrurIWUIP8ZDW
cZnbGHYez1zaQxId1fzN+ddZVctBmrM+81L0/h1NkB9rkEW8mbKbJo/6PHIxBf8g
jcANfcxEAHqBkuyTZXSgoPz5S5bTlXDCY2kLGAUnc7FDn/92Fnvqymyn1w5GwpJg
IT76CysO650TcwjKTqcm+JqVvzWZj/i1ZF2iMo4ILoNp2sFEHyYTJHU3oNFyXiXa
oT9/6zFcAsAswyNrX7ZP+sSG06LrVKYy7hEuD25fPRfuQwlpVZ+GOS1nWnkrMrrA
nwmB4Xhol3bLigU+lZV13V3YDnsbcAJhAo3QRZ9RFOJeTVjDhGTYyyD5vhVxIQYu
dWeY2sFqRh9FTWqo7irbLWHSOwUleZGv3Y+xKYEvoY5TRDKa/zwtjAV+vApkN6Pg
KRL/sVBQcPEoqYEakwK6al01ahDcsLyof3y3Bk4bhNHdrXqE290DupjvZT38Qchy
4Wlv8hrjz944EFqu1QJ63Um8TXK0Ooa02LWrGLRFAHtBFLN6Gep6CcwxnJ9VuWdm
3tB2sYn/rldinzgvUuFr83Vz05cEap5gPBW07qn7ffiNvLSsOqI6HHl/AKAp+2yW
JJ3i5fxTnxNaPtpKdzn+x5JjqMj4x0dv/tQQzMcA34R2SPdK5ItGmYtpLj8XcSMQ
mZYLqdJ++wB1Y7Ui00eKkCSQoEBJ7n6eot96CMPChgKdxO9ONkkq1XgF22cOyfg9
dqrB55QJTl/f5Azdk0/zi+W3/uOFXvEB0UkrLQo9iybenfPdgdO/C1sT3LjMXWe3
xvQlC7zM6wt6yWRYbpTParT1stmlxNWQgZwLVNVygAFnG26Wj1oiOXO0a6Un0/Zh
jWNC/rlsmkuY3ngDTQTi2bm9XS2NXoLzjFVOtT91C4/dBOY3CAzUF0TZPN+lwyS1
dMFyQ+gjwZc48Buc/2UM96Nd8lB0J1tpasGfLdGyMbbZJma5CLLVxAjs/Oh1WbyY
Hzo/x2V7KR+jrC1Z2kM0rWyg/e+AXYlFu/oZZaxWdeakw3RDu/eDgst0vW7VV0o3
bTag4WX95tEfqqxJTWUXVN6H6ERBTM/JClTFPXPbGXiPf18sIpmAPATDnrBWuTWD
3YHahcpKI8O2u3qjH72RPpr2lXIM015dMQM0FFXBCip/YVm2jKnF31i1pOVWkvx0
oG8xom5ETWMhi2wueanM126W1jSraBd2FteR6y1vYfXkg6ciqXnCitNCEOT/oWv7
KyMSSKYRXOI/uuA3cPfMi01rJ/FWWjxBgFGjmZAZtVthtIUHgmnsNe6YK2t8Rzjj
hMaOWNIlKFSI5WCMqSJLtBAnptjWsVr6KP76HvrpjqrCq5Sth9fINNG01pQe6d+d
5aYeVwmOHuaypyXsulXTHObCrPlsUwFT0ex2LjnvmoRi1Z4GD/Fqhz9hJZ2D+YwZ
7GVVloQBUu50LQDKFsp+tH7zbpmBgsMhExeDCFcfOQ0zbUj2CAtDgrSbX/FeR/Wy
04PZ6htXNWwjU0EpTyO4H0YkTml0SdIwyPagn/l6J/dWO2CxBVTP17RbDbcOBT/s
pFX49FO3KXL2sbXnmZ4wxALOX0VDVcmys3oYxCx8jPae+U+RCvX77YcumFrhYF+n
bGNn9y37tnXdPa79AO4vlPFlgGjYTwCVO5UUaZzcX2OYKkTE7L7RgLVVbyQrZO0r
eewWBRIwnzcLoK3iE61qB104AoCsWSVHkBWhbfd7meaZjA+NNeG/0BNT/FP+t2Xb
zkTPXYn/3ToJ7epU3Ock9P7oEfIT3JoV1tzueRQWJ7OCL/hEIWK12TfuAuIjOAmJ
0VbG06m3Jpa+aB3/sQsdA44Qepr/ZFoUzgcNIoPnGNGCK2HHfVHwD8rd6Xq3noJt
PL1HOMZ6Wiv7acZkkAMGAodznlBDSCsoQU9hWBUn6L4hvt16UxIhHnwJlzbP5hqT
v8h4nPrSVvWF1c5hK0BGS8gJGojKb9zl97n8vwa8yXV/nF0GioWr97fEEGcxcz9P
o/4tzrkb8NGCzDwcxprgK5FOqdrfXXfs1UILgq83qXBb6iEEjsaCacy9FPwQXkrt
9s5nmz+7qajBdLFXgwFz3xqQF69S/4+CGSVIuVlgQReZZlUeHPJpvo36qF8JjsLy
pO2DhID9pa7shFxLMilZbOFRT4fJaNjEwSc04Pp6X+cGHKW1m9zJFWrDqlyoyyRy
6jd8HbWfFJ+uqOfi/Z7W48gapO8HpogY5TWaQ09IGwinlJfo0SLZcybTw6JBWmp3
N5UiyXyAVHaLDQIh33sozjr/5LCckpZJaJ78hMNzSJj2b2gDI4uoCDgO06qDekbf
V6aPzsxii+emjm2ElQGZarI76kJMnNrlVSTGF/8jG+nzCy3c9wV2kdFBvtM5DO33
yVu1j3Jq2VE6txKZDN7ABFMUf4sdj+Z2CszyvXm++UsZ2/ZYygoxV7hXJjqLGpJv
UHNXacdbjMaVcG88gKj3kJFHFpayKOMoqFNqvcDH3zdHUjzX80Xc2pF5q7/D9HFf
NXEMWVlz+XzhsK+BMtzp177tKHkNkgLOTR5efyyPP/4inEGWR/rHgOn8NdH7L870
9ezvzsvin750o5s68YjqXhU98UWzmQ9/jyCoph3j5Ha/z4ARInxlEW1ylO/q/b8o
mvT7kY1LLw3h/ui0A6QwI/LWfolXBeEXWwRX/cZ92a9EX15uDV/tgeJmfHdr6TUM
2Qs3ct8ZHme2Vq9nU59lg4yUPbjw3x4cp1Mp6IeMqxyYWbVmI5oHaPJz4b8r1RZY
fQIyQe8UWiFvQL6Tu2ZuNyvXwJsv511oIWtofGau7qzm+/P3PkhQZVvZrVxq3ESg
ihEEnoZ0v2JEb48fXI3Qvn9LGloyP0A/b9EAEqh5uWEJwIArH/D+O1h89+DigX2c
o+RY9dvU/Q6I1Ngo8TDfN4TTKZFHF9fuZyg7o8FR6ZZfrnbcsiTf1lRlh89/HuVS
U93PDFIeD5YDHXSm0ne7kU6On5VcbnnSMC6FzLI+NKx3O4jRlwENr7+9zqoNpMjr
qoVNk4iII1vGZOlRj7GsVhfSjgt1FiDgAtUJr+9Xi0ek+opbBaFlUjTYe11FKPmR
+2Fe0thT9TrYhhpl/cwvNngvU+EZnhphAdApRmHq0jw9q8c88Vg9l7RpW6li9uiA
jHrztnbH2y5xPUMZI+6puNVWgu729hOZ7Gaoej04ioEEG0OV7ql+WIxuA/cMEhpY
4VA7sB7neknhWkywlv4QYn6VVypPVDcUxHBwP7knGW5185JlKHMo8mY5dt4z+xk1
hLqOrByKKevqFkQeymSGhtdzAPkb7fKaEaCXF3DMor+xPws719DhSZ+uX7Q14/3u
p9D2eDxztwFX338uHc+USPtv2q9UnjeQCW5dSYyOU2LnPuuRvyja6bTggBqylmCO
TxbCYFsRD/pg87L9FikkKv82VvE0fDjGWjZ+ziHDRwtP1OO68SInB3y73PPXP84h
6Z+dRLF+3ZnCIscjqssICQyUWMKLe4mya7Q0UL+waq5ZqFwl8ZD8mPXN1EEeZSUW
8gWlFow145b/Zwp73VCY2TyGDqCSBPPKOJrzjwSmVyX27k5QFu7yvYld4pjmeXe2
13fWuxSiq89XgLef0kmiPhjASjYj5IZ5ABMEpEQA/xSplvgh+m//b9SRkhR/1l4J
h3je5WQkzoigzCYZKhHqhIzXIppzvrp5euVG5NJl5Y9sbLWljPTSciVWNkRjkc9i
Zz+FL5l/gdWBZOJ0sb6FpJr3aPXfSMj1lbguO9RovMwkBEars/SAoVzbj9J1ICjN
GuaryPtjKEIp0wRN2RtFFBacpVJsCND45I6mC4Lx+E41r2y5uKDyNieJJyNXjs+q
F5OoflTyowuzUyCl1Db8u63pjrHvOmadpvkwqSgczkkFDUYNpTGLSeobj4LMOZZ1
FmOJg5HpKmwMFE/OLi0YCbZ0zFmZ+mrPD41i14O4WR8EsC6B7Z3i7vMGk9d3ISJi
CQbbi+jWPQKg1gK2CdS8BFKcU3k3BVQtn7EHhJq9rUtqT46i7NzM1wKoxKftN1OM
KSG3CE8gAmvx9fALHvTQnpUlOa3gZ1rEVGDg5uK3eOjnfxwv/otMxzn9EAnZKQR3
J2QeUBBt1melMuCGQfRREe96Dmg5EzUjY/ozzWqcXFmHzYSQ/w3iuy+x6YKAPrBj
SViXPn7fm4aIEl4d6ata98pqmK7Gi+VOhLa7valigxNVLh5lVOS8qgl7bQ7LWpg4
IoQ+ZihjSa6jZuGXMQZjAa6DJnTD9tChKLcV9PbV/5G+ildlXv+HRbprHJ0TJhuP
OG/QsY/3VxR7eCZyFCwHcGhkmV9fYBM1kjjqVNUtPd9QeRQ1ieTQ37Y2uoQQfzXM
kZ3emvYw57QTz6JXBhwiAIj2GUe5PK35oc2J9EjsLlVDsYGiGHZ0ZIkQ9zkrj7MX
AvitJjCBzZMk3nNWFyuUygYqljoE60mZ80Nbf7vf1LvAKYeJCTVaavuOYPQBEXTn
V/g2/TqeeW+dV/U8fEfhUmNnibzAMwSnuMw6Lo/7+QNetqVO0mRO11omSCwl+Vkz
BM3yeDkEdmcg9sTt/EEo46fpgQj0wIsAkZ6FhIzqzHcK5N0ccelsc/vD7kxN2iHH
2ApZtqDqqKrbLsQIVDnXhXt0HXIkjrpY9rRwLZYdecyW9RBJA73J6tyHqSzxQWGS
IxPceZtzBvLgjsOhxIPmUgKgL2nKCSmiKHE+QrYd8YZ7sPkDARAwyNR+4wCXWeu+
C4pluafeNIbdmZAy/r8I8lovA0MhB37eY/bYWlNa93LXNsI6ekTmUhsn8bN4swQx
9SXsnR7UyuTKqPDrrZPyhJ3eB8ocBBAmy6x5RNwPaDSTgjJbOFwgKYHAIUu5HzGW
FMsMAbyMA3EARhp8FW/Qc4CNyJDcOzX+uy6Su7G51apTVMEZ04urSCLkiOE99gq7
8RUfe0r4W7xGETwzkZV2ml1o4WUEjy8wdoOv7EfMpptRpprfT9J6Gu/tafqP2nFq
HBWAJy60jh/nULg6W9IdpPW3JQToPl6jaGqlg8zTZEwAe+0xbQzgG9AbyhPXPxdU
PEPgCPdrfFI90/BgxbtniPwf0JlXKjiIL3g6RCIpCNF9nZvTgJ3L+iz/xASsW1DI
RWrbL0xkUcFDMuMZ59q6flcrzev2bB8VEUYb4QNjBbKMGa3waY/AasDz/ZLomqob
W8IP1N6d610WiDipNmrz7WaV/5lJCZZq8v3kGmZIL1U77qRlXd/7AJuJwNpNJJvY
eoSnXyrkn2/Yip6NeE1z3ss/cPNlZTiJwd9LD/XL2h2tzdNnmiDS1NboBEocoA1f
ZyyKn3PNcsf+JzfDLMCQKoPZ4D9ONodJ0uUIY++vSBzwRgsb1r2G0G8qzGf4P9Y8
BKmj4OuXXEUnPR0ksdRSx034wUv+goT/cDMxaXqFqFh1B5xlZebyMWqc6VJNAGcO
o3Ebdg2nzUmrvZOQcho64rQLg8oJRXfI2Tvamp96rv61SXpvlBK5ru+K6HHu4feI
a857cC5TKnzKrh6ksbjaHZLW7NnDYTlUAcwqcSLhMtETCE7o3MU7ohEt6g/pOhd2
OdIZEvuRFpgdhyuAMVp83itkNRRX8LiVNcV8mXHC/vMjgPx8OWrc1/wxUGNuG+AE
Zb/EmQuFkt99ZwD12DRKMbzFepa7hnkpb3qx52zlWzCzUuGs0nb1QE8CamGHs6RA
FA1C+7g8My0zP6qleYUodIvV1MKKczvR4ZMtcux32DJzB2Gstsnb5BaJMzmJG/h5
6tLatP3Bxd3M3KIDfzsrLrJwGYhQevBfs6BpI8+vzvoV0XLfbvzdms7EZvCbGOd8
NxcCmYeuvG24enlKN7P9ZGA5MqI9l7FU1IHwot5c254UOfd5ycPPyhObAzqkr/P9
BzRczzeHPkcfBYCmE/+DY6NwcOxG/LW1Zdz49vCCMXmPqmF/FsXXAkLgrGFGpf9f
UQo5SAV6J+XgapUBvazxyv3zAOO6kVdUoXkKeXIGLugEp7tNtbgvpbWeNp3Od3x7
IYMmWc+JToKOBWs6P6X7ep/+ZKufJb85TTAVUYCZGkjJRWXt1kn9pp9TlTSCOeT7
qv8XRU6UPz0rY6IwXI0QEZ+EeU2z68Pt2QH1+Xg8494sqsohW58frdpXLrZQoY4E
2UW/Fs1kkX6rx4EdGZ3ERle2m8PZ2rAh0ut/yTpN+5+YrLV9sAoQwsuKg2a0mg6V
PymbPkjKnF8VMmXla+GOK/zsA6r4MuOqrqIqQVujQ8hKkgxcWhodEg1aSdicOul8
mSAqn0wYnTCMEQbSEYfb8a8iB0NfjMA9+gSADd3E98V+XZbbU3CHIhnomYZe2JBr
OvKBRQQDKrXULuMPMExpSvvs+tLdnGnf+JClRMLd0PsNNuaUB78Lg8vm58b0CE9N
5RHoxqGpfLTF7NzGHVa/x+7m2kzfAqfAZOvvrTt6dOaxqojzSfn9ppuuYCQXsObq
HVTgmKBns2ndsyLVdEFWD5mNuhbAmQUY/Hq8uPTwBS7MGKlPrp9q3pzbR2AcQKbP
rb+mj2vBAlgMgwf6/0muJItYOJEhuo1XwQ7kB7UPHogKFirY1os3anuLAz//pLa7
1r1X7098unIjRxHXJDN5WkW4QX4I1NLHzA1yocR6nv23DG6a6Rt6Q96BFq25LJ0I
KV/jW8h2r2vkaZJ8EB6oPjLUkewvkSQSI3+/JH6lAVYiVJZnp9a6mhSd6CndXtL4
LNwEpdJGXqQ8AKnugm9rw756Q8jS16Ge5quOzy7RApT6tepl3Pwj7Bs7FUZRzYMh
gV1wZasasDwjf6w9C1D/u6vzPil97Wu/utHrPVMQ5UdGow7EAK3qVXFF4lXDE84i
gmoQxpL/qzthitlewrXQA2i+XLJuBg1KhGWGx+wQEQY49eNnEjjVV4KxglevLyJG
AtG6Dj8u+RC3ExO/gwiq23k4oJTmfwhWJBFaKIECgL4yMDgCp502oeFobAmOu3j/
iHxAhEnS+Zugsc/Wam/7rNvlSF6hHcNxUC47+Qw/bV6wGDpw0lR3Qu3YvC37XQrA
4HqlXxDnV1SANn/EE1y9EY2gb6ApizJgj+12XXn+WnXX5i2HXdBFSyUCZh125MuB
Awp7wd9cjKj77gddmFgeY/mfMw21UJMGGOF5Bauu26bd67XFtDgrnM3sNRsqOYfM
4GCR5Flp/inkO9MoFGYSFKhnkcw5ILFFJ2DaCtz420GCuJqlt7aZISYBwbd/lUwo
SJHI9poQM+GVt2uuFMc8q2OYp09iNJZBpzlE3H4iktfQnpyR9hIKxqIs7AZ/3pnu
azOtcSlL5U4ssbKMfZ7gwuP9+iEPJrXqRMlyINEBnTEjpeNBYKIO82ha0CkM26wt
hBNDp7A+mO6xwiPrsvSC+SkhYNMSKA1vOaqnonEPQ3D/9HWda/zuSXe8aGf+pU0v
WkdMxZ3wra9EUQs2wGYGPrhgHeA0EC1/JA6OlLidcInLfiOYHAbrknJzBVQoElcU
si6mxjzRKkFR362SqI3nU/sa3KjnpztjintJaZueJGZ+PHS3Nh5+uyULziZEiS9B
8j2EXpy5rkHDSB08mtpdgyWGVRXHtKXnKe2Fh+TTlTOUNeBJLKFjPis9Y5Y3Gbd9
CYbRhQuyVNReaKO6NV9RF3W4W8KkcTnE7lu8ifVZZn6DRdnx4tNRscN6Mb96M5ua
gEYL8HBjN21UskPr6FpKWkSIVxxEh5TA+5uVdHVIO9/BU4W55f/EenQZrwzh9YIu
PE0yXO0J/xjx15A09mAkOZ+WuSZIPoGBAS8V4qlilri4h5Qpa1rvY02xuZKVPTXW
V2JLYYiQQxGSZ/fD8mabA+VEcmqYSKchhJ7ll75lUy9XNh3PleywEJXmVGUVdkq1
bYweMDqxsGMFz5Ng8kYKb90O+1qUjtF0k1viNg0PtwHJB6AGu268A6+TslvcZT4K
rovBAoY1qJknVDVBCizJU7AsXGvu+6SsmPRSRlJCOCOBirbnllkmhvx3CHTMKj5I
Hslnqg6srwQVpfgvgyI/4xnfdB/5K1UdXSztjmv8pye10FlF7C6HLi8oR82lcXRc
65LbHMUutY1tHeH5wWIvXS/QQA9OOnzR0Q5DqrKALuD7YqPMBl4BDcHmYP+VmhLM
1tn223VxA+ke+7H366gQ8KTMP9ac3gTlrCPeOAsS1tUHUvs1btYQRU9AgjWN9B2A
6h86T7K90t4GQ6Q94VJtKWsu9bdj11WwVsPwAeS+2/PBa9JYmiG6A0ebyfD83RZN
XGyR4lLZqaVcp+ZIghMegRj7/oPOfNkyW9ufRf0cYbp4bfb5cfztSbI2z1LfWrmD
ooYiY6nd8psyLSlDkAZX1Mmyn/YtYjCdyf2DDi7OExSJWjOI/pRmTY61q1MrF2yB
YyWvFxmHEJBrer2/d2/BmZWunhmsGZjMYcEf/aPQIdfo2YMMrf5MO2DE6fZcKqnq
OjG9p2zR/KYXp2DYTjj1X2pTjTqhJPV2Qord9Uyfv97lQQAcEQFjT8ieyEnjA/kV
owj4kG7ltJq/GIAjS0SiZQFYR0JOZUIHb2Kj+Hoi2yrIzNMAOe/MT0ToBaDz4TI7
de5qHDiyVFcz6jJsCwh/8Fj8OTaVb06huyOkQHNAo9wVmzErWmSua5Cvv7dqC9c/
U6UYfV3VTMNdYBmqaN7RwV8XgwJkkNQ5zRb947x/OYwE38IlrSZjEI3dAGjOuBte
GhSHThn+wIlTzW+pOqOiHaS4RMX7F9aFBdA1I4KXieFIXPYVRev4yKux4ka3b0p7
+sRzOTcGpMugySPYYUjZcFH1ONQv05401f/bMLHIbVmv0MGBAYxPgHYNT4AWlJ1M
uX0pkKHUyScM0PINX3enaePpqe3LVdIC0H+cMfco1ATkPWGzLehm9O5BogIORxO3
NHNHgHSwmXrd+WCcw7bChlnSSUx9DRfxRJqp0YEdkGA01b10Spex0GdoRMsV03J3
sROUyn5dcK6ZbeU3QpIv+qfVSyilhfN/cWqPEjj1L+lit55cWrfjbfxAxEAYaNb+
I0I4ElshveUEvkYpbVtc/gNIeROgw/0kJwz9cLMptgzt5vrhWItjlsSJ87a5InWE
h+577RJd0g0howiKxynBj7cnXSd6maxZaTybk7re4L0xxMycP/esumC0KgbPgs1W
JsICIYpJLmIVISbdZauw+/JEQLeUwrGrUH/x6SjvBBiIZH0bVY5SoeU/Q7lomhIf
EzL4PfJ9KC2wi3BSNU42r7g2ktbxVMwOg+KcpbWEJ4Y41uJ9ykLBKVHDIVRK14mV
tNyhI8fivxRubMBx2ChAEAjvW3z/18V+1BuWWvQxHdIsSlZqbrs3U7PRYDLevAHQ
58ZcFjsFBFfaKPdKQvmRycjjekyV70LuFcEHMqzInKEoDvwveKdRLK1bz7qamW4R
+jFiKroWMrK/Mr158MmhrCv6RePBI63Es/V9//47UGHY+3P25OECMIt4HHn/GpNP
YnV0j8MwRl4pahXoUZuIqLMAY3uazu+NJQSjhpCkQCWsov2SJg5zv9NCOgeQ0afL
bMoxYVHgdRLjvm1dKR3Bc5BisF6kBIVbwyQR6ZvrOJ3MrA1+bdsFfmayaArcDPY9
Mb6NGgkIQ+rCzKjK2d91A7cNd5v13PKkt1rtfnbQpRbILYIBbYeBTs6SaITGQScf
52hPoA/c0yvQF4OBdHYXjtfaWHGnL9mVivQIebTEO77Jj11KbN7fND84ql9GWPar
TQZ87i6a7z9gwL61O1kypaDXkc4X3ZBUA4JUxKdmgiHODx23Sn6d1ry14D9gsRn7
mE5sLVvdjqpwc545r5QI2bN8miaeZCHadIhbm912RagTqsfzpANB7q4JtsoYaTFo
msdAVDuLIy/id7yy/CjkU15QpyUd+v96DDE2S3FfMyZzK9I2rs9rfcFCd3t4DyjJ
GTBhlIfPThwni5QSbLQklKvzz8mZNCUW32xe2fHWBDWanDDIpNe2FAR7YcGS2Waj
2j3dUA1x7MO6uxR1rEDevHTCYO80pdE6ddBB8k1P7MpokbMGa//Zk9MFRIqZQiyr
OvZYN8mTo7ELS01RmPHun7ZNr0m8bCGC6Znm5O6hzjlLBqBAiR+fFdSQsRjUt0BV
UQkzh7L/z+vmOGEPM3t/oTbwRCoVdOpd17DFamwN8Jo+cyesNCnBGx7bBvdOfzXW
Zg+Te+lOVVoOOVz/Ssjy2NIbB8FYsziIfYjp6j0sM+gXMvOX3UJywZXXs3yqEYn8
Gji/5CNx2Rfo1RdLNaunQG+mUt8Z3TBk0L+WF6yFmNbIr+51UwKBUxvW1sFsLeFa
jE77SdZRBhG+gYoXlc5JyF6i2ucM7znASNMankwiPkRgkDN2BLH0D/5zTcQ5zWDK
gYRhw3bX+rsKXkR/yvZ6Xbr0kecR3Ox4ocles6zIEa+qRGKNU4+ozC4cjgG76P2d
IDLvtH/39qrAM3u7rKw1A4evt60ZHzVYBqVcqmBWPdLCPKh8iYBYeW1E9lDGTdD3
RvpV30KGAr6OYSE76GYI6xXONpD9m1W4PTTMI5LElxeZtNBnZAY9ZXED5g7AD5/v
RWKVvq8PjdDs9Y1lH/8zrceVMuXKa9a/zaICDyx1T9qyVOKEKNKhbOqxGZ6EVev4
GPFprV5qfcfqREXz0Pdmvzb/OTt/25ZXAItXRAS87wH0TgEh2RSLF8B72wR3o5f4
CYckntme10hmvgEXpnKBEuLYdtXBhoQpUMnsptaYu6IebbxIVGW0rmgR+PUfc7ea
bbKdk3PVg9EgsEdYG5nH9PPt8HiHvpaAfUmjRXIJn5NKlsuj29uo+Uv2EdfgfYhf
z28thQCikL9+jQX/x/45NqDKDp5jOqnx1Pr/eRcE5K5EMwu/Ss2hDRqYTqiitMrF
Bx9uZZnZhRlMysjBHZjL+oL+W2drgrn1c3uOZLTZ0yI4NKQBBSNgzssPEtEKvxEj
GHSD82bg6VlzRm35j0w2Z8iIN19Q5Z9fGeebYosg4I+6EsOtZYPkz/RVO3IgX0og
IZ26Xj97yny0BWzjoh0RSVlCEcfwE+4qSttUfamVQ7dE/5992PIObyx0uWhnPPNH
EF+SjQnKLi5J4YmMsmIWgJbDw5NkGHW5XQb3DFQllx0K/SBen2tuwWYhDSGOPRP9
7Ev/ZI7wAtq6cN1r9uzfP1gZVsh/4qnIgf4rzKcKt+0DuQdx/3TlxR95yRmb1rR4
MVcLD2L9nnhMVHXV4cvbx2GzVtfPmX2aTigm+XNcORfY14dlcocT/XRxIU+80ofu
JfcvY1HLNi9Z3qdIf1/pgsOlnHM2WTSMg46cgmwtzFzacOHN9mx0dBTbOcGCFXZf
ndP1zaiWcNqqPBxP4LEKXl6IgRzDYVfFyrzZXv/LMKijBXLn0RvVNwaBKt7DXxwY
l0kbOqDh/Woc4rEqveGY7cRrNoH9EV86FsjrM3z0VQrSWj0YBX2rCbWD40dVdq8x
s8mmj21cWqqf4rKsitMklbMxiRDHknZetswczF8Jafhxyw8IA2yhiwOvLTXBdiz1
ecFUGTVjX1h5Ye4zZCEyXjoTBM+eJEBbMJm8H72/YymVyxcyqlTMaOKTki+hOxrZ
tmOBzyecZopYJyEiaDg6JDqQ/31xKTEMR6zQhwHKyL+WgUHvcuJaY8lspTTUNbS2
Xwd+6aAu/76tgHrKx+42+CYzGgamDxvhoaedxAHI0tMHMaQMHKCV5NHcZvVpf0Jw
MAycjCHHOsxCLD0vUtVUzqmiHxZDt3vScDPGgHO7WptMCzYI75cDaxUDg60TlODx
bV4E45Nq/Zi+1eeiA/6yHrYrfV5Gvbllrw0sZ2LSEP9jKr28DmdPrf9YWcN1qZb9
vyd5u3LaZmZsDX0WQNAbp3qv0/XJwV3T8k1LtlRg0i+iNr9UMm+KOiIcX8B/BAVO
iUAUTXjNEkzd6nU2KoNh9GC2A7SpuB9g91ZSX0T1Qi8VNNsyuiom0rlL0leiUoY/
FuMCbYQnchY8FOFnIKDnlZbr0AzTa6EspxyYMMmG+P23D2eTDr9Lure4BP1zbGvs
uTPwE+phjXhuao31haFmnrALoQ6cdIsg5PwUK3tiVKxt3WuOIekKNGwG2b51cPMA
+skfzsDaOGqwkopdoJIaKUjFGCIGII6+ddMbdxzCRk0vLzw1WfvwnHrzNNlj8OrT
C2jolr5zRqT9WBs4uEe0Rs3fzs+zDiXi3IPyIVmojDLiDfl2o9i0wPa0QHyHcSpw
RZ35JBroSE75tH+R9nF/BbXa9i9PhyYUBpDQmuzKI+nXCfeMWtlOI/IeysX2WOSv
mAcC0hx7KtVsPxL996C44Cr/G6d/1uKV5spaYYlqVfC8U9Xn9FalJiU4kP78JFlp
7bl1+Asf0Gm0MHWaL7+5RuaoI5AsMxSXYu6N3nMHwkyHZ0NjGe6rtFJun/YFA8Tm
4fcq/pWAAGjiPuUhq7rubhAaaq4ZoYi7tQRdLuQhJxc0yA2b+4vJszqBrMs/AOEN
JpjwL33AcCHEng8ZD5DOZ5V5eWHLdguLQQdKbYrLuFPtlXyE8ggSZ5P1slBxePge
1zuJ1/jn4VJ0j8LrZXMiHUVrjuwfTVZ5sm3tyu5/WeEFF1s/SuTrsD66ZXsGjCVt
zwI8HOQIq/oMxqlzOQN46q5vT1QBogB28WpD3yD10WDnOfol/ruPm+r2saXNE6bk
rqAYF8Tq+UWV4wX5i4SSFb4P3Q4TDrlbSXjcfGmYzX50cAIq4d636xj5HAbgqs38
Nnd4TjsenHbUlvn7+blExsZcu1+TgyuU3QhhYKwFUFAzHkHcFdcDdt47gEGZ8CzR
AFdRoiXJWWZlK/7y3l3Ce1inJS7czYkUfEM2u7oLIWl4Bwfo3vhSLQBuL+TRKyyL
EC8mdaaXIbibRzwwtVAzSt2WHEIh0Dn0UimMgybAppr+arM2yxy4kPWFDC7BsdX2
BpvgSx6xsqttgOR2jOm0MIjElDOlQEHwWNQdqhU45iSm/wxypwiDFXxwnepzRyss
SVZHV+XsjkV0S+aQxNyx/2yS88u5L3/jw/bVz9OE5w7pqp8cqWKmcX6vzYcM4Ltv
Q5uyJABvXt0djgHe2xGA8vyG61NxUwxgxfIHwKMEwV6hSrg/0Cbr+aliqOwvWTgY
6bPTX74l/KanWgZfykGKPo07hxBomPztQCxZvyJl0Ozpf8gV5BH+CaRz6Vhu2Eeq
bQ3DNyef35XQRCflLqNcxrUOXVYiSkjnJoC/k2ovd/S1Vo+Yh+cbRU4EchouaAPN
MMR1mGLvjdCoECULs74MoRnugQXBwLCHxUiKA/oRKR24jxO3mTW1Oc2Xx6Zqmcrb
DpoGEjPArYetW9JDTamfHzQZMR2yYe6YfxoNq1Z1qF35dbYlcAI2h2cnVCIQ9z7O
i2xG9X4UWKphoYoG9uphi1OmGgvT+EEzDbxrl5PpcOUcJ/JHUGKx1hN8bV+sLb2j
cjrDhf1ndjKNYettVX0SUwa4MrzOr7sMuCkIsl8RS+6CAF3H/WxIa/++IEfEmgBE
rDijpzh9KLuLGN83r4RF+o0LUYgNUW1RWF1SoWkb+HlcGGgo/mBOp8DC8TBZkLSF
+XHb2FYAj0p2696hsJ1NP5EVTTwCfR13txucQ4+/gJIjz6drSEjy3iaOwfpkQAVD
KVFW2zBsEYsEHmtKt6AYxs8+9dNldJ9OU96qdRzpalOZyPBk7/C7Eq7yCMOBAAdZ
LkJDKZQXo6lQKs4mqs15NxsoaxhyM3B6iLI6VnNPKkxj6EnHb/iN7xSC8xlAkZlO
3X+EM6nBqoYoaOMz3L83yzqOwbF5FtDIRrIhm5xtx0q2+UKn+JGAec4+1oRTlann
rWWDWi+2KpXp4R2kOAVLi2qFTxLO2/eFimoK7k7h6/1AsoWub1sDULoeIjFsLbYC
gNx+IMnGDRJQb/HJqhv8CJqt2VImc4h5C0WYqeJXLTdw77TFxzGWRbdbXcFeWMIv
js9g4OHv3LSsWdwJhUzeTA1v/assbuiwttdp1F1SenwFK5vTctRsOx6KS9Ic4UtD
IGAJj9NmFpxoDgXYJ+juktQq+1noDordj5Mrgq6ZFN6WgJ/B7hSlYiS0Ezy8fkWm
i5P4GujVvcsIsSkOUJLxAhwE89EDlzfulzvLlR5Pa3zd02MYayLrAXj798fxJhEw
eS8z+Xx03QuYj4ATndlAhQI+1BeyUB+q5heMfgvgwPjouXM7WPGcgQ+iWLEFLIKp
QUI70ZVx8uKwIgHt9MJ1RufHv74YaXm0qPSbMLoO2ZVb/tYptFzhbDM0K02qRbPX
ycMhwBILMmilMYR9193ypPQTuy430gDJ63zBcuepbPkhMbGplaI0eU07VRlmvOS/
sWSh6D88YVPpG466+D75meV9BGoA+zmS/MAvMiloqFsdZDCQGF3gr4GuOD+RaCdp
ML/uv5pk9oZWMIsRFht9TN0+Svn5KYWGL80TrYUHUZ8hO5U3LP07FvVA6lEG11df
uzdHDJIiKaomdWrvCjRk1cESeMWGYUzOhH6Sg5cLjlFsguCmROJx9jzjouB5saWb
3hNkoyZeEG+ESAgMp2HFwln3UOC5t84DVKv2Gj6S92/OWYQzw/M5PHDnooZM4UTK
D1wPWdKIrPZqndsSm0PaiyIIv+TQ11qnMSYefCnwXxth1lu4TTWigl0dm9/kF0H0
PgCDL6gnCDzvkVCge1S9g7tUbKREbY4fPqWKmNi2fI0HaMV48xVfkfV1f/BMrNWZ
KPgn8rdlcwWiHgcG6Bggizjhm1IhHkZg/PDCOpzjj2FSZwtAB8OGvB31WQ2QZ8K4
5Iap8gGVdKfjedKNkjU+fhcDmVlvsoa4wMxFYf6+Nx/JRs8xJLV2PgG0IkjMx51S
uZNoPrkHUuapiHIyx2jetxZ4AXUgum0SAJFHhDjXhQF6L4cGtnB8SkScn7P+g2/b
CvSpGKF2OiaEGeZxRpCNI0dVEKD/dOtIPB5qJE1BX2y6FeOYaQ8u38+1wyo2uMpn
8gcWqbRGww61ytBAvGHBX/BG/1LHxwv4+zOO3PdnBEwsQ7BZbyuGf671XKZkUKtE
ezIETpiLOVBH1b3/XZeGzbu6+KIsc+llYs4iVmsDgPJAnMmmDMhlPL91933ck64w
z3OFiWhZO1dDnAzBOsLFfSZLO42tcqme9TzCrpCCcRQlGL0pmHAgTgZadpwsj+ya
KAV6oBXGRVNQOLUO4phhHCrIGVwCXVrk10k9jvHjaIfkLJvS9Em7UetE4/oW1LA5
+poYhVsvyKiwWx3oHiPlO6+frwRePKlT0iwaY3XWldxvtQ8aUca7Kp2FGy/Waao4
qGb/LTl7Yi1b15TBvSdBtfeE07tJg5CF/j6OkWK+tdgAD/Qvq7Q56DyZAwAGSbMs
SDamFrH7WrMoSAJxR9OVcd96IUREy6hfBesmJGSKBtQT7QU5tPa7blzdL4D9v33n
1BWzQWnbiWm02Pji8R9D9d/bmLzDMRpUXyBVaFH31qmxBiVKrsODk6Nd1TfZbTSE
2oUi+Q1ADrXFIAX03y6B1FrJvl9Jggl0hAPsoHLZMamyNrAHiDDdskpPxj862Bin
3wNonVI/Ym6Qkade6N9CBsSayayKYUS2lEwHlMGzZerFZP7nU4cSFwHc0VhV8iEg
exc6gR/g1lm6PPc213UbhNwfZjTLwpf9XTkNaxMfDcchoSKglbFJeuVXi9MENuo0
KvCMuyR4sdjAn/rkwCfwAQ7D4DJ3FN6Bhtkad3DumoXOlHJZ43dWoUcc43FisDZ5
1C9y868J2zEd8uyoj44aHwJSxnNNt8KfO/rBxn2lZUSXeN3Anv7l/8sfMRmvVgA9
0iTXi0Qjuc0gZSkh4aBm0Kd/22JMwUmaLnldjDXzebpbSXp+9fTUWs+F0SjKOmQj
JSqQPgLwoj3DSbZddABlWyZONs05Doc/3tXaqC3adTJ83YCT3eulOc2PnZHD1Xfs
zZsgOaLZzp69psAdpliE4LK9GrAjklEM7E3JVvHlGHIFgpLo4G5QLnByPcqpwXiO
C0SxdiP2bZFRySzQcy0lax5ZEMi2Rhhf0iNnnomjRmDibacXt65qrvxUSZZAxAtX
NwkClFWnL3dX+rxwVQZ8vzbnEwp4+eo4SFfLE/ISqbI+OIaRi2ZUn8rfN7BzpcIB
o5XpdWFBuzXzHonT44tT+QJhNlWnb7ayq404eo20KjjGYo1WqHHPmlETbYrkho6B
MJifSMJDdHh0HshQTZlMrnDH9MgRrip8r0sxNJyzs3Wafp2q0zDFddQtXljfjDxJ
bZcqlBfaOjjstSgiZiGBZp2Vo8+FQiCvvvnyVrlbMxuPfvpKAn5IFWEzUiNSQ0md
VpAmwb6DsPPOc0KrXoTImAFYFigIknd+qHK+tIHpcAM4Q8AekX3W7iAs3fXiih9O
5eGPEnYuYx9ThGoClsgudJ1ij66lP2SVvb0VMr28ekI64T7nF5gaT/I76CsuUuTL
wW5BBycvsVrECTEf8odJsjuecOdfrRVa28/nKf1uqleOZqjNFvxcRLmGTQ1bjTg4
VgKYDDCEVqnjdjjz6Eefr/V+KX3WVY8gxgv7bEhnFCa5B1qLQtK0ofJFwQzMOQQu
cr75WztalJh88Rnbb5Js1KYSoOz7TR6+BiyxCiagu7LZFR0mYst1QZIkB04V8cdk
d+ZlHSKOIjCKq9QS7KFneo/+ubVGR4LeqQ7zH3IlHVxxO8sUgjgfKtkqYHeyTNYK
lIsbODumypL1pYh+n/RFRlSMbxOv20b74JbX9hq1d1AWSU4zT+1gYU912bGTp14Z
pBbjxORRKX4/ijGZYxhebF9rjGftTluF67gbmbdm8dXLTnd8qjvDzJ1WRI3FYAGu
XEqgV2VzRoPZE17/Npy1UFXZ07N1aCH+TIOsdJ++df5ZK2icsfHv8C9K64n1gIuy
Wz/NpwJK5sQu1RnbRn0Sqf6FFjlFASutFPAWRJRXewTFtEUlL0K116if61cAngFA
xfGeB/hZUM5Mt7ZXhJY9uVUHdP+h1RuseeMHTjxkAj9Ua+lVKaJl9fY7COrtjewC
fk5cIqr52ZqWmkXorKpCDivDRZcqSv9X889k+XXTiIpXPEBBC25BZCJOq3o/iBtS
e73RDuwMxisb5jkiOjXL9+lv5Pip6QWqm/UXbp+HCVy937byZw0RIu1OlC/koOR0
iTLULa+mjF9/LU2Lvv+bY3UcbZSIXWaAyiHnTqsPPhLNOJuZ57PXBLIrSlGjyR9Q
a8DgugwoRKM/ypRySEffnnUZwrONERrwPe9ftiJZL281ioHrnvQFbioFNx6ujJ6I
VHnumKMge5H6RF01O5SHOkz+IyiNUY27VusCnEZkJeK6Z1HJYrnF0Tdk+RprmvEY
S2riYBw+xjJpV0EsiiyOMjPxhzzj5m8gf1dSkxAzbD+VNoELA6565qRB5RhcIuQh
N85Lvb8ErV7Os/JHMsufuYpkNiaM5cQpByb6BInTUEWAvlvKIkoiehLBRUaslcBG
Q6fFfg1qv/EfN2M7qCDVg2nq131ESRUBCvYOGbpTmHYPOa3ZCKhQenLTlWa0MOSu
RXNJY9sdvQxna6xpPg1gY44jd8xocNr3WsAVThWZgniHid+ZJQJCnYnRL/bfgbYO
XufjcHQ/kPYIrL/I0OWiqLYqZNTnnh0TO2ojPE9zD2LvJVH9QoDSZYbjAiDHF/uh
PWYMj0YWwkt1nLYMA39XRPCIYBe4PldL3BRY76oBhMVt+oSfLDC+sQqkkSPjHfHI
OLttfdiWHt65KjI/tlQNKOO/ta9KYyLHopes8b8B4eBr67IPPbLT79n2/6ya/Tut
CYo4xh9ekMtchLnGlX8bOvz+gli+iE46nHwRaucOzdWEnUTu68CBdKqKKxZ5GCaJ
X+9KO/GjkTZHW9VFLChE72KuETzaWqc+6z3xr7gHvIcIw6GRLLrKein3d459Uqm6
YpTVhvSUD99BH+7d8tlVej+v/cZxagC83kWfv0qrdkVTDi0HrYK7QntXrszPA0f8
FExyIWf3J04p8owdte7nyeGaq5UfHdleyLRt8DnIW9UYLcfV5akgWKYR73eZ50GS
RXpo6T8W0xJYiQ8+sM7L6tIWfay+GYnN5RBFhCyCJVaT3cchoR31Fs8o7I2EHBm7
1vlY6nF/O2ZDemZ+baqzO+o5YYrf9+EnTaWboRYMbqw1m9X64OeVAdqVQdyXxKI+
6QXQRRjwZ+XFs4TbYwxsvv6Ee6TWmwhGbyrZSsrA3tLHlS31MllB/EftJmffbxwC
f+5Vu0wKYr+bGDyCz7lLqcn/J6a9ztrMhH+odfxMwwao0MN8uG2hkYI4D30feM16
ubI3yJK6FJvbf0QSlj8c39qBxMwrR+Rz8EMBpxzLa7+O6kVEkjVpd7EURTJaRrBH
v0ajZWFAElZ9n3NgBeFmzIc4d0H8uR3LyZ7hkUdE0lLaF7FOM3jJPIyqk1f0orp2
FoU+AMQe+GXYTNtP5mZb6VP4cmwGsfKPNtpYrJx/hlcXI2Md7J5O2uymeFMPi3fg
hX77cUYtNDVYAkRqvmS2daO9zUIRiFtS5l8AMzvEQ+BXRQ7lbKwZAIr+fHl1B1tZ
Dhr3hywxsXm5HHTj7NOp2YyWJ6MiZum1PFTL/a15nTEMBFk4abgc7+CxcEACEVw6
bNfaTZ3dQ5iY32UNsW6DRGBxjFTdtiTHteffuOZmfBaK4/brS9V4TOdi/G1XFUbX
dIivuGQx2/HD7+1unQaBw0oCyc6RmJ1BeA34x0ipKf36pny2DoVKYd7u601+C2ip
1oRLN50AJ8XA/yd5k5ESASOc4BMgH53TbhB38k/mXr35WROHhgmzUbG08AZnqjyD
lGe/yppvpAwmlmDFo9YS/9M6qd95wJqQe7/qMAPhNV3dnonMKUHpoHH4r8hRffP5
kxNU8WHuq/7CgMXp+fgclDoLUaElp0W1/aOhaBSYuxeJdjXjHl18qxdWVpTcXlAN
7lrTWpKKoyA5bVjzcX+kLFRwiIMSgEKNR9HZdgyocuq9iqjVOZ/3wf2EeSmUlgWU
Vc+JNZSlxO+D+/mLDsid/MOsxD2LAWn/VqrQ6Dzm7MSUWKYJaSrcRb9lNllQ6qFD
DK3WeJLSWe1aGvAwiAttL05fHiNGVQc8XO+YUSVkccBCrbHHLAyD9jfk33T+hr+E
OHUdGX6hx1kVKvePDoP4IQmnkn2z4S9W46KeFTjMzIJD6jY9bY5u5PNpqC9zbX+A
/d9lizfhZ2J2P6hMrwueQoOiZWk6CXFwTMdkNgZpfZrmcKpNYeIYbB7P5MVLryo4
6kBvxbY1CUuZICg1a77MGHvbVOhY4L5A5uK0SslyETjpQk36vWtQZDJexPLuPXoP
bpW9DeevOm725+wKOrm4BKICmcKfzdbysIE0DMdq/FA8+N5s++EOzB2M4N1azCFh
zpT2qio8nX4oAqy13b471L5gDluRN8Dx3xh9GAN5NjxZA58k3KfBdmU3j6RnRROd
caZVguorNoy7PVGmvWJ19qpFTmsmtN3/X+0sJ2Esb4/uQCsNaqbabqSmeBUQqYQD
WC8AWw8Xco01/RyR5OxzJY/JFG/3bsJUJwT2TxBA81Kl4GCVkccsrzvTLcmyGkto
GNB+NJR9xpWOZ66yjYaMa+pEHMo9iPZobQ14JZ3olAOPT0P/RQRuUT1dek5Duayf
e6j0vKQAu+3iyV/fuMrU7zjA/0NFHLxF6uePmbeINrUNaDBHdndgWLDR6Ol/0Fnx
LwWigInH8qT2gJ0wcFZx6rhuGp49qDJpjePz0fOD94eBH+b0QIOD4eu1BL3qCqpA
V749HnPfGtl6knwsbj08u2Ocj5c5nTlBuYVC21Z3pXiWQG/dCep/zMFey8iR1u+W
iVz5e16aLELXxINjmGxQ6gNMc+b1awHzTaZBdECqkk7DCc7nllrh2+HVe1vPtHAq
8f3+V0ctPekwpKMylz9eH5NKYw7pluwnp37AC5GBfsn5SA5mjC8gEItWKD7jhfaU
4WeUHzRhAHuoO6CboqIiq1pcm3Fv+6y97FlUikCRwdQwdSjVNo5bNVW5+gILksD7
vIiJrMccUR6oVSvHkHcJ6X5BtrdJp5vjCCVEyKsDfb8ogkzDcErwV5skv4efFh/p
cnXlIIKFayNqMOyrQC7c7+rR0a6icjpjnJkZK8wOKExUkCe5LqM/KCf7DksDDV5m
/Bou7N/iAGAIBUGq7CPzq7XpVwkeVlYGELZ8i9/FBaTPDrscgFk4YhuwL+WYZK80
xf5bYmahUPON70I5U4k1Xkg4o/vmErQjXZSgjTpQeyoWjbLGX/gE6hP4f2RMBgqM
4GBWr68HqRzVRH6xRTFL446HG40XMl00pgqRYaEaELzqHmhyfBhEwCbG/VrpmN3B
ggD2UB6F9/WB9YuEWiPzDxLgTfrnt5RNrBNfiZgi7rz54NM4Af5PbNe5SC4W36Zc
6mFr4mANhFY9PY7ln8HqdDeNe3bJuYEQ8Q2Zmx76tykHfHn3O+Q3W/nt2+dUE9zb
WK471GOASSiaU2xrS4fPYYcEAnBQo3wlBXw19j3mk3SA4NYn6ctHd+c0lNVjSlOO
AQlJrVZ2Sd6jtwyazEwRLLa9RuYUK7cmbapaIARZIh+Z8bGZvQDlvne9HMoArkvB
cDzt2CK637cYr4YSvHwlrDYcQCmaTQrKluYzXqDJfbzBv1qIGDxL5/pYgsWnKAoz
aGwO+4eyER7Fchoq1D/1703VeJj3MZuhAMQOGRTD2uF3ZxYq/ZiJaHMRR1hqlW+k
vOteWq+qR4RusEBzukZttsnWnbd6dhLy6WdvFaAOLjEq/eZvtS3//mzmKJAmyD/d
kDROSlEVgrod773P5pnkohjrYNVwePWzg25mLxZfaGI2s1rnlhWOyY/9Xe5gGkwu
hKAlRYvtRXOP6YikJl+0eBwnPD3+JhxLMOD54S26Fgwv3A6gFFZR37l/gf44ApsL
sPPJd6RSSa0CyGLvwAEXdQ/QtgRZwdZeV2kaSlIS9Dnjh2QM59WmvU2XIpSwesHo
OjkAN8PUvjN5U4xeyq8i+Je3mxTcYaLffaeW2t+c847nY8m95i0MAV37dV94TJAj
+vI477hFWaL6pCi2peEPqPShk5JcWsDJPRjYSmYQMMM6S87MSKWOdYZEW6SwnaPz
RLEcpj/JvWAcYVNseAfNR/lz4x43+BrNcpZ4pF2N8XH1qQZm0hwOlH9SLSHGBuS4
87RyI4bORew+OIjxSttyBExjgw/k7OR2s9hvvaACkH2yPECzw8/XhxGuMadAjD5x
tpqB3ZmH+NnmIS1JSzgHF+76UfKt/0FHKS6Aq04YdJLRhGjOktcaDsqezY7yH1F7
/aE3fdCUwC5ozxatCU4kWu6+YY2Kx36YQ22Ao3GS2SQFM8uE51f4PSsZVNFgOc2T
kKTFwmjKhC1OiZA2h5MOf/LBwboiCOZ1WFbWUOV97tFH6UJo40jX8bc0gx2Fl8eU
HYUQU1pjGvwScUbrHzenFUX8EFH0lhCJj2OPtMqV4Q0OsijfUN5C+yYbno1Ie8oy
THCcf0VV29shxig5gewhjpOU4xpzjWtenmFrNaSmgJQ4pUhaXRLBs2a68EKsaloN
UwOQ4VtYTJJgbP7D1RXslbDa1MoMkXuFhaMef6YDHKrzV0oIsl16tlkK2R0mkmza
IKvM9RIwv5o4ws4QSfoesUp1b1CErqUC2SMiRlz/jHtNKrxY2A7NGMgBW06zc3s5
+UlqpJBZbwZZVqFjSpvEtOXkioKexdgR5nAE4jZPfb1rXBklEzGqpN/RYB02ltES
W3Yof9Ey0gj9haFUxepeERf22z9pVHjkoMaBB+v6zKo8mhEJdeWDHC+sx7iPA8Gu
LQQvqDtH9xjBRiDAIVxHSKNmTwSR7Z+vKxDRqX3uH4M7LEK5b8AiNniT8N4HMapQ
vE6KLrZYGrHGtyZBHjrpvIT4TjT1I+bnH82tt9znqMZnz+AVy6ndpkDxK2Vj2Dki
iju+cUiJ3TfP4BC2B9R+gO6F7/H1sPwfXZ49Mq675QSy4ca1ueCxjPsJcbjIYEku
vVAwYe3gLYIS22IwVYcviDCB7YF3G4+MYBX6xAExEL77WyHnnAMa+u58Ur2DTb6Y
4gUwc3XKo4t4t3lPkahRXaX+Q8vrdBsJ06TvYByCClAUHmRUlDHR+1Thcj72nxB4
+kDPLtgN8D65zDe4UQxef6Zdp50kRyVVG/dl6JSEMHaIiauzWr7V2LUkSpQN1XNS
o6scLxy0uLvPKHVJ+aP8OO5GrDfdw4hYHtP5C9mCleP+iS3m1QB+MIq3QDmNtwOt
2n+rxS4HwU4j0qY3YXeaf1FsmV4xoU4fNgzsXZwyxO7Q9P9t1C7a7PGObSEbPzXT
7bMXWsfCvYZb9h1A4pupHGK+nGMPClDOsTMkaPTKNa654N0RHzKfAynlL0TNQmOI
wLfTLts/6BR6oEU2NRtV3aAcNH9ORDJi4mh5amk1dTKZhxDWSzdRmsNr1rfz1VTx
bdvEb0EkgXFNsyFwMzjp1bDsNbyi1gs65ZMYjN9B+vi/aZdk/C3SvPfoJ8+/2ah6
GHSNEHUWmCojf88DgvosH/ThjH3QjudtoRadns7ICOWIF3ic72FGemQw7Nef6gUO
ytTlq+gls6UEf59UPb6wc9gIPVqhqTaNo3OE30jW/2Ab4dU51M6gvOSODYxaLseH
uR8V/akfsySOiId58sZEccijJtiPp0K5lsWUl1Da4TDHEkteeoUm1T9g1p2+jMS+
3sbZdL+yO/hx9a7Vh4gCShHsDIItaZYPP+ctj/90A/oT7Nz09ETIOBoIO4MgO2MT
Mapv6DXPk3SKJEqRn06jE2jA6mdeDPNjd93Z/QjYGmJyw0++Jyd/GAhWKicUO09h
jS8Jeo6tDO8kwPu3OzWyzxHYSeELZg2oFrymm76q+3RCoCdNRAG2HUrI6MNFWO7a
FZ9CMmvUjeRnC7FDFHeJV98RBlNZ21f6WHYeULqOZ88o4TqP6mjhaGa5J0FKY9EE
y5spLf4DOhzWwjJ7Pa55flgvmnN1bLMYxNqVm7UnWFNyH77VR5QVVqCKjV52lwen
86EghRAVm1aeiIeEJtMHga25EoErC5/FRAZ65+HqUxSFwkeFnNjwPoiIa72Ytc2K
fqY3Bbxxv507bMzIThWF2jTN/z5ta4zvwmkREKbSvDQJGbaVzxPvCNesr4HEE6BY
qEzWfjzWAR8bdtJvBb3IPAUYg0GvPybtS/zS6cVCBk8SCQRohndi/GRe04DURMUO
kNEVeMFgg+DFup8eQxcvYcz85FXAvOQbqf7Q7CV12jOPKmQMVZYEcQbhFPzckOs+
Qkj9TYutwMtYdEhlm+Vr5syy6a4X7Idt1KRSYZl0OWdJlKByapLDjuzmULKQ62x1
ZzGCtjoJhOOcKAMqeIXb/Uu5VRkwu//09XizT8Tbr4BN4vbBx67Jtdbb3yUHSgtF
ofnDIumhqZNZsBDLdymRDjvxsay4c48aUtk6W454I9Rn4a/m/H2nxrDRZBbjhd4j
C04CXvzxKMQOfl7uvjWxHksZN9sQKU2HE2swSPdtCtnwQO6g49J2EPKtY/g03okh
QbXGv/I6rTywRPAW+Fr/tBQcv2nwXgMtjTkmsUQ0AawLjgOu8Z1nZvANgvPftt+8
xgUlYdPzP8Lv8Cqcqe9NRAzDJBfW3Y4+Kkvn+XOOCr2P8RZtkxVTdW480l00g4Fp
mwS2ImpN1z7163gf4vlVXrbAt/KPirNm1TZjqy5YI3Mu9pBCVVFDpipgMgdRlc+p
sqGleYOqj4HVeuOhkCCdy4bH895idQacfR13Qlkz3dTmIjBTqej75kSsHgKrWUzc
/6GXHLHHIpbR/W2PVigLXe6ytRI/7tg5J8T0N9i8smfzwL11Y38jypsgpUOt7c/G
1tofV7p86ebk+71Qni6khFvbjWbViM9OMWyCRBhQA2BS+d+DvJT2peJpVf6XS9JS
ZTNzfkbVJMsJkpx6Q8Q74+bJeq7QGR3CYkrkPuYVVATiGooAOO2kno06Gnp/oR5h
uPuMVYJ+jvTVo4I0AABbWJ8W2vJhccZkUy+Mf2TaocwnTTM2ciW4/M9NCcCl1e1k
BjuIeYFA5NSWz0AXIcQTDZ+SgRSKHfASEM6sg1+M4gQhai6UaaELDYz3YY1mxM6G
X1J7Y2/2govn1oN5jmDoZFz5JDy4YEEMmP9xzxP/m1cDMdw4KteOaPu2aXN1+xst
O2VCDIaMzNT4GL3yWfvr7Y/JFletOQwIDbhHZEK1LA5X86vwuUO7bhyVRKPV/S+b
qHF9Lv6v+/C0IcmPhoLG8fFxVBej058f0J6UxrTNgXbv2a6T27JTnYUHqSaFPiBT
75SmObu8DgHrCsm9LtQNaZHKeX7Ore2x3hZNxTB9PQi9i6fU130GpTl1zQGUh6uO
AZytuN3Y8mRgkFgMM/O/zQNGZSfdZeJsVzQfb2XSXLWCWQWFPzhz4YApYoezVxMA
gmEAhdX+BhiWO7nzB8NQxpZhoKVObC624qWeQndFMOEnI3q+trI+ZmGIIfYYC+CD
MNL8tQzZQ1+J7vWIay3GPkOGgPdgAuFN2thsY4IDJdgInfTlg0qkETviL59OWnTm
yRm2L7jfNMvuoUOkGmYVFsba/GzS5ePnC3kkgRMF1p8uux2LVAmPc9C/PvFSG48O
MFtK2TLE4UWFEnsWrN1+dioSwfEVa+q2EYr048baWU0VHLHC7tae80VsyLP6PUL8
oEOelQjTWayVaGy/mzQdmaGPihLoWu779A9/F19tF+gfF8o977FVRdt9tVBybcII
xZNpb3iEzr7IkyQUUfQx4Lm+5iGUx0A5NWET83cdnFl07ChWzNDvICxEwI2XC1Vq
HF1K8bg4tSN0/7SVuK/OrWl6hgVf98FsL9qn+z6CQchSEQm+P/xD+WU3rvveLee0
0UbUR/bzmy0PvTUaXqUAavM+ywdzoIIonPWBCN8LtQ+HV5HGi7Mzit6FJuG3bmFW
VoCM0AsGneH1hlmfWMp3JQsvWzQsxelasftr/QxAHnvqfwvPeYhV+BDguWtsaxhl
HrH6AqX/xG7RB6kU2ehe5O/DxkWosMbCyWXooSYNEy1GkBh+vD0V33ekPYZCj0yT
SRh+nPQ5gqkdaoRh7f7V9Ypc6AQZRocdkagHm9SbA3uoiNV4hS08HZOKwCq3CnXW
Ewr5RXnWeGMydtT2KhGMNEy2rRNM58NRzmOCbvnnB9guuwbqXV6WOL7mKtl+2pZR
fY8r83hZzX/+Ww1PGci1XjGr4XfF8kAresVandEvI76Q+sx2JvJKb+EPoCsrgNYp
e6kEPBU7EX+OhvxslcxEzcmAZEL4enzfQ8HjODECYYldw99ik5MdBJZ4brJyQBuI
QOIpRGBku35ArAaeXFWof09DckSwaqQUB2r6kwT8qAdaOTDQgG1DGGjJo6M9GdLQ
AI047v7xSq6JfGrgB7O181qhlHMo5lPh+qj8nMBuhlD2HinBxYw1DtRj4HOWsqwD
a4a6rlW+wffidx55pyPoolAbCyq41Q1B2JtFEabow9Ee8gx8eulgwqNFtoqhrx60
TKWOMlYP8eXy/fc0atRu5nqB6AHtsG4IrCdNAeRGM2gKP9hPsIDcToTPTuifdNgS
OFKc3PUmM6/2GrLJkssoIk5ZeRN1INQ89aLa+Mv6Bml+iVSsisD6J1h1a2axgu/v
FD33RgN0SgdulBSI8DLWpHvSWB3lXhUOBYET+BCzcZmg4KegKA8eSz9vwTJdGfpk
GZ2paIqKnfFIRpxtwjHpPT/BgmRJUmqxiU5QknHcn66refjOOOGSkgo09/3FBN1H
Gk2ONpVNZvgnnZGb589qhe7lRkRtD/xSu9Sd4MtI31rsqZ0TgHCSDTB4mTPIoZPC
q3KCAg7FOoAtNsfugezAXiTbNBQV5066nDGaB2fjBlB+ngMqtDuer0AJxKyCOyAa
FI9xLK3+caEEYG346OLo28aEOHtiUbfkwBrbh5lmF/TZVY7PlqUOmEH5hdjRO44/
kh2qhWVRbjM216iJJ3u3lgRWx8Hy4n1N9wB8Co2TCVPJDMEhfD+sFljnigccr3mk
LTM7JzS621/pNUasbKRePWtM8XH+4VEXYTT09yyxyJ0rPlfvzz8UnE8Qzyj6zRzK
U7pd7wn9G6C3uRKTZKJ3oCjHHR6LJI5CeaE1ZRBP813ryY8BoOSQqRyG14LWKFtp
Vfn9WkixEkn0KJPST0lKwnBXEhZBjdsbb7qpqCbToF1SCD3zq52/U0kOK+OaxI+m
HJpCnp9P8LvH/EhgdarCQZUZW+YXbUrYrCSaN228sO629bmxAkkzJXTTe8Mu0H2c
k/HZMYvI0W1vaHg74QkCeQwOsMZsq+qHSxqU1ZsMqGSWCuRqfORZBFPTP2YuR1YC
qioDLbne55HQB6Ui1zlqPyXcxm+El1sjRSGdPZO/TfkUsx1S00yp5+6KCRAVgCAb
nzR8hPS2yDrNgGxq/Z62T6lF+z1Cs7h90jFCKxhPno/mgTwT1C+ubKlBTffg6Et8
4u4I9kztljHEDIibvamrz49Xsgx1e4iYXUPKQlcMYUnC8GpdKvjwzhWf9nuT1ZmC
uqeihst3H3mYlozJQFWwfpshknU7dDHycNIjHz3OTlwf9/rdNy8cNzI6sIFLn9eL
ipqpfGBC0ly026bZoGmOZyqPc/NJiFF0F+80qDi7xkmWwZaEZuQZB7TvUeZ0po6n
KHfRiWlvo7D+Bss1WbkffFAR8MKemzTSzJEU08WjI/MsNT6jSIx2DsH8SJ2turyr
DD1CWC/ZQxndXEIlqYsLcrDHl8BkuVUHyi6R4lY0ODBxDMJN6ttAGm/Wxq94ZuDD
rBjJb/m0UdbTXvctAHCTPd7Keiu81C7auDbuyukE79hJbkBGxneIP73iC+O4z4Cg
Dl+sLbYEZbsdrs6+A8krh5mpuOc1K5GzfbtLUEWWnAlRWtjJvMsEvVBRuKY68DCO
+npX1OQzFwLFzDb8jrbeuX6uEpig7zs1bOwUcdgLHNTfeI8001YePC/TSCSObfMY
KyPlYT9PhfiEOldHwccAvEZ2DWTomYFPqQ9994q19/IMGLMrL2I0sj6vmxOm4KfR
BWDrCu6+bYfgccmZkEmGLa4z+Knk9U8z50uKNYh7jCg7OjLNf9ylTAscHhDwx4Qm
lZZ0y5KSejF5F8dFSrJZGn4zIa+rOxeD06ogY8EyT+0tbaPtJnIpXJZH/E1uVeuB
DEhBZefkgsHFEWCNIxrUlv92CvJ8n/aXzoVjuNVS/9j/tpjJJi4nqfnJQtHEzgpn
/cK8JQlhnaer7TPz3keZ6W2R9TvbchjNirkCxZn9u44ngev/NtQ6JfVrtoF2DdH4
A34XA5wbXgsByDWGhJDj6f0p0A0W0VmMSwZE0zrcD73M7SWD9HHRUHkm4BvJvaTc
hchEjbgTN5zpDx64eC5h7i8Cm+jlUyyn++GYY7Es6GCgUJ9sN4EzfZ5HoOMGg5o8
D7pbFF5v13Qqe8NMKpMo4Lz2q8etoMGzvb0tnnYrsbIecPlvFdkLimOqGpckOiK0
ZAsyATZIi1BjKPG+8XQRsVrKDghAsq/X8Qm3IPzLDmuLLB0Kf2H2TVksg/e9KS95
+/xfSgB3rYSd/aVCaJA6hVzSJts/Ex+FWvaUo1cStUX801AKFeTKQGTugNy1UdWf
gk5Ju+S4t0rSvTUsjHmFv3osrwPvhh4nHLfl6wJE01jZjrPo+Gg/hYJVhVWbPjb2
bRsnhzb+q+aWFmJiS3QTwhW8ih4i6uWLJL2oQgUhN/sp6zJqTaRL3W60I4kkWQ01
NIkHd4WbdLjCGy7+7EhvOWQG3g8Qsg63jWSw9wQBi2KAfPQXWHMvGuiURSl/0vqP
tnsQNWxoqu1ypl8nhWx8LS9ak9efoKznP2yUrLQAjhOINbr9c2M5TnzyakT1Vg0I
y0m0jq+xvGiFFIGpnsPko2aRtS8PT9nBUNQj+1LBPcIgQKSqKd8WsU4NNeN2owmH
sBQxyEklzeT2xAKwBX0xlD5DMEXeIpzFtQz1KBGynyRLpjy9jcwewLA+wXa05c+N
g6szBab9qBK7eoRQGWn4i/rPyejgxmlX5N5eVyvlB7VAxSxi2VdQpqLIQIorGhcT
mxdmBRxhn0Gz2MZJbGjz/GoIYxbTiSIE9rCFJCSEV2hRkweE4Tkb/4qBuq/IhjWn
CMQoKEWMmtjzZoYOpAXc8B57EuhluXaP46vEL4i0V9GZvanKpvHVqdQtqqaDFjYO
FJX1Xz7ZBkVUlKKyQJhs29SSu0DMh4nykJzwouE57R2kBe3pIeJD0zPKZvXlh3gb
2sNjcdJtQBASqED+hzzcBx89tQbdkLDol1d9byM9XlcCDp07rYYY+Z0p/mEPodGM
2IWQtNJQqzJg5jmIvO+Y3I7VwfX0uKwua0P5r4MMKUkUvRI+2ecxrwJID2/kN081
x+GeE7sXX+AkHTf/u6h9/jtkLeMwG6fXCc5gu4K/G3Gq0kmW7BPgX1Q/xsw0NLXd
m/oIF87wbxzS8QTr6q7NhZ1eNOWFc4Z0oDKYUwBq4yGoml6rbj9gmt2oF1RcdF7F
uTQAvP5ruMR8fHDQRg77q/ci3MEWwI1azqVbf+sl4/hWPAKv+hOjnMEi7EUMiLBj
ChmiKQvFbXi8khpQfF4/DzBPC7w9XOiWwpH6DhQC0X9n6xrJ+C1UDTafaPIdS/NV
HaMoqYRkIOrL0nPiPuHHK/uM5jVeyDDgnvbSj77+3iZjg5+BINn+riVCfqIyPoDA
e+PoSDc2bFLf3BLIyKS7oWsahd3WxQkNQbbcwvQHA55/9swaekTVS5qW8jhC7Ld5
hrtzasT7YQNx85b493Yu9/Rvr3CtPl/R/78egIlM3smMtgGFkce2923n1kQ73i7c
o/vL3hM+HRleUHErEOoiD9/Jiy2qhj1tPWHVcNOfnRBOdf0zXfL8oXVLy35ZSAuF
W3QQSxrZ24qweLIZzy4fTPMJQZ43lYJG1ZS/vKZxdcSpnQvTiZxTH7xe3F99yZZ0
5I10fJan30iNfMCxTSdTBvquVFYnjgfY3Vzme5JZB146FRs89vouCaWKh32mqSxR
+f71/GXs6d8z7EHEbpmWj/Xa6NZEgWBKHrTJCkv5LRPX4X4Zku5UY4UdEcexqWXZ
ObcC5uRcR59pQyoWAHYmaGuVznWQn789gs4LnJIHU0vq6ZlFN9JOqLq4Hy6yMDki
YQkoEzCgH8fL8OSSNc65IjfmyDAtWkeLH9uErqRrFeb5jyj5IGHQxl0xM9KXJeNy
2ej1VOUmuO0ac93ektcLJyRigGGy4R6Gf04TOuFeH1AZBOSrScNHJXQGsXHbwjaQ
c5KCIu5Mh7Ppn7GNo9MKniyysxF2YJJ2NUs26PT0iGBM5dEjP7IOfgEcP/JooDDe
Osyi6WoNPNiYliXHnXdMf7lbcbodzzlzVWvKsUgK60Q3KOrMHJifKxjLS+1QpuDl
xDuD1H0cWdhFphkkrhY2Vp4cvZGK8lpvYBW9h3UlvhaEXigLdcevZZkCH8fXyFW+
JjgbNs/HVxSHZr97k+d+owvtqlTvBbZ9f8kHAX3MBpIRcAZtmWzstKE/nTdc0ziy
9Ucgej1SfFdLLYFu26QDqssApsBCQRonk628PfS5Vgjd7npQJDF+EaQS5ezQho0f
Uj9+qRd9LqifstHDLB26NN44lgMJsQLGp9/XBLggjt5jPAs8MHz2zbGmavVSj+SQ
FvqBJg7mALhOVdzCvKTrj24XoyndJ14rLmnBlghL4ypwz38KHEi3iW8gq+VKsLa5
kzTCie9cCanOxHCozjvaEXtEGfv8EceXq2rOTxT1uqt1gqbt1bKHButiciiCKq4C
Gj19VsOzV3YVzoTbQxesfwXVy7JZkz7n5+dhxLEHpaCEVeU+VBDAeVNJQw28fqrT
AkcXG8Zl3MGAkDnB6kq2UWtJ47E2tLN8YLfokZQSxzk/DHAU4ywtrEfR3C91mVfx
psvRKdYZefwUp6A+hpcbFxkd7K4wOdWTUywuUMazIlpNGzaqJHW2zVYJehvAIMxm
3V1lrMN6XjSv6i9n4ScpRz0PKupe8aByHsmz+xN17x4rolaViGVQL66tBEYC5un7
kLhdBoU2wc33kPn5CuTYeBrHw5XxhCRvI3rsrTDRZfXtU4gMdvoiUiVM7GjVW3oJ
Xk7QMZv5CCDaNYFMwvPd9bTuylPcTkVg4Azafn/pEVlCm1Nx3Lbbw1/nzlTudZbI
nBRuSIET00LxsuonrtudvfPHzPN/etG/NqBxd/tZpQ5zvQfnNhGKxeh8AXD4kPla
5d7tZVQmBc9XCi8yCA9Rq+oZcTtmf8/y8JqF6TcPooDVQU6hTrvbpcI08t9hVcHA
8i+8dup0v0GEAn5CcCYQ7ul6vjkM17BipRCuwvMhxEpRUmbzqKnCbKoIdY+2gNq2
CcxRjdyiQfrsj2hnHo7+bddOH0LJJZp6wQp00MGEL6vn6mnvT4NMT1O6GTu54F8K
Bs+ylBXIgpl+qzDl1CjAV2bFot7sVl/r8bAV092d8DagCA0eyhcBT8EXshIvwUNA
8cwJWFHmynoR0ujizN/vzyNLuayHj2rux+Ksg+ejhHXJenC1J/wwS8p0f/ZgmCG0
SuvdjawdJ1XDMnL0QwSy4Gg/XBddQKnBS9RFZiwvhMCWX+vnrN8CrFYnZWzhMmNJ
E22FEdsy7j0MXO6k23Q+V2HvaOgxOpamnJoEautxD98i3IpwwzIyOBFBbMNxyCCJ
7qSbiOHX5eNzkDrsXTDznYUyS4jAsx8XKkKOQmo8G/M529VLKnR4uOCSlTE3HWQd
UbUn3g2nXxaYldpo9UjhqDNsW8FTGByFPbsp2JG4A6jCt0baQmcXlX9qC/3SN+mb
YcIlhYdcJvFnClUZcD0DQfjbptsPRZAWlGoVdOHf5i0QAuzXezr1JygC+lSIFSKx
xHvtwjb4WsYD+jzYRlPzQpWtVple7hlBqEOs/qHe6Hxogfnmo44oZNZ44s6IRIDh
tT1bWK4dlFBTrthF75Fy3DUYWoQQg3zMKK6CM0RQ4gyUc9xnGBYk3K52+LOPQX8v
jtP/mLq28PD5qAvt2Xrcn5gqEkt0vRCYJZ/ThjVqC2+7dlawoRxbHEEq7apovT1Z
nrg1WNbDRjyM5z3JvZt80HJhPe33+yU2EFma6T6E4pT21c7ev/tHkbRVHFbE4Ubu
3vkOVTAusKqAlEj8AvoEREDKEtndZhB240zUSD+E9RRf/04PkSpuv9JqltYaB25v
8MIjBB7A2FtruUn2+pgqGbbFxJNdpBwR+BTQoRIFSC3Oxxc/Zyy03Dvg3cwoVJzZ
0mG9zcN3B3d6KKWvB1JYz3JGPSpb3XZfK9dV3LSZPftIgK1iJVsTHCsYsSYu+HRV
V6t4o69WJkUn0fMS9vDx84vIVNieEVdx/EfuQgnrPVR8bzmYiKGQV3hDfVfuhEBj
qgUQ67S2aU8FU9i4lC4TGgx5bNxSQHJOYtdhB6h010wJYbCpWk41Mpzt8lelOeJx
rhcOCM8z2jE6JnRKSUdDFpRgYL66yk4BMTScFmQFS4EPf6lsB39K2uDoLHoI7FLf
XpK883E1Q3rOurQgtqny9qeO8+6dWW+hcNTQNC26PoWQhW4HuykuNPcmemhJn+xQ
AL6fXRIv5XcpoyRYST0dyBhlW1FeDXK0cyO2l8+d3XM6EovGRueb7S8VtJ22PEFs
znLoDZPC4Ayu/INclmsQJIfQy5/3mNie7HA9VTDSK7Eln8WmEqb/Qo4h/Qjo8G+e
/RLukh9zr99Q4wxREKHZ/PDYvrT/aT1jtze3BejRZF6zJeyP2Y+W50M1erG/skgs
qEOTpg0v0OC3yIwPqfMfLbdw+iFL2cWMbHajg4StvY9sIpELbnHOhzcuJ+w4WMB3
/XIg15NVidCHYVLteYsUB6KR+UUcereOq+SucwbUKFiCPReOhQkKKs9MsHFjlUHC
Q+5RAKkeU4g48Rz4vXLqvf6zjuiLGfSxmTRrchibZ4JftqzfIXK0phZIur4K1ie+
g3jfdm0lCBwTkc0iMpCmzzGkGyfr2kaE/cd+wAzHdAtUqt8ojobzxUueqzs734uP
9QyCjW7bQpgNiqH76mG0Z7xOjIyal26N0U1XLx7WzAnEEZhZv+ws5QxECFscm0LK
Ka0E17G0qmhJX9O64vpJXaSuOtHMPO6dRfyDV0OGS/+pqLsMWbh/dxggD465f5HC
Qi/MRfwp2ZMnARvEIu2UahLgzibj1fPilFNaJ5YqboDLDwGAQmMN+utoStE7nIxG
QmVA7sJIeayMEebjDfulgCamyPjawT38foHwsl8EI1nh+z1cOFaRzddiKBppGb5i
5RawqlFAX4M6iG8+rNYH7Y1jq+QlaYQMourSixUUHHalWH50vWc9X4vhm6Y5CR6x
5oXgHEoP1vcNo8ykEcxHjXG5GxtWwZHkZy4VSKfYIZ3nRPoCfOLEXXbMLjhlPyD2
mlKnLcP5A+ETDEn6vzPJjlOcK5g+UZYg5CrgcqGqjRZfZHrsInbKlf9+idKzY8Z/
T22VMJAQFhQNqphq8rNC36xq8Ug0kImctl4Ql4PIwxjsc0O5ZCZUpp09r4vI0KPV
VxSdv6GkEbzsjqS/Dl14eKcghjgp3XjN7gpCP0pe49E0HkK0xpJaKGgFXjcK6f4J
aKOB8ReBbtee9ZZhFh1pk0zpl375gczayYyIATJZ8oseu4IQM5Z1BQF2wPwJtjZv
Mi6IbSqd+isE2mBeM41ZoBHgJKW8kWfCbP4yAr/03ZgGS+rvYaS3+XPBWcXGKDxW
kzujc8jVMCZJb7r29p8wVHOgU4i7VceFv/rVIrjRlmYli3OKNGEKxBE/GF1V5r9W
eeEW1pMnmBt1kiBmrwtzUuRRMd+KP0Zy5x/Fn++xwt7c2M/ITCG9L1xJvyHmQSlv
2xkAfHp/uXVdEZJIQs23r8i5v3VTi9n/QX9rAYgSVjhrnLXSs5lAr26H8weoC+t4
mFGNUzakv+uyrqwx74VoubqdidATd3Ku9xqobejP0yiWmaNx1bdWp+IH11ceAfxg
63Wim0kiVJGkj7axIDFFBBvOIytvQx/e3vokEFuqG5D9N+lbzl1Hsf8G2C9ij7rX
YDYUiSSAXIDmoPf9hdmW48SOnSQTL7tgeevUgpie0UPSvw533SP55P7E+vcDlzZ6
V96fDvtwkS3RRIUgkD4J8G9tyNAiCuMW4D6/BB4sNBpGJzjo4xcIxM97RkM5FP28
ofFyZw57K1ITkYRS+J81ihaGgMCSxbN9JTa+44liRFGKVzxt9wdlgUBma2B5cRPY
xx1kKp2NBJXl7zmQz7fG6gmWmu5neJh8UfYbQP2Tj169V1P62nqkw16F73MA7VX4
poIo7tsP58m79tZQp4N7GNdzE+okJGL+Zba/UvFs2VbIeWK+LIcgUH/G4yomTqfj
RkaHRQToE5VtCL2ckKRKaeEu/n1upDcmASe0wi/XW0qfvlGJutneHN4SSLRh0rJX
F3/raDmbPTlx/Kinuo9ijmHx6BMSE69DdShGmKnk+GUz4cZNymG1m7U3SF+FQDYk
3XLzDriVTRqd393KyjJi3MCTRqmlbDmBb5zcXWHB5JsJeh/Qq0IAWSEIhEbjwzcu
uu6uq/yEZgA6fHmYEuOt9lrvUUcYRIOMAF1l7KjbKkLe9Zv07/Jw4oQAe/qpiY6l
drQzt/5vpJjJReEoGkl1ByLwCgSk7NH6sx4xGiX7HDRV3mBQmVhTgwFtAzQSr/m0
IY5EXn4D2PraXIfzn2S4d6zvw2KopfOEpTdkppnMpA4QYNbZmsL8WIr9eTE7JBSf
QspF8KAUJ8za1Ur7oMikReq2D0Wvo4HpgbgGPLiI84aZ6qyqXfugJ/uz8BQJPMPi
3ZB6RN4AVHF6naeVgsYbFtFcQLahFgnfhOmNz+SB08idY0uj1uHcfOUJNqnhGT9D
I66Eq0XlYGpbHcfjp8F29l58jjbMKH3jak3Wo/xTSOeW0L3so55AS7ZjlGMBJu1H
VG8MUBcSs08h7yQh71OaqyTvXMsTs8EkcKoULEqcVCuyohKbT+LzrGrbR/A+hyw/
kGcXvlGaUl2FRk+iWV+4R7NFwIBb6ABWYc6jsDFjH7iMwg/JZNwu7dg6y8V6y7Au
NExCLubHzI0mOlBB1jiJ470jtq/2cbacar3zcZxGZUbGx2wR+BAroGdC6z3KgOnN
8PPHSDGqhWomG9+RhI+mYDWbhFU6ktwwpni+nHYv0Bg0s6liwe7mw4blN7be/OZL
vY/+enEnL+YTkIUT+KnfUwiqOrCELf+AiTJ4bRUA/d8dQbtlAX+Ut1cYKIH36Q7m
dBGE5EMXeGOOKSZuQ2dZLMaP6HYS3MzCoDazbKZusBEZK18OO9bUkgnwA/sOzLDy
pLZDhi/9QLln1TNujAUR3+RPQy+UAxzMfJ/KB21B+U41abo+WhCh/DbkQQmS5SyF
qnk5EdLJ0aidiR3yd5issv2vXiTBSLbJ+lo2zRsGcPrsQ19ITD3JjUvCCTP2zpvt
0cmHy+AjcBNmZicQchf5CzVC5BZc68HvGgTcU4xCZnUFxDtvrZEH47Ac9hWjZ+pk
sZuTtvVELu8Hv0yrqJQmdM7dJo/azKgQPFo8TYp4d5Z4Hcf33twkSfQGfHiXyL5C
3rJ++Hr+DPinwWcUXqy33Ks/zWmQ0g/PXYwIebBqdltHegXld4m2dEt60VFJrF9S
lp9xAH8Fp/d2uhuGSx1fOt5rj0H6vJPDMBnM4eenvr1OpPXOQfSV3Tb7NRUUG50c
qXThpDiX4p/HvZCjU60qPtznm7qkHWVTs0DEAly/XHnWoRWkcRKb5+S7Mdp2ADFs
aaRRJqprETidd9nzrwqy0yEGAChR/bPCaGJbjJEhVtD9HItNelMcDPQNaOkyndXs
GXGIDdZhIqiM/mApNftSEI4a+QBHg7z1b/CkJDntEx0fJBHlhNKlDhN3H9bI1SFh
eCz2BRwdNfRsbDjV1mU5fDJcT2hy7ZjfRC4aLVls7rWhDiQ8/yXzWzCsnGlR6e2V
TN3IcaAh2koiBjbMYCu0zVWjw27vhDUr9SDwtl4xf3P17sEmgBHz/yZqQ9Jdb1wT
OiGjeiaYPjmGzF2Ii4M/5QdhxbPiaFyMuxDwCLXfyJi6zFOwls9VMbo3zxh5JbAl
oRISasBEb2LDDfBmWqU6V6QCcHnCYqcaz098Fm6vFRWX+nPn8ydc5F3YaTZCnc6K
dOwj1SyrlO+Sqa9y6XYITPtR6xy65ZP88ZQsMvrb6vovdWivP4BiitMgN4Dyd1Jt
3nCrhfPIHpUFHlwOK12Kztp73ZQeuRsylQ4l3JgLYKtplodk5AetH36nR6aEE/R2
EjbavIiqaQ4cIN4pg+yeabaNHuz9dGsgonK+kNFPtwFiBxgFnShpzfrWaOjmsA+7
qJk+W3JGqwFO8pFQX15Npue6n5ZAhsrUZkBtOKQE3JMcOJP3oUgLt//pM4ErYfst
HOKs4kFAXC0+mAjewP0vBSHCNPL9QSpEhrKTyASp/0n/NXSjxjmesp8P/CF7WPh0
kW3DGBMYrfwMraod5aaOKJ8onOAm6n3RQO9XgI0QJCTS89yfF46U1dMD6O7q6Th7
SZTuGMrCTUJ8aVOjB6rZnh7V7p9k6ESxZMxGh+wV1diHwWQTX5CtkDeXxjgr3JHK
GiRuvsMdusGTZk8c9aEjyY1Oa0tsTslgnZlII4Xg47Uo4b7ODzHm0zq7L7BM5uNk
NI3f4KPy7He+TjvksDzms0l7mcQhv1cw02ZJDOIDHm50jHHvNo+5Kd5tfTbKuXKA
3S5823KP4QglG5lMbx52zdJRqhFVPBQYnf64Hlt8ahbjFaz+QozD8+ES/SDXkCfY
ZwOYxV+IsCO5iykEMjHnQxjVPECYki2XXNv2CKxdvQnj8TVQDGn1wq7rxFJ/hgoZ
pVVnnA/JuOL3AJW51Z4H9idXpc9gQy52jIDhcvrtBNyn5go6QmISAjwtHKvx+Y/l
S3jvOYx8uA52U/dITXO4PnWLWNY0Taa5oRIMzkWCJiiPFjoWTWHJgSNgkr8wx3PW
W69Uop6R5kAP2MP1ueTv9025HmsGFvvTdrZhGRji1LlzF0uGRQeWTNzV5BbPG0Qi
WqIWJA8SbFUICvUoYZVuVsbrdPCEq/55AIa0wge4/QttZc/yFHK0F2zV2s7t/wIE
OeSGl/IdXCoSnA/gzUwTBg7lUxOJ4JA6Q3vjPD8WW3ox4gEokpcd2A0dnIeckyYF
QCyI4QM2j0W10QFiDL3IUY1AAufOW5PU38EGuQ3Iaf4VzFr5yd+IOvX2RGy5DxUf
Xrotwyz8s4aZ4jlsGu5oH1bYteBtVU9z38z2x9aXamHrCyLMpATHWssJOs/9XOp3
CZON/bqwGfuz9skEaOOYnUk96jA2XlwsV4MQz+46xauTELOGIRfF20gypjvQHojO
xzlIGGCI7BN83M/oMN6te05PEJzUy+60d/5cD20Ya3jEKCZDzoobX6dVtYV4dCQ2
tkiR+uQ7v70DCGRMRZSZIHtB0QBB4FOq3buFQSvmW4ThMvSLjk/QBJ/tl4UZ6DOn
5ATszxhRVPiK28MFWZ0eqmZseJ1igehozbqp1tnc7Dooej9kgZYxIZG9Hi7uPFJt
lCQzMKS6sMZBBzif8eugKSKS5dtnpk0R1NAePj1r9obqdN+ca+5u5B5rytDRIav8
+CeyT79GGF2JiWaEPOo8CcIQ12xyyTUTGUBIYCllihig6lmspYsEDtoLzDhOFpJW
o5gJbwVo4Wmuqe+DZLMpPiIzIKNvBSJ6dJAhx3xtzyolAoLdivaHvkjmhpvDsD/V
8Xc30MHawcYoERO443vehtF4T2tkmu0/bv//+X+9eftWl5rtapqK6s91jmIEF8Am
h0UGztLmzTnzwoAhDjmyKf8s91HEBg/DbsDryvoBSeSIToVyYWIks/zqyCGBfcu+
1z2E31fXKYqoTm/7HVds6RSa3K5hrupl/+QUJAY3pvg4GeoZvOUysV1Jbv8+Qj9j
1jMZBNsD6wWmGq5WCYSekt3nUlvQB4ovJ2Cf9y9Vewc/1KsqotGU06z4T3zmK09z
tfMO2EyqFSme4DXeON+aZvQcbLk9/ceYf7P7lWv7JjiNi2kleX5OcPyFxnaUDUPp
/ooMSVVRSEc1QONF0jfNlqHrpz1gKQPieOYDnvxQ3gVhrAVP8bjw3gMMhsXDHlqO
rXdVpboWK6/wNc+CVScc5ZkTO/OyuGZIjGH3GviTMrp1/ndUVk0LHSqGRvNFlTfY
3CUu7NbWGLpaf5fZCUUXmxFj5c3l4AiMYjGWXWDh8m7cAyeS6t13yDyC/8Pu0TGe
r+nMNf8eb0IusLhW6TIifn1kEBHbKD4u7AyoX9f7dykfR/bkLtYIT44iyAldTZR5
4e/z/1Ba+oeTiYXPi+u7s0YqYq0CX6oBeNN1UezZexdnscCJLg3M1XSLpCVg0aNV
eWMesU4c0Vr2U52AB9WtqH8z/kzj61NbxMIfCGVCnDRTbQHancoSXHI+TVXnnIsq
qUl+5GJZy5uR2AHBdVN92It1bm/+4+2hPYf5a6E8LweO5M6sxyUluRGmsVUSZHXy
TMVtCuXhTrcVWlbUyoRbBK5FMvRa9DBMxOoayolXt9fP8DtIzouWbQQvMWvLcilU
jvZaCVNAFLTRJjJGi6vy5bmnppa57fxKU0sh/lbcH2MzclrTO+VVK/lwQlb+s4fE
Y7q6EeUvZPTOO95AruIcksgDNdhhZhtQfNORDZgAqV6REgq63+0ZwJdK/A9Qzsiv
cANaaQLYYHbn3I/E8R2pCk5lh+n3sFm/75ZXrD+vgdNQfZ2WgL8IUU4rt1Yo+EiF
6bRIId4n2kRt2d/3zzvL8JB/wrCjVSPsGre/dRo/6GKS+iSTdVqS/5Jm8uBevTtL
0WWy5wik9q7thG2OeYVDGEmYn1vg00zy5W13pWIb+Kgv09EBJHF+0oKZZbPRFx3V
l0xecf8sFwC6ss9AE4IEMu/Ik6Aaa/Hr3Uz4sIYiWHr9ZlYRX02kppUeDBVwUwqb
1zl3hK4JMzHVMUORrZaaJxXwZxhXvTFUqQ6Uz6Yci3QRNRjNTPIq/Se4GOEKsOVA
PumFwSkkV3Y7fgyGtxxSqmRPgyAGIX9RylZQOvM5fo0lctyYyYtVyKMG3Wn3KGV/
+OHjGa5s9q80T8Xp4g517E1jQHCxtDSVTPFR/fo60k6IvLDLQg+xHJG4bsR6v9UI
XvhHe20s4EFhrD8zFpxw1a3ISDhfwpHVCOffEF2ysKQpiuKmwWA/HpfP5TqcuNQU
/liqgGfmyngCcmvv8iklqh8WSi6BW8NEBTIPv1/wBfvkJy2v+Ys0oOUGUDHxlMcQ
2Sg52AHqaDfZ7Q0PS7l2DQZTlp0/BJuzAqEGXJpUpmbgIfh+1k7q0VhoWYhtN5Zm
LawN+hfqNmhBuvXjfZI7YoXJ5vZMO3LDxHxTWQjxfu9TsYJf6gZ92NBkske5vJHL
Sx75ZHTTAjUdRAu3Y1XjZf8SHo9W+4kK+C1Vn0YVNfSIbLamGIvnXhlCZIAcVC9+
8KWAKW+4ARQMjyw5TLL81hM1iIABBKozwk+EboPZe8RTGfGOPhaA+xGAQlqcrM00
HOluAVksOFB+AVXjOtDdKy7XpMymlfPYNQSKJca/k1vKaKWtV1rUKKJ1gsBqbjzK
PgMHZr0rwzXU7abFTovn66so3/xGmC00UAIMYcBQC6P90NpPxSwcglHo8MWgAGbo
LvQ/TbomkhRz+apBtsq2ryZllbm07nqffonZtD4hnu0MrH8EEPBJoSTLDtgLnAhP
pHtO9+71OfnPtqrPGGzgv5kWH9ECpkRMINHYii1odRluxAJfepISZlMo5mP91DG0
Pe346A0IH4b/rTnJY1f0zFOl8KW8+0dJAa+SrfGUKFF7sE1ZpOTu1mEqljiWMkJa
0X/55wI6jaZXFOzPVKjroHXXxQJMY7hGlrkxMaJwp5VShpSWUlEyICg8iOrF9AWL
d4SsqzdKXVCsUQHRP/jBW6GGzNqJsuRsOup5AMo5JHED4yPvZf5/JcIFVHtMKpBO
XH+JKW5gGfzplEwyWZAasa/6D0UINIHL+48JRbfdUwncb+UPT44Ez5i+NsbgmNIR
RPoj/vRkj+j6p7v20fYW/i/FmrNpNluwTk1dQ5PZj5L2w2kp2rFSFE6wUJsEXHDO
gdMSIr0w2hh5F/8gOVR5G7iCdwXWKRqr5mu/zxQ+ELKW7EFdpzRuBABraxJwuLHk
duCTCIqNs23UfC4XF4ahiWEHsVpsbhd0Ja5Eb43uuO101J1CyXPXfVyt/kmHUkxW
cmVgV4ymoQmMuVJ1sq5m5+t3MV9bvWT+PPJRPXKtsLDz+WI3eP0vTi7qifjpD5j3
kv8ztIkt9+eazLr6LOKVCV8RTO0poRbFAfJnGSLG3/xSBH2Qaqe3LyQq5XyAIGHR
p/xscS1BejEn4VfheQ4M1rhGIzQAnXHxuB8ZWWEvcFjag/i8halhi7NoqbYgtA1x
YGBFgkRTU9jngKVR5bnXmjHP9OgizxrNLJIrkfQCRi34gX7PSHE0hokjhSn3ZOZo
Kb9p7nzJ2WUSiRnIYUJ6LyIUzNjxc2HIK6Ro5RWByMxhMFe1f9qaoUlPovshm+Wq
g5TgIfayY69iKR+V1JqiO5zJwFzbZJIS3QeDPwUJmknSoIb8kJaNq1Rmla0qDxRt
0jM+KX12EbC5hXrtZvAhhU8EcZH9UCpOTd9mv4X+nnlfwQ2nqmV19BWN4mnnc0P2
B1KzDWHM1kKDh6eIg7VDnXUMWhZQgDnNzvwv4/m8UfZGjkV/r4yWxvm9YDE6LEow
NnV5B5XrfdPaejRLw5Fy35HYDtYGH2xPL/xg/yTN+PKE1lE2Tmj1XZ9MzwgLshVC
lxGDzJMIgenQ2tbb5O4Z63qE33q91g38/g/GJ0DY9wTIz/kMjfKxAflCgeDtESNt
fqS6tnp3osT7y7OrgvkJPj0V8bDxWK1wqpc0OBOK3NJomvFjZAjXnRFE4j1iKWwC
/KwU97fiEvkirDZjHm/SBWqd7NbHsdrOd+RLJBeSKoCuvbkYVsJ/0BuGmKCkJoeX
bSk8TrlU9Je3K1Xc17JSqjSSNVxSs1Ug2drj7c/WciPfeHiZA/2ez/IhyzISlWaS
z3reqx8yerXU5e0IcCw+BgoXsWuYa44myXeP8ILn07Isti80eJW/AcNv5lOlZBG4
/vLzOlIwdKNh/fMmfZ0oxU0ZcfsNy591BABvvp6f2YlcOuffohfNebXjEXtsHO3O
3M/130ob1QAaHDsyPx7ljKn9rKGHazuZgRupNqgMwwvbyK9SrleF5zYnQJY10huO
obHu/XPuJyBLOZRFVYDXWsPbZM/FCHAE47qWWMFLF31pcmvZt590vd0//HfsOBE3
q2LHeTArFFUE6RIU6erRFjN5fg2ddT53J0KnHKq2mOs55WwQIPxQqiMGlpsGXk7x
BLS41KUpnNrag2hCmbNWogT77akQcTlEdz5AVAWQ0NmDR4nrURX8hIz69DJzhdT3
r/Mw601SKRjRXZ8bim1ZFGEzN3p7mVjWgjRNGYn5gdo/t0NLLP8LsuX56xNNeudb
Ko9fDutjQ9TOKyFRxtA8XjeCD5hdH9W81+QB+ovFQ1OJYVXjfPHWmmxnbtEcZ1Tx
A33TmWfrCfbMJjpddsMTNH3euJ059OqLsTbHiNZDk2rEBwInpdBwlEGbZbSagx7i
4+CW3wiqgVGlsbbX6p4j6o9NZEUayuxhgnvPb9hqB5gaJtROPmcfZXDFpDelier2
0IKXIZLP7GIeA8CLXkQCEXlrOrgp0loR+iNm1jTwQozO8azjdzP1dw5e9y1+Blox
srlvcGeWEK+kYrxw4p7HnQD9zfgtxrGmcLkKcAGATf5HS3VUGgsVUlDw1qgEC3Yq
FZuHgHwZsWkk2gx8ipWZ8Ccw4mNnb6WvX8WaLXBsSskIMDu88Sh6w+0coQ7pRUVB
GNhT8IMFP0ECwoMc7nKpHQbqhBeE4H+ilCdWktemQve/I7BYDyfLvVZfpW6KTkmB
6J5yPEVMz4W0SVsCjjMLK3Vo/t+rKzW4LXu/2vQfvCAVVpnCoMXnyzJwzC27bWSL
5fNX95Jj5jFR1KmXz6WNs551FstVYCnF4zaxiXX/nKdYSpmF92ZnBz23puxnFHR4
bV90O7sFhpc+YX/2jxznVwX+7iWob1RnbZShrUxDOr5aJ88DUc9jR0tuy4V1pDQV
CkdLpK8TkXhFhojxeuc+XsO+BehUJ/OTTgsKGpKFJMmDHnxCKQPudAG4/GufSBeR
c630G6eB5UHC8+oh3gc0BCryoUjD7rMks6AXuLcq3YOxk1ZHPuuG+iQ8OrytODvH
hq6q389H5aUxAiC5XJq2I8EMbnOGorOMkpuy8sdhzqXK+u99B8VK+NfvEJxVw/IZ
ryh8qwr9RG+FAKYnpAYXdP8bP9jqidgJUZwAB5QOVKKVvxZnQ/ODx9TXiQ9w4Z6M
bKAhmeDP9DJnO8O+XnLbEycZX8KFom0wJRJpFfsmcVSa2Wo1DQdT2WyoHCxbgj+v
ngL+pPMrRmh+dRSws2FBKbC26YZRCyP2KbMXS3BJmSCBNIHDP7VM1u3j3nPMIrlt
gvfK77vIoU1A89Kx+AGTMVKxYOV+R40Pk9mitTyB5ds7hE5kgISquFp3GPWO/84P
TQ8YUqcIATBpZmwZx1OfM72ooJqHvJ72bvVUrQgfx1Uw3YKAVUVXwjCLVUcu2RCI
oUBSNDlBKP4Q68GMCtX1Yp7HkX0kILGgIPzIr8W0X5Y+jcY2D5xIpNJtjAyzqYME
pe7yoBMj0xh7ce+PrmgdoJQA55LmTs+SNFHm8c5VHuC7qGwWzXUJyVJZ7CbGEyWM
Y/z4caJr2kP/CT7qxicT+HBkWgcjkfpP9S6Cfwg0ixM8oQNX5phzQnrodrupsq4A
WFgU+h1WyNAdkjy1uGjqPzWl+EobBNAWInwmpVjGYrn2UYN/4arML/efOBdRqE5k
Pp/JtZwq3+pSqQ2w0s2ZHZfx2zW6mufIOgCa/fGvEtydRyH6PubcgnR+XoRHdWtw
7Hh6xZ5xmKxGphgOCoI8brmvRG0dTSH7PIedUDeSc8xBmfoVNNnfEqZ2uOPgDwkD
5y23+OiW5mC2RFTT/Utn+4Tf21MCiBVcOHsKsCJ9uD6RWxQmgkZqliaH1wpTrEGd
KGDqHJxsZw9tWUALIUHXsQF+kMx7dBK99kigGhlcKgXK/IXgASlh96Cr34ymGOs8
EZRuu2SGKWdAoZOGjQCGEj6tQ2GPeVVp8bL7uCnRLpUB2LzjkkZvzJlN4rssFFwG
F+r2QVWtMS0zhg9RT2J9RZrsqdpDuuuD2LDn9eHuTyVygXc8c6+5Dd6GaSBRpgAu
DaS0UjGFj5W0AXBhXdtgkjxfxdSXX/7Ynze1+P2U+PsXcHhAV8Q0fpSTSqafBKYH
ru4brTigljr7f1v5AwIQ9kd5iqeZGu0FDN/9QJlJMcFd3kSLZRjhXjt9FKBScfaq
TJRnR5CobL5C4Zn+KyXQs1/15qTJL2flGRP4Rgsfkil0IhtKIQDrEqjlX6hBgi3e
kcP/127L8PUxIS0BobPPupm422UNAluRL6EHI19JOmjnAQ0CUR69TWKWbz7521MT
7FLQ94GydbRLBMTHOQNtPr6IELHrBhFTzykNZ7/9GNbrBmbUOfBsmO3I2ZvqNstV
st43fcXyeJdVII4KYjsxn+YLovAAu0SPfxHxZLRzJWgCIPTk9Kx8Ve9gNIIwUYXG
iGW+6UpTgEqIzXnPLsJJGBrnS7VgN/1oP3DuKDREbe+tNDWenfnlrkWrlFQKn7M8
dB1E30UrNNGL2NC4+/B5NdvFujitJMeE2PW71ALrDnzNh2frABC/VCvP814U62gE
7Z/SVpbibimNnuRSQFgHFXUX/+XXMDh2S7X3kViA1X4wn/UaMgE+ypBjp0STAUNV
awQnCgFosmsZ3SUPq492rZRtzEevbePVjz2ZyPnF6CR90+RepQkpRWAPo1Fph4V0
y8rut94HjhOUDOEKqtesj9beOeUcJBvsC36KSbTn+1YRIdxtsmrIEWoihwbQ/EVQ
pN+JNTlIYn60tw/D/9WG2Q9Z10GJJSbMrxC08elwKsATm8VfO8OmKBCy509aGEbI
b9hwcN9KXVRwXQk4txNaSuDeWLjgHKcYWaMqvVkEbCxfJUk3v+EcWPKJFi4MEJv7
fNOWeOJ9MV6JScIRnZL8zuRhnHFPnuNkPCckUJLNeiDlDwNei1mVGb/BciCg0puC
/td93wspwVQFmjPu8boAHub7l2+tEjzpAG9WAwf81pMczhTYbDbe3FD664dKjPyp
w7y/OYhVMmR3zy6UzDSZXlPmPP6hoC92PFuB4LisMtKPYVrrNCeOQtC5QsWcnuT3
MUt4N6y+fwcxjT7a/9qie0NlYQ2o/wodF48DnPWI6y4Lpv90xS8Oq27anxNp9kkU
gvIUbhS8lrSfVfM+20AzxdSxLDJR6ynSIVlUPEZ9uBvIxG4M/3euBe9zAvh9ECbN
34Q/qBepOgVvI/tb7fL63buwTG+wsFMZnuzaIoqcGRAQ5V2C2ihIkffCMWz8Spe8
oklEPNvko3hF6WQZZ2aobjUAu3g2WKZRjIppeLTxb2laNFffUFE0OV7ZojNB+ALd
1Pc7qMvLC7z8JgYXRe49s5PrJeYh5f4DtSnaQqUp4onD5N5NMqBwKubmdJX3l2bP
RxzMXE7uxisIP0r4MCA0tugE+pQaFqQBTWBJDOS+qDBtF4/u0Po2x8d6+V65evxM
KL8rp+VlAq4J/E5loEXOQNf0A+igRfTnXB+1dFq7WWwuWwO5O6l8hYcOSdigubSI
B6uIYPa8zQ4RuYwdScYfXEyGNgCtVWd37T1hL3i5t4jvzgX/KUjKCua5Tpr80VeR
8BSt2S+GWzwWtr7izYwNb+W4LGrx2cm9F2CxFOkFi8MibLo+PwPjg/WYmsKVymwJ
494XU7yg8Jp3fee/4JR5e8VRriTohKvgHrclw7SSq/+lwM7oZJKGmxPbaYp1/kEe
E8vwvACAMaqRW46o5uqBiIZc/KELEesiDFqmqz8nzQayW7uW1xe6KaIozSWS+8dP
BREyG7NbguymR3O97WAJEOpx4riLb9QptIqRmszzT4Fiq9qcezDKX6Ia0Q8amHaP
SZ+sY2+pCn/KeBVln/u0Jm2w6gQ3WBnrgmRyOQhzd5eTjyja6Nr3wwNtdPFq1ILo
5i/wQ/SWTMwIFjAcc75QqL/7BMKozm+WrbbC+WYf2pocjHOTeyPfemfhsTBCh/By
E9l8TT4c8VZ2qoXyyGKzpIwI5CjeqHHVG57/++/YlmZn2w8MmbZHmv9X8Hji7kX9
L2gRnZ318OCSxHtthZSvsC2d1YiCRch6U6DWNa4yLBt2Kmi2sSB40brklbXlbQuH
azdDp1j3T4+0of1BDHZrZyRsuqPLD6zUMhPTHtj2/IMpax39QCAlsaAUNJEJFovD
kR3RANolnUYlq7nYd3+nYWKszKbQ6p/qKgd6CyLmSleiUzyf8IXGmrlSKVFnCw2G
UB69phet1AjPdxn5n53ZpUZ3Iy3//LMOUY/piPu9XVV0IZs4FkGvsUXi2OMvvovD
b/Z5uzPMkwfueFxmYhJUAXGCHvf1MUnPJH9DzfmzLUKgjOJ6cz94ccFCZxGKD+zS
ctWodi8QXm7Tn/qwzArhwMtp4DBQA78d/Dh2ps2i1W6I0vZdr+VGn0CYu6haHtgz
dF1SfkYkb6CCBaPG3mSY/3lCkl6EGcff3TKzxyfRbT4Nt9L2E94uZNkCcO9l27Dl
E26ktBQvXXqCD18QaovDILStoUUQSBth3SsK6aaOes/ADH8eDD5EPVhKj4tiqCmA
ZnS+j4XrSz4RCA+SpURVGf6uPFfoZ9K/Od/j7g5OP2KYhyvzf0D+ZiyPMqh93Q18
JqFQJKc+LyC0HjBXoikKLOiQybdPlUkvsxzhYPLiuQdB/gipX8hd0wnpcOU+TSOx
ADqXM90fGBzK3B9NNR8EGjkTNZEmiadu7bN/pKP2Jui4d5gfyrAT6IW5Mxnza7Yi
C6YEW/uyvL6B7q42Ok4AVH2kNA/1VKDqCqyCulou8KKW2p8/DtRVltnBuWiGlTnj
Z4GV/U//O5MaJ9DmhiT9QSP32IkszKNyAb81Qd7L3VYL8YcuJcpKHFMNVOvN67V/
OevafCSLGCZV1Cr1K5XuTBCTXfFDd6Z91eWp+EvVCZeWEtLW4v2rFk3gKSiMW/x0
fyCtoaLsvqRwmLUoWKMgiX5e7gzHAHWuBA/UVk7E+kEZUX79BZvtsg3wZafP7myX
TBNJWR0K8anitnHuGans/zDnOV2gaXmZp5oh+ltquZT6kKNNmnxaDGrU7By+WIO0
GrHxeZy/ThSElbdTOw/NoV5eKlZPzmYpQCKkU47CPZukS5LvU1BztfRKAbT0XqzS
t2SS2usgu+4JjF/J83QIEP/WSenBklse8Z8PFVD8h5OBLy4l022cUVzq3xcfd2yz
1QlciJ595CtfRlT/pi+w7KvSxmUBUhCvh2ob4khFN2cBS5A4h5jGTL8v/hGc2WoE
G9PjASucwobeEF1kUNB2vYffmxVLDh9bJgu62Htoy8HzT1rqiI/oFwla932d2aAL
CL7NUcsJXJttKFyobGgVe6hY6xgkYXxabddQE0Vb3rkHJNkzhsEct1pt6Zz3+ixX
z0lpgJm4gb8fSsZ70nru31WjLbelTIIhC3emyki3Mtbq7bmKENkSfN7KuRAnbwcE
2I167UFv9BXBhtAClJaq9QhFcMi0chbxDdPJH6Gv4WFJf4jssfkrpM2LlfH1uzwc
2LJgYF2wIHfrf7Y25Q2+wYX1G4/TOavMWjXRBlSP8hBOvsvnU1ooKOcyl2czIuXE
VASCRl/8jPYl49vqB9iReGW7LV9m5tI3w/JNNKZsEACK/Cau45wZkFvYCk42LDUA
kBmCWDLMx/Lgy2bEruac0CdvjIAsLWnN74nwwczXBn4wLrLxhaYLuEm4cQG9yj9j
3lnUn51P9oMz7u40eiZypvIAIWsrtkwrXqjgL3mpqYoftBfSoro4tk/q02t06doF
FD2n9FXPmIPIn37ooMIHhx2e6J0AZmBgzSBXy3lyoE96Xgk1QFOl/ntUglKqqe22
7jd1VzJxLUjjORyDbOR3XT08KAwCuPmGm75TeOZZFmbREFOQlC1xfL11OYKHxb5O
aYlszO9iixpj6vAwOCDH2kmvb7v4NRfykWqaxS5P3HhCG6B+DPnmvYaB2dibO2Jc
+IGrHITY/et7jbAHVMiEgxUEi//a8X1zx89moVCYPUDLT91BH2drAxRA+eQWWRGI
ugIU4rWFUG3sZ9vL32r6hPiXJKdP1LZsV1ZTUnRq8Q13YpqC9+cyM/hpKRSWAP85
ylPCa3U0BIzndncj2wT5+VjQEJTqhrDHI407Rm8TujxgC+YB48SBv19YNeGwp0PW
0F/3G/QJvvktrJ8B2K9cLXSZf8BFIumnHFdZwOAhuKnwTGdybiNaETCgJr274Tfp
afIhhXdJDHS5XC0yD8Ftj5hw1hfLywcAuh58kRWyZ/KVzkuyuIO2UC7MTUwy5IC/
J5EBDdLzxAtl0Y5PGeMNUuAfbeso7nzkjZwfCFlu1jHsm82t+Ffea89o2Q4jZ9BD
yWHAC8RU8ypaBChZWx5sabLJ1RWtRXDZC20ViblTtaO2muER0/vhLqb5eqIQa8WV
jtfRbZ6XZCzUjghDxUNw8T8mp541/jykAekXq1/pweZ2h9PMJC4iEKhUp54xIwXD
FZ95QbXeZuwNgx+T2Mpl0bJkxEYWh8ryI7HTHDV63w2yyTbGvMfjhKsz89+4GfNm
WgclHFxlGN10qvFKRV1l976zSCjV0ieG0L1FMGOVtjiUYvpG6TGrad1FBBdsFS55
usAjGr7vOAjckX9njDYjTewAIpoR4s1mHcnZZcUdYG+rCukct7nf0Nylg/C0H45l
f/BjtU3lO5mpiFW4zSyYr/6gmz5Pesl4VYoy7NyjxN+Og5hgf/key1whSlMQpuZb
V6g+cidR5VEvHpCxEYReUqzFzkym30+twYB0Aoxqom0/Y+d3B3bAgo02K0p/TDkk
OR1K+htFz2J2ANxAJGSdBjAHkjhpi3Cy9ePYb2sehr95sQUJDRUqDBufYhBLxsWw
V9p/eeahCxelt0i9SfQ6JZfryvM4ZFpecqip2OS9Feo+vidJZ8VcJ+3JIp4N7JzC
fJat18UE+kv2cE79Q8Dv4uLCuOOEzliptgjLLQEvRF25/Hh7E97YeOSwrglcFGeN
uSUHGKns1SF/oCETJKNKzeMlm8DLrqAT6kaS3zzk0DWCtlAYqZA7xyg0f6MfoDwA
Lyf3QGvl+FJhX7mxAHMQzjSIT2rrvRO9nwZ+VzSTlLtQGOZRj+djyuYSHPtPlecf
uzYKzyZGRxVAh5lGU8IhvCNCQ6ivAe+d6vp+nXIgOa8Szo2ijRxKf2EK3EFEZoOJ
ipFvpgvyNDu+nQfeLmXqJl04IpbBXeJFplVxcrIZ0QTUJ5zWne3/7wP4PLU35Wyf
oghwVc6PDqVF633CzJOoWtffyMygiz7mpfa1PrJKMcnxLKrOZyGK831OedzAlOFW
bRBjYGHLZ85+KdNyHcXDO136ZUKzw6i5Bump202Dg8RL7NhfTO4m2vfENnt77C7Z
S5cn4cAsbasQz88c5BqJDBIzzqdDp+dCCsqJI1e5iB1Yd8HdcJJQs4VDap9xAHpY
r+ZoQoQOXLDRRuk/7kqb3k8b/ESkxAWRkuYRcE1Ehozlqw1qznyZvBhxMAa7Fazo
2C0V3WrPoeb+KkkVBWEmnarKxRMxZhSJrDQj4C/qPGG6mklUhWNV4VEAwV0iAG45
OUbjlgQ8qvz3H0KZKkhIZdqzkANetW7JjX+8/TC7CD0JdjbszXfFGVmOU8v1/7OT
1VstzqVM7PmTHJPCMy04oWr6hKkHKTZHI9HacRmdXAwUGihU2kx5Ek93txpK8bEG
LI4kbW7CC0iXxjPsZSD4H2VnNCJxti+HnsbCZ+p2zx6xLBHh7DiYqRs2kbS1AmIF
iPJlyggXujgucznnufLPWnYdTG/EOLHJhKKmPFHH1acgsswF9G8HQI6HuXwjg1AA
D1/oLPkOwgBkqQFhvoqB3qX/2fWjs8HiVngyYqXo/V4QoxWV9YrBJjvQioKQjonq
78aSyw5iGzFRKCY0FgObCvOK4Vzkf3LW1UyyuspmTjHBh33sk3r4iAwTrwb7Diws
aFbWy4HQmpie19YJUTGIRJdY/HTBAq37p1NSeZULrtoBv0TpNcI6KDPlWMgHyYMJ
BznbLltbOLzGlRAb3oaOs1tf8pSd61v+aSC4V4aG7RvsDXdqCdsGGAw6Pty5Kexi
xc+RKTNlSMTRDiBQ60lU5qF0LDHpivRzglU4Vfo+ORV7pim26iu2s8ZkdhsLzk+g
10XlffdEtn7ULOVCVbVZSueM8ryw2FqGBOnPuWHjIJ/IkyLjiSWowMOVUqB4mRI5
D/sNAoojtsnDfrfgMt75TxCLTk+O9dORMQg9W3R5yRcjh9HitrZHbkLx/gOH5d8c
37kEerWaME64uxzHSdK0dqrb8qcwjfYEoU3a2S3Ltb2i5QXBmYFEpr9I6R82kSU0
igxmKQYvFzAUZNN51kjZ3Az4sSs9BqKOMxi4CIbJWz6p/15fRoJ3b11vzWRlimwi
Ighzvu+iZKGhH6qE+AictSkeu4SE9DZWwfd5t9HcqRxRk9rSlfaoz64Ryzw5Bg2O
sz+lrat6QtYZt+kIbDdJUM/QUzf5H/cfVedhxKLO5imw1cYHHhkEde693bPeMHQU
n2aX08xseCpLw9zpRXmby+/oAFhYWhjjcYcBfmapEx1SJh583xk/F6niyRrQxVSD
h2xlWcFHGWC7fsd5ZC//RiV8FowG/gel0VGyBxfiEqPKHn30lJaK+JuZulkYffoJ
c23siVEVZx812St1ZCqTLEbfJQ/09XpLYaE6MEvB4MnNkffeDwL0S93YIYc8vKS0
Chw/ulk/LMgzDEzrDENDsCyx/LPgwaZQiLBgQD1nsKb6LZYZMQwscYkawZ98Vrhc
vefhn+s2xveLR2LMUsRlj6exiCI60CdP1ykQ24672EwJoIgkSs4WL7v0AxOVdwsD
YaTNuar38jc+V+1FXEFb4Pm75ByCUV4nf0wBr8nSd1JYuhmPp+zSBNTXX559aBkV
NkKO1zWjg24XH1AECmZjY6RwOrdRckW2tTXryEBRc43p2gCEzS7UfJUgUsMPZSrh
w/JQNwRpbAqThyzLFdaEICZVbCn9l21q1X3lJCs6UllLEMVflwDbA8OdsDaEuw8+
tqFpLU6VNLNgDvTsb8akxTnXZRqmbZ+ni29Y0t8ioZ/kO26NTu1HG1ypPxNyoimU
YR8TwvspRY+yU1wsDN94YDUlg0xQfS/qoptCUQ5gLj9AmaMNO05ZixNEkksik5gB
uTmO9yZbYhnpXl/bIusebfqgXjMffe3EaZ9mESNvJXqh93NXH/yX/3iqygMrYkX/
R66C0OT+/j6N+MDzP7VSJqNNY343n39hsWk+QiWg5syAek9LnHjCljEh2ZmHp1pw
onvJINZEEV1619yibg18wJGURnbV+LzYNpE/oQvL3CTCxmiIFzGvXMF1UeaS/Gwe
07DSzspdqRkXZsW2TX3T2mFKfGT6JXLAu8crXsEAmfUo7seslhSqON8MLo/5EXbM
5vn7mZNyOxCmRjo4BcKRneAmxwNlSFz/eytFdimkbyY2nFMa9VQSvt9aynJbBXTl
CjBkMyA5XuJZfMB95wUpJxXPJ2tA6NX6GU+ELbBaTzoA6PACs+qczCd3xajCC6xu
DAh+h9XwV/+3coBGYM7Eg3ur0eAYaa9oh+tgUwcVhBpfOGVIVUdW+fJlKzE2CCFo
+uda2N6PFImZ2LBeUPiFlh4CDwJdnXYzdaEzuWq63apS3hvqtasSM/jrtsefHDHp
DK62t+BXFcqXwD9rgGb8b4wUOtJ3mq55V7Ut9wwFKtFUpjuThLMrLdyNNm5R3uCW
BdAuoNtudtWSQyxQYvEvVPNmhmLxm1iOziHb0PjtHqd5BP1iKTMJNITi4kwNAPaI
Tbc+HcJTJJ9Q50G7a9EFmK1gkoOh4/iipxz5LOvlXPnnxf8ShMDeUvsAFCe/LD6e
wRIwxngYciX+w9TgqufbpQvxMzpuge9oPVt0mj7aH36z1mDOjXTO05vMCJQesVhM
1RtQq+vfipm9KjxR9+KmwpIeY0ZteA5rxMTNMeysw52jMyH7r7TSkhsDp4vsgTpG
D7W+6wP/qtv9Nthy/IpQxg3/m+QU98ssX3vt1ZHOiz24noyiokWMau1fF52jpYUz
u9Q0kS/UUnGcn8qRb9G2Yw5XDys6+J1UZCNaWdy2j7+dQers0d/STcfnLgQyAWcZ
TOXUhWLm5TGVm7jIjeiqD3XrC/6YHmgFsvgEbSB+y9cMNNcxoH7udCQYyLM2vUc1
jPlG4rtnbHxa+buHWz1eZ5exShOgx3bCBafwrMOvKjg6iFdeiWhK/xGr58SZ8wvR
vcwyZsu87OsU+3tVegkNG6n7dG7fakyrRcdyCIoKsnqVKgicfdsMAeP78ZdtTfu2
01IFoWuN5eYg55e/+3Nl8dxBP5UDiBquNYRQS8lNU1QKtgpRimtJ2lZPtwkK8Ifn
aeJpnyssthGLu5Y9Q76fuHVOn+vEB2FG8ZQd0bGJ6gSKJvNRWNiKvDcAZqGpETPf
8aYuhGJMwydJpSqgVltBOdYoG/3rFI9XHx4vs5KuAixbUHIMFzjztyUBLvxa+Zsq
vDNr2INjJrolNo9N7MJVm9ThNQdIkMBT/KuVswaJckrlj5yg8uyaHCVuoKlXqtQh
IEFkg3XWVEPoyhBbdi8ZWFpl6u1Z/M/3OVUEqY1ATozbegxels6woGGJAbpshE8A
zXkDHbc7PLXfdFTt2ssUZmyn6U5E7RlH4yCtP69PW5clTcw9BuCQlfkHjOw0VGWc
5Sjy/iMOPxDC2O29EYa7TvIK9gvDNoJQfZ1z5tYYKoXCOPO8rIZjN6JIkXNKOT4p
WM0vDvtikfGvMsRq3H23B9P9KJ6mt+GKTcPhOuxv65FrcriGHZVPk2/bBZzGxTY9
5GApaauTbuLjbg/8Hjfm7H5pQETQxBwrqXhNgcyafMZ3v1kkd6Eqac/cM9weDzT/
Q4lg3XLPJNhghWXqgJa5nfOA7Oaya5yLtpsxq0Y+0RkFViL1sF3Eg5kLVVErY5cx
NAGic1lWOFzY/rG3AxgrRVu5CEPxVMfcFBH+yq+hKSklnsxvf8NRYXDyA/7oMSPQ
oOIEK/i2cM6tfRfzpDLzboiARsYHlkI9rnZj2nFhcHfccqAUMd5y1M1CQkkKx5Xi
8K3oxFfhuDiCVMw8aGtGMXFBjE7lukyrEtM0W4P4xKQLCd4CU9VeiZZApGtRu+6t
cm7lzxwXzdtQZ9uY/0SF/zBjDGqMzwQjKWfo/TC9b3mSt9UGPgmhLb+KnARNI0Ag
FjyPFEBZcS4atkMDV5b79obyIHDJZ8Me0O3pKV6liJoRloiWE3D9XXee+qaZnQbP
kPg+O3OgBn/z37Q3mGvYDya3ncO8RJbWgG3fpnqkdBsd4C646EQiXzan9hIOimXQ
Z+Xmn6P8athC6GngnhQelYAI3KIT6UFQeNGkkGjgedjV6+gj4uKAl/DW9wuiY1Lx
AXsHYbOG+/FnJk8YezomftYYpaPh4a+vEgn7oiMMioZxQKSNDPacIFVch1zo37ey
jZ1uHM8vJ8B3RPyuu1TaUR0dfdC+qFBmICYkcIjnHtQsTP+xY/JSYUq1uITdoGHl
sZz7KntPL/pGq4Q4f5/wvs46vd/DvT/RMX8oDaURkAUo85hLnG1YtBI3HWbyMcvM
BGQ8/rWilo4tyTqQNnlgI+l6n5rZSTpnyb1ZvuFpAt85dZWaTf4bHYIWYzqb7c7I
jaMzphu5ZqFh6KsR8lbXKUG76obJzZA/d+QTruzUxAT1SRtMtN+07p6rxHg8B0W6
efXlr92HcEqQzPal+uOJUzOoTROBnBLXvy+DlWLVPoBdHZN3wnf9i/xozkepPQqY
AJZL+Z/BC6fjcCLdmwW/vxJ8dyVgEjN+njl8u74QQaJ3kMwtBXS6/4UYFoc80qWP
Y+Z/fqzaAvvblcJXk8QeeHS6QPVvCrdlWq2znqwddlZ2HVX1fsDeB8FzPhf2sTSI
Bz8JPGKg4lB9n1lZUAHpYLDUIUWvMKQbmqPS5+aPgTmUdNu+WyfkK1XdJYMbg1er
nbGS8FShhKxfX6jYxhsVMDEsAXP3hjPXA9b6tc7mv6Hz4fbxrGNcjtCP2ayJPykr
gIykB9oNr0TCub+bH9w+EetLhXHl5jGNqOl3H8XgPrg3046NhlO0xwN/GjOk/TJv
rhGfxTpAm3yTezxVUOd4ZUbfbluxXG0czUzlYnH4jnFy6uxPq4F0zl9JRJAp/hTo
jwqPhn+KxpdfeXF2Jk7pkxG6WcxeO/PcKz6e88LxGcZaWtTOXSCswIWYPGnU4RCU
oCI75ffBDtSIuw5rJNHdmwR/QOOYy6GKyueT5X6YNpc8LYWLbwGk0/RJQRkGGQYm
Fc1uvlr4XYY0m+yWdIzdzWt3ptyEajBCLpWPaYO0HMXxvFSEe0lYnh4wr/dz8pO6
KoK5dlfIeB+QYDdwUMD0Q9DDa0jKOcC+INrun4Sxp/UUt81bQ0+gjanKkkcwXlCW
DRB079v9Cd72bSQXsgCGK1OljtePuEgQyrse/4xkdv5Cdq6kpiubPpG08YWBlyjd
dYgRDeQAx3DyPqRjVSiiiY7OCvbkh+rO6WrnX95dluFcIQYVAck4MnNKxFvnnxNG
mZZnMd0JaCMEbKuG2APe4pmpq769jzxpm5RII+xkFLi1De00bXtqxFplJpVu/TLy
xZmx7wNMBw+Ab2W3YTEQ0m2thDeCYyjwRObCudMZBbLzYwbKuBBI33z5uPrR9XO2
ox4j/uwzeRrHIJswwBIByX36+/Q5NJ3izYWTleGnXuhsZC7H1xwd6ybA93oC4KHG
QpyHeV75Btt+mhe3xJZA5fLnXMDkuGc1wxdTxeKK0NzP4YS+Xks3YLPxMcJtaPoR
9MxR4E7YAEvcCb6nUJxwj9tHVb79TrOyAqOlb3bFkXqX4oy78k5jCaa9hTZTgUAM
SI/8AdNtUCkjzoq/AwMyZvDZn1ds8/ZmJAPOeKCcow27vMzG5lQ0HVxxhwojFukb
bMvf80BRmR+UdMQZ1SI1HygD393xTI6f7Z3DAqxKfmovIj+oIZsOcGn6fREPzYRA
waFONQuwC/w1mXRYYPl4k5Yap0AB1mZMxHYQuEFDcqFmwQD0H0xco1oCnPKAcn5o
kq8dLv5/EdPDJ9jx5ZHjT06RcwdqKQMxB4g4YyhASffMBn2HzSjO3v53QU8l+4rJ
BJA1f8/XMF/sk5YS6aXpQc+DCtwYuA6By481zMF2VPT25vt6r//rjKWArrJ3RM3F
jBHY0PzRtkFTiVTLQdSMxuK1/wHkMRDvtg+zXS0N7R5Y2m5oCnDVi+W5kO9cSn3O
JogrnQ/uyyhYDbBY+uTdRjoH5OuRjm1YoGGf1VAAMuh8a8R5osMp6f+H1H3k9EzT
1giHNPWa6GMpId2YyQyciuShtZjiunTHtgD75Ghm1ABT/vgW0cCcBBir64uab3yu
B2CirA3jSYte8WWFGU8kqeps2MX6XH+2F//d4DMgQ8s4HKJkdwffWWHsVnR4tDZl
Ml8AccHMI8xA1vEajTMy9yBOpdEwRLMJ9frTkG7c7I2UjvHrSpgwyZDfSambi6eC
/RtoTWqJk+W8pfaxU3IGLh0cj4Nlvlf19hp3YaMNASX+rtPx0hWOq+j5xaMZ2Iow
3VYPxhlze9ZNTW5eysGT+MNAkXiX8CucaxvqZ/kXsjDR1ENEO+u7rKW3nzH17s1/
GSs+/1NimkKUzNdCj9BcC64HGeqpX7rNAigC0oCuoAGoBptN7cQh9TLx4ySUAarz
gcqIw14rFVQiM3J0Q32YH1RlBLuRDd6uKBiZmOVZaHID8EgDwGeKYwa3dUakRbFa
W+uyAeEzJxUMGzGfOGhvtEgC07tWBPJz5BHy5ACiNDTe5RFGxWA1tk/E3jBZLIrH
olBa7LcKsiOdR5oFNpRUgQnfVz8P1B5DxIfr9+Q9sC2atat80nJ3RsLlNIjYLR+u
s5BfGcepgzdVWp6JdD0dKgC8Nd2nhsEHH2lATMItNRtOD1kvrrc21hwcAzfaeBZV
FjTOHIqvwo5cRMQCSpAXhkPokfCYArmVtMIxuA0C9WX5AG+6ly87tgDoDRUkjRQ7
8kec8f6o+AyojD7Zya3kbXJVAI60cRrcXGMm0Dsb0aVXaoORZ2ahCa3DVUADRUk6
kXo/vVYaMK7CEVNfXazHNS6EYHPJ+GDIXY0OZhlc2w3LnIybq3Fe99fUppWMjqCP
YUZ2jORWZ5tqmH9k7ssENWiNWTHK5frtz8IcxlHFmzgw3u+F+8oPE/bQlCioiZpl
DRHOqcV0p8MK+S/PJ8QjqqqY+2goErI/LANATqEZ9V3a6kjfwydWhEHAP4xWtrFO
Nxi4/Se5c6Z2DUGjD0JHKO4oEJcjBvJNZP/JuDU0C4SBsmrHxBLT9tx2zIItfJU+
SM9wFGYw83B5EkHrqO9iLl2Q206Qf3Og/tjF7J2tzbtuyw2IcqkV5pQx5JCAC9Ho
GASfHURNNVyRmeRZbRQWZavgluyeE4n+aDVbTJGqgb9OvYBlDhN5bSjWdq05q/fO
t/uz1iGK5rUG9q5fo/iFbbkca8ifAKg216GxJQzrqZGErbp3qEERse6+TsciAdXC
IqbN7GTWYao0AczT2OhTxORHCpAW7AWeo4j7iLPfZQCej24Nx4+rWG9lVNMUXfGU
h5yZS94FijF62AMV7wt12njanCtr+iVb+IGDsB0hkQBT0I3vLHReRxHkW0aJcWA9
WGX1/yFWrIwrTD/Dwhi+lKZ3ZTjZhp/TcrAGrWRcAuM4Jzw2qwS5D0utgalCw2J1
1+Vl+aoqiPeKbhM4aT2M7ZJHvnWytG/hsyhF4jo7DopSA2YzRM2G6otGqJnBSeSG
TtBTSYkRAgAuHmieGuOK6fsLHi3wSoHELmLI0yJwu8KBWtQO3hGu3CcgyT7xrL2z
2kOUvxyQafbJ4i1I6Aiio/3DlLVmZCTtaTFdINEx3VfStLDtJSfL6LfS0MZ8ihbI
40jIItW863yV+zuXBvG4NblKFwGMkvnMoSucRpJxkUcn412dBStwftEBNVBZ9+PX
RCPprE439ARtKhpoCjMG1Nbxk8TUcdGODmkbJn3fekyfvKmbqrWfKHgcE59GWZ+c
1MoeDSoxnLIPOSiGGAxgrZZDvsXigwnbHuJiK+c14lqhX7PwJq5Qx8TqHjTl7yCg
m/dhWxrFb1RD0Z2tZpXvpKs2OHAlazvlEFDe7rfvsSV6/NPpwu9xlgtOzKjgdwdA
uaHbql9Ess+QCAkr4LojI/WllSJb7uqwfry8PVRQKPwgaUAj0IeY7R8lo0t6Vvn6
u5DR2u9BT0lo97+XL8D0vh0w5J1eEt6y4gXGMsr2FCQbS08zyJnC9LQZiZgcmHAL
nLbwPyOJxvhYFGwT9NUR98KKzNNgAnRZHK+CoImfxraDwzZX6toeLPEBjqnzYl5b
d/i3Mr8/AJ4AobvQiVpoFjS5Z4bmEVhhtVUXNVOjWaKOQcXmsBMJSXhWWTJmkIPW
tOMvj66LQ3R1S071nIBc/zzCHlEJwcd/oXqMEqhPmS1oVGJJ0X/rXKcxyhF3rsPS
yyDMMCHU9WX3W/XsJgswQ94rAdzn5k0UrVU535S3HwfIkR7UyW2A94DEQEjKwdVp
228rkfxOlls5bXxpYwiTRGeAjNPdP94V+cIwxeuRWTIxZyky2+nwwd6mJpfMD6KN
k/LAlmIi9eAYo+lQ1T9fRkzfPuoM69+KdfvAkkr+Q6n/785ky0InqQkDay1iyhWH
Cdxwp0O6QOFu93MIxyzpl0DS2OZhsOq0aecf3xpsiNde8ZV/XVDGc8hH99I0nZmo
nKvSjveLD6YC1L6tmBO9l+WrC5XZBIoONyhNBoCC7ZJZFk1DbWL0VsgoNfs6T4d8
N1qcOFiWH4BPs6bIL1I96MvxeFZ1z/VX7qTNBYJ+7BWyMZ01zS/X3JbnXPE5Q3Xj
K7Wjo9qh16pymchEUxAZ5KLmZo1X87J6f4JTWZGLxR0oD0ZUn3u1Lzw9Nd4saxJW
lF9eVOlHzfnTI8P9q8xPMKOWiL8oBtXE4AFWt9w7LKRJCkwR3P5W9nyY0HUHZz6R
vb42X9GCGsNR5AIdq25XfIADv/NIhH9pz8Z+2KHQgeQhbWbyfqa/Rxg/W/EzoPR/
kenG0m4eOoRUrSfbZzAVKMG7+1F/cBPo/u4tJOO2fLnv7mup++EShxktDTicIt62
oDkXxHlCOhg8fssWUxGHptChtXR7l5/O+1uz2lLJu2voorfhCEf4DOwcvD89kBTP
2J7/rVwUIBlUMNbaZ3xginY4iDFK2YmQuOphqM2b+v+Vaj1ikqLlG8TDwA3mXkTF
vbDrfBBd2eAmU6moPt9r1QRwb696mIHdjizdkMOMOZqr0Rwrvf9xUg9fk4qXFYdB
cWPP7iZjXUo+10f4U3Tr+VqABv68cwqjcR/oohOBs7Jw4s3f53JiDdqYVClaVnOV
Clm6ZyexhtF9/ONKvgGAnEC45isnQk07f/xpe2QeWjbSwuPUJQcmpod+6oBcQr8L
EGtCNsIpMkuNEq7IO0VRXZD0VF8dGd2ZTsWBAD3A0JCQsIFgD8K3ksILVxum9/T5
XVwj+pi5R1o2F3wn9lyOKBCahGXWYwdjvF20ffPNlc5HxKY7DS3Cce5/qAx7GhGU
DuQ14r0Sk4LL2FAhhubNpGA+cf6+0uwXIZGI3MP5q5VOgjUyloDEJ/gKWfU2qab8
OBSSUye9GFOTWONE45WYpgC2zY9AJSH0CDOSox0+/s3yqHjFOii9b6tDkmSyEUcW
Qo8mCUleD93B5+TrVdTQupAJLaSOXassWgg0SPunQCnHp0gDglKAUFn9EZKZK6yn
Erui+kdqGML1fC0QBIXLE1y2fZqhUWRV9GtshesyvuDtHba7RDqVyfPWi8zSatz2
6a/dzE8E2qwvdgkBa6Z+O0xJ2od89JkyZo9b4jVlGPOX8MKmW4eLMRSQrJUy6ZEX
uddtULTbefGqSZQlY2X8QebY/6vP9KcTz6xFTzBkATO5+/cAQfFisJKb84PzVox+
fIGKmyzKKCF2F2a0ix5q57Erzfmq8R64vRokh0RZNPAkKRhIze5Sl3cHBXVGW9JF
TsdWBBhHjBISmSJ83DLK7cDB2ZnNQl+yCYWEHHq0Kd6MaVlyqLht+ZQ3C7M0K/kv
sLfedEY3Tg3tIW3E7dk6w3PKDdFFMYhLl1qKiFUSWEM8Br6HIK5/zJXkWVMT8lVT
4at5bfe5GyIUiflyNfyvObhAo2BPQmmzYjU4CjsMGFbcxsN8eosIrvVc9UKwZk8P
5mFQQ1dcPSuJn/uI7wwRsG6N/Wx0INGiDjKWHnugTwzuQebWAMfSue0ERf0iWDpc
aZryoRvpVU4/417GLvIvY/DPyDK2uVvO6K38o68BpLrKTjwod4jjd2kgkYTgbSmj
HZXclfTDVQCvAUlhMVkwQnzXmjeFXJV05AC0rNeC3/T1xN5cuUSAwlFmwzKAxZda
6M09gqSsmNYBSLcLBuvkhmg8DyaX9qf6WdVavI8jNu/VnHh/bToUTSQHGIKcBjdm
JkIWrHQPG3JuMFcQ7mSiUKZbC7CxqOTEAdizOs3N4+8zuAN2YQhQ8ROeohLH7xAb
h80u5FGjc37U4XGAAzsJFU5Df4FSZRNNldDPIMwXoIzGMZqdv4erY38K4/V16cFP
YBH3bxLtkc9XyDjBYs+zQ8D0xAW+19mawYzlORVhfK9PpGLezYXGGd1WsOmWyLZ3
Dh89KWFTx+1JxrddiJQAxDG40BBdnEgaizSs9zemi6nI236xVwF3FHBva7XdDSV4
yPMAvZVJihp/vv6SbdetNMTEHSbaSdn4di1dBFlkl3Psn2HYVWzWn484d8rV11EF
lqLTt+3qNLhN/FPGPoj8KyclOXKiXAtb9LEG6+vtZh1MwGPp8RquFbaTDlxy1yvN
Idb0DDXVOPwosKHcm7QCrLBihHisTsvAxT9GS1ADSdlmqfIyG7nbgSUcv5U/Jr+x
iOjAbsMBf9aW7J0dOMNp08+jQ4rcjZFyhslpdB9Xf3OyMaGiegEHzvvtfAcmUXQ/
oF5y/jE0PPvv9N2k2fEnRfpz75VaMiwOBVw/hzdlPIG7c6rg8mWTdsSqKtECC66j
Ocgt9/AMTBuMQnvo4s0d7PTOvIkXVMNx1B8JRfJlb+YmxlP1BUnRvMnDBqc/lKo9
7dzdQz6HB3dAi14u3NR/CRNDBuaY7VKa95nv3Kp/pJa1PbGzb6Qv6mjJ7HG5DHdp
FkKTfOgz0jujtL2BSSWM1W2DjHR076DqGWvSdqT3ldybow63bmsSwL/PxJWuyOCg
79nJu0mZ8jYoxDRhkG6s9q5fQ/byHuzEpV14lThaIRekVzi+RZwVCegLgfQHrvBe
6aRgQvMgRzkfBEi0LAOLvRDyfk96GkgNQCi2JAaZMnvTSwgt2hK2LLN12MhJi+WQ
+QnNq9wgNO8EZJTQoyGGQKSVxdDOjxVDaIWKqre0rlsEJnFjeg4YR1z2EZuK2eo8
/exF0LOQ5n1QOUGaaWxo7HutXnUaQTBcrlG+OzZ2acjVcnVXyk7bgjBtxhp8mi3J
E6Oa36DdUpuW5zHvOd85eN2wxwcw6WAqEw1J9lq/ms556Fa1GFZnrR76R3F8dAl+
dnh0OJaReq6yAyJWr/2gI9aEyPNmyiTNk0MeUw0kXwSNX445sRCFw+ImDk/+9PeT
ZHiSzO009WPoI9aQ8agE52nG38wquGBmWuo4uSdrocE2sDEzrvJvZ8cgSL+bIcsh
BtJN0zJ7pAzq5u/N8bDvVEr8rOo2zOMOniXMsDaCj2lFJoEsKn9WrimAE97j4PRv
LL2VzCzQ1YC+7WGeN+1mNGZYoi8rfM/GctUyp1WsJWMQKX75S02o0r7/sbSXE3F5
+jKawbeHSCOCr68qbUr7PU8DUry13x+PVTuhqpjXWxvcM/XuI5tSxh0mwVt+tGFl
NTPqBxS63xtRmITh3M5SFgGZ6o9bVHbED4edu0csUWmn3rAsEYQuAlMk0jMHXA53
nDSoUfvLInQaGpA1b3IbcnT2RJb2vdbxklbxBFWWr7TO6ZFYRoVZolcRzUV5LQaI
ButTfOyJ6bQEr/mZ/Ch/DD4J6h/V14yZUDlfSRD5eVyHQlIKp7o7GSQ1YLyxvCRC
EPQPDmLFTpnBiOjJKn5PlnSab3gXerKBRqArWhWpXY0Y1IxrXKj/5DdU5xn77M4I
SUVuAw1tFAgGElohVP7vEZRcuboHrxTHH1TWGxaeBBy72I4c6L7IAz5HUYrQ3yFf
56Tysf0NSu7urLjpzyQoy8iWSc4xADNudXCXsjOcjRDhap2eKX2/6KFSz+OE6Y6B
qbQhXzyAeftRemRXi18iIC+aGkrsgsw+z9mhLOMmEug1ctr8ur5RwYAlRK1laClD
8wPYqn85qd8ZZJhd3ySUONAGjyvKru1LtPAI6DTy7obLpB7slFXQlU5ydCu9E7ss
/Ye6gfcpP9SsRIOjLneEzUk+Oi5xt30YHme6+ovn0OM5INuAUF1Tx4BpJ645Y/dV
u2m4sVJGNEsn3K7IGEEC2J7fb7HLCHTe7krA/eJcarlM5ef/foRFMVzdFBUDHh5e
UJLZmqH9ABUNGm2VFFwuQSSQijFNMKp5D0b6yLSHz+E0OJFWb4EquqkLMLwng/1U
RSMUjdYo6qAxsY7j9zLQI5vfPNeAvFh2SOZm857OfhzecUHvLVcpgDpCnzIUSVXl
1TLlvpxpfI6OSzswm1yTX+awuWxv9W/C4aYSFKWLDnvUxHc/zZOt0NiOkQlG3tcF
wlPFexj5RQR9+0LdFYZYfORcQMe3AavVn8z4vxxO813TdVb/ux+HB0K6IWum1Q5j
L4XKCwSGgJS8FmZdGgtsMkfkEaxBh2O0qI9Egge282MdjgJzCYHMAGVvzQ1NJUi2
ADme5YI9Nf5F72VJbAvjF3Vb7j6EVfhxakRfGsTGOW8XAzL/xO0Kzvw6KgOSvBcn
IjAy8K/zJajUur0dQadsQQ+/H1/UShdIHpZNK0OafSl+rBgFsBCK63bvrCpjL1PC
XMbnu8uzX4s+NrQHXgOfT6TPDdDY5AL0bRGdgB8zqlHTd0ihSR8zVCtVhSzUDNOU
6BbEWbyuPUg+u9AfQM7KRfY8PUnHlamveLgC4MsnUa7jdDfFa9eP6zqbLeSuzDLM
O3AQeVfffdYvLtQ/3+YzQtBA5HGLIe056dk4UEcK+iqncR0l8cs+bf/5ph/ZrTDJ
izKEZ12wfECb7XrzniHInrgXNxLzqy/b3Rbt9RzT5W2l16OZbyryhJ/EMl2ShVdR
ZTqNWRUztpsYQmFuq2RgfT5JYOKRcJBqKBDiPyU+odu9spWpw52KpZTpCL4RPYcT
ya+8LNfsGjHKij+XBfZEbXZING9BEd8hPhg3WKxdnKRoG9imeNT3xQWjYXbXd6rs
M9tqEaes2nTHxfGUXhex8QmhGWdjSV7jBjEbr8u3A6uM0Kyy9OtzjhEOBcA34DH9
f0U4ZOnrCLbFRuciaV4dTppbJvwQEqAuwKjbFGxTzNZuCzjZTS1WSHWIknk1Vu3x
LAH7TkGrVPzfEzN0p4t6E0307fdXR9pbT5ZGmoepT9u003bnw2MHg9WuT07UNadG
REJEjFxIyh3S3Jc/idDROfxDwziLtpUnpOQ9IX0apiSxQW3/CvMJTc1KvvTPaH+3
sGrHdGo5eKWQk+/paYKsInG6nftEYzBjkBnSnQOv/JyIy7JjGSS9YfnTyPuBM0QU
xiLmEXpb7l+I3wwu5jxpv9yYsyzmDfjsh87Tkz9AC/fRpuKRLpdGzARySk5iVbiv
Ibx3bKXlc2bcZReF9D5pq6ugThMYWuylZk498A/kOTk3GqfyNf9uHYdy8IrkPFHp
TKIqAL6JfyKC4QkLbk8fYRr/wvar79ldFcFoT2EY7aik6/joSh2U49HItpP0s4U3
+Xt7TXUYRwoiiXEflGW/ArraOKC4XscmjqOzeEKqhsCEhzX1F7MfFrLEVUEtADpm
W+k9U2uXdEWoiv0TZvcQwmYU8XvWUnnpH4nL+ttAysCgVNbdnbB/qGSaZq63IJTm
sJifn6f+hjTmiN/j9FIzH0i5Z4UvLXgNzlaWTrlzFXYWjO2+Bw/Hb258BW/lROcE
zI/UxKii6qBt3KL4OtZf/zX5JhBlLBs96SrYSudtTY7X02VdLZXNzsPWtTi/3rBl
4HdjljSLh8BwzCohEsGhHF/Mz0MT7hQWhieqfX4pWpDr8BUrHPz5qa1hRGGxF9pD
mXrwEyGt/97dFUAEbRWOf2zW4BCiFmW6w41EFURdP3fU8t9hQ3AXjldG6hZ3rGLN
Eds6dMXIhSvDL5vDADV+4HG82HEZG6UYmFAFHLVA+Ug0lmhy1nwLkBw3CHue+bRt
XH8EQlr6FB1RVMgyPGQCA+5Eq4yf4/9vKm12Cce/FsinKwW1UaxeOJDEGOYpA3M5
IlGigsbqO250AV0wTFIpovZLmAcBZYPWEWfv+qhiTFhJbE/u3W2lg9nsV8SQ0tzX
Q1ZTAJEkVnt+2lNk8McPiQ5OQRAY6I++lUX44nmqdGXOlVenG2A4OOW4Qe00jtvb
+cWA9U0rAPN7niES1V8oLSrvm4pbGNG2BGti8XpsbWfqYelbmBXIdZdjTM5q98xO
/o4dY76lwMaY12Vh2unuZDC4O5fQAYaCQiFMimSvpE4q7KBdHea2kafun10Pz96i
aweZtafAvmoPJTJFCammm2QZahVQbfOsumcPVj4ZykM7+ObrVLD8BG4KIc4Copo6
KZuUvZ6UWDgx2g7TxtnOBw2/gUTCn+lInGclyTU9qiRYYLz8ayFzp3r5nVwbA/VC
bg/AlUioWoJyrKlKMJf//SQMeIJwxznisFqXPMeIzbiT2IRn8SFgIpWQKVfCwEtN
TNn6/XQsW6BitN/MPOSt9UHhX+1DmojEPyZj/YwyPr7Qc643w8wBUXEPXrMhIxtT
UCSXOYRU/2m1E+6xnOI6tV4Wo0xrIMN/MVyTpdcu37pEDrihZzBD/rqR06RapNqD
nhz1vcvvgqRKeR4PxSs6RrY0Ost7DgoZjLphTINDOJRYqjNBQudAnknUfzKxsX4Q
ZB40MoClE45wG4z/gCuPHysXPTzSJXw/xge7ySl3mTgL8p6aB9I7mzSqLqudLG00
CgR1YKQaoMX1sXYCHVjQgCaij0P7cufaFxQfWcBEMKIhMxtmNjYeS2QfNAbgXvdi
Wse4yK3BNh7gYpJ+QJ4M4Iu0eM85G5CF/Iomb1O+qaap/gwYwlWOEqL8+BCGdBAZ
eU8+MQdMvMocqLqOf8tmZ1pHnaXV0sE+BRiMuF2jAEX7+pyxB3dpMeckkeGASlGp
7665WAA8KZKKjfYizejWDx/cRykJ9/+u8RFRrN2R+otoFT4ctOOrZrnWxwuVQwh5
tdhuujJLvDbXO22wjN6CzrU3gNmdiltcbMfUwmZyVE3io5NYA3CgAnQfbw/XkS5b
RyHumKZ1na3JR7XUcFKP55pctcSdAQqd3JeKLWqpFabJkkKc5TXBKJa5WbPn/vNi
yASjMHB7jYJ7r6/bUu2i7JPoAW1DHX2Ke12NHZZPpLwJvfH57CVOIDRh884+qmPV
w9wg+w8ECNA53N6ktMUrSqwe7/4f73hySYwxeBEusuCp4ju19U2cvFeINHSK4Tn8
YNY4JDKnNdc0D/hIsXTErBveabDLWB6EITCoKRMP444TP/zGMnky90Ysi2BbRtWP
C6D8uFCl76KyY9T9+sS8OAa0IsW2hdLni3jq6tHmP5qkJDj/yXzeAcmTYE4MGh7y
6phNDek4XrOEp9IB3ZC4+1mmRhfAGE+87YgOsIdS+XSEXZccp9aYTuz2CP0hLJVM
TPz1zGLLFUlYVSzeDS0wUqr99IIUea7YgechCGYwZogWyq6SZZFYRZnxoJsHjkLB
UswFpcy5inr44oq8TsdyfAdkK9FrIUUsp4R9zVeUjM2laxCS5vggsyLwOd2aomNF
dM5AiyKcLNa2NWIhugbJ90meWkPSI2Gg7olT1x+b6U5nebWj5kUFbaC7C8e7KgQq
FvuqqVrwV4ovXqWf6XcuKcyPZBH0rsBjohN44AE0okFYMccrWoP70iM7xpa+ZSZH
syTvClox7LkssmxYHgwnLjw7TYaJgLESycLZl/NX3cMnWcqPrkRMN1STmUi5+YF8
VEc3jNs2Y+wcGmUdrdUu0rEnPHiwxT092Y6mhZshbDDzPmR8g+ibu6sBXNvqZOxs
Z4IXnXCdiMVoPwfXkP6vRyzq1wh4+erRrUKCGa061iIgnqCiiBgnA/VFdtlE7+26
5CPLlxBamqOGS3VK5PAPLHkq3eMHRHnJs6tdTvLNjfiZKY+hJ33QLp4+Dgi30kWR
SBuoG977GrUfq9SO3fwcpViGM+JkUOtAc7BscIeGsr23sAt0rzf9hVdTVrC/sIYs
Ww5ZJhPT5Wi5xsUFtj6Quic931/D4uC2yXL7Hh9397YVLyEaJAQXfHwfRXW2/cQF
bcx2UyAPmYnUYnAaJTAIxqQodHvxNqbtvb/CLyZM94yjmozL/takj0a2fcURNrd0
lGmkILFnLUHlf4lOPuJqRPcjlrwoX5QjRojAnUXS/VD4eCn7e91NDqmsbE0hGuo/
T04NhA9BL6S4OBZCo/1XtSH7msC39cYauEDj31gtjaUD7vFlq0wBr1zmIZsqoDWc
sFgEgXa5LC/9T0wz9JC/+3EQbQS1pmkIGtwM9xcjLuCxa3VYuCXIQWNhFanS7N95
O5KE3yTEBDWLQgEf0J+Rbl6pidaQcpBzeOr2EP+35Ywfx0MzkSpudQQz7D3PbJia
BblrP6B0R6Nwlc0kTOqtfgVNUW/xjOB4Ztnr89MGz/nLvp34VccvhwvLmpfRa9Zv
J1EWMaDJ9jgNhsk7G3m8sk3niTC/07chETULwsmaMc/xLAXdZJ1SZTUU4ksLOhl9
w1P1GDthlUNpACuZEfA7um2HhSysZ/jqORhwggydyQlLagtFD8vvaUhTz2Q+w1z0
5L5DWvII3ltfTwNh/45LRLv2rsgAjI7WYi7yPQH/vJXJEj5a8tHAak5/L6BnAjnS
uPjShsSYOayeU6l3lnfD27GrT4DFLrK+6CO8wH714BGzFcDGSgPMJnO2vr1HBw3d
FtB9ooPyllvV0Mh/k2B7QoLxXaFqMwWQAfHLx86881LpRVxBi94zCjSY2+0KldPT
lTazd52xXxgXLec/0DYAxf05+UeN87JExDzzBBi92T5c/mrPgWgg/JrHE1zSZDTs
x8war45KtxcRVXduDVT0I4PkSmQ7e7qb9VpPbDzhJd3DGyvyr9rPpKpX/xVouksg
LqxQTRItHUivzrNVRQbUcU8OfS2lNiwsZk9YhONaaJMduX8622Zq3CO+CjdXJ2ep
g9xXvxRYcb+sDb7CrO94IpM1P8AM06xHBB6mF/CGMeDoH0Flpxh5CiK17X1dmuYF
P4nFJfn88v4leAq9zgOvTGl0F1oIlWKi2zaEjsiE3jRk68k+5Glp4cLSiXEZsKgi
OCrrxT2irnz3jxoM5sK973hPMpxhB7nQG4m/FJXvtQuCSltUOcOD6HuAKGQVq+4c
LAxckk6E/OTOuYId4lG2ObGJLikdfsVaOY/rAcnlfLD8WD5dNNbaLzNnBhVALTKg
tzM4KjUG6qTIGXFuMXNsVifTHPCyCmmEaK1naC+WL1RxPL92E6Ylf4EnqLkcEyOZ
/6pkAcN40FxIoHJVYip6uqjQJx7VSIFGpMFfMZHrkKm8OP0hwQj6usIyvrDDxj/C
pmKm0HDfALqPEiFhNlWybL3ULbYyZaXjzE9DI3JKUSQdfuFZTaukbJGfAX1Cj7N6
u/f15diK4xzdDBIKwxPU7xGWww18wVq4NXIYNq949YoPjH57nKn8tkMfoWed/2l6
EmA3JIYav2YeZg7eEbgGYz/pxNm+4/6Mt+Yw31wjKKgpsuwkKwF9d5QqEqkrPEsu
vRZYILfaz0gbrn7zQDxpHRdHsFckPKDKGHVcrmiRGDDZ4uhmmryviVAJVJQ6sTwd
ZxvHw+tQHWAGdIUdeZZ7JnA59jBLPfkTFXJFCYh16q6hjQM8AT8NCMpl6aGo5ct1
ZOu65MgyoizXX4Aqsht2E0z31IjjPDBh7NSa2eMuAaIxTYAW3rXdD0GqIEk8eRQ4
nB4tXq+8joUB4a1ZEDrDbGcPq7ug7e8EEFBW/SK9xFdibA+AmeVyACP3lbCVtcBn
SfbmdGEmh+iDUD59URvGyPsOYv4kxI0QLaQWtrLUWdlZuvO8cjrSveHgC7n4FBmz
FqpwH0lv73+Zk2O/eP08zaXxcytJ7qMYGB11HtlhvxHiEsL0Oa7aqVPEP1G/6iyR
4yqp+P1Bm2eSTaiw5VaAWMCyi0icqw0Gs7I1e6RlhecW/AADoLFqeZIl1jiGNGki
YO5dFqMnmOmTiVZAQKl6Quq+7ctPUNwRE15+neTJ3T+UZlcriLuzi/jXg2+g8b8z
lmyvWqTU1ZxS9xafU4SI+Tybaennf0YH+zda4eqvTk01JSgrNYPOtp9ssIc6gWpB
liGPz3nDF9oTodnrfq2upOaVkFFADXS9+zr5m1/MmG+sViT6kOHsdbotRk7BZbbY
Rpj4qS+gw3Ucy6mfGabuyapvSNwAQ0FgLEy8bnv4tIbj5vvjFkpqnRMVOTVjxmtw
or9N+B1JwTn2VWBL7gGeGS0C095cf5aLRyzpfPJIu5YRcfoteXX7wdLXkIynnOqU
iEz5X0362xywQX3SCdWzRoYSoVwQUqVDeK3PJfjzxGdbCaon7ZKQZ15iBNcITp19
/Yv4IVjvxuZE/ie1L6ks+6m6UbpTHaSlY8Wqo/lRtW0ZEu0GNgfTQ+w5eIcbZ1jY
Wdm9PkNNHhZPM7pMd9qdO/MymYHa/ggMGxg996BRGHqI0y8y1+jyrJMD5V7EpO8n
O0YFGuFq8S3Rk7h/qgImWkP2DQ2ar+3hwNL7xyRB2uvfkmPh+7ZJML7Q6V1VBbH/
xBLEBQtAPZLaDtIEB98v7EkG8sHur1NU8uiasSSsJOr2mkW0/lLt2SSokr1HxVP1
QmIxXr25vMaWFxGvaon6s70VV/UulohHIeHOAWJzodWHihRf+oGBaFDaPIVCy1uQ
5wSoOUNa1xakB07+UPsxiSDR/AU11KwniY1x/0x+URx3Fk4heDwd7jFbeEfE36dX
Z7BQHytYErFzlvAlekVc/Xjvdrf+PYTBhBGTpKCMp9rTE38PhWzUwB7lXDxqOq0n
EniHpVkD7op3WFyVnKxfPFIBI/YQ+SZQnngvIewM2BR9APS6ZV83rvE2Bd4mJ/oD
yQEmxqaxR6LXNuo7U5zGfEuA0vKYT0/RHQEQuMNZTMbBfCj+inMo0C9AtHXLtUEt
fA8DpFMYUKw7gAVrtWkLgQzqZ9JiUMLAci6X00m9Edl6fa5jFHBViGi717VkYUI1
IenU95zn9NsSq91EA9xWmy9ZbBpfC/WspqxQGxv7rZBK7gxoSdTQlxbkfffQWLad
rwSfHJScD5aecY6mJjn7dgcYiPQjHIclH2lRiGmSUUMfZ8HpXNJuoff7kzlH3VoA
r9vRUtjwiHOkSMmFU6RjsL2kiparCbNf+evf+gXf8By3uygEUHuFKOAjEznF/T7C
6uVlzABS7JGxPIBi8VI1UcCNpFm037+yalrbBfOOiEX3fqRIJ7axGt3cxwvc0WxD
I+20rzRU1xWfUmjF2N8ITih6cFrNSSoF4SeOoji5GidYjkuOWJ5a82MECTDCPboq
t/94xhHMcha6M3kLMM4nCkPQXhkgHj3DwuZjrgxWCddk03avRhJpkWdGw2uFU8u7
uge9YG1+JpONobG+FhSxnoz3qMTAOyhxk7t0l2YWa3e7zcq9lr9A8+/lUJyeSmZm
ZvAeBfnAj8fjAupdhRXzcafaACblOBuCpxgJnhzxfAkIkFSe8aI9Z19rU6WgHqV4
VYRFX0T/vpKz8cTQn6/r+HTx4wllEQQy2hUhQOf/aBdLiOeRA77yNckzcbfcu94w
SYZCzWgBYgpjdUmZ9rscM9iWwa1YJiIOqJRzxZufBpLOkes3Pb4jBV5t+LXaAAhl
m6U+vOfiZy31WJMYPI/79BnPG8zc+M2KCAnSJnkrgDfVrsdphWgdJgr6+DQjEFrJ
4WzR4CS/KINp+zFL0kO0aSN2ngGbxYfINabvSnpvHZCtcXqXyYMRJYwOo7i62yaX
Sa3GwkZmJjadMHA2GkAcW5VLrbS+W9kIV/sDHO/iP/By6v8y/FW4QUxF/GQads1h
mSkMu46Qw3OhCA6NQnQEcbV+wJUlw2N09jJBow43PieyJBAnYLlTRvXm2jrf/8Op
J+L9UL/jmvcPH7hVog8tdiDRqdiVxlYrHUPGsg5JZYgTk/mwNyTmekcnXn53w4ld
Q2tpjp5ZjAi46BAiuOU/AUoGn5lIGbhX3GYlYnaG+6l+GuiNacAonegIjou+kSSa
RVLx9EiE4KO5W6scAn/kHOz7uREWrcFIuGIM7BXi4OaqPZT5z9keOsWqHNlhuZwf
TIA8tNr+s6Z0Cnl4KpTWvQio+czldqiVwQ74FhNQFiyb7kEdIdmlkU6Mse/+hYcR
oeN+4oO3GVYwyIhkM1gQhhwo89EDu6ASA9I67C6d74VRj5d0ET+6OLqOZjHTYPoU
BBrH8llL1iTYYBvJeV4t9k0UwB2vDF31lrROt01GzWlWdnwQ4+XO8OH0p+O5BCyp
RvFoR41L+bRevwllgDitCPzS54f/pbafYTphH78lxZAh2qfAA+lg2+SlBXegLEJk
4GVKW77wpp0vhS0SItbUqU5VThsoB4QYwloE2uwGUjFhCiOX6TzT5lg0X3hvU5ZE
xZr/ssUCfMXC55aOyd3VtBLhbncXfLHQi9D3M/0qy605Swz4Ga0JOEkgDt5NXjHR
VCEbhrQ6ify+adULmxRcRGJSg6yWV00vdWmtryAebjzaocM7OQoZ7WXIK+CiP3gt
eoO/CVqUkMF+GLLjj0Dgt7z0Hft6L1dyrLatrpSsKIkM6ScPfvEep9MpPlZE9DOR
E3QJ8PsAqNd9bK1FfW5chE+BVhMK6g9f7Ramzay+E6HRCXVFNZTfvgm0JCvZn47x
VohP2aDbOZKmwqTbEJUfpOzv9ca0EiKz/dcAKTfDHWWtONP217PeE/tyw6dMswFI
15AfiqNXNmrmWXuN4892LonsK5wGo5UyBWRUOPaRsmExylSNa46IsE6D6+37cQ8U
ug2QIXkI88YkxiSdFrOhQ5KAVq4dABW3iQ6P58NzOIgQWZGunEH/NOTGdCTgIp8w
LxqHsIuoEFnuPKno7+MZyeXA0+xZJe50sewAXFbSqRmAGEpB8GuVcNZ3zRq80XpQ
L/50CnEgit30zqtAQYElji5aLSoQLWS5Hfc+bGxsWPEWSzICt6F10zUCJsuNTCO8
dbsR7ano4nicfXu9OFVylDlWn19+WRCBGr4ayBIcwy55TMbhgsM23oNJkKsZiX+E
9kAzyfLKQKKNnWzF4r/V4znGc9ce7N6+Keu4bj8X7czUIfWIItVLo38N32+OIUAR
6ABEuHnR1z9JkoB1j+d5SQBdXZmh1v9ZvAdi6DokMIRTiiPUX38tgquiCR8UxMnc
pdG/lo86nA9Wxahy/EDJ+KiM446GO7Y/la2GQW58Mcy4uJmmKHwIyVh9n9Fel9oe
SimtaYLZLn1uy0UDVDTnHG5CgeEunWbP85c41WKlKepaThnST8RL295EV64XGt2Q
3A/nyfW3zr6GEED/P1IlJ0GVYrMYABO0o62n3CtKYvM24CNOq3O1Cla/bzQcW6UK
Jt5c1xiZXU/uARgMm2GZPPEreIyhpdGIa/ZqF9hPVT2thxEMzmItFm/DlI0D/Lqp
r7hCrztb1VmyXyjP8f65a0xG031jZXTRLpb1XI4q53tnG3lbzi0eLkD2dL1YI5jw
2h7MLtL4053YVsMjcn2f1RS71ukrfDMUJIwPP1qK46Z8PxDFFtMk1SYEQu8UU19f
pwj4Q92w8ovmjhzW3fqJ7pZMZh2b2UexcaxPDvbtSwvX2Msv7cylD5ACH7K8mpdF
GQ5q3L6dxvb/6fTwQ18BkINy6MAV1ZklrjC+shuR7g8u59ng2tMEtCmS8ZtEREQg
TRHs8TZkyMhGOqnl+98c16Pst0sjpLjPQwGisYjtNTT/ihX7rXZQm58VYKu81OlL
+Jrrgr0V+HSXCxwzmr2brtAjkDsS+353zaBQJz4FzaAuKAsl2wFTihVv1B3OZpzT
ljp383rnAQXktp/gT2Z7aHdwtDQ622abUKYRimtoHbk4w3080wOE6h6SsotoqLzE
RETihR5gcsHGhkybcU5kBPqhEZoHluhH5JkcpApSpP2DsJdzgD2AdYJBnB8YGsvG
fC4UkT44Hd7YJ67wsIzMbAvu/65EUrYudvx6rMWjwcK6Fibl4TAtDIUK31VnLiGx
3Rmj0LXBLDaZXD9fTQzrGMgY17DxAyksYJHIXLe3SUE8wwsv9W55ORr41Pdh2wN6
L6fEIkFvKHfT+lPFaXVFPGqsviDEiPmIUglIr6TA/1V5MPrOBoIyS9MoALFEoL0k
ozs+ioza+lUC9sSazu+fuFjpD5kbV+61mPkpu9XJpBU1r8dsg5/z38PUIt3NKWwt
ivoW9V3dwtm4WUXva8PEQqvznkuExbJqd0+s81tfrk5ZHjgvLFubzA1/+zCAJmCu
h+IqYq9H+gTOIKXv2QEmFS1UaYKuVKDtVGXeoZYiGvpOxG/Hi3KZxvhGl3rH96lY
tUv+TWJUZggt6ybohwoq1Nc6oM5R94H4znTCFAm1u/tBLt4zkl7nnXzEpFJ63mxF
UAYhWdMe7nHaECFL8FB7v/5VzD5q/JERACNoPZxe09KIbj5fKQBs0G43OfHAgBnR
h98ptdQS2y1e/HKbvYOMnztGg5xzss9yu1HqE9DSe2N0YO0XMhVFMy86oC+4nMpC
QRsii5rJLuFrBKkrr8IjsblnhGPqhVyhkef3oAgjBX0KjaCb9L05ZQJT8y4owX2P
IeisJSI0Oh/4VCITC5LiOQYh9BlrmyNdvEnoyzAnt9RV46iNyWB0gNDQH4y9qmld
chMZ6O5kBWPQy2VfIaobAABEnuL/XJFukhf7yrTximqmRHkK3RSoL8tk/jJra8w8
62OXuQ0ig7m7vX6iuKbBnHadRboRFZgnPnpbxEhw2pCvKpNDmV/WMwiGuloxZatR
8Ig81zO7a6nXAeVlUkGOffiqSfEJ6OgbW/VJh1NiVyQJplg9g53nrCKEAql5MDuA
+iFRxBbfUGwIAqdB4Bs/KupwigvDCM5sstbeDR5WzJCje27u5x7p90HLeUrpWfai
tVOaqpsUZN9+NB+DsLCSk8/amDbPBIc4vsYQbvZR/LtQN1NrhAyEHtu2slm/Tb2G
lLiifv9+K5gozpe52wNQEm3vl7KeFFRWLIPuekHtM8TTQVrP6AkxawOC8ucusar5
HIVrcUiPPvnKhWm+FHNHl5xX8bx+V/SU/DX6E2vsvRvC+CZIvowqCAPRl8K+VTAd
cz/2JS90a/DQHFVDYaJOj7BtjRfL41g1HCX5tCzAjaMK+YBdQ+2btmQ4GwdRAdr7
nJ8iMwyf7jAaXv8XQTiHjnie/EsfJEhq7Y5SDBkAwQQ1lkoRdjUqxKKvkwIJ36qH
G4y1zkoExu/SNJVz0sAY7AWaLozqAA5ZQlXz87LnwwPutJR9/x9F1kDuJpzOgLdt
22zpsPwy2CH79NNV0ISdy1YrALlpJyH2SIhGtEgTUJrpptv+DxwLoWoL5+5ABGcG
gmAESKR99gqsFF0bWhmiH5vUsS7afK5rWwkSFLhp0RRqqstHGu0ZF1YmbF+UwRyx
lpV209uY16t13+W2+dgrXbZKlx2ibAvBB0i5QxBPtZF4sZu1Hm5Bpm+9U/5Kqp5h
Wk/1GM25GGbdauhQjzUFrZ64NnHKJ4qhBtcKs4bvvkA6ZaUdg/TjpmA1CDD1P2Oj
05ntBUdjM5EeFYmH6O9FPUAtpjLzqxqr58K4vMFWu5vvHaFzsTc+rgspfe1ChgXo
lUpwwLrIkZ2Qc1O61+Y/Rxa3AhsjkeQoNc/piqXmlP0eUMvDzorsyjKMHgen7F8f
+KBuxQr3Bt/A/NA0AlPCppusvIc30z8OjrJlWd+zoqUH3e6BX/HQRqN88JSHaV97
+Bt3Wj48VZUJ0FTatjJOK3X2IFgdV1uKStFpPpZQtSaNa54SyhfLbaNyEOeciW9J
oWtsjvzhVczJN9nZ9AOpcKb+7O7BTH3TlYha6o3i8A1tIv7TkjqW8JdQusukcBFR
ugKH4TbYZpGZaY6g2MYw4X58V/04Gra9T6bt4ZvEqmKSmOqDf00YQQdNfVn9moQd
fJARJlzL49Voap6R1A1p3RZ+9pUhQZnsFhm/5TJ2ZmVCnTnGL5gb0w5rLXwtFss8
niQijJVdgVRxqIwDr91/A/gbmRyIf9OmsX3An8lrjFVCt5L6IcyD3Kg6NGja1267
BSLKq/fhd00ablXaW3nDjZVc2kCiNVSo6Vc9Dhj+eN2VFCZAmDO18gN8kdQYPlD1
xr9GaBFwODXu/nyP6FVyVEdt56TUbZDQGYQt5oSQPkz3OBmksRrEVpKAe/J6YC2Y
1neVKN9zUhDPd9xLVX6RmU9K0CKh9u7PKBzMB+O89/i0vjGggxKhj2dVpZzCXmDU
zv0pL3K9yhPtxKeWRm8MCLxXfG3/OmiCnA/3HhlK2ZjpIvyxOfb2jq20G2SeM1Fh
0fAml210xZFN07wTg+5KTLfia5tOB+RsXzkmbAeB8iQrTV/92iOxfifSwCzN3ryh
SF8jxLqdoPjRC3Zvv0F17D9guKD1zsU1gsIGqFeTJc79uF6icvk/znn/HadSrL4G
1eebP0k3Ad0PLIVGdMx9y5xzhMh6plfCgdMpxN7628kDlbWZi+avY0eB1OKR6DH6
xwo4Xj52SYogOeEPiyR1QWvGNpJyuTWGnbELKJJhEqqIS4PtnD59I2+eTxDZbJnd
5y/ywRuLkrYIaG+XIpM8rFSrmRsG/hAVdGrEnH5pFTCtoFqOX/QRuYZ8428QiJo8
3klRct+w+ONH4VxnCEgARAByS3Hyasz2R2gbcUMEbLs5zT1ECfAMH6jNBq/2FFWl
NHN9tUQKT/8g3cJMbOKy1dEYrSvnP3z6NOFyXovmJeDaWQ/ZMaL9F64jyCoSSPvt
rqIVbAdR4xgdJQEGz06HOzEqFuAFAl6a6OsCs2JIHsTrvI4wJlp5uZC89x1OwLU+
sgdsRFDFtisiai60MB0zZtoYTxY8nkAvEazl5YaKNHdcKTymXRUwtwUw3iGTbiiz
/F/srfM58/7ZJvyxqk1CKzjDOe+3GJMKb2pKwJDgcs4Yy67ZwjiwB3pTajYLAZ0r
+sw9TSq2/qrFak+1fLdbnsV9BCcFqUPI9GDoKZdV5sJHzYsSHJZRUpz1c4x87KOY
pBAmK+rmX8K5XumM+7Bl8/YHtXc3N+yJ+FmYeaWLGqytLneOj5bosMnO5e4ZcGE4
18XdburNtrc7m0Yt3p9d/pB4lAhXyeCPooaBH2CTYg/qM2n2fAngdjHJyJt4gKky
if2WsL6RrmrK99IpibjvJRMmBoCyZbH6GFKk0OHfYTr43VSg0teWdRl3OTpfxdjM
zGfm7xKQcln/rzYj40L8lidQmwjlyjZ5NrDTZqDMv16/9T9OWllKmVVmcyu5+iiC
wbZmo9t7p0JwXhMpmcwL/qNSCN0f5aYM+psdchHsO/rBz57x8rcTeJmkbJ0eNQO+
xCCXoBbvSIb5j9IMKXu5DLrR06qZbiXFQ58y9PLycSKh54vu2KGT/g4lnvepoR6O
2e4k6Rgxmc66mOMRj+U1BzqKjpd2CFmtSylcbXn07lM905PzNhevZ3EgpVAU4Hsp
0yitutq+Z2fOg6DVuIZjHL8PDV8tGOnZRBVPToRJYRJS7Tbjfgpc3RMLlO7jH9e3
EjMtcqKgPdk554zL8+I6fguAQqG9zAa60m0DW4HUln+D3Y/SCixE5fV6MgcLuShs
ZITzg8zCZ3q+GNHZJFzym4kDbk5k2lDP35rC/odobaLyWcKwdW6QtB/+4Ze8PF6q
ps1PC4xn88HXwOtsRXy4D2aqg7jyMIlmpb6hSwUhJOz8mRD//hSi2LcXH3Cmk+Id
0WF/g18WpmEpuPhPimOpn9v6QzrPnR7/lQqLE7UlSUZHaLCkiofGxShhShR2o5YC
WWHIyo4Qa65Mtu/Iu8b30rrgmM8NtXYnxSVfY3cVlK2oJwQGFwqvXMKraULNKDgp
ihqsWAxhHyeB9xs9QAkJTB9N6EifH0oSjKcevFnJazPramoJUOjKcOrRwRrhR61E
ZWKYEFaq6mP7YtZ+ZI+7K8aPf8lnFAPTWxpAgZzOFiW+sc4NGM8txSRxBWuoYXRY
EGyM6qQVmrCykmmd10RZpGOBGd2PP0XGhxHAJFbXuX9C/AygwQ+pRdCkscDT98By
ZX1u1LSBTy6RRUO/1pdGa61K2wssfPgY5llT8WxCQUHzge3XHAZoJiJy7+qhq3YT
iq8AEgm+i/FsrwvNoBWI5UFsExMJ3gXn82vUnFJroQNWj2S8aY4PrM8t19lAiCxF
a2/2rIdAhpF9/KJu1KmD+duNtvGnjVefAIKs6FxF0WZbeJPagNIVAcdALw5ognWK
H+ESBszQRsQfWVZK9a2o53+iiyzI/M9n5RiofbXB5LXV5EeVGj3W4qzbR0idvMkv
AlnsrqzOaKCI/Iq4vQX7hLxQ358PLVIHfz5bqlCpRPlaMqmWcvfBgBGjXvKmYXA5
VwwwS/q09MZTJkUmytvxtYoAxBBA1xiEkAYCOx5XpobscVaJ1tX1iAoWS+a4vXzC
R6Qv6+B/DxlBUfmNGrb04VJaLGloc3K+IXVf4cO6ZnJKej+ChMS2SPUe8DxCgWpF
0ARel6Jkr7Bq3pO0D4p8kYrrHvU5lppejAUSTxyb2jCSsVMHQDqXZ7MP5Q4h4PBr
cBa+C73wDj5NY3f5XhWPx2h7AVFoEzVy8cPaT3s9CkvMZ6gFdaY+FwdI0Nh8eBTP
yVoV5aYbNwNfCloKuSaAnSSu3OzmkYxuCrrl0yXViZwPbDh3Yww8j1cKl4cbJ24b
6SNgXcdpuMZ03CcgtNQSEUgyR78Btg1IW+A48cTNWt+bCta3xPjBJEXNxIBbXGRk
aaQ2gVqGX4461gDsm+UArBUpmh6KcZ3FyqiGU3jQ0OXcmrCnw9ACtwatNBAN9FtD
3MPBxRm7AEFBU6/McG/12V+A4QAigKBgVs5P/x3vl4qmRSnHyXQ6DhCU4UzlZ3Qu
XdbiiPvNvYoVaihXEvi39ZaUvP34C3mzKyPp5dWDZz2+tyM8MzzZ81/S9xx3wcWr
gF9z6BMOg6ayBGH3d5T/CAqd0g8n0LoVWKwoUwvZTOvNFzquuGx38OIR/yh7imAV
+yE1KosAOfCEVrFH9KpOQnOw0OtMG2IDDWnM/yhzY2uGuFF+r1GFu0LW0FVphDz7
OR0MtaCDfUUBG/PpV42IebAXpISMj9Qqzx7AWSwh0j7G5vqA7cJw1wbf98cJizxT
jvYpgnt/WadS5XI2v695wYEASsk88RN+YtBPensQaPXqEKLQDNSBMtLwQ4v+Uxkr
RowQrLyks0MpimkJV4++Q/s3mPZPBBdOQTNNBI9vUp2UnkvlmqTeQIW5P26RWAWV
vOnXvBYWXJ6DtkTs/PuB3+wZmJ+4OyXk+C/Ruz8El4zbmC3w9m2aC1hdJ/Aw/7SP
ZezxrUviTed2TP7SiMmyckFE/EcHeA+6feaG9VJjXi17EUXxF0pGNsaatG34wlPG
9Z6MyAxrSkTADfjkf7R1aDSML2UIzu242VHobaYwT4px/00qahlzvhsgMTU6VGI+
pcS5CUbmty0e1tPvDAKew0nxSEHFDYWaon3i8oSeYoSeBDx7FTZfodpDdXQ5yt4U
+JfjrMnIRt61ZhzA2XYuy9IlpnrUEaMbAXqrQoP954ylkR72VX5RqfkrNwtDe+Gq
ROJ1/0WFggVXguvEMGNtsdfNIt+WRoz5ct/HqfQf8015MMlxezV+oRgQcZeDQiXM
LlOzZRaa3wIWEB2JI2A9JUpXQ3yIBnhiwLZJGhVcjVXMTxLjKRGHG+jQN83W9UxS
aC6iuPYrdcn4foQ+m/3jsFVxWq9MnTL6nNgPQkCw+Hv6vlMtNVRc8ZRWaKVbZhWC
obZSkFsOLvwUd+RUKvkD+mce/VMDjG5YArMuVf5RWnbEjUJlBcp1/zRq/17z2Nr6
Ez0Ox9xzh9I4gs3+38fa6b2n1PcBIsJb0LMK7AoU1u+6hU67AWAct0kf1NdJ+XEe
5S9C9nJPIkcxGI86TUDKr9oEmHWn8+Rw3lcV9gPjXukFnpIyyF8Irrvaxoofw2Rl
/jSnkyltXDSPTJzsALWRGGfQVlTQldEqskV6qtr/nqry6cgaTmq/kvRH/TLzYCGP
WK3xYB6h1TCRwF3nQ67E/419ip+R9CkLIooURYc3cfcrQoPxG6opH8aDKWs2Zx4l
aI5P/XQBBgXeOmepU9jsC6uNFFSc8W7xFeNshg3aGnLRpCcRUWmP0rw6tiAue69e
YUycrO86nbFwqjDRrTnzNWbE8HaKDDfcPAJuXtcVULcZ8os5rNUXF5RhFBNbqDCg
bKJP3GuYUWkq/2bYMVSvNvZZ1Wn25yhtp/nCnDd9AkK69RJH0UKVTrVnwyHTvLQq
DiW4gOYznSN7kGl0QRBAqe0HgzmU+IVCJp/RC1iKIDQzHUUq6nwaflhcdr0kMZJh
0IvmXllqMjS6rhoQFOXcR4I7ZsYoNHsRp8yD/+iJ03vbo/652WDx+SYzybz+KUZ9
r6ooWpPTVVOmDoETuXzFAEb6i5bOFgJ3xiWCBjLcfV0u3CIE/NEV+TKGoWitXuIb
YJPt2PekVt/ws0em6ueqxJ87O6aa2CbHNx5quqLNzq5FcvM1UHOUwsWZZvxuuTZ8
80NLb4r31t1q1YUxRQPGTR3eV6qdvpGTMKS6+s7IdjQy12zzWh+a/v10P6AvCDGF
0PvZFgIZ6YpBgcln3jlTMgWbmUNxmNMdzPaOKahUCtGDs3iJV2prth6jQQGzFZPZ
NYRKekTu7mfY0LfiUpXYak8ZLvudTbRYYBVGYQPZR6G3q8J18FF697ifrl3vA8M3
EKjZMnZrpw+HAcHbp9k1F0AoLFjx7Ce7wAUF8tDAoTjb/gFnHbbdqscpiTmXuf9c
I8BYSP9knaxoexSmxYF4WGl0FTiYRUnOudScqZnxmPHMbxj/dEzrI7djo/9BCvOj
A1Ku4sQ6mtMQBolBWnx79FtVEmbzaY/EjnVEJlXaOt7Mh4FaFSlRzJxN13McI7nf
5rx8SRR5czQ2P62raP+p5EcYNMha0n9vhKu0vn0nhJOS3bKDgD6azLnFYOWaTXsJ
aQCMmjKDCfbnUuGyNee6w0TYfCT8SYF3r2+4Fi1z770VbJ35Uk9VU0oiHwi+Ipwv
qR1dggaBvQHzNS+jA1zAhOfC/Y/u4Mh69L5TAVOc4RqFrrbQY2hQE9IdBhZAs4vb
dvz4IfHqs2Lm/tSjFlHAHmhF05BsWRvHLxTKDBdknwZ3uKw5wHFfXN/6pTEzR6P+
YpxWO7TZWxTsGuAwHd52OdChChnJkn9gnFUVrhJEj2sXI45D1GMt+Nq0CVx0SvjU
5CGjaxF6eHgi5/RQQqf4fzDzORkcQaNop7D/HHodvEPDc1cmG0LjVfjT4gz792YX
e1G4C7BsnIbQtWDVcMMbB3hLPGjGXPEJGeFO2VapFVWdGmH+TvsewS2AXocES9D9
5MbudwNQ/FEuEFMrR12uKvw/q+SWS85xaDgBiqm0ep2bG8PcCmyus/rfnR3hx2b5
xLqwu52EUj0lpSrY9YH2+hpn6+F6Fz1WTCLkY5t9JXymWfBU5cuU4gx6MjPIXLBx
NS7/zPpJSeumO/U8OjtGGnDpwMNVg+YylIFWFvwQ1EyZT1SPaZ28ncj9m8YKvgEd
H1ViRIVgg6eWXrJvh+88iX1d1FixEU6cOhaaNlDqDPIbAR2RVsII/yq1q0L8jWhy
RAOIreCNn6WRwoXYokw3QrAD5ldnz/kXm7qMDlzX1VhyUd7WnmOFO/06/4QGvBTx
xsVzTxHmrsQtjsNW9YF3kY2KPfa22Rm7Xu5W91ahIpDOggPtVb91L3sWWZdLeGYS
h0c9Hb6mSTP43MqfnPIRA8Kh739KbJqaI2Ja7XJgbuaq5YANyn9T/WQvpkTsDAVM
h9Qlitu2hShfvfShMLn3jQHbGf5RqsxGlo9ngZ6ClKqcYxCDF1c9aVmCqi/Zsvwp
M3SYV612akkWsJGffG4+K84Lr6WI4VCzIMWT0j2+lMzWJRnpQvPK8YJ/oOfVQird
Enecut/FI3n/APG3HvvYw358f61suPDNEB9Mf4jE4ylnU8+7/3fietF1M9hGO/mB
5Ysh6fhDGXqBiCyywsqw2PuqIoksuohDaSutUQOVa+BO+BvDnDFNwjjGHaz+nkQz
rU3Z/W5sQKM5m/YMtIu2cyupNnY6L05EuAA36Bj6E+jkEmovDwIjLVkDYZZl0kG1
bBPuR3ARS4RH4hiy/Y8DjPIfshcnDy/83fYVpEl+0GbkCNHcBNVvULXL8I/4H9np
Zddyg9iV2pdJTh2qJ48D/hOx7sG+a1wWUWb9EnGkmohiDks3pU7vkOPNLzr+oVrk
ah2DByceXv8N1cxwZJxrFLSS4fOMCUj77wxYrg3lbrLpjLnTGwwZe3o2/f5zelaU
kbqCzpx8zWpxM4t/rGQLVpN6kqWRQV5Xy45EuS7Vv2l7vwDnqFM//YMgB5CWgRk3
fO6gg0le9BZx7wIDc8eBVes3RB2DbR6iMhJj3WcY2L1sQROXNql+tVCLiRYUFdJc
QyhKEJ+iA+KOYCjlKli/H9JNGKR6jK4GbfBVaAlBIc+3ipi/03CHiNZrH5KuV+Nf
KVxieEch+OoWBDp9e1O3zJiZw00dek1974Qz+WamdiaOlD9uk/td7q1HjUzLHLcU
l4hrwT+nSS9lE0gnojwFnVIYQ0mmdzptGcD64sxutkKLy0GTTIS9wVbChnJMWxDO
UhDZyDhLHwUzneOadYWclQswfxQO7TPUQqXXne0D1fNhvDbMeGiMD0eYQReijf1Q
vh/cBdvSQbRPZfHPq4uHMZe4Iw68aS+5j4IY2WzA4B6qM2JXGUxTMngmlEM9vjCu
QxIeSjwN+jF9YWqSHhc+0j7C8x3+NX0AdtUZfpqQNYZ/qe54oBm4IawE25kLCy+v
rnbCzRwUDW+8+kiF8Hw1HrCk9AfmM3Fc61sc52EkfsAVPiu4POpl1zvz6RZJfFSk
aFiUL7jcutk0L/xMakP1YUbL66WyDVdszAR2JTzPfGThNfiRHvJZ07sv13PLX5cj
7Fhj/bLeQUL8hW0HsebqRc6+RVnCv5rbRfbkbLpcowHH0rDDSICWGu1yoGcBP4ba
qSsVQE02lTf3hFjlRJwc2XgXFoyD1iIy2DHKRgnLypQhA/0ZP87KIfBzaVtJl/+M
olxck3YUmdcFVd/4wHDXiuE6/4uoBekzl6/ic4AXG7iMs05s3264hsFXnryzmjcd
aeQsGo5SIQ1ez41ZDIfgLAvW/+kxEIHS2UNKSJqSwN6Lawm1lZDHnji+1NSNElDD
jzfeF/nXKy7yRcBWFdJzxxVzfwDAwUPlMwX+oZLK5uBWKMqtUxVqYTweVh7rfD2Y
s1hwsX4Scc7kycyi8r3hQLU3MlyfQglb93isrXitxuj32TGvVFqAEijciPdFL8CR
E9jAFNrhrcvbOZXU2E0Q9nJxng6QToy3F6O35bTigjXVf/ztm+JyVIECh9anIoUy
Ywqcw6zjp/m5Cqdnv9y44brzoSOU/MGx7xsVb/RXDigOndxy0El382gAQvf0yC78
2mZKb3xbwUJQpMCKj/IeV/m/PdvHuJZ/S4nOxF33RvwJ95hSiu9LZPyd6hS//JgX
a+rKHFQXcvncx+YxabL4TCJ19ZWUv0pxyMWnGU4K6zKGllnU2CFXRGQ2/O7iRynu
B5SVnUn8CYu3bqayXVtfstfjCV9/NgwojGrLZFbBoHtSDgZMkoKI9Ds5LpGt8OdE
DlGSsbaGoJL75qZRrEnywmYM70yNnfP+GcH9fDCPyGgvtdsM/mh2+6DE0mR4Nrqq
qlk5AneHHfzDLMjQQndrwtqFox7WQTED1Ah7GMsRYslNC2MPG7D4d3svZ4PS4Qz0
Wkbk7FLthlT1vRqetYmr8f5zXlkG1F2t47RkVhbeCQdzsVbn1PxtbmvLsyCfC5c0
b7Ar8sMlKspAX7TAvQt4qJXXofEP8Gxr4toa0Q98rx1jeUHBBvs97kdFZ3PFjNJ5
BlLNOfQ0T5e+DfSf0FblRmtThrTTxyUW4nviZEBzNOMX1gSSC0I0Z5rjg75uhv/c
CJVfh7MvavC75m+pkKPnpAMnVMV/uiNaSuSdCdHh2yt1y4av39Odx18h5bnmcoz6
jdy4d3tiI7K/q3rZsF1pYtGC3jj9UIazt2Z7gsCZcdBVHKisnMcMkacXNrrTI6Y8
Od3vkdehC2njDYHzbn4CNl+zisXc+h6n6CLcbB+H/dbfHORN7R8tn5EHsqMlyQUD
FlEHYX+KBWIe/dALJLRJTZYpedy0BH/x0RzAd8EntGJJPQuOxYvjYy3jlYUIoxnL
SAHq/LXFldleUTwno1J2pTUIiyFX6lWnnCjbj3KwEeWYTVCpofv7bwC1xs+N8sOh
QbMZLD3L29vy82ZrJC1hiMSYv055sMGddc4Iv3zU85AFhwtjLr0RC8BWrmIKan5c
QUPx2v4oI6HQ9m474gjMdlXOo40hRLVlGGEGfW+q/b4bO8j2HlYCnn/3/2e7mCR5
x8QlJ2crxoSZrf5OEjSKpz29MclYPQBo9PJHGRCkrFkAni3i8lYuPbmQnZS48Mjp
jno7V+CyJj6civ7UeqkwS1LYAngxcB2B+nd4VVeo+NHhRce39mOXRxzBg46nsVAe
WxWXCOEuOgETM6glTbXtiHVO/mF5iUaGWqCre+7kqVtUwAzHeB+jhWzoWmonqDMq
3ZC+eNmMJJY5UxDwh2jfEExa4k22i1rOUeZ7rDZ9OWMmiLvtZZP6LpYNQIlZXLhh
aSmjBLN0JYTYK8cVzYcm0UCJW0xN43KKDoFI57WFVF/YJ+CHKwr54yWHZYjQGEEv
eIO8jfenUt/nLOlVtqGjHqggLJ9o/OK/71z/YYVnBWdug9BVTqJQNSQarWtuatFX
niIQ1GAMQTnfQCYP1X/zNpaBF4+XY0jghxsyN/F2KA5hBf4/P8xtU1waUc9CgVxk
cTHF+cFFGvua+11NT1fRThLpmp9QX71K2rrq+6ldxcho9PjzWD2DzPqXrzuBRDlb
93vXT8+uJ/ttkO7WxgLWBIm+BjeO3k0kSH1wlTjnAl2pl2Nx+r5t9n8S1qOfC68c
HdlSHFYDYjxcrmVtNK3MgREukNYBTeyQISttxBFFLZ//ISC6ZfBydxKUg1JBh5oq
oYXcsMFzNh3qdXxYtyUhMPlkwP1sUJgKhtFIVk8iIQY3CnjfY67fHkOKfjFvpzKX
rkvmdID4/bCIg0kn6Iw2RNSOiZ0leu3WGD1MxVhHQrt0mjztv5Lu0jvg/Z+X9ita
R0SEm0ZhhRKFI98Li5kz5uhVFs9tmDSwAleV6Yr9os8xMoat3Q60boj/KrZUnY5i
+X5w+wtxo3luU9+55oAEketaQzMKMDdZDNzRKiX8KNa4E33G/HDplQH/8cBmVJWI
57YDCviZ8YCHUWmT3Rgoj+nSkmjUv7HehwH83oH+epgLXMdURU5L5Pb/jR8YgJBY
bkEYllSyo7FrRX7tkaOrg6gu0a5XIMJdyDsHxWjXANbtwBqU3bwLzeAegvlhcBs9
+B4tFUqZu4S78qbH2v2lCGpxG0A9b/ODQ/PAfSriN/UyKQ7/1iyelxOMiVdSX3LE
3LYdd54AJ5niLME7dKCfsEWarfD8E8cJMhwOT7IkndEqzRIrIGBWLZDYmEHzNGKv
oCX/7H1hIE3a2rN7Dq8mhP84ws3xWWR//cOBJboMmQ8fc5/NakJ4br82tyVu50Ay
fW+ppnuQWGcZRbf9vSAKm65xM/Fi45ZFnNfqHPaLm5zlYTOXf24N8x6TiMPN1XUm
kJYAfD0IJi8rEJ4PJFb/CV+lIA+6rAIsFS4UVkf5bI5Xe6Z/WBEDUTgUb/mbnyo6
K0oYNTprbZinG2vGIPXDJKliyE39+15njxZjrL9BjF/6RO/0D2v+H4d33rop68Rk
uPg+/w+gK7nUB6hhGCu1sl4YtVm6Y/VEi3RMauTpSgm6t/Uf8qAIxH5n28DWbqR1
+D6gDkVxfYvV3MuWr41jE2b5Uao3Tysjn5WTIIvJGdqMaUakytit3U8HzW2hc99A
FhAghFmHSABWDUcraZqqj+rOiw7T6x6wTWag0y6cJrpGGLW9FPTIT5/lKBSY6oY1
TBjKf/RiA9HlTWjwyiZxATAU0FKZnRXrAl1puBHB+kq2sNO2iJZirgJ2u5bmGuUS
IMui/08jGypOuX/GH+mHVh8mGawULOLZU781YcoSiyqlpEKi9m3s0u59i9oi7KcP
RvG3Y6iZBRMCIokurqjREe6sdH/mZrX9Juu+qUJ51xCere0iojtSd8fBQqmQ+tba
2cIwjPmT979KRjYQyvx3nAaoI2Bc72F1nF4s1TwM1qBNgmEBBZ3G1dKxuhddEUvw
7txIZghKoxIhQ97pdJsqRZ/vcTsDow8Tl9WkbdUP0Vjczdzhd/CMnNgP4dR/ztbw
mqRNEKH8Y/XX0qWU9b7UTFVhJY3j+zM8GaoaLeVvmeY1NIr3R2pgwxJ3TbMZcsPJ
gTfXvsygzAKXn4JKaRNtIyQr1cZ+4jZXKh6zTE1tE5QUrpBigfoAds8ARBgr1yCV
FImcSTGpZmQcjPBtOfUqgL6WzbPQYeGkY1G4G4QmxC3cA7L8cod8icmGMuHC5lt9
Tfc4rMZi52QXlwWAuMGwoizmL+LtSjwsGU0pLhORyXng6JWUEHukdBaKayI9ueu3
sU1R0ed7FPIV6/T96axeiJu6iu7liKRmCqk3O/3mR6k7LFEntKcGzjuR1aTjQytK
x+hxdDWpqb2Beq6RUkuPNK6ZVmL2d5a6TWH+zWTk2D3bMe1rlvdHx+mtC5JDiJVn
Ljpx7pEdZ/z9FuJeSt6AkyF8suHi10fUuG71yX/yeB7Y/4U4jCFIhJuiIbIY8/ZA
l761JD/HU/oo7vWtmzyIeERpEQhq5WrgBjn2qjr8fPKyq0VANSWQeWxp6BMQKl34
h7TM3G1XKZq5rERovMxmml9bSPsHxqmpoSSD/WcKMKHt1puNrQ3cOxXYpm7Fg+MR
zlBwwI0fNpVLHCHvgBScTW2OGMGjOIY4o6DLWkO8egI0NG1dG0U0DZX2vSHcHiAg
dBAya/D+1CwCHHe2rtOFryjmIn+CxGbEKyASTsZlxzi1rbnxe3vaZtVqFk30uTgQ
ZXyxY9UDPZQkxJ4SrT9jUMeYQxFNrYn2pyt8m0s5aMfFKXXI0hppi3PYBsNWtFce
ammpyT83vKyMBMglBmqCmX1Ke1sABud177XQoHE1gMde8WEI/KhZWV3+J8F9g8WS
Hpp3EZOG1Yf/cNo26pI5rHLAOxM0GP4q4RAtbm6FFNbvIUiclrpJy2gCQl/fjK76
4XJychUNX5c6lTv0lRcj8plQwhCVEB6LRRGfO5/tpudCQMKpB1GCAHGTly4zL/1Z
O8aStzjnbhSZx7lkg12x9WlHNZsQAATsYhh9u6B1YrOa90LGgBQVR+O0jsd2ifk8
54n/Bpsii0E3sMkKgU9IUxKbNbaKtlms39U7ev7SGaXJLWgGk6ZnPnGYCQIY7595
4PKPZGdq5Crzfk/TijsRoW2yGj/UUzAe/NqA7nD5E6W4iiUciJNxV13LxEv7z76a
vzdUgGsatYy6voVpFz7fuY17rnMwgA9V6WB30FeJUTbCpg6Fo5OK+w6AW/zaHPbe
2MEwsrVcAFIrSo4seM+L5VDyw8UNpvcQjnmHX3PdHt1u+1L06SeqA/F9tmNTjfwe
9lzj+whsGbAekYhtM7pRW/z0eqhxjpVIE7OR1s72YyyPk3EvOvUsQIIfTbv7ihEr
yPN+ia03siY4laQrOLVAX2tduB5MAWQmghcO12/7pnksmcG2ssDsC4eGmnEqhCqt
5uLR4J/xMpIx7wij217qDf24CaUtbHkDSz9+hD3i1WZF/McWnUeu3iAbqqJv8DeK
FK2E1HD+S+2jIicNw7anMjXgmTzUIA/FGs9jmQlsA4RoYTtvivOljx5koW/KjToG
rW5UVflb8dMCZXFOnOhqECXILEU4heIut+x4BqGiAGbheM+c9MlnxARYTwaWdpT0
i2kVWVvwMEIXUkUmQEeq10WDqOVq8dJ7o7S9Zpm6ZEHBDaDFfZ1UxDmRtsGNFH+p
1vR8ps/DXtssDTrdxQK5XdYJu5UMf+yo3wXom77CcjhSR90FVxPUK8ed5vfgwm9y
SoOUKYok1co/Wiu21rgB3Cmgl+v11ve5caQJ0OXOHj1owWQ0NUVKm3spEJZTAKEN
5x1X0puoGVMXn6b2z7GbmEH+ymOxCFVVawRskdhLe8XFUXQH3UDMxbLy+jUTRUVZ
rz+iKnMhqrFOesrBewkmcyQfG0tLCqaxkJDvStxjtDGkBEHiPjAru4sZH4S2q+2J
JdSOB1woTwqpuoIgditls+RERP4kS0M00NMUTbHgA1wWQEnn8mWKmqrIVMKB/XsP
k2F1GjKiUlAPXjjtAbHEnuERrABz68Vjds00OAxfWXCHYcefYKXBPjA2cCV4ZyU4
4bT7kpOCPGZE14Ijj+oCLuC4Oh6+So+pFC7IVA8+U8fwliNpVN3INhIj2r+0tqmW
rPqClpvnKfeMoS4w6VimFqpU2IjGXodD4oY33ziMDF9ykxhn3fJjtmOKC5CQBwqT
l3eKJw+QqPNIpt29Zq+iGJR0KOScbkjsUTnQ4+N3vCujL5DBNDP+Y0V9hjyXbK4m
fnC6GkizjfUVMXwA7UUl7uMLYdpCM3wFx8nEeZ0HKsVMjhcaDncuwuJupHtXNaPJ
kQtMkTq0Cu5RjwJRyiolOFJSFv7luyPGG6h1fJmtJ24xptBPAq1Bye+EnndG7plt
d2uu9XyH2gdGp5RDZbfNar2mVpWVhASA3TZ3irEIcSSRfQd51kio3lCmmw0Lg1Ea
EKKxL6RIWcILHcosKl27lhD30Cg0k0h4biOPIqCBNI2hOZA7cTP6WLfjBVvnECJ2
rQsoihH2X0q7wyNCQlr4C9LH1m2gdd1hN213CqxdNAm471UEFTn9S5S6/gFG4cdg
zSp42TRN7WbzG6UPqLbzBmucNrrrkyiVudTNeIHiYoE9q8rHifv4fvLP8VNIJuM3
FGw4zY199mLunr4aUp0X6mz5DxI9Zw0AdeVPym2rbJj0dMhheLz/oaTAOH7gT7yd
3FmPPLgWToq1HGpDItbDHRUdmzslPsiKZlTkZjOlMnCrC42Q/eUoGQtddhEoJZoV
JFdmQr/eaT8C5/IMSahRjLBS3MKkDgGXkNBQsLyGDL/irQM4K+HxIWOAjppMZWiU
3Sk6p0nBGCsQhJdnbokGl6jteW6zXAzQ3WR+l5dwFa4OQZzJ4klutag8O0TWAHd7
Z3YhIhk6ipd5UNAnUnyu2vV1Ypqp9B9KTwUNVzZWKOQUI3ug9vosM3wJbvLcJ2wl
myGG/soB00b+MZji1xj0PYzkMf3BQwZqEnQnegPYiAANgxuIInoX3tzuB/Ui7DKG
Fh/ChaQPfU+KXVYB9zYq4ehNA4Lao9ON2pGVebjG4eGOx/oXfwB8viAoIwofZqo3
++dzFEfBZbWyv4nAjqCzqcElqXvKgvSMx3zNzine0XRK8CB4sw4Suz8yA/zZ0zcL
WxuW2HidVGBxn9nGlflP6kVz/AdSk4xeWWOShsU2ErRfmoYpdjW9X3L7JikOnzmz
ZXrSZycioyCzDPTAfEnGrm+rxP2eNXgbpDzPuV1soaqJbDHwZLKJga1Up2ZevfyN
dM7YeOCO27iDDhr0JFtFD2swyGr+Z6m0w895fdzlHLWOOoGE5tht6D5sdGrNnWQY
fbNAyrfQaB8BJsYKbG29UMGQh+31Kf/8KtmfcggRhawCduhNAYpc7L0aONpGb1aA
6oTaIaUk/Rx31jZAL3/CPBHVWqeMBH26n4aKmD+vSMo0izH/ykSBY6p+7aRbvKsr
F4dCudlVnnPUGYpDK7vX4goXu76MaK4GKTRxlVGYlDDa/6wcvIjTXs1W9IqlZYua
kqRCRPrj+jltpLR0DgBrQVsYzqY5Rp3LeTNTNC5JLmx+/oA51WRxCFldU+6kLij3
bXt7WsB5sYAJ6/VxYUfJ3VANcJ7Tz+nbqpDwIebB3k2gpsLvKKIDutXzTY+8RFyY
Bur8m44rlhw39BhjecCkBFbeELUlmoPmzK2Otm0F90b+TfeBEGcyWpOLdLhlFqRN
NH+h7dcwuYPWBfWdWFXiUEvfH6M1neeCzpaFYfudh6IQ5oX7hPu/axLGTU9FFLTl
hVw4i/6k4t4anzYAmxXJdbGeTF2f9vWJ/SEXjuwNxrsuAuVnWuVqTz+eX1u8krII
77GYsaw3F5BfPEItbEhogwix9+DFVYnx7b+oyyOtaAG4+Pmdx1sYPt9D7ceSELxa
rjGMRJYWZQt2nLQT1nXLO2aZk96Y7Z4hGJplMEs5ChazP8wf5+pOp+M9SHS/5G4U
r+dJEpJvUp1kn0TyCducondQJx+VO2SP234NK1N1hayMVOLP83L1CRtqU7l58G1A
0lDR9sQuTSg1iq5u1ZA4ZulvwQ34d574fXFk1Dj8t3lvo33jTWs+2uvUAPUXZtfk
FV/B1tYF/wVCqebe4pPKSzmmi51jzjgz/AXAhOc6ZqjeraGeybaEUIBEqhKKT1If
SAgbEwmAnD4JQz7VlyFQAReNUKefYix0vgEXrrJ1Qf8gKZI65OR5N6EaDQjwv9Id
MQ5hZ0Df4GSwOiLZ32iMctEDshUUpgDUdtYfEqirk4rZTSOqdkl1/W0C/kNeBvZo
QwarezJFDmHDxvmFMO1oc/DkHCSNw7xU+Nbkuu7hoXSuXj1mjXcZkqPJctrHRWT1
k16jGbFw1+NVhaA9JUBroralAuWIpdG3ZY5L/d6/40p7lgp+99VIgA3i3lQe1Re1
zAkfJC40I0Q8mkRYSVPj3jJkcOBQEPbLnEnu+RWBwDhfCieMANPFWRCAi+UDJ4gy
FulgaSmUoyRmoV9njSS9IRNsLsVovxTwkJKXMQ/ZvC3hu+b2vFf6F0u5EiF8R3Oj
sJlYSxG9hNNcq0xn/nWOvOLbBWrXE1KV29ErzzDR8NGUmGNpydzcjOCrAeg6py/S
JHnoZrkJlT8ze+S8/vKnAzOPwffguGI8aEkL2QfmBztOYuAcCmhrGkLbzRDFlUOF
ObFWTspuP2hrr/mJ9+JFwn1oE/Hn+oZov5Vn+ds1x88ezTggwjbuM+yuoxQoENw2
K7uYMRi8Vh07KQkAVCEVIDKXrEYyVY/zGDtWBNP5IvO7M0aR1zBgLXiOvG0dal5b
vOKRQMoyS3JNbVs1hLhTaCJrjsENC9+rnkm+ANpPdDLJa8MIGh3w4TzFWbthTa9p
g2k5L9kr75VJ4qBKRYZk+h5x9pAUbvMo4LGxjn79O5Gp4bP6Xs8dz3a9Gqq1smVg
TjocMOR/2Z7Dw6Wz5iSPUpVjI0HJe+CS3aF194uMhwOVxAhB3ebQkvwoETTkgM1d
PN4x94dV7xWvDyroMc331+rlzAWx/qn02DtzQPugNteotVRAzqgVl86CQ0Snu1SV
J88sqE4mgyj6OrSq60yJCFPTiyrivBL9pcHxfY8O/rubMtIjAldsazzX6S45hBW6
zr92LN+gQyFWRf/d03luVTjt2MIJKHC7pX1qPF3MsnGfFP/RT89fIQI4y2nUyy6Y
v4aEWXDsrEefyUxxwyQDloHRZNytNFr0Y2EvQHTqPMO59Hzz/SNp7q49elYT2UVp
RtxmJl2TFz0MKTDbwcHVpfpIHsvQ2SPLyZn+pKCyeVyX/XaV3/r5fiPUxZp1RaZC
Gi6P+Cc3q+7V0e94JM3mM7QsDXcn8q8ApWdpBfwagRE/EV2gFwYzcEwby+cP0hGZ
YxJmPwtkXF4dcqiVRs6AivkAPJKncF0OE9l9nRbs4zfFOcnurL9iDMGPa1Hdxz8p
XvQ0fmp2UQRn1hQS15Q/BFkSlNQySqWW0RZzgnHKR4ftLXtxIqPM5sBzg4XSCIB6
5r6pm/b9d/FzGhF8iPWUQUQF2vpZaByedck+Zv0pk3JcElpZ2K6b7eps5kNN/QVV
ttU2jP2oBmoIUoLYpmSSTRPv41aeK+gixO3Gc6ov27rERWttg5lA3ZfSWXvIsqv3
YkSpYARmfVv40z/C4ym4/w109aryc9d+jKo7xPFE8lvcpkiIN8bO79dabkI7ovnR
F0ArK6dW7RNFuWVbFKGCg1IhUxh8IwCpkMLqpOAO10q2Ef/oQ58G/QOPuOPB5jhF
psuNtHxC8RfoJVabNT/TP2AqbMHfOnK1o4mXOs/GD7MsCCtC1k3B86m9GSnQr8Fn
5uDOy++FB/WQUYYxu9vfHpuC5dONJwS5DpA6FePnhT3TVYSEVzMG16N3zD3eSuMV
ScZPViBV8QP5djnL9+3ZcBW6luFbXFH/4hqJBfud5H369U2yh2wJj/ySQ7MPOO9T
YTOImxydQKMDfyFB27FcglwKVRbpP4Ep9DYpxgWy5e6Nd9tPaXV8oJee+qGtII8G
95j9JhFYPfuV0wTIyzXg9YVB1KyehKGAakqBUCa/wixGAoZ44n/o302Lqr8JRLbg
qW4SCWaOzmAm2LhvtZBmTMGTdowJQn7RsW3q8U/vnxdyXH0v7qvk3ySPHaP0k2hh
fxUdMKoQVKPao8I/oc54axKPxBPa+5YzEcbwZNae0Cn5b4q6P+CqI7K1n4enVT0k
hiTbLvmsB9/jZR6NmxGw5qKajAZKt5KsCrxSeCHGyxx2YprwSkfgEoBfkwFpJ/te
L4gaUKHT8GFtO584h4Zy1IzRVwYJ5rhtGhwH6EBfsF00Bu/jXHcQEmmhseDoJbqx
mw2FtywHYiKLZci1NwaFbSIDdAkXGxkqIYL3F3YrvauRLkzAIOBbCNxU+KrNLKzT
VZzQE18Twm8JhZXlO+JLbS8KkugAjelawJM0sHPTTK+iPOY84nPfBrzvKTEUsYAw
Zjrbzfilu+uIM1QE7YoQvp8B+Hr5PbaPUYulDACowQ/UAw/s83OnDmsF2aJ8UysT
RYjnMhKLkVOoeRSsgt0YwoT2Y8w+qUpaepqM8r0t0QJp2G3Iqg9/+3rc5M9EauNd
ynKyFp/gSEfkB5HUoj9HdE/9YTTt/f8lvc2T0kh68vvIvuZyue2ssMy28DUVrHD1
nVnSouMwS9LWqm6iFVVRYoZwH/6XTGRvWeQpDnAhAxrlYGwq65aO2xtQohPFSTjA
z0ex+Vz8Q67udQimawgUuNidSnkeoOUE5usugGh/pW0zslWmzprsY0luhIjPzHj7
/Ff3Yd5bttb0XZxcSDw7vYWsXH6HBh1lWMB7QZgIQ3Ubx5RH7lhE23umZx9KjHw2
7r3EeYVFbFQ6P6RrKJREF1dmqt6ez7ISmDTY60wj4EVEjMcA6JkfqjEd5FJ39eyt
nwekEPBwQOZLqc1TdC/lVdWBlgO/Vjku6KHBJlcISNbUpqvJavufgLHbeAlA43qP
yVygIITEYjBfBEg17ArXlWq3wCs8dnsdQJ2Uej12MW6Seyl/ZUlyJaWflg1ed2/E
0s7wofFfVZ0J5Gw+YngSinwDBlt7iKAo0PXooyNTs4z8CKDrSYVSv6SlnZmmb6u7
ZIu6Te8y6xdJDPgVvJDZS2BoEkuuBGo7Vab+BEIxbjU93X1fVAsv7bUmwdNbi/p7
4U++oWOS63Myz8wYnI3ahPHsj56VkZtpOpeVF9uZ06/Vcd6+YHpcDPT8RbOIg8ou
sT2DdV25SJlmcS4Q/GBv7wyH22UuJFfXo6d9MZleUt3rxsETETnvFBIAUtuzAXuy
yt6w8zt3SZJgNy0S7iQj0Pn4uBk6AKZxeAWinDHg4vmmiwcgkGz25JY5AtksVLgJ
EqvhLgKuH8HVqQsIgLiOXkk2CIc1Cku7HhR0jNUKIfo5964jGarCAEbfw+ySDWke
CdwOW9eh1OLDJjpnZWI+dXxpKKAN2AYScte/HEdj0zVE2eEDwRtp1kEwwa3ps97C
+8gMbk9YAF14vm7JJ7cvm7SCtNrpYav26c0EHENnk1TvChMx2tRUr/kRYv8cossM
TdxNUld/ehmFHPLckQ+7FOjUlsJ994Iof+UCnA9mO2WwUN9lNMIx/QyDDrIwDigh
G+THyG6bI9HiltS1pRpwS6MkS1mYwStK2aqIsQq9/kOrNoHfVk0qw19QzYit9E2/
YXTFOrw2geDNrh1s8GRH6mejRk2lxNkNByqphJFZRDC2hXyNKnsWNKd+/0dqJTty
gSLkM7r2cAO+xhwjX1BrDS2zc7bN1wWSF7vdvrGx9x8YeUTEiH3Ekd+lj8Oo4rU3
3FSQsw6vPY06KQSrm8X/ZbIjLbSXLVQmm2sfeCeRj9+hgESYZbZjEm9aQCoUVmir
BFegTitwPpWDJWF/kdxSmHg+b8LeLX4CY9z4ziFaZYmmz/0PaXQksWmeio5z7uHv
LFKcI+AkZwwhHldbuyZH6DsFjlD0ponyB0rjERXgewSYjRaqfEvFdpv/GLJqHXUn
iOoDw3ctWdw0PGPXjqASzZAsAD9/Vfy1ALRfhl0/1fDsNDhIh/dnApLvKOJGL3OV
/VfxStaLuNPSWz3lXCJAYEXrAK+VmFmAbnB8v/dyQ5tw5pUjVkV42YS/4WOX63Q3
sOdqOAUmqarUoHtRH71leSxwWcXzMNLjyNdYlIdFD0+lDHkBjCKsl8oxuivYxXvw
pt9IAmuA/Xts/8WAteaLZTjhzi1+AcmJtquBlCavAn9MKzJ+cSMqhMOY+uxMYzSs
4ICVz4hsaqplahyFkZ92t23KGPhW107EzITCLTqkLSRp9bZ47UHaBFNFWoQDNdrE
d6LUEabaTwhYqHgwLDzY5EDPqq92koJLuoMb2wRQg0KnrIwNydJ5XDbARSEXwQR/
VDSdP6Cj8KMffsAEWHiPhiJMow6xFJqNaOI7ftEBdHRBTRsY792zbbGWwFXbk2av
CLOOnE2oyGT8Zhg+UaotCuuKkf/qqIOgeqqA8xlJv6nLVDm+pRYKpHBMryRtGJd3
lrBX8MOu1pGA0WpikvUYy+2RNXCDeXrR1CkpdEtvhYJfP2wTsBg6hnskAJ28JCsI
cQGeyqyLLp3XgKxHM3pKF3TI2ojCduxVLU5sjKgItSPsXYtFAaiBOjX4GFcdeUZx
R6j43jsZdqVK2s8eQkGFzD5NCSi0VmvASC4HRxF077U5JFnF1PqqbDQ8tk8BTRq2
257ifQbGF/0BsuzPS43ODyf1NOQpBkn/yH6SrLjfmfsh6cs8lA9ADzwyaVyDyx8N
1EvrFfh4yyrvN+VjjYdSxP2cJ/iU8NfyjeWUjBFSuAQLMgK8dBkxBaPgvqBReYYi
towKCRJ1OevtZ/zgcnZXryGctYXozmWE0o19fw5c8wzUowd+UHApUJzfyTKo24eX
mmkQNEWCUYt56z+iOVKuLW9A/XlSdrOzJxIuZTIVegnFRVa0ZcxeHaVdP+TFMyHC
c22uU1zsrdkBprXOaRfrGdO7odoFbPK36WdRtLaQKtj2l0QHZZ/3C1RnNrOKT4r6
ogojQ+ONamrp6yTjYydkehNt1YY+YUtcwMsAwWGIb6p4USfeTN8bKQmFYIKx3Bab
08pNw/56//+DRiHfpCuiQklJcCrSH6e8Uv/SxT8Ac0Le12ESQexZbVjruoPTF3ad
K+5dbhtNfw6q9mD42uT/e6aLZHRufW6W6qQn4cyLsNVtuZdXa6sV5tCaONXg/gDY
hcTLY0G2fSijS1bliacQrhb7DNoA0SgFf9hKu/0BqSkfy555nnKgpfTY2YE+7rZj
D+ISro+eD5BK+Tfwlauf1sknfQda0fivgimfBmNndgDiwTl/MZustYY9hk+AmyIE
ff+ARB2l+xzyaK0LtLBA+bLBJLn58JPlPygrIaVDxm25k62OQQnjDzTcdqZXY2i3
PtOpDN5v40KX3KccezkAZoW+DHPS5vA2A0/JHCOdjAK3tmH0oosTPOeE9jFAkWdC
Lb//suLTNwvRYNEJFU4pksg0g/VpMrOzenxh1B7VkriPstY8xXTfcY/eEFNKonhe
rqq8QczuTBM1qCnfM4lZ9m8rXYcMLpvPhNzHon9nm+vUFrGlyu2ikKXFpz9dBV0J
ZzGIaW+m4h3NClV3N0AQf21UKWTUvoog7pXiytvaeJJKUqeTobXJK2VlBwJipGYC
O6F0dFxpIVPXJfdQfCJx46YinVApCWRhjWdZo8BlRBixZM7Tyg6gcNYqNM0y4ydi
jQqjz+vxA4fU2abqVCWcuSvYDWQ4dxWdAMZfAldLSmP84POxdYZDyuGgguN6Us5P
qUnl9dqjL9SSe7PpggOtcEf30INCL6e2rCES5mqOcN5cBoLzqmL69E9vBUPZHp+3
NhCkixoXTrWj+hD0YlXS6k9xKhDlaoOwL3AWmn23Z+rDsEtzOl/1SDKCrq08camj
gEf5OZddvrjUAyQzHF1xCKbvf44KbhP80ZanW0n5q9fmJhvmpvVDJ5IlxVjTK2Xf
4fJL1B0abdDC/hkzXZh6lCFnJCSPg0q4YVHSTczN6Nf4zlkoClMvuL2HqDDT0rDx
oW7rjmP77hJ+VyoP+QZSA4y2xLk3Qv6A2LgtryY2hk/2vq6gDft/JQxPjYBnke3S
CjCubn0UZF/Aub0sOrLHsEPlL0DLUh+dt2PJ5K53H5pUebopFEmipKEGvx5ojSyc
/YgTRPKmRactwrmG5wz/3ZVoGEoa9Z86VIXlcpbLPCnpKo5hA89p+G62hMuqUURU
CrCMcqEvgklNcr/fkBkAyiUwxj0yPoFdhgr/DYLIyGQUfUgxJCtCucYZVbNsXBUR
dHRU11LskCDmSTWcauCXXorDsCkC+VB3e4EoolU7FQx/0/b7jZzREcydVZKoJcPj
n1QotpNeR526Eb80xfQzfbyjbmIiQ4Fg6geMvr0dTtIArKRW3xdd+6+tYvxbbug1
74MJzBFKqB2kIjl2YLQvHzOOrbGB5tv1roDO6y2Z73e7WmeYdaOPNfr/aJuWcUSS
qOLPQC+sKfaE2AWtO/QSsOHbwbrzcvl+oylnqr4WKubd3vDOIxMAU335HR8fUK2x
noTpiwg58UadrZKGu17Kxzow/WR8reobELTTXj8kj/1B07Xpb5HUVmD4xY0BrnZH
LZsL00Ybaz3WYMd/KX43LtdfC+VDgd2iaxt3AIf2kZZjoew1fwVXYxargJ1sq5US
8Gux6S2eBSAUv/5UoL7jq19WoUJvEulKhxZWhoa88cWYGLaet30h6soNxVpJQONb
321iDuggoT3W2KeLDN4Rhz8QNnCIAXZ4TAF+WJePdc+6Tc5aUemXMowAZQaMIQgV
9oKCvIcNTFqwm/K4MAo76WO6iBBrh0PBON+2qj9UjCuGXTdLow7pA8KGUBLAYoLU
0eBud1QpQz8lyKj95t4QSaDF6t1bORiQNTQsJnLrDqE2yP8Z6/hOnpN4yJgsYAcb
Uypopz/S6PC8ADnZoXZtZtMLnQCt6SIKmqjfwVlqTwjps+8UoejvPJpz8FRbB0ro
LacLAyVFYgnSJNb1FdhToJ/iUi9Hc2RcBMhZF9fwLRCm+AlpUEugwwAzO0BQ1Ar4
X+1gm22s7OO1AMb2c3YYXH0eXHj2MztBGnGmIi12P8zzL7HMliXioqxS7ykNa2ym
FgqZbK/ruRRNhzo2Dr13xX3hwYcAffb/P/6iCP6vSI5FwunWNH0a7V21ZATgcjW/
nmKzfeJUZQUkjgLUtdhZAUcBCMH7x+qC53qojtmevhTuE+jWU3epRyaFeqfW/UZv
eXnv3gcNHodLQL1k1M0RYgm0ZlPnif+bUyLlx8AdkdgikHVTsEmkVYGU+QAKU26g
O8/1LzTYvdzn703gIpP7TWrgST3mqG6vi/Er57W6n5cIUPhXmO9N04pu6YVWcHfA
8ptFAaFqpm90DB1YzsapIlort9KhynNTMVdck7czJ6rXgU3PkcQfwNBqdMwsclQR
xMZXt7znlNJ/qhGHuODOCVv8WlnxNcWeb1hzlWUZW1MBWJBJRNTRDbcaL9BYnQi7
syrKWkTwYQf5N8RkqGQPKf7jWH2p6s8TKcWU24uGmlFMh/BjPvmZRSJrN8jhfJl9
7qZ7p5tNZXFuKx5Y6TBTFFYSE+3NRK70ow25OAhGwuVSwqWH6RCO49lXFwJfWOhP
z2LhKDBpLReaSjHUeBjvzrDLQH683djdLYDthMU5pZE3IaqJWFeCId9XFN3brGQZ
WPbvTazj3wYy8AiLq6KUoXgDWoLvwQLgm4flVM5fRxw1Sg14dW9bOf+dQzxWBO1D
JUC5QzFHw2vUK8AW0xMygPMz2jexR082Wm87sernSdi0Pxb9LpWER0VjAPy8+Ly4
mqg4/GuKEgInyOo2HKsBF/enAcfdFVvQxT+KSM2OCcfhzyZlN9N/NJ7qzM+MhAIu
UWu2YlmArBrg8mn42LBkBWYOTBrvgkPSxJRD/l8+UIFgQpaRjc6cOXy8cZQ7hUfN
htZdl82CcpKmLy4RhoRzqDVV+qfEjPxQoCj+03TeX+h5GEbFMSYUCUo7teRlP3hC
kzR5FuDqIMoWukYt7OAEmeOvD2JIKB1zeEtPo0BWG9O8pRYtv+PfGyd1KJC2ATum
JaaXmWjtJEBOpwk/xkayi4ikgL8fgCxaOLfFlv/b+S69PaZ/YENfNhgnKaJgi8qi
FI/ghzPQgNzLy5yjW8Vl4qrxc9fr316zryZhGvrgnJHNqM5AvnUt4tWIVPiNBD/o
VYB5m/ohi/NTCt0nUG0w2iVlpbm+KxZpAJOVs+UDMsOlTbvtr/Ds0TZlU7e15I16
RT7j+PupMpRBIZlCfn13fnvwJHo90IDYC8wmSh+gTlzmtB0XNtrTTuTKo/KOsZmp
5Wll9Rklr9ZHpcbCPflqmWjv20M+Vu15Lz0ERdXYvKXJLDXX/DmlZNdTeY3lWCfr
I44uXQrB33t2zEb/T15EotUwfYC4ELFUHIqEpHWDa61aViq7rlqj03eClR19j/zs
zNaUCJQuCE9KDFo0AQMOzts456qB47/BmDpYFO336oSD8niuLeEIoLv5810LkV/9
gRVl+QGmxZuZ7qhMYcBwkK5S9dDgniB/iy2NNkbjS9h1LAcOrK/LbrN/9q1hipg+
164xWVNmMT1vccLS8K5ITdMT9gbE5k9pCNfhtEvH+cuPZSygM9U/f0kz8e6OSUUE
pzFfqBQSHim3W2Yv3Fjr+oKl834f+8NR/++5NLBAG+dyCH0uzwegWmJ0VnXo1Zjp
5xuPMJdtZIZ+bU2g/Br73r86D24xWnaZ0btOx74hf/8Shu57yEIYlH8CqeRg4VcE
hFjPbvBrf00pydHsDCcletaIpAtdaVaviJ+ksLJvxiIoy1MQH/pHjruoJgQBqhG4
bEnh4kHMV6qvB9gphEFlTwSjXP/V+MAthlxNVMkZBnYRSEm41Ed94Py0DUnQWvg2
CDDANpDcstX2S/cVU37oq5W2BKKsV7L3/ApcDgEzbpSx71lDhueRUp/fXEIhUAVX
You67OMw3SmABBmoaDMjzGusaj5IyRZQzbdOxfrB4AATEHdxrRfdLrthTHL5YZgi
8NUWSopKgGFjjCkLxdCusUMkDq3A6gPxzVL2J2gBxC6+jOmfnLuEO6I8lWC56xoC
A3es2gHHsNb135k0MP+drxDg/doBxF5wjiAAKhZOFjmLk0tFjaoEGdz9Gat6kk4J
3ZNTsv3E12QlQSS+xCDtio/aHBjXbal6nHCh50L3Rv4U7reZSI0qAbKmiLeMtAMW
8HJYs2lGzuHO8Xte5qa7PHi/7kfRd93wq8Xt2raFFXdXCRrZ7zFtMCKdWXRNvMws
1rFSr7vTKMDfR9Wr1dVgBivqs5zUG6+LYF6qpJ4o8dv5tXWLh00ESPv2kO0PdVBw
fDmp6ptCPn55uoZCX37pt2wYD1H2dQSknedytRvyPP7b/ZVJuA5Hl/7PkGkeqDP/
xi7K1daNkKeSyBqBjOZDlr9/aE5OhcLnGEIS/Ci1i0OgcSrpErVZvY/x1OOnIc2K
zTQVq0CC7puEWJL2VyJZxEl3CDuiqyXP9gbJCKA2oz50naPaH+h5NISqPeLMV0Go
6qvP5OU0UpwKbwgtfj4PKqTLVgRcw4lOyB3RkR2m100HUxhxa4HR8PDfn0cTcnUW
ba6VnnY+xhcE6/xKg55C2CveyeRL1CwVfz1BDkE6XybMBVAN/LzLAEY1Vs164K7m
VGQZ1MIPOHoHrDfSVhq+Jl62uXQ3l43KTd1qyRpuUoJIzHVVlKe4XQcgLlGuRTuI
oLmaarmteGfDwY0sXCsz5EwWXu8IPhOAFKUkZRbb4sXkOyjjAM4paA6ItBJ3WgK5
OFO30ZnysWeuS5OUV3gWolzrbiy8ofWDZTvYLWF4QlCSTgCiQpJsWpfaK6mvbREB
vLE6pZga3QK11GLx9xEAoYDAdj/e4hy5cU+ivImJcG43xvnLwnKbBpxIDsrXXBTS
erdXj2GfsfA7qoo0T2AhyCHQk+GXI7UfkZBZyV4yccN/zNDNSQKcyB0e5h9E0FwN
3rhi65/OL8SwHtP01bYVZR+h02+sdXrDQzsTF/OiLGl6lqYK4eoQjGJsP3AGfP8G
hv2PrPx0fXqtTPjcxYUx0N/ZMh/CYz3AVLbTz9xTWW43yAUsn9QRfO00XcyQNvHt
AVNAaYyq7KiW7PBV9Bv9GW+Sh30HTE3O30+pDNT5jELFkr8lTBF4+7ACQP7sl0uD
xcIyps38r0JVXUzN91IopLNnEK3Ar8FoGm9VS4OmAZIFdQZ7npbd/yIjd8JdiHZ9
1vQmTgdk5VoZyyU894AUpqazBP9r+D1RB2hB2jRVyILxJU0GpJOJ39YxEkrekhaA
pwIbuO3H4P2rVhybymfpZ8eyzQ855SjuSJ/pvsOzgxABJS+TTXMn0CMf5xnVUfa/
6XxXLWhI8SJUWv2mo1KkTCayzlq8SHA/oeIB1bGzzWs6mE+vb7gsd28Ps5Q1H5EP
h367pUnPT1qCY7aAao4S/FhKfDxiJSMhGVGuEtXW8IBjJQgOeYtfdMad4QpuaPPD
clbbRR3VLoh/F4t4Xqb4NauBKaX7FKGbolHFfDvFsJPgO4DbUvc8YBmI8NDnMPNC
qua9QG3E1glraE6np2R1QfnfV9I0lI19MF5IXeOLUoltT2taYwXNIP5uEZ2mswuD
UflsGZXpJKR6dMIHHHTZZ5k8//KwUIYNVk6idphmILzs7c8FwNUrtm8DOKb2qZx2
6Ez/7xFuI1NDgRfhl3sokTzwu7eg6okpSCgNk9PG+NB7Iy8SerANwwVkD9pEtHEy
a0ySJDKMwTQdt+E9wGNZMUmaRiLVV9u0lZYKXtmBf2nFQNt6QX2noYeDP161Dx9n
zsgXrNH1v7oHF7OXAWBHxeK4/YDCvLfv8SKALx8eOQB/udcbGf52LnScWi9bFQC/
R1A26pjuhyTN6FwPOdyW+u5fX9Jb/SXVXydCDKse2IVw+Nj3ShA3uVtAvFFLtbER
ZdRx+nZuu8fS1jDWW3Q/67nuVcVOeCSwv9lXD7K2auHVxYC6kqRad4wSGbzIuv4p
Tv6+qihIAtwT1h+T82xMagh0k13Eke9ggjIaDdTbshgjLA0DAdiEwiMYpEoHhPoJ
rbQo5tqIsbiCvIzYOgIkUQCaGegbV6HBiTdAobmlMoFMPvHr64/3pA3dUN85qREB
6QI4yk7+/lPIgBUR0nAkNvzoYBY7FoeTWNYEWAZ95dnSufEgWvyo4LTYfr86/Def
Uoj8n0ob6t+1Q+lnvyBRan28TQIbjqo0iVmgx5h6fQUmCyhkPYWkKmA2xNlHqg6k
fTZd+hDPc6hH0uZbt0ESEkpk5sG5fcv/TxXopGSaJQpEj4B52qVgM10IXR/wS7my
rR/FPTlyNQzphbB7ght8OQf83+QVtFRJDvaG0N1hhp50vUZ5ZCW4eJHKdVjqHqo0
0c4zaK8PC/IWo+umCgK4ITFYdd46pj3BkcRNrAN7a3iYSCiy/rMmaaDmzPxmjMav
+n1CPfr2AQ8kllPZ1ya437SyypBL9oEx9PPgs7Hp7E8yXfVRncfhtfDRNbUixnqn
KZZD4dRDHVBglTTxndoUVKlIEZbSybCeiVTwJxK5LoN9gyJwhxhR0Bbwsh3Z0ZnN
UHnzUgUkfzTIK4i/j0EjqRsGdGkrEQm+cxgL/vBcEu71sVRCiPrk13c6PnHzWO7f
r/khoeJ6JX7woVLugAjRMXtHjigPaxODPwHVBjF3B+DwvVEdHbU23efJXBobqlsZ
ZyDT2gSwjRsmQ/4Ib5Z/cVHjVXJfhPZv2tP9ra8rCBB7ECRLxYr9A9nCemq9g8ba
41+ty1rUSeqQlrUpAJ964KhlAob5cOBLGCjLxXIZ/JkSfJ0aT0eMyDTVMQbParyj
4RFIk3chxHwavgR7zD5/Nun/re7XFkA5Aq3M4EXa6m5VrLpdbxr+IuGMGWLbVIU9
rhsIcbIP7MwBMAhzbmDKBFwCgIB/CNfwMl1I80erM3DiOJFiiB0HM5rK+FSRIq9Z
hwzyOePIJofkEcc+I3oOzqQNOjmam1Kk9zjMbxPBCcXJDSwFKbiw94Pa8cGqGrDm
PJa2p1VlxjzrjtcGMekewVn9l3/EmdR/U6tm0V85ifiKN2905cVklVOtZ8oabjGr
FT0OlX0lXyrz905aEEZHq2ctm0iDezXsbi3FrpD3ZfeJ+WRwTPE1s3pqodM70BdG
KQF0VFd8wtiocQvq/StKk1suqbDX30Wc4Lz99qY9GuSejAOoG/bfFH549pnRzL2Q
tmfFeix4gIz41ZAaLKTJeMdXYJ7H423mzgF3+q4vgXs4u/jn53p/QSnWkgAIfmNK
okfLBJrgk07Ho5pEIhW3/kM6gNrQlX/584hD07YLL+NSTi+9+1lkiDK7zbo1pBtb
sjcgHAuyh6cBmX2J91wtUmrbRh3aVIlyzHRPUgvXqWm3y7euwQ2hkIAvqCVflGSx
mNe5J0mqrjfJwMZO9s+7p6UtAfPTuwjmvfs5zm9LBLTBdrYfehQH8wyg7Nqi+iZ5
GKxyq6ahrIbzviKTIEPW5gUVyVNVc/4WuxWrfj7vfJ6PTYZWIPBMHBfIw8xvRgl3
F7rDkBY2RWnFhMPJLObxJ1xFmSL6b3IMvyX/ZKxz27i1iD7wJIfD4Kol+pyDYiPL
7m7rlzc9VydxUgShS7Or5tc0Bae7tZXan2/NOqIIC+xfJxh9jvtb3mgCrdZ75Wzk
F79aQ4y9ndCP05zfkXwhO5p4Akw5FdnFYb9TAA0Q41m6HjyxkhsKsl+M4/nQeEpr
eaYmouTBUAV0kfi234ap8CmtklcGlyCH5haEHXWhEHjqLzUZvgl7yJtN7ivz3xvG
gFMF1PKX72WNcyAPY/wFwouEybr2mpKA1iKxHcyvCEmSXRaFmvwFN9yAMg5AFJBi
IiXS2M246foxdNLxMb9q6nWbl6WyYwlf5Gd1NF1TMzThsEs1DMwUYu6mojXzgrdu
Yik0mQptIg1AKVBcuDe/bCkswRaEhp33F97IzuiYWFCUCYyNzyf70qPBsMXww6Xn
7IYB3D6Yr0jXfBM/GtLKsdaudXVAallrq+8EPNNHnv9ebo4qp8MCe/gZoyAgD1Uh
E9OkBlVHIWIsG1ARpYmUTtK6uMlc/9J7S1c89huCnTlu2jrMWNhXisbwnnoMMiyt
wsT0x6MmeYK0GU5xYNAYa4t/7DB/s/+6BgpzyjQFtFcFPMHIan2Eu0+32Ap5Rw8w
lOzEjcfj4k4oKpAs5GQmEDcNrvauOn5JXCv6NJQJOD8lqhnP0+ZFtgcleJfa+x/K
isl+uORYegm0uOIhCxV4srdUYL9XE/RCgsrRTBCmM+U+kCYx4TnJQjrpxvnSqB3f
zg9eY0eNfeB5Tjt8odcS5ksOJpuGuOuv2iqltltbNggVZCBWHdb9SN/hEDs7WhTo
ZGyfY12Rw2MExxj0PCQVvgBud7wgyeqc9YeR/P5D6KITz9rCGAxktbpyOeNtH4aZ
htWAS1le+eRlE/c7ZipPBqjeAvdRjti8bBC08/IR6RxDDX6VVxRfddk/V7upwOkW
EyWxow1+m2MaBwBc5xPqVU9+JyHpol191i08cdp/LfVVzrzh6NhrRdq+sC7tcoTU
/88xNG/sa28nlU0QSRDrK8Hz6Qv6zv8VNPnsJs9uWsm6NoBHpo4ocXlUwO7GAEUd
JKNJqJ/vuKlQH7grikSnrejNi6Utcz+mYNE3Ss6sZIsBNYyV2THWLx4xudRYzUEl
4sxQr92+PnwY+HwPjEGvw6/avoa4t+oJClJTyTHR0eZlYZgiWEkBv/sekHIpMxnm
4bQwteOeiiz2vbK+6t2t89S10nb6qycSk8JikIJrTpKaZK8u68oSu42uUdpswEJj
IaBGYP7UmGwiEDOV3ygNRON931N7Uxwg/6O02KvgLHbhYms2kGzokDWslp8QUHcz
dFlcIR+Jl7lasD7wE/7R2/Ny54rJlPIlI+vhFBPbPITIlsqW8cje6vArTY+nJKly
PX4QOpyqoenPnnbEq7dOICJpvxEp5AMQBDNsj1OTzkCsJJy7A2xehSfI2Nb8WF0A
o8jJcMrekGMZBS0jJW5IdzpKYNroWK1esrwd5TxqJNJ2eGv0tq0YgSWhiY3iaFOL
MVoHWNOc+rkysLt+9MuCfFrDbPyG7exi1DdkFk0DrLK4b9giyA7pb4Ir5f+m2fAB
BEI8nD3CWoQWkRljMNlWQTAUIXtsCYXkCAyYo44bnrW1WnRC34eglYYG7WwGE4t5
RS9ivd7Z2ZhRQ4eJmKj63i9r/EegJ7zdztlwZaYLXktIysQz5Kp1aleawhacOgYj
CwJwE3W+3/EMqRF3HgoDdVnx+aLTfkKbIzfr+RZz2wFw51b7m3RAsYDLpswTVK91
rUHOO6KLF0iMBbfefZNR2XNyCyUu6/Nfn5OShtMyDF4x+7TUl50ourlxg/qvSSTX
ZpYaJahiUyTDcH9O0miSPJLqdWoZOCNWhpvVATef7K9373liaBhVxaLNFodp1QSn
ol9sE6CQo19Z82MURRMb7EXZOvAjdkKVwJbgsm4vseb3lVx6LabxOFA+qFDPqzXL
OvZyDkkl6X6czEZKF4TmDbKERqaOv6Xwxf/1mD3ZydprvY3jXgKIuYZFklY0RCLB
M1idZQD4WXptiwbfPtksN1IOIVcktgP+RbE1bIITYOasUk8yhMKsIoOuFhgz10tF
yToYsRnT6JyfPKaTpvvN063E97JmBiIsa2WegOBkCltKHOtBwyBjtd2DGw4zBGqw
1WAhSs8Ywk+3VDaxQcNqcsT0nZA1zBD93fwEBEJN9xJop5UdZLAxrGIfO2I+ZGGo
+nGgiYPIZ1S9+8ykLU3y/6pHoE6DZpccSLXyVItlr0kLWEKZovk28k11EuO1PPp3
V82HE5q7SHDkliroyr6UQid63+XTG6oTrocWU9dCdCEEpRWS9vLYuP3dlKiyB+7Q
w0YgjkKRWDqVfC9Z7AWhCHgWbWs8fu4IhX/EfeBuxv7sqIxUWXhJs7nY41YY45ik
1QgXybAh7M+tLgyt6LzqQf9rEk1tzKWZ81msG6Yq2dYLnDqsIJswq7j7aPqz/+H9
/T3w47CbaLuG82RZXZpixSHgFSODd3SfHLQTBgJ0v0xAyCrtpppIxhGdKyEX2Av/
QklLJ9bKqk9kRh0d007c2X2tbHUyd0ScNevPtoN2KNwdSApU0SRfDpelKmnn1jV/
eQfrNwlb2PEZ26PMJ4DC8e8aavM2ztX75D9Jo6SbedmhNZSGQy4YNPh4K3fqRMni
nfDaSI3XImStksWjuxEwal+ZDpuT7FAD8PkeJZfnDnkRJ4eCqvAlDC8L/XIRyOq7
JuCmBDAVWeO2p/IVBfq2+jB3/PCfe9xxYpei5A0VYfD4M3cVBE1Bp3fW1aUG3L/p
AVpKo1326hruKpZgSd6VhKDcu2mA1mLmjsDq92yHOS1RkC9U4HOsHttlOOQsuzAB
qaZrIXK8foTEf4Lpp0i0o9lOTI+hDYCxHvboFq0jq5HHJHJPJMOZIbJogs/ZNF2j
BThcIjVxkLYDm2rlxKxjotioXbGkBVGlj4NxyunXv7gJoXYh5p1aapeKR95jXtSb
eiaJHZ8EUCQ49p3ijmc1Wtdgw+AEGdZbpjqtMIeJgOiREYzn5F18OyByr6II2tNC
GjR/fTa1FMzKwTG0lvCgdzU2P4Vbj2r9r/LFIRXSKv1KOOTQFdvIv6nZNGjaG4tT
9mbYrx6SiXwCsL9+mXMknLUOt4dUg9aEY+agbAGHZ9IPqttCD6Ir2j/t0jBiFefR
Is8+RJn7DwVqBZazY/QCRyt2OEey+t8acxiIzddD+Pdxz7zeJrdasFGBMT+EIROO
QDbeWeQOUuzuLPSGvLn53VBuAaXkLfjnbTg97fjdilw4kzch0kRi3xpvN+zd0XQ+
/BooFxP/+3BycSfbmtrei0a3otMK11IXhWMdgtkQ0kUpVJtQHfLDBRKFhJ2svXDC
RRXcnjmeYJLesph33M4GEUkSIg7zc0wUet353lQ5xCuKXmEWdAJOTgaHqHj3VtvZ
LSdORCfMy+BQmXtezmol8OoKz+BE6ARnBV5zQhbgPwkhdj3w/jWf7KLNdfDL+VFT
lAERfBl2w2Lrj865HI4eZNsLp9SaRvsFGDa/3viiMGi07ahAbJKMwYhHhA4A/1Lx
Or2qqrjn/xwt0cZvguVrB452fggAVb2kQTgy9EBHdpJgwNqPVd5gecfXiYhGXxij
yqGPHyJogvJ07PIP6/hrk9xEoMaAvjwypHFOMLqHjm5dBaWFVCnAGE/P30HZIPtC
rfS5H0kSgGLEq7D2w8z4+6rOBMpOG3VxnhDRKZsHiEvRZE2eEqJUOkslZW2WK6sn
MULyShRU8FZ4HthDOTWFIyZ8LAmmw+xbMc4l/xolMr0kL0eCC0Zjrocy/oL0+Yp9
hBsF5Pq0Im2Uf710r1ogEKSwr5qNxTkoIAW0s1H+Cuvvu1SsX1l1c8qMWsRXo922
LaUBueK8qNEBGw6uu1/2oMzM5amFTHDdwFi/KYRpBl/Z4lfwcEnnlBvFS5XHUGgK
soUTIGqVSjpbV2elk3RD7gE8zRho+I91zDIFedYf58eb1lEyqMx9Qznkb6Yn9JAD
4ozoJN1hFLXFe2odM6jVE6rJ2sjFpHjJr3m1xNg5U/yKJY/LftZqWwc4rxsVTsrL
LPxU8rDFmnjgwqwXbNT9Gu6N1cgNc4ZyOUE+RkfMN9et+TeitVQAAmrqaegRe2Yi
qNomwsIxpsnkvlQ8MfaX2GqlnkJc3Lz7SX6wY9hJo2nEUjwXVLehPKgEa36NrEYl
SCWDm5SMvTMxpLJh57eoaL1BiCkrHyC1YSrFh9w9XRCmoWmCHc6EKT15197TYfye
lDoSOdMUd8vmkb+hpmLXQciv4s5j7zTUovnq5w+KHkoi87JayPyCsFQi6p4Pi/rP
VPbix3TJZf6LwG8crZWn8DmclrghOVsCI4jBkBO8iM2oViwTbr0OhyK7giH4ymKi
1WQDyp0p5yPrLLhq81LwheBEmJeOyW842HWr029cDR5mtBXyo4LtTGw4oIf+ZFNn
7Rj3oo8WIfVcutPzmG+VuQZtyiDqC9ssczjmwd9rfkj7VGm7A+AdobRSx5E4UnHr
mRALLzBKOG6hUxkp3bpY30ZoZG0oIKf20zvlZbAiD8fNmWx1p2dmS1f/XV42vyBH
XMuqiaimQCVm/Q2OKkQBuWDJVGr0mPmMWWAvCEAkVxW6bMMyLn+/7POEKv43mYp1
paoRPn2liqetfMbwURQrpznhZwe+XVHybahyqfDDfG/9GDUn8mbpyYhhMKZ5F4JH
BQDC/dk4FQlmlN2aG+EllYr+/kH+25XcByrWV/Vh0GIGBHzBEA73ZoMU2DT/XYa3
cn1OO98ERBlnUDvHVqZW3x28K78T3eDB4A40fI9a8LsGQ96le69H8eegeifmXTFn
5q4lcc0g4AuI/Yw3plh1lnNsFQUnCr7xolbC+D+akQnncdq2dlwNuHx/AC+2dGMl
uGxRtbGPqzCbmVBHIIvDRkQaj6s1oTAgDD45mxhiBFhTSgECr8KE1BGVdMo34Uq+
gTxWc7EWfZvtdoC/Qce+jIL6mCrsFfK1c1CmIoOMy8kHeHqUMzTpFbFwTAmG0fqH
BWeMGBw7ve9rigee6DWHcYnkzxupH9TY/86Zadbd2BDZD0VOR0W/HU9NuCwxxhfX
8DVpsWFkPHOFZTdutYgI4AW8U5KVq/OfgHu0lWbOWvXgZVWs1T75j5ZdPfVoAV4r
FNQ4hKBJWo9MqGhl6U6G7P0sYAjk/iKDJdTpNvqyaaWgKcKWqdEkW/EoriVxxNRK
b9J48tGC0fvcbXIb0tYPRMkcMPT+2xSc2xVyk+l65tUvXGTtw4yNZe/nn7DbmcM/
zkP9vy+91plZfoVCRYr2K5vlg3ya1zEr17mF+2KfylHB03CkO5kJdziRr3RmKyX8
+doX4UfdvKb9MnDYOJtHoIOo/P7oyYp3irIWQ9iEIWrMayBT6w3RGe1irhh8OTKY
WWrfncsjGG2Srub+unQUolF5UfyGrpTyYeHp3qGJNXBetGRfbG2CDTCrX219J+x7
1vFJIIv/35vO3g8kBgcwbqRhUNMR6znptshu8cZvDJB6Yh3mdBLdnFJ4+EbHyF8Z
F9+fKEpot174738ZmdQUhoFgERH22uE8HAslKHLHe6cB1RH5bQc4JPRZ5P5tGeO1
efNdE9M6yz6wsTDxL78RCWImdGEo1nBuf8u2JZGR/LTt6AplZyq/8TOFIXjskb1Q
zGrj1lhIwDoi3l6jKAWkXhujCDQb06IOKJ+VYcNjTzdsz3bXot3BW3nuW/u5VJbt
W3zHIXLriJnZDt/S3P3T7THaX9CmUuzLvaAGMaRJZZhwH7xKhKEOV8UK0yV2YQX6
nprMDxKuddsk7hqF1XLAlJ3H4yoNan+NQid+1eN/dKvpZJPVmqXiTuC1s8k7aP4O
kx58Qgx/gZzh/KeMJ672E0JtlkZlwUHfsSuK00oQQavgkL28S2v0+UcNkYbMaHi/
MZVYZoiliQ1cWy3gHsm2g74ptbssXB5lzVV50liagvd+vws0AghonfSBndGuDkK4
EbN5rxBNAoixNzUGTcI/8XXRzgtGTZQhmgOVgsoTocvjP3xOc+1+FyfkM3TpekKx
5oKrInawAFgOPrYMlN7xOHEhmY8lTD7DcIq4Xm6LJj/kKwJIyZBlF2tqOGNg85am
ArSFBcol7UE7y86ABBiBJEWHlcDdiUdvuRkVmb8xZzJTi/jtvqwAHNdC9L9w1nSo
N9IW81Jm9QMqJwpQvQbspsvys7hABKZhuzC71jyLnEvT0D3jz8WToiy78vYtf2et
6Cy1GsCzKUSPhZ6CMOAfRRAluO7cW6KQeiEwYX7QvLyboDJcu0dmgQFRTI7AaVEF
x9L+0OXzgSTPnWNkk8yEF9caGk7UvUozxFttVc9pHgDqQo06voNph2SOJhneBNNl
cBX2T6Njgo1+5ZJfUYkJqxKX4Z/E1BnCKX3LVAR4IxrP1tjeTCLz3UuIMx3K4Iby
jZZVqcj86mPzAHZ0Jjee80oCZenmYsSgcV69dsMCQlGUahtpT+LHZuc79YUaLwzw
udTDmXyzg8uc9hLVOPTVHCbS1azoZgKKnBa2MVoO/glfC/vEvY4WQHgk6dZYiijl
tchmdzQBp4w4RW4AhbEhJA60T1OcvMV5mZHQU75r4JRmtMu7X0NXg3lFr0s3flXU
5PSD4OqzqR+vb205wNYFsS0GvOWK10GYrsWIx5pgkV6nSczNT2fuPCO1uOLR/5Gg
3QECNuznBDn6RtGw1eDjBLsumFvrm9ShYWyL89zs0RiJekIA2sId6F5t0328vqFY
qryx+Z+auSF20lwlpauh6Aat9SUNfXO+sW3hGdzGS9IfdmvmXp9zJMv1XMHnPPmC
QLOnv5Mi7P3f07mv02Ca1N2Seti3EUwrO4rijZbRJRyoQVp7NhzhqUp9qmfYzgcC
zX2uTq9bMSZm+6qGghErkxd0A092xxg1fqAtQow5AXn6KiYBSZ2qBDSUZLENNltt
/5hs0bNfEacLz6EzWnYuhkCz+kdsYeaUsJnQ/ltNMKV5610t1rhaquqy1FvFkREV
DHqQU62sk1XCUrCwCr5nC65Fc+KwnQvpQZtzQwe/0y8DpzAYwm7LluuiSUotkNBE
trmfpn9vVERGJwX6rtdXYfO3MlocCaSZfjk6GQOuHxIbbc6x5LjZ61Ny9qgGrP0M
0XjZRvfuY6Jk/P7gzt0kBUv95Ojf46lkto20zQX14vmH77rri1SVXR9hdP+NC14C
anOyij6h4VVPm1EzD1lNh7VHxY+7sTBsO4ZoHyrvOMhbwDxPW4lNDUUXgCtsVnVI
EtYPkPYzguaS64qMW8u4/M2vmbiZejWkL2a4omPALOlxmE9oJaTOW3hPf0z9c+li
TnWEU/8m++xedI0ndX7OwQ4j/7xh411Vawyfq9QA2HrAhmL5I38n0J/KmTRtIkDD
5p+NEdzBOg5Hrd0Y4iO8ewbnZPqy+FmI+zBFtHDe+TTL//03VYKmu/gXFc/Sx/1V
oXytbdhj7NC9B8CxgE4BsoPuwKq5K4tpOAe47WZKrYCzLZ+cFJK4jqUWg7L1qy1C
37PPzRHbevU3JNLbOFYNEsrQd5wcjL0S3orMEYzeJCExjAe+n0SDZEPfgpSJiaax
nKjpucx1hgqMlg708h4fNsLU9ePI4ZO69EC/ixHYiY+dCMF0hDtCqNpvB9/sOxWT
KmrNAbIMPWOMlfZIvuU3EVPgu9Wba40hXuTfzWEUHyv9dpkfOWFoatVL4nQ3IZUv
gc5K1Kd3wFf2ki2cGpVdLmT/TZ5z9g70wMMvowFVMvcGnJJ5HnyZwMUq0N4TLvI5
7jGw/DGb0eL51r6HvqZ+RmrD9LlqIGkxKsbjZvw4AYHwfi2gefd+XL+yb/wTbFXW
47NjRTNLRBVSpx3vPCGxcdWs8XMeS59tu6o9zhYbDANeT7nfjbXl3k8A55ftwEs5
bUh2J00ve4+TZpeGWes5D2MmV1ny5JW5nqU5wVbhW0qyPIx5AGgkObSNao2zywsP
q6sPMWvAnCr0DUuwcua4ILuGsyI5Y1+cvwaqyMMRmHFSeI0RtJOiw1VdLpLIYRWJ
dPlbLUg1aDmvLZu7RhWmjTwqfTmcs46j8dDDR81rlpyGubaRc5sD0YUlvr6qVUBg
c17V33QF3rYra7NCPlhuV1MaOuR1dzOZf5o+NkuyZwqVFCNr+cHDtbPiQTc4hwJH
PenAg1cJl7OTYLwTQjN+DZES7LBOqfU8D9gWVhmZXbTH1v87AHolDVc2A1RyfBXz
IcGC1WT4Cwnn2OwbnlfOvtMZWlgiSJUxP7O6Wax3yNvApMSZThCw9oucKwIZFiZz
dnuJDRpkeEJzwOHkOw+qCWEOu3+wjhRziuubrIK+e0q2paxeE5T15cTI7fHVKz1S
fm2s7MDjx+sFNQqi3m+IMMUvKyFghe75l2UxLBJCGBRna4IfBqytgyCzBxJRT/xj
U5vkAugyk9nwHaJe2sM1zbxA87ZEC/eahXW8LIu/Lh3JfCe4+k0z4R4J8GSBgZGP
5GZqcxH0ytwhU6w599+rG4FOzI8wnJy4gEshGVnZytORoSM33tCzK67Ou/TlghaY
eEtH3OUqoOI8yCSv+OkyJab/lQsWoYPtWwDNb2gHYLJRegjJRBCrb/ddBxqAZkZi
cvhPgA1s25vpRTU6DiM5qfNbiY9B3AmHr8gVVUN5VkEgJvoOSQfZQIdH60Mae9D9
YOYjA0EMkJOQNsLXSKCs+z8Fxm77sS8TLdobV+rO+HrMflMhMLXDiY9GMoKsimvi
aHVcD5jAaPZIIcYHreWRBrTNm3fFxwI3dSYbBpr5pDfyd4EGa0vWeTFyQOcPlt7r
SY+XBfN73azrg1JuMXTzR0j4A8v9BkPbBxZuAU4uL8VMzCMWtgbO6qHRA46BFqwI
oa5Ott8pwfplmEPGdutYiGrZ2aJp8zwA5Qd6pShgN8NFEu7QN7keF8ME1xSqVahB
YwMy06Gqh/5qYKyL8FMCzsPBnPfk9e7FSMbv7U0E/PaCZehk2dygKnlYY2w8i8xI
7j1+I6mDxncEWUwzo/521N7E35Qd3xc0++byc5sYjuZmVArnrqPW1NQKj3I80U/D
tNHAX61KxbNQAR1Tv8R1bd/NdSVKPVQIYsZNeDMHab59hv565Xzc63bdeQxFQSt4
r6dzq4j6lcoQDrTjMQTZlfUJamNMmCy1z8x+lin1jhtLUvJPQ5p/7Wvv1ChkXrU/
W7dYn7Dwu3bYElSDwDg4wX+urNj8Og4I7cWm4WDhZJt4+1jlqoeF5XNgGr8EJZos
1DPSbwlMUgYIutxcvtS6MF8YJpIfqJLiKCC/CIBNKdDXOLpLP4Uw+HMJVbwTqpxr
NCKz3tB1Z4iGnVPoqYInDW5wqfhJIgvUPNVH/bU87xv9Lw5cDDna0pAH/xVBu4I6
bqErqqXrRB9HVpuZk0Sa20CjaGjTj47Gxfiea9K+/C0ChYwvbvnxEpHkejBq7sem
q/qYvJg54xdNwafD5E6Y3OK/LySafbckDU0qasqyx6mKCL+oMebn/cyogqlS2Q5d
1eU6WqkFj7uRVk2QR0ydSpGJZEuoodVje0nJRV8siD5+/OXxYXkrbDYWca/rY+am
z32/eXlyRDBCqikvR79pZlq2h5Xq49DhYfsFH1T8b/7BQwvENLJRi0RfbwhfOTUS
CPcHA7tYcx7gIV0ZaeF3edu68bMqRQ0ZgAvWbCPDQmwSN9ZCjkPJCFV7q8v6Vbmt
WIUUCipk/7MhcOM5LmOreQ7hThbLp9i8isL9LSPcz6111MkC7/O0x6hkq1Qq3d9a
Jh284szki9He7tcbmxNeVyPwHgNoHunmnAFuLdht45heQyRBFYSj0IekovqrAbpR
myXWFPNTmXjnRi9vfeFUo/7AWwTi17Du98FwEePxmjtMl7n/5jA5vmQ6ymwzqO+x
aLBxhpS8QwPVF9nXKXjWbwmITPKt7F4FBPAFCtOGmGEiwS645ll/Issrr2oz1LGi
IOxP55wmt5qVfISe7piErTzuKV7anOIl5enwUY18qFg/iCg5X7M60rw5/9j7pX8H
3Epf8EGwGX1UKJsjWRQDoI6UkIcR4gmgPlaTIqO52V+XrNSnQVVVMn3pFlX5NwmM
3GJ/opYFkwlMZXH55cpVaRwykp9qU7ubPSVq7O/0HIpqswjbvLeW4iW0YTbGmpdA
U1FZ186flQI5OCbkHUJuKyZx4ZdJRcd1O5ldQtbFKl3q6P3rR9NQqmGIuZgvbUfb
WRSS8zjMQNeQr/Z7Mn3x/fmU+AjWt8x+bMGNg9ZjCy2OLyBWzhEUhLnf+uOKgw18
ND/UE3YIFNtflfX1tTfAKHsiNYtIrd9oqKSTpakw5PAYUScXnFgyGECVnPQMlJQg
KHX9Dj2glP0uXIgPktJxjTb9mFhF2EWqIwNaBbg2EeNc8w+Qaf4aEQllsfhG0md9
MYj+Lxrte+CBLeSPJIiyeG6Uq36FmFGxaOoQ8Sf79smMDo2/uH2Tk20abREMJSVh
WiPS1e2XMX53jqJHpoZfnBrQEBv2ZV4/n3FP4FVfMtWWC/Gc8Y+rCfVa5ZNHxmlr
MZq8+xFq616dqPm7mcn6zDoXyI3LPRdE2zjJ4wkv6C+SZ/cxdEJOzeDftEN6BAWo
Pe0F/05EJp4kr/t533UyC3iWuznBnHaj08b56QQP4X3fPlGnLlqvAJ3hZ9T6qro1
8ZgnWvm7+W7UCvHjSkvs7KnvcjUtRQlcu1RQWngsmCuxyVaKMQ2SlGqrNejOS4JL
aaX1xCT1DBj4OYIHF0HAnfB+T8b5tvi5r480jqQPNLM4nWMS9HYGvNhP8eCmhoS0
RsoWO28HIzvhO6eiEA/yRg2Rn4h4gbSeRjQ6qNuAKX046bXap6JkNidsMxKx7PUs
vagZn1qrGUv+J8puMd1lHJb97dAA3SzZAp3MP5Mip4mygwXxh8xdLUcTWMmARMBH
e4o5YEpM096Ik6IzCs7nztm9EGSFUsnSUXkG8ocoVNhIuHPBy+qW2B0o3yHyZ2MX
lKMqKtLK1Ty9CwfnGNM1es7verfJtsurvPA3ZgahLI4x/25N6SmR+LDYNUZexLXR
GPQEdJXmjgDEqwkEL7rBV3PPA2Cgb35mv4IwSUX9SNZ5GqQw09jry+NJ3eWmqadX
jI5p5v+y7A4LDXKtMqQHpvtYEVwBRf3mi1G7miIMpkvXvaV0d7tcjWby1KxzswC0
S16jRe5j/tDqtt/zS/8YvkppQrsEYtvhVI6O6PGYbEHTVoYa5/fIsPTBTbt4jPbx
EEpK2+z3veBuROl5iXUgj4LZUBiQwrrsV5dkxIk2mkQswqILnBVj8K5tB/Z7ksGl
2uRCo4/iF11RaRgpiPB5cKNum9UKPIbb1TPJPCxRG/uvgBKZTJr8bFuACa2xTO/J
qZkz70US7ub8haqAMB8tLPbWOBPmAAdA/VT6s6IgwyT+VPFcC6iNkZ7NvVX5m6B4
hLkVhVfNk6bzbqQWJTlVRUoxKAF2nz/OIv+I0e4B+SeopFHnr+hjNTfpXVGvXw+K
HGC8Qijc9Atd4aUo4tHOql72IX34uVdkCTmx+1pauEdlnmZNJHR6hPbOWBIXLZdj
2fb/2cbUYD+122llqJYB+jucU/QolfmT3BBK/ek0KQIzdd9cTI30HiJMF+TAv2Nc
rboqR1Ct9SwkruyCHhn26SzFwt28S9sr694Z9hDPEWRnun+06E0DcZZx6FMA6qyQ
q5OAXGi+cM+wgCytSTHLeetQOUILDxRvc9RCDtKeOBCSmw1FH4ANHVUCbV2ACKhX
AADBj4QnwioHu4UnMbxzLnjIDRXBFy02awwzUp/aF7+VA8qhVpfWLAPGvRTVYUnn
I4bWW5H+yQeOEW+B5X7Y5YrQKYgt/e2E7CruOm9zBdcpimz6Jdq8S0aGi8oIVoOr
o9S+k+tJbbKnLXI/INFY/BFSD+OtS4n2LfXw5Mw8vAPzjXZ74A6/sWOTmw0rtjva
tPBxdh4Oa4ZnyGx1mZv/JxMFsyFacnxWnSZiYwB+NqxUZn0sEEu/6IB8VRNGNflg
ytgXV6v3M6rFc7iMSsbfyumBsaompl+GLY8eGiOr9Ba9jR23Afd0WfiFhhxx2x7a
decV3vcjv3s1ew4RXEJOsYcoPHgif/S5w+YeDREcRASRk7/X9dQkLuzh8104aDzM
91VQY1L6+p6EePRBbL68GX6W5PL9ZtAB/5bjiyGy+iRzcL31vvx5EfPTBaB7bBUI
xkNLi9ZCA2U8iH+zdlULaikP7N3TXaEIuhC/Ju7A7PHwxh3+h6R1rqC48rzwpJ4C
7A/haR2XIAKMRzF+XoBwUux/85vNIzRz9bryTFq22slHjuE+tu8vCVwyMH0RDFpJ
uWYzfhpdpd5TTZQS2HvRCOT5BaWKbWr8j0mPCP9MLuqzUlhvnKo5iNoRkP+pj0oJ
wnlK6j4h+e3Aap6b60o8emZ56qBBB6GNt+tAdCK3ISKGf/o3mh/kNp179eA/evNm
lvBSBSTqcsdxMGjzN9wM7nQxB9Sbs+cS94zlwwD3DAvkfoYAn93DWzOOXBiNHXiZ
OkxYbSDf0DDgLmYnBVRlHw+DcMPVX23uKpiPRGA5wX+f8rVaCxEwC98DuaF+/gbQ
R8kNgMwfmMrrJErjS9w17uZ2cSpp2GvR9c0Y0doXDqr5SdGA2wLZwYonuGwp379v
z3JhUc7K73XslTx6frc+abVGvOgWW0dSCl7Sr3z9c4VJDSb+i1G7eEWReUGrd5Ia
Q4XG3YTpBW2dcKXzId57IotMYJyJ+0I8I6DWhwq56gK/J7Nb9z/Uu1r+nXZC/YmE
Dnd9nUzaxY8vIbwQYv9iCOo8IxJuJZSApz1jbZJEheyxbOH04VLsvsEa8WH9nVDj
pTAmCCkHq5iOOiKLsybfCz04wIvyuzr0aYLCqHJKVH+yWjLTjBjpDCTWN++pD1SU
GRs0Zz2Un/rBEtzxgFDZJFwKW/Sh6bzb4EmfxKdip5KYbuS8YsToCqd/aA6L7x5e
m5Lqo7W2PPZDuoGUtL0gBfktixfEA2p5emcwbOrSwOc7ilHo3kn1BhGws3ayaDGM
vIi5fKTdA3kNRZqNeEd2UJCz9O2SlWEPdSZz/MvHHvRKLhPxYUi3U+ey9DZUtnpx
2ganJuaf7F6+AFMBXCv9DDBLS1lZGAViqHawga99OyB7ot/TPPfO+Z817g//DoRC
X2I20pceZ3cxcAEPguYrj9j7NfI7dS2hjJoq2BPPsbERWlOXNTR5ROeVK9M3kWuG
ajAt6YuyQU2OHLwFg0meQKQ9ejj2MGu6Hag0yYMQ9FVpBdZwq6pZ+xhxNl+T28Cs
CbTJ+AFMPdHiDB61p2szu6De7qCaU2c2Bm1f7K2dAV376KVoatw3sb5407x7PEpA
uJVSGpC0/IA/RE8VnNJqjX7O2QA8G1Z+bAOpEUyo6NLm+ZezjCLA9wYaT+tn+H4e
e/D0AMFX4FzAhkJ4E4Ny5kQuNqgvTqeTBAfwTqOk9Oq6GyBhKUo+F5EeWu4pue+O
ccuaUWbZQoVIhIKTzX9VNqdDRoFpNOnvo9pCMnxLRkxAhpxtEP9M0RwYR4KVGil4
i437oQ/ESkymiYRXaP35ypnccw/+wTcci5/xbWwa1/vcTQlFlF6ND46wFXa/slXd
OYQLE2EHnU2dPQLrYQkqeF0QFhIP5Lw3nme3Nc4vBHgQYv0DFdwZ40Alkg5ogidn
0DSBTBQUJe9kkefohRW2sBjozAXlzUVhDJDJ+egJWgbgQPdJOfOXfD+ZlwDQvH3p
w62OeIcj/Y2mu8OljMQ/bPHUNdrI3iQ98tVx0IrLL1VkRVQIEgbmjnTVFr0Mn2s0
TYUr4o4u8J6mnlRAe2zAVu2AQGynvOUd6TTmdENLxDFi38RzYcvaVb97Nr4KwrO6
nCJ+VgeBwhZehx2C0uqyyAFP5sLmaXEAzfFSMeXBm4TRmjzPpgVOxzYem/28TeuY
bADGoO1yxu2pjn6p9cAigU+0Vq5GMH+Krt2MK0yp5VIYklDxADngR8DcSCykUBC9
grecpfBOg20U3w5y70CbHaNr1VYi/soNxGnD+uXtUEKj90rKQsaIchQVWuSG3B0P
QGPWghHV9OFqJ4ijKq/olMkraT1GLm5qPF3XU2KNVUjwm9GGyMVVq1h0vi6cy5Hd
XrK9k3ktqJ1luOwoFKDah9TctzLNYXx6WajK6Q1HfJJ04Gt6RFHDq6eiAYxc3cYs
2AbjzgpXKFO1LiiXY+CPQL5e4pdKuuB2Eq8ahvhpDO/hJlSa4PoZ1opUuuXbned/
wDwcPh7h2pyOVngfHia1pgI+4t30JKLwsjBsNnZE5N9Yqh5JkekxXczX580oX73I
6Iv9ldO3zolDu7m7Vn9A1CzPmalnLV7daUAn5zkCPqyuMUF3/M5kqi8ZKLc76Ge+
ArJ5Hy2px55g0epHu1dzaDlj26JqIh2YioFGi34n+gEdNdwyCu1gwgPPEMZggi9H
KX6NIlvLtJYNfUQVcY2L4XFe8e2LJyYlzWD0yQzLxxHQTBATNKP92FP3IvXpb77h
Kfl40Gc6sP29WPmG2q0n2dt9RiBH60tnDRjfiOVfTprZE8nN6qv4y4JCooziMFCU
Vqn6WezhxREjhqiN0cPZ9+B4rvNx/yG3jGC35LhbztmldYj+OvzrZwc+ynENKXKD
6+yaP+HNUdnT4we2s/P2W1Y8xsRAQGw1xiuNW5DwcdN+VjdjeiWEUZohYQfUqMAr
5S7kL094wdq5u95DO507gsUPwYUa44X7prHX433XhmA1CrGBpAWXjxfWD1Tz6yeb
BwpnXH4nqvz94kitn+r3HMDT/nCy8TFyd912MjqhFJfrsKLxQyoWd3HP+n/3PQA0
L9I+V/q1RwtFI9bfbGPSwajnPO4jHZMaq+gHfvOKuEJShkAfFaqVuNj4j68V3KQg
0/JfF2b0Du7CmaNvUa/XtQOiZ2IpP5a1Ettga9JKluv5sMfhQu/q8mwtZF2d2k22
YkIbn/3Hxan9TDa1Fiz4OKV6ek1g6gwbsqS4Mybkd/c/Sn24lqPhWjOebnEMG3Q9
Ec4ybD//BW1CAgQ6wcFBPINsXUxL7eBrniownZsWeu/JLc3dImtR4sH+6R62y1IQ
g5G1/eaHit5IocB06rf5e1ldNNAEkvef8epG0tUlacMkIDfJK5FSgn1iuUUs+Jbd
NT/TeOAsbRD0g62j/ugh8U0ZB9/xm/fj6BABUSkjB5rnO8Q+tdI11GSQIJr3Puaw
u+4ykbXg5LFF3x/WLQ1q/ejmPovOccJBTmpYRQdejFR6D0kFKf9VABcHPIneVhfz
ks3/UPIlJGfZsmlNCMVPNrF1ZGrbXZa/z+oVa/W87JYRBfyfk2WkTj0/R02AlOex
H2RcGAmZncWV2nwxGJZTpJ6Dk5HOgAAudQ6QPbeLFRWVx4saO56heWdeZKKZIT6B
veP1tcrXEKVPWJhsiNLOU5xHcFRy7we5nLWzhe6RAON+NDASNGWToWY4IN+t4baN
9E6I6o+V2Ym5Pkqnx6D4tYp7klDs4G8Qg0cpfpXeV52ToCrPV9UwJy4pPf6cb0hU
PKaeD3Boens5Y0WOK+tXDKGB6XKdk6tS6Rj2ApoLE4MTSwdML57VEFX1IDCMLAX7
D12N8EY6DgBBn4TCDiWS26bjyFmxrM9GRV2bBXBvtdbo0WnW0a2LaRty22tlkbW0
QupKv9FobMVGKRnc3Zouj4f8tlPfNo00lRqbJSBH8RVkzeFw6GwTMqzQ51oo8dNJ
WL5q1DWQTJ20aUobkpQEkRP7jyaQBLkDR4nAMUeh0Q0SzSBV5FAzIXsSebFCQwHY
B2N+62CNPD4kckMUo+GmZdJK1VFGNtR43ODLHP5ctxX9MF6BX6aPtpQDvb+aFO05
qTRaPXRKtWfto6E6PAsxROzgPQEDW5m6S5ls+ItOXBvbWL9WHAT7g+uJv15BHrFi
MQjypO982kiwpIWVXZbky9wVcyEE9UD9ef6tyBkjoOtVtH4v9FCtLIeJ0H7uhJuc
Lcb+c+JlqikdlTzosi/gz11j4g4SMNUCZe+o/s5rnOL9SH47FcgToI57wViNxvlb
wo494uE2+7o2bAHgS6saofCiOOmL/kDy4UnO8wajAYXg5Z/uOdRehuQBOThSqZba
W/MlWLC2cVi+SXdrAbUurXs6DvbI/XKk7TQUQ8c1G/em3qWNuv4Vyw5/QOuNgNSB
L0AcrNy9z9eN+KnlMR2iJJWPpCtFP2FHqzUxCiJUDGwo558C9Lkp6D1cx4cmosyX
JRmLUQ/TDXt96o53x30RlN1U2wSrmQnyMh9b7kGledk12Mvuydyxn0I9EBpuAUxV
mRe7QzcwgnYhvWgWlqnL7pewbod67bsXqyEJBP4INUq5CBl5pjapfkQGK5lLkV80
9M/fLGDs1Hu7OO60dOilPOsRC2/ic00Prv7z9FkBVMq0+LHwQi5udjpHCEvi57bS
Am0G+g7kJDmL0l5itTQrhAZv3o7uIjWq+ARP9T9Vi43bg6X4er/sAHRZ1b2mIXf4
NV63x1r5y0Fb4GuTJmJuHkuNsUlQ6o5q13PeHGbl+xECxtz1LRsAqoBJND5Ercs7
GiLe2hbU0ybHbG37Un05vnffWVsROZ1cEJRYTTWEwt0MscGw0fgu7azqCWqhnl2M
RlI+GnVbvrYkZoSmq6nVBehbFUeDIh0uKASx5NOefvrhrXRQ8AMzoyWIRrjnQtdl
lOja0gUaY8c63GUgNJG/IOggG9Qc92NiRyC3QJOB6jf0JyC0iw/SonfPvCALW6dQ
+LVOVcT2b1q1ODQl5g5gkoX9PALMyRRRbGJ/iIxJhJoCF8GZtnhbBhxuoiZcN9Vk
Q5x3EJk2oJB61b8SEuhiN3Xm3oclalrskn/eMu2L7R16JJQe90lz0GBpWYVLpAy5
84d4SLTs/RUpjtlTkRb9Qf1dDpbdeUTzjioEtFyH6bqzw9180vbF4n0tOHJGigii
sv8P6z+Dx/Yrl/Q3BXOGgPLQFW1EtUMXHMUxPN8ZGzhCp4ysd0+16Oc/CAhlKX3v
3UXADZzCWXcoY2e5BJ9uT/IJK78f820jKYN40yIpbwzgW1OqIe++HnONw6pwfPvn
t5XOcWUTYTSj0cwbV0tqhtfKGyXrKMh/K8kwq6ZGxFf70nNEsLXKMef6iTIkWTd3
4sW8aMpw0ry9yScLykAGAjhAgO9OIzfPB6L2RMvUdvcCINPor8YoA3VTWY3Og0Sy
KUFrvGHQiaR7NX/bcy1VBibBaShhJp+ymM0mTIwYpRGOMTcEXPzra7v47X8d/WvO
YUk24mXhGQY0TwDObX/LSvcknhfc4FPVoWTvZseQGd4RTe+KVm1aMiMpeWYewd+P
LbDeosp1Q6TRrDh2cshdZvZCT4y7thkQkqSLi8XXbBdrhStBEAn71eLNZBcoeKiV
rb9HZT2yZkSrNO8nsSAfsQCPdAQcEpRvd7ZFtlsyY8HBMG13E+9JOKakztnjcIDF
darCQSoJ5omoTtHfu6EDqNHAwqxbCA1Sp7FFOTkx8VJZUWtG1FLOC4oWkDxnTg+n
LC6i9t6qpcB31VaNiUzudowGgJEPX2lZx2vS7bIKdbOJ1KybowzCHWqWAtLE/s2H
FhbViBcyw/TQBQ8NfNgi7StoIv66NeVkm5swalywN8UbpHdpJ+uY7E7HbFHiw50Z
2WAezAoNC/7xH7HvTVey8b66D7vzdkXyt7xH77UTf8zwMuGobk06g1gv8Dx5d22h
058tXEy5vHcMLMT3Nz3n61E0xbqZPlJjYD8Amcipf1Draq4J9ph1lUtOCvtvLx9E
3lQ6EI01le+LocVQfN559PEjQrnG3A4vtE6eBPwJdnvMez0lp8tyZMzww03bYBtJ
DMmwdw8DWn1hYd6RZ6CQ3m5bQLnIKoBUboYg8U6SZjE/1Z0OAHt4MGx2uXOmA2Pm
qrjl3/RCwdWhm5OnbXmKO4lhQK/yFNuFsnVDg4sKbcozXdtz5KdrWh2RJN8rOmLT
nM54CBSV066yDLYqj3gkgTTG3CBwk2wnIxXzJCWUWdaESJ3FtJUxytHx3bt4qk8x
EP7NN4tGOyHtgsp5XDVvSYZRMfvCHzr2IN3C6N73j52is2E1klWgz1bqqkoglMyw
4mVCIzAOmyDXSBwcgwr8x08F9+OiTRSZUeFdxSowktgXrqLVyVn6Sb6ZLsrrDMCo
lwZXISFa5QzlqpB6FTe9PmjjWb8DdQxmN9f6Yaxy+Q25N15pBhJGIojKrdnWaT7k
9Ii62nNq3AU6vGG64r8CQFYkA/JULszq6gZE27pryrdsvhxkvDLpF3Sl/ou47qFi
GEFG/Ny6i4xnjtCHwX0gRFlmNc6hc85wHYHfxmMUUQxT4AsWOIfAPKOycT8OH5r4
ZNXIfzoz1vZ/+hEjrRkroKMWMH1Plvv2G9i+U134urS8IRIi/MZorv5HA6+WyP9m
oRmiuFQURD+QeYRwssqrkaxKdUNCYc6/I2gkfMFn3q/BcVVGQZtoVAPqb3gm+zuJ
GD212fgeBuq2MaYAWw/jgTjaCdoT36TX3QRUJH1eNhdKkQsTkCuu+bhgmHkiFKRz
ZT2oo87k5KQ/+xbRxGQ/RqQzT7Y8h3OLjNzle/QTCEDKQAiB0oDWQw0r6gcxqrVD
FVB5yHlPxSY2GhlV/SHnSUvE42lyo89hfWRjyJFs9su4B0V4MGm0kgf/D5nmuMPW
idX9KNujbhn8uXslb6CW32v1eOtMf8dSw+tdeoR4gVnyyznT8BdAv0CHIaX1rZDx
qPT564lBHfXg4yXePpHjYEUqoNvHR4iDFrz47aE2SlPpZkxGnmhggZfqdJ0BqRvk
SeI/cNXronOTBWfuocdJuHjx6+b/wN3FZqbqP96Sa6hNKWJAZfNIiOdn2Osj2xNo
kHRUQ+IkqFd7Nmf8yqtY+1rLlTTAKRy/GqVaHEC6AWVbUHCJlkl4s9MfHMWyB254
glZoU43Wgot0CBQcUNoxhb+BuhS/n0jJ3KDVnwlOWyVLm957Xb7bLqtHKBWXcghi
7ly7lV7xYBjcwgQXf9HeLP3Qe9hu5UDkC9GGHkKUumCuQ2o4leRggV2v/HeQ+nd6
XOl9QGFH2HSjcMgxb3pURRIifZ7BNo1QfuNllYILNWHGlw0yglZm5AOZBg6LglCw
OmEzkNezSSsXlmZr2ouD8YaPKsjy8N5K0r1NZaAS9nx61COjvAH9cnjGVsjljd62
RC9D42M4/qc+wAZ8UBBMMNP3NFnZVBPlBv6nWQJC5GRuFMrqUL7YTY8S0zRbM7+x
NNpjsUjHTD6Ye1TWmifQ8KPC+du+08rYgcKzZrBazVttb4leLuWqfROjGapqR1F8
rapmWTbZMmlh0BE9eFvQyfI94mjsOTxXx3OCcOyhG7YK2zq54lzasfLK8ymmTyrG
+/ev5CWA4cmX9y6nD/R6nnSjepQFwX8zVFpiUG7mtLHv7mfoEkScJvABWTG4pNCU
pRoqTwBzQ9Z3migkp4JwFFIxhwE2bndnVo0Tyh38uFJ5/7CDP5yPykSebjF334Dl
C12wkbDohtx+UCzGX606ZDJDzH2oMIFz1+JB5v7tvsSvzrwCFaletQD7qCbLU2fJ
EPG/4lQ6KdDCJipC5M5x0bNQUKgCsy/t+8Lx8rL3wWBfA+qEVFPJNlpaiBxfOHt3
3CisS5OqquouiMOicul68w73uJEcxPrMY2Sg5ePcGj2roQxeLjMYsIsA8gV8nA45
+Op9vVKcGw7yBF+b1RiWiS5PIU8MCLd5qw2gjH7VloIc9fkTuHTPLd+hM42BtG8U
eLvZReYCUtzVZeIOY9IMg4qXKsEfLFaduYqm2h24+dKSzV7GtySla91Q3jox4uIu
F4aIqh5W9FRn2jz4u6h/kbS+onBnb5+BSAYoTyYp8nnH3wPBQajF1GMSVqmbUnUW
Wqw2iLULD0hbo1WjF6Rmrm9b/oYUrDLUH3x9BtA6W3/MY6nEO/z7t0+9bgFCqIUM
C1todCd+ouiddFeRKeRuHVy71qAvI/dCfcIo3WkGFSY+/G6ahZMDHuVRW6smp8Ug
eCOkvuCjh5J07Ktmf21wrVfqb/NkvkIaef5vOkXGW88duwrMcDByOw5uXzVtZtKQ
gCHm6sLPigP0BmyDVkYtcJM0DnV5ydkmOya5ujZtUsK1YHaToVEhf0aGfOBT6dM3
mFgEQeEPa7HYOdnrWHntOKOKk7FSfRO1bRWuCjBBVkNqrfFMQrueE9RlXd2mMq4q
N3+6PiojGslIOdDHHvT0CPVUo4z22kgpP9ql/B9v6LmkZIQ1uoPBzdwA5giyw1YY
Cq7Ko8Z+szSdpzVaEsx5DoG45Gjr5mTNcqpBUqFjToYlHlNsrUhzA6q5l+OHhwwh
4RLKNQZxijwdolaioOoFuCaoAN1JNk+vN0HBte80IYT2ceSgRRZObB0gbPKbaVdA
LlmUkvAXvGthHkkjN9FJq0LXGWrUi/2B73LcUn6tnXqLnvMaUptvTxnQxyCTfgb9
XBmh6W3VAaBHxNGfTHnUPCB0clR2lWLbpHNBfYsqHusUVIdkOpDMR5riwDOcc2vT
6iEXd/naukIydiNxCEgblrWY4HUzU2xuyj00iVp5wMZloR9bIA/KfWMyvyChGdMT
ZjVSBRRnlTJDnjSJ6QkxJG/C82tISQHXr+wrIn39xdWrZ5nJChdB6JLH3XCSFjlO
/6bLgi+TNi5T2QmqWo3J33MAAhJHVk6aNt1P+/TJx9vjbesirIyG2hyMiVi7EpDA
NllVsRe5liPLXJZ58VwST8rUEeGBuOkhDAHmBCLDa+JhSqV1apxWtqZYntkudDHs
VPTtK0Xjukeg9aCAFvNVOF8pB4KT3irAGen9xxhiboSgKQtT8mE0EI33YJCUuNk7
g9woZIIUnB1s3H+YrDw/SfF9YfiQ9tIOCqyPwliZ+G5DffTsCZAZeWBmPj2miIpG
pBjJaVY82o5YO9OvebTf4oFdfpsN4xPEHCq90AMO189kzU0NRlMkdkN1orFF+W6+
95Ac8fX4vwO6/AjpBeziRwQDeVe4jzpAMsolUlpV5OUuBQrM4N0jA94nNO62TdOY
Nb5P4FbQe/J628KrVRQ/RFhbVsbTyQS7m3PQOEFgEK6lQms5rNYKnY8EqJRYsV6S
0iYXIZr3sXHMpJehJYhnp4Sq2DqKLhG2u4FnxArAjazNwYDiSlQ9fBs/U8Ecd813
QxS1v0IRBRRzdD86hPb/HSJdzz8iw8g83PK7OvPmT+TiBWil1+lwI8wDcWnwHvZl
PK4pYOgMGe4B22oiSBLJbH3oKwrTUrv7GMB+TQR+y58mHh7/hMRBoAq3qanoEoTz
L/WHTNnjJBqnGiMTIsF7HD8n5FB9QdLyfI0eUyp9yS+ymWCUH/+vwNstoxwuPMUS
Q0V4M364tbCXaOZI4vaEFQnPZzNDV7qKLEkTMukuV1sHu+Jme48iG6Jh7NmD6WjY
2i57wk27GId8aNs14fFrG6CJGdiZJLzLzwGByASkEdKe+KY4erPAUxj6bsxBp+r0
yiw2vP/wpqSFbf4hkUwj/A8I55gJoaV5sCCluoJUq8dgvV7MWxXHukSv+GkDE386
5Pu25mL0GSra3z92kjIMHFipXzZv60WX8jfB9fPxN1HhsZU9INZHHvUJKZN/xoXg
kZtHBLwET3DAzYfe0W6vQ8qtzL5ttBArSTJEQsqYNn9h8ayyyV5bI1Ou2SoDnYQj
d5qyxFNgba83iEIlo5rdmaY22q/TB7ZcjUWORPRWG++mWEsnIxmdMa/APiKKl8+2
S6QwYoXvPd0CW1pAr6nJpXl1/uijypOQtIat1Olye/S4gsB3NSs30KVNd3QF9R0j
gRXb7ImWWWShNyh+N43B/OoITIwsSBI9tF2KdRsUpvW+O0G1GDORzNUd4fSQIfGU
9+qSm94IgTkZs2FS74lyqob6rJZ4x06rIkpWLyqdjVtie6FVgCHh6w2XrTjbLJgJ
X2o28ZJVTfe/wCMaDLw7rdqMfsaaWNre9Rp8lOWvWgY12/iNmkxZ9y2FHobBkmQ6
etJ/xxE0LT46BPp9rBhFyccopLx+RqXAyM+8DMbtxa8x9etalhvSh3HpJ4asLx2h
x08Epvzmll1f3n+0/AxdV4TzPmNpmlUh1VcZwJjTB7anUSiQIRrczl2vFuFUjkKG
57fY7mwSPOxgmX9pbewEVMPuDdOYcbvkGeSkKEDqT+QnwJ8dnRLJu4efPTAI8P4x
gtsOs4JNA7YE3PzDpRxdWi9EcDAusl6fnJn1yKC0OYTMa4li2LPbVraoJfF6AOQz
FCcxv8iGtbv8usHnLG49XEMb4dhPZ0tirKQQn0OQ59MHC9d7J33SnDJLmwDiYrWW
2Lu8Boe09TS+NMauvzz3+Gzf+AWYJNcN9bR2KZJYFD3fLj7Wx9YkqAqZVVF5kQYl
S3cd2CeM+tCV2nYktZN8VvMPyBNc2Lx9zCl3hxY/m2a8ejfqNQUBcmCHOG+AGUyV
Mp2i9FqoHgZt9pbYjUYJ0YHcdOABSLNJ03qhp7pheGOrujcVLw91ENSCedamL7Qs
+BcMl0P9UfuKrpn03UHqrvpWtmyf8naSwgRQiPC6G2FdLfQgwF02eIPUOTUT3cag
CIx10yZzj7bGk/II/3cHu1nLa1W8x2k7WTU0vR2D0NMcZI/xX/612LoRrgMLlZD1
GnfOFMcOCXRrtjoFJqsxhK7chz4zxpOWdvy325QbcJj5jvkgTR3Gw3fIVvWmrkY2
Ix95+0VEg2+/4Xx75ItMS7MHeGj2ouJz5KbJ4euHuJ4NoqmmSq9ToIOssH/F0pC/
03lGCGLab4L0OF6NCxu1PkhR1NeBVrnHkgBOXXlP1YFN4Qgfn9fKFaoR3+H4VTWn
imLqRN7b7/qoFReL4sTFKK3+l5NsGnFeEwrRAsto9Ov7VWZ8Fd6RfJytwyvjPW7o
youuwdvNXjAZkyrft7lgbOGeCZlm3aQk6/psEdeyNz3NpXyE0wR0INEv9GiaA5/K
afTpvEucWMKSgzILLt+uXnPJ/NdCy6cOPEHivTz/aWt6eXWQJHj5SNhfLMxvGXO7
yVVziU66JNSJYj2NdxIP7z2kWc5Zkb0ca+GY1N2eojNqbqzlNv3s4M0vQPHFR3ae
/Lix9H8YW6t+sobBVc+P1VQD+3hg0u6P9qNh6FNT6ltRtuiJmkoC+3z+polCmdUm
INW8he4bLl2DxJVR1bJoHSB3wm5BzhVi/bqIQ55P6EAspgGv+ItjCfpq43CmGgZ4
njCoPVWp9a8w7OyJmPELpY1OC0wUk2TP07nNnC85QZFdP6I90xefjItTAfX5DCIq
mSd1SCM0us9iLLCe0D5q8wuTeR6DGD4utkSb9PWM5WbwN/5RFpacXi72Ms2HDOu/
7J51u4jGtDx1TyuNudJUYOYo12t/Jj9Asd+qgi3ltQT7xGd9jDdMc6T6j7cBRpvw
add/8ObCIDUJ4fUhlfMmL8f3Yoskas2/XTguzmVDze5oyWXE7spowNsXynM5KyY/
FwAXTaHqQcX8sgz/hmzYN3b4wfmFF7WJLsnm/VyvexBoh9/c/kMJrlXKEjKF06tR
8Hk4cgYDon08QcE83Cf1TmjJ8yTB5xowVRc7ZzKvmLodskIbNG4Wf6LSoK6afxXu
VciFNpafTlEh8iMex6Z1dqdt+A3wNxWQCwx+Nhk2NDCvdWOjKFWl6JcYAB4fkjVH
1++5jPhKCylahdhYE7xW93DmfZQv/0/6YKDx4plRLeKtdLGR7PS0hkfhpPLoVEuF
w5PAohOoi/sG3YZEfkIvhkdVTFTIdXCDe2aZBT9vuoQIOiAJcx7e59OAIkG/mjAu
oey2GdpMOvEb4wAVD/xFsAkbfT9IVN0p3OAb0xEKQESySdpbZ4i1KwsZrm9BQHZB
WSebZGppgkbWquxyhL52AflFuDVuQUfgXKXqZJUxa+V5mLb4r6fvDjuzO8Noo2fI
z1/6QZNRG91VWazB7mAyky26PBg9FSzwUgmEGeIzZkZwgxsDV6lTjSnPO5eY6ndB
xomFhrNkcmNrhKagk2Sc7ZJ93qNz8UWDWd+WCwOTspqK0DG9jtHIXHu+pJCkc8wY
dfLY6QTgEOLZonD5etMM0C7Zu9TTRV51hL2svyyuk3s/3Drl6FDwzIwHZ7UFJ8Ws
BpQdW9lYSmQ0BB43DsfYEkxh8UjGRNF0z6PHX9PNHSqlVQIa1gUeXqY2chM4KG2g
2u7wohEHoHWgoHVJuYXNRfxCuOg9ztoru2gKGv7mBFwWX0JfdB/PzTN4ckBZtsiN
emP+ftiaa24QLk4XxHDtF9RFJYRBizkkXTq11Yhpqr2JY6SN/QVg46tEyHXKMegN
Y7JPKs/9Brf8XxwN/Ntsgwb3Y/Q2DFW4fkr6tphtVQjFBjR/8TmgT6ZEabI1PxPi
DBL5EGtZgAHJuiEZ7I0b4LYVKFtI/Cegi5NrZnksGrYlI8MAuutOmS9Mna7tAtUb
3J9nhEtyf0S5OSL/o6V4iFteC1wSKRS6ZQXnKO6N48J1A4C4QO6orkHeVN6nrokQ
anxvXYO2A1gdGniBx8stO56yTKUHYV6uwobVGavkVwM62frS1TGW8DAQx0v0LUwF
gFF0xi095bs5I9JQPL+HbkZskhiABHlqFEaYT1TUZRNy2zG9iXzAbqMK93x9rk+1
3+ZNlkzexPKR2ly8e9cEkVL+EQzThSxsLuMuLXC1XtqoSWVKgyaURS3TrN0PQO9Q
c+IPJX1jBYEVoy14xo/Bf/q6ZMf7EwyHhje0UT6YwUo36/gsK5oqzIiytp0ooEhx
mvpyokqC/SLZItvzJiGNw6QoZV26MaUeQkjnhIGCcaBv00NilPomJkHGP/5v9qZX
0cwtheMsSPHkZs2RIinfHENkIAg5CRa/y8p8PqEAw3iCQPi0XaZ5xYk1vLw5LUUX
Ab4ev8nIq4pQpk1/+Z2l9eyJLRwnJPQ+KhOghpYobZr45M6L6THck0MXlpqv4TX8
u8+tz/R063gVBv0xfYDzzY/C0SkvykrTIuYOlLBeaUHs/Nm61eaBUjiI4gD/qZfB
fY1BwdG5Y60GYRyHpJeY27iIV1uZeaZAUCB4D80TcvvvB4/gA6aBHkab+OgRTE5c
L4qAkWZonTVkXtdHi6zQvqY5eQRuj1gQcTzjwmycrzFLIp2QVQkojhUpzQOVMTSu
oIYfp7g/sc/9NKxDkwOlqe3Rc3Py5XIJgQ2deRROa+kQEaoegn+XWwlBY41ApFQG
BY0nec7PnjKXDEJWF4f3lcCkf+VROBhlSAEPp8PZ38tqpAdu5E+t/aSLKN1y9dIP
ei3QfykUC7jXVqIaZEmd76sii38x3lB+pnxTVhIn3Kd62JBFeKXQhgSPv5h29qW7
bkuus/wChg1+OR6ZQmhZuCN5/WdKAFiXfVehejdQ09gLjU/9u0TTEAgWo2OUFvOA
6nuCjQoWW8cqX37SkoOd16egOBQnVBpzn6bJCphO4S1a9fg2XvM0o0PTW4i+BXCl
WPljmIe830TlOp66Ho0raSC9BtkGTmIj4VRoXbi0u1yXC0EjydhHK2gUFbG7fWig
E3UB0dZeHlTSdYSAlzIzqEWa7pRNuWmnHUbaMAZdWd9f/jmjqfP3vB+J/+u4plY3
bOEY+focfNVtCfH9X6Mg6DzT1ZsYQ5EkhAslwwKwBhLSm09QJuDpJrmI+PiT35lk
pxNGwjDOOMt0eTQcy6NZdRI3f0XlPfn4DppiU5+hhZCvrGjDiKX4jMs+TxFn22vv
W4tNioJMOmvTnQzGnTNxyuAOm6bXrONd9RX3Ny3lywZcdAI98RbL/IQ+6c9elq43
8H/roBTKTspeC7nNzsZFxZ9eOE1XiOvBKEURTaC5T4deYml5MgirdW2e2qEDj5vY
xoeilMPLNoKuhdG5ALnZ/IHYdLFRZMb9YWJ26305GFgLVEBHpUSTOPfbPrR7TN6i
X0EM5GaN/emEfSeRCxC21ufQIiPbLxnLKhQsxXiUQJgQOCJcxhXlD8qAf0fRRTCX
MJp2+d8oSFbgsJJeSjMnQFL82/5vtxNFXEMcZfohxQv1XK/T3hzhk8I+YH4ZwBli
E1anV4kteW4RAUXvJvgVIao6RdEfsBaKwB3Ei2iKy3evnag1xDLS+3EEMfRl7vqf
DhaKPkMhrNZoNplnT4WnoU1a7xbmx9KaEZ9QrbegKRLir/YERsI/+LI4WJfqBivQ
lQAD3mdFlPqTn9mE0QG3SEeX2XEXrgEbpOKkkFH1GuFqIm4wHgFyNmkAnjtdAfF3
A5Vrzrzsf8RIDp2v1VHugddNx4Rtrq5dS0oNhTUIzf7kWJmyEsxSYNGlnhtzoUVI
S08l7MT+VwVYLfNku0EgTuIT7WEDkUfD0PtWr0DciHXR19x4KukR0W1bSY04iC/z
WQTGRWayct1NwwB7hhuLd5my/h2vPaWKYvY6gNs/LXqpQTpzMEiNdmINvNPvsQ+4
7yvrt5KOvrYh5+dg6A9pAfc4kD6yAXa0Hly5nfeUA0Uey6Su3RT3H1dffxjZELc0
22Cy9xFGdXfc0tro8RtnfGhVxdCmnUlDQEV48RzjQwlQ/roFHgDAb2XWjargeaE6
jXMOdWuPv8DzQibpEX+vUgmJi4yMIT5qx/DVQPwRCBpMDNx3Kaq82Lrfwq9WQIgN
Qm0UEGQ7W5Ouk9i3vHS+PFdIB3vhohOqBJim2SE+ILT6RMidEMMqF52u+Dmp9pX7
tWt6Bz4JmoL1hROiBgFyb71lneMa7Fy+Onnn+2ZryHHnrNTvt9y4m1vzyk7BXG0y
tPmCmvn5SqlIEycqghroad3ZS8dT4vtI+eKxSMWaosow1J2nDyLdZMz6d30WlsbI
JU3vTak0GkqC3e+gsch8I6IUOXRFXkE00lZC5NuJNPjwwktWqILpRYiDD2RekHK5
AlPg3CsfJnPrEN8p9JYt9yw/AEVivndXRGJ/8ihIWGqoCHn/EgKOa9VqkaC2loCd
F9NrLqsYZQ3SM0HvqLno8oaR4Nx9lWNyCp5tdMyIvg5g7rT3szJoKfz4wj1+inCY
+i3xa5A2x/HwVtWDIunwutZlZL2zHcNt6xYvL69oEKD1PbII3nVm7LY5wfwfcx/n
iTEUeSbrjHzRixpHit+eg1o2uYDo7NbErAPZ/AZr3wEfkbRH8YGfvcvyO7gFycgL
TOC1vPMX3Iu31tIAA/4EZamceREqvAqk8vy7Je7yx6xlrI2pkROTlmPJfLy+0THA
+yj2fa6kHZvAk5URzrpJ+KjfI6lw7N5ECd6Sv26dSclkqz9m3xdaK89gPVdtk70t
q8BiZM/BVmEC4cufR+fL5LVFxcJ1b68FIzAPas+cNByApkFOEkX8Zet8QgBXOZZj
UdyIgcZOZI6oQ69IaGPHJ8MM5o47N7ANBBJg0j/blIrCxft/EMk85qRpHjKqnBIR
y7zCVwIeQu+MmAK+BOzG69y+87LmJMxHHLhq4G7irPeQwmwO+/itLYb/Rok3x0yC
wZgbJJJF9r8sMJK6/wtbRfWYVF+d3/AcjggakLx7b8VbWssV3kbmZDf2TOAih5N/
CtJsksscyTqLFbPwYEJqTYXH1tSOJqYp2UNy7Qgmpm8MnbgEmS6zYr3KgU1XZFJp
1z9xq7tAxu+gHlXXNnGTW8lsVJcrT+H3beBWiYibZW8+5bQaAAABaY5+SIcRlhMZ
C+fG05eX2AUE/5+WQ6loRKLl7vJa/lTAxpf0bSWo8mxQoWKifcIGU8QjI57MwtYs
SeOqazY0Sn5jPjIWjgq+3yFyOyfte951QW2m28Zrmy5lwCwuG3dGcudBqHNE4Ekf
+Q4nY7cEFvbtlY60VPHL00+LCCJs8OEZ+hiWObUGlF+W0H8gwnsGkIxWywOx1VCR
rYN5ge+z0BTj23zQiJ1xz5E8gx9xPFEEM+JP0w3lO5lePNE1w2Ix6kmrIp2E9N6F
f5Q53xWqGlUh8z8G3QxednT1ydQ+xqEIheBhQrzBKf020BI9gLVMmN33GsBb2wGf
JjwnhvNMJ8quRl9R/Mc50wVczAPJJ5FLUPD+SMAlvJNFmQE8vXaZm81e0poFPQUG
sKaT2iZg1mV5m4O174+hmLd3Ed0vqD8Fv0IgpY4EFHbKtquC2Er4IRVGls+G+uw5
JxMLsZK0X0rzo90aefo8rtyLn79iD0KmsSPT19hfizV9w2zxnxhlAN4k249I5qeI
t6ce8+xDdy8fxSD8heQLXK15ywA+2ZxwITTQJwXwHtvlS/A0jNg5g99dM7o6L7z5
1XEBZUHBxoMBXM3hRfDcxyQ/lGCQecoSzREXOrU/pRQmfn2WjWC9vKw+8gXKvcmw
TKgyJkKy1+pQOAxxmNyVJN5CrkUjCZDOc/gou7V0iADaW8dsbLQfFX4q58qdlWpV
RWA17JJ6SIVu+mHjCM1UtwRgkcR5UzDCVijJ/i9A8DqRaGabyCUymrkgmf/cuWb0
hbLT3UHuz4xI9zGo1dcS3m4c0lfZHQgSjoHOP5fPQT1w7q/MfoCRNWSjF3aPt2fT
PHwC2H0cGSwS3w0DxXM5KoWxsHsSV9fYIPtP2WQWg2ycTQ2XOLwfx1cA+SRn9zMq
GVrKCQuR7uTP8tyPWDO1dm8G5irmxPurRSHxxM65mF8f7Orc0uMatuxPAsBd59IQ
Ucx8iSojee8lhvVsrd2MO08fXK4nHRHLPwhjgf4UiMk2haEHwX5LAVLXmEHklDJJ
t78B7ksgRIf1Xu+SCnvTkGqPVJjYlca9gmT28dZUVgXIZ8ZLxg3NPps+eCCSrUmQ
VDja0O+xAEVNiOSsDsTdxYmdy/3FdtUQPaoapt4PnclSECdQ/mpoM/sUpxzB36m3
FOKzlofGWpkR88h71qXaJGJmVMqTRb+Q6rAT21wSPkoPZKWgDhd7jWM6aUrw/CJo
p382XWDx31WxKT8/vKZfiBqu5v8PWqekh1vXDXYF4rVS579aQKCbhEfwHxdOhWqu
iMizJ6zNf/XM5D9w165IF2b7fS8fIBO0ZwgDFCH/KmE0MGBaD7dRpYtBVOIizEVx
8dwlbvkBYMHBnRRtRsHA6mP1NoK9iP2L3lR28f58cXHSDGlKc5YEyT6JBANvqiKx
3r7bvZ7Rs0nI1Ujz3SiHGjSyMCFeKN/fmYokcIwwErMMMhY1yCPEFQQX8vEPy20H
n/FOqWiMDqDSRvYnEaZFLOi3NN3Sr+dr8+BfMdfmmcz+ms+629eQUfVwUPTaYWJA
u9muaiUG2lyhPwNnnWf7/xffYMh1GfNXyFD07hQA1s6DDUupiEZ6wDKUf78KeayY
W6GLZ0JtfWvKsNMrvOrqbVLD/no6Fpq/QGwfvGhFD1tljWy8UH8f6GbAOzlCWxZ/
XcwRIEWGvV075ejMTMnJ2nLaPhZygn9FKneR/GIw+eGs8ZEXfyK/wHAmg+oQtgMX
VT0bDYgnLl96ZkabTw7qG6NAvPIMuVhNA8V74sIS0SM2BsfD722yNK4XZV91XN+D
Y2p5PHMh62koQj6NL+fK0KPVumOjhWNGyO4WbJ7dX4kb2HhAWAIKKGgv6sNYyUXu
I6c+grXjWTsgaCW+AA8fGRv4U6Wta4AwTi+mnF5FMLxQpkSXo8j3P3Q+wfGltM21
Xjfbf7W5s2v2zLvF0MIzWdmjmXpuPVuJgDo9AG/A4RROu5iTDzx02aDHHcCAJeBN
CP1a9rBBGkwV7bIUjkm6mqJldeVIPCmBQ6iH+6M75bF4BGBMFbDxeKHLyMNXwYtI
JMFcJnCPdyQIwzLojdZOr1GzLVRBQUAC0sgDhxT+jKDtzn5lBLofm3m6bfmWacSY
wRlGINcNZ7ixzQ7ud/M/Y84iGWWmb7xpdFwBn+ami9GjKgYyiAH+B/mZlrp3Sa3J
57uZ3xN5R1zKVDNCZyYoQjLa6r2Io8K+tAworvuXZbgfCaj88aFlOL2z7ga3Dqow
Fw8Ypqj5GnDkPdcebtAb7i2ZIJ2/hZufSsHsjUVyt6Md11eXu+17C6Bd4eDcDz6O
VGo2usRy/1N60h9Tdz+/hDnzJGmZL66ntlYpcCugBGVpXu7B1md6PW8YLtwDBzgS
TvHRZFBiqs+sdjfR1MazrKYOcFVnmisid+5j4DgDLH4OYhq5ETq1IeGjOV7fzSud
7Y1rLFQzMndGQb1Hu9oU+EmIEXUVdoc6yti8r7YzIA+S0hyKORPQvThwQoKc28lP
RKilns7WyqNG91SeSgizW1TrctkTa9OiafULwrQ7EBcvhB4yTXB7TVFSFWnzAJOT
MJiry3xUUttZS1Qri1uKyIltnIRTV5d+BovWoChryvDrKK1Qn/WdsqKLk8M8mJ2r
KkrbGAjmfgLZ8EcRu37TShnkEyBteJ1xtmaHbNd/JRopHnV+oOjQBmtO6OWIJ7Ha
RnV6uWccNMpunyOgWnmDCpnf5xPEWkhOHSPBoKHwRtHf2QntaOKmTXsEcOoQSWJE
YNEqOO+wCczZCOYmlqvGA0EujAC5dFjxs0DhyYCjlNrQOR04X6nqHhw7GIFLeiqy
ZhC6mHZTUOHS/epZZ9GJcbGW1aOoQQPxXEqp0BSV8FKNG/LIcrqoiFzFeOOMl38+
GKVimIcLRB6galLoNv218ttXlSA4dF2SV8Nktfkc2hBe/p24dptqPR1W91Y8qdGb
YgULKQByeD8ao6Dm29TbBYBCjkOArVLvdrwkujKLsqSmre2V4obmLK78ANv/fauO
arl/BS/If40s+znTRtcRGSPpv+IWnVT3864qZH4ykOP4qL1lm9idiNIUg7bmgwsc
GlzisYbroNX3MKVDrCdSe0Me1PqdTPsj01D316lrIOacJUoxurlHERHw0/l7MIgW
Xf8mKWi0cYCBXtha5y6wfTxGNPrQOnCtV65fMx4TtUon26fyvBx6/shvWN2d1juX
M2H4nhBBv5NnENm9Q3NgniftoLqHTLzff/D3UxA8MTHIsB3m/2g/0MGq8KdGJSPT
9cX8bLlhu1YH9szDoTjgtiTn5rZ6Fan+SAPuWTCpQLY0yxFF1g0e6RBhJ83fbKnq
fOwPhZVUlWzcRrd0+6QO8MDDwW8sHtrA4YZ3KzABXeU4d5c+XCSe/aVVmEcNnyCd
3ZqswYVWGCAL6UMPIMMpYhs999O2DIaVnaRTtQrc0IDj119esZvVjFJCbYdgb1y4
15z/vf5QBoTssKz+CEZctv2+J9uPwM5+aJ5TpzlYasWU3pQEhJm2yhhnZZfzaRmR
sCQYF+Zgi9aGRD7041U0GgppLxpvyLdZIhED1Y3qOTzmsD7SUyRTfTTdqeVAJeLU
K7oauRu6qnrSwl7Kpx9YztjYGFeC4+GEytX17LLzG2fKxRhJ0Brl6tb53OaacY6z
tONWqV8iek0YRlkH4NNIjCWIbd0RCyPAaOubLHhTovQXxjdHFWMByuyc+MW6paUs
vKPQjevtjVPA8FQ07bQyf0AnkrdtReu0Hu656DEtSh6P04bH4tlks6II4lP9Hodp
Rs4XeFDLhFGhMsg21GiJhxw8T7kzxAQJ0YtfyyoUQkEID7XgVOqTX1Ilfx17KwI0
xJo1N7dVQ8CPeLZ0VHjgDfWy2R2YSqh+cZhXP4QH4Du2gMqqD6jX+UH3WPgAsYBg
RgNI4DkUeqwvizJYb8zY98MDREbXWsBEmlypcxIsj6iGCp7EsCUtug7UOvwORwyK
Ck+9JyVGX/fZT7VoGSISndexZ0hJSBrffSmzQutRg2poe55J+YSDOGZlh3aG77Fa
raKD1FLHboKO4q78FMi+FosoSC3AfKs6VJqLjBf5xcyCbgElaqRVXJfuN0JVWSHe
tIU78hqGM94fFAKt+VVbjqyZAVEFOfn9qsAi34Ybj45DdZzOw+yqwUmwFykcacPD
J59RoV3Fs0T1am1slj7hDLAZkTbqm2li0lC1XNDaexqS9668pCKXTbm3w1mM99jo
yxrOx4iRQ0LiYLV8HQvO755ci99na/gdvdcamBofPDioi+LiTey8FY+18vNOeGyP
jJJE7KKn9mPkGwLdkABblPZxoaI6vJQrhZlt2Q7bRT32LkdRnPlI1OkGuu3u8iL1
RhIbOnNksLlkNt9hpVCL2A/T8xdhOrNfLtXD8G8dRD5X9S8OcN+Kveajk537qK+j
29JoJP7yG3BcI6M96JFSIRz+WR6kjMlYF+vUoLroQPf9gkZmsOWTDDYmPx1hKhAw
XqD/Nasnu1ifSdEfcQZbYnlS7rogkHV8Nla9mgrto64djPGSdYnUyokbHETtmwH9
5+njCuILyMpChx6erzP1ZaYQ6MQluNytQldyXnpQ0dEk+NJ2pECOuQ8d4r82Nis0
z/PdmpSDyT+pjj5C/tq8brqFVZl0jSdTXtyr2rwxhmiC15QX0ykp6qidAEin7jww
0enQQPhuj832bOKejBA1PyMrAMjxSyEj5Sp29BQRRv6mtYlhNTU4M78TuZjrpWTs
3CXG6PRmLguOkbbce5Sz5DEc4lan2s3Z9CVOqsFWYu+hdbcV4/Q+N8a8DHLYxF5z
9yGgotPWbRV5zYPjA7FGKkuNym7s4vwCZd4TcyMUrfqP3sXGQbGO/YbZC/Sd7ECU
cjBp8oG5llsvDGebiHJZNqRTIom1Rq7RnHiGq+ovPJC6pcUsnvp9b+7k8H+tvm+l
9DyKd9bM0BEAzUW6pLXHTWJjUfb78Xop+kdwyAXLq++oZcZYjCBR2CBHnLmNxUVp
O9fBmjtw4QjeZqxllSlVtUjlI7kO5laYD1vXrkEnnT/A0wOMcfWURQePlhZm7Bv7
NmASNVRp8cJV8t/Dd6h13oPWNBN+Tg8wfCQCMQoBDHaoSwUPgkg2RmkLIccs1e++
N7WpXa54D4C5SPeS+qyU4UDx7QqtuLW2TZeBZ+ceFmyh1ssTFvvbKr7yyoY5vSs0
L4sOo2QkZFs3Sah8IFqnVCaWmFCXfjjGltxYca8WmKrK2F1Zfsv0sAWfUnXoPwNC
aHeokfUFfFgK8PudNL1JSvSFU13I2uBN6pdcTH0O9L4U1Z29I9l3Sv0XlH7AbJEg
JCvek8TN2Qty5XsSiAHUZiE6XQWAMdxfN1xoQJxoalkpmqmO92NrrIfQZeIC5Pce
b61Gl5myLxtTFgeZQrdA9+lPLuxwFvtWB2lArLR4HdjCKljXvGuycr3AckcA9gqE
Xza6LCZdNvWUCM/i0VqM778xsMIn4Kpfzc40glOjM1qtVj5ESM5lMgCTTS/juGjL
z1ckQQ2DtlhU0+P/5h83a0t+AHz1npMqsxC5+U3jK6cVVSojKTRPwWUN+DOCkQlq
xQLk0+0VHbxSqvd9w77F54Wt8ZRVcjIWJeVcA7Jt6Y15wQgQeJMp25OgR/r3D0nk
UBwkv4+BHZDKKu96wYvNtrUvFu/RJhmNW2N4Qau/FyPlHQm2r6m4Mi6T6p/uGDe7
U0Vx1u9988OaRDDFvz8FGnngo0VFywDGAzgJ3zmUf428DLvnMmUTRGTDLa3I8GIm
kSFRpLGwuzV8RjUf/J5zwoUA6F8uNHEQygLdwZAKDtnbNnY8JhWF2P6tl3GMKhPm
8TxxskxW1ZVqZxRFRS7JdVxdMPGgidzFqpI9WiPjy8CBzPjvyqpciXpi8LPcqO/C
woJiHQUXOjYRkWkcpxu4MlM9jT3p5CS33E8F+mS/ytyp3lubfeOk4Ydrf7Emi6g0
r+6aq+OtuF3KxhQ/BFrwonePP79IwwQ5sPfn2swhKh7YARNZQGzBSGWTHW7KCSNv
do3vZSgr5yvfAAlzOGKCZlVH8CF1LLIzQ+z5XpDniQRd6QYepQvSxm9k9NnvDD2a
GlF8yD+iUlTSOGgUXbcikIxEKR9ZnuDRINBLo0wNm8QsBf0kXpyX2UF5Of15BdKE
6UXYXh14GLYOWmBDuvqJt0bUBvvtZM/bIHymlAiY5MB63l5ta58L19jek0rBLyBP
fWT+pfzdPzeBqK8j5ddlSlZ/O/981/ikuDoq9fCImm02h8/9JMzZyFfU7Pl6IT4Y
7dlfncgwkL/R5jcuUn5b6QZocYtVgrMYJDEFkn4NK2LD2wsRJ3eQBKqIoYaZtiAL
f9iA3hjSwCEqCdzO5hp6Ss4ejVvEYMHwiLqJ2Qm4h+HiyJCQFprz0H6uTNYnFNx3
MWbL5MlFKAFO5tFRdyLQQdDcl26eHer3RpsQ+fTYIUJbaERJMOrURYbNF5rXEUwi
iHMy+D0b+hYXhWr+M9aRENEgn0N89RsPCl6I5odMpDKxOl17XgllFb3DZVHC0fin
7khAK0KFcoCeBM14Ehhqsx7qh34sHxeC/MSCprvNoj/A//dS7d/OWjeaHYOChxih
H773JqO/h/nN8I9zLsr6+4EYjCJt6XNiv9rt5pF11/ZjJ4QXSoAhaFvCJlNN5xV1
BgKXemdNTLqQ6HlIPZaSlWuDRRheIavC63dX7l+zFzlSJcrB/pg2lKow8cK2l97m
ahCxwnRW21rOCarWuxIjQggYg/1WgAlwXMiLy8MMV7gU05n6bHXANUkLR3hBDCJM
rcJJFsEWIIXQcG1DKYqT67r0RFS2UERVNSyNDtMnfDSAGd7ZlOj2dUGvkuUOevww
pJwiqc73hIQNA/w7sjOKxaI9zMOFPO0zTAiWLSNVdR/tSAA8qgySudEfG2dkMkGb
fW5uB7ubkCIEaaUMTJNGiNxyFBOtzi+ZFZ2iwWR2hleZKneE/cMQgPOslz0679Y4
V+OmdbAuMKt8FpC7QZeQpIDPnZRHuW8AajXSH6lZafEQ0Ti6sKx1lCOsx4arKnsV
j6w/WC9lLX6nxMZoEBJhl4EcYJOvswGevT8sTnL5KGXWOzmzRMV4VE8J2iSIG/GC
H/X0ENxEYM5i7k0sApesZbyK6UzBBQl6Kf7W+ZL+zxnvZU4R8EjiTNNpM0/ANgNR
3JMVtU3bcPPABkrLYHYgwzT3ejH4jb5DZp4uT58NRHi7U03HdYEq0BgAwlfGpYsT
Ykj7+wrk3xutN5UFa5Hp5Rz7LayJVJbo9t21gH5gF5OaDG7mJKCNJuZ1vslotvUN
X4XQMuBCSj7hPluKatyyqCfjvrXdpOZ1G8ZypY9n2JAX94M8U4QmI78vGEY0XEI4
upPuLyZFahqTpFQsVjHtKR8EiTtcZz+4ExWW+G+txigE4ur5oRmVERhLe3OmYKmk
+9wd30fZLdStidGLGsyAhHSNpBM2ntiVPQR5fqqNZYspDBNUKQZyF3E3MLa53++d
NXrkPSzipmTUyv7EjZJ8r7OYAdkrBdZYk/WZJHeimWOGPfKPgOUpco6mzVI7gzkE
b3wqpxx3T46yZDUL8wfiT4m3LMWvR7yyLTGg80yywCEMlTnebCrUcZRGHkphamzP
rByolzjctiBGuFIVJ5kuBwPKNpcemyfTrKxe9OUbRNRo8Vq4/RI8Sr2yFwOY/hcH
T5xkr7b/+AAtWq0AhDM/NNW4w03QuJKLqts6LrO/SBuS6IYV3ZnTj2S7aepQOIij
pN1fDu43hMceuroEJbYLMgmFsUTZ+wxgmphRSIzno28nUhREpPTmL/R4DDscB2sI
ZxF2l1pg3rFAnwpvtyGZnE4v8BrD62TBhvA0tqiwiY2bQJlty9nSOP32FamrbE2C
cQpXNbqVtQ4RKRQ1cEKggbOOwhXQk5JXxPfMakhQu0ZKikMpHKULKSbnsOkTwvMd
muGTwRWDrrNc361U+lE9sABhmsa3Z/SUvfNTO4HF/Aul30jDnL5PboakdXUm9+C+
kDW6l/E/4vaX2j3RQ28dJFhEZ9Df8kaWoGCDNnSJJ+h79CxKsTnGcebzUdN4apP5
UMPLx3x2kHIQAa08RP8jZSDywFXk4kd6qp4pV747tonnMUkOfgfY6g1gxjSsg1x+
CaEzl7Tn6VFvrRDjuDr/Q05RqzNXQj/Q2/1gw33MJU0PVuVRHGwb8VFXNwqDjCqN
jeIVdX/G68GS1X1qsNuDoIZrUsSbp/076jnEKV6KybO/r0gu+P2qlorDsTv8LLU7
Fu3Ivt13sndhlYBbBMORl/wkox58TFXSZRqKK82uawy0KbBgMTIvzRE+iFsMneQG
F7+crfLb/mX2JZ+kPbbL2PoktOULQOcMYlz+w4Q/rpLvwdDNyqx8+HhW6Lgx20F+
sagjiNhbmZ29TnbaXHpu+h0YxyuqfaZxp5iX0i+XD7Rq2YqHLypQakJBlBlHoL0W
3KqKOWbdhrgiPxFQopFen6HCFEJfTtdnejRWXVIXj+DnOQ0uXlndbE24v0kxchf8
MVNtzLhJ5yuAtp0mpim8rS0Ps94dyPMlJ97NIQ96oNbkltnRNhWPGFbjvZ8k61iE
AtpLVFmQ1+HGPN2HDYLaEV84DLzV47tmva//gBwmeYnGgMXsMm67QlGLNXARh4FT
UO1D88YJKhqG308DJznLUUpdchMfUsbc5ghMIBq4+8mK8qHuevFZaMFaL6a84S98
qj5IUjA19ZMuNHr6Xz/AhNwO7QnKuxF7EcKmNcG+1ClJ2Eqt98Ebk8xe/50EyT0f
Gm5fyMpLQMlCeCJZ5d6UHRQCK7oG/zu6nFgFrWHdiQbb3iCtT8jEFZc3bkJnoc6O
Gt+0wNdmyKgP1+o/O7KGjaq0cVtwyow/VF2jFtm0toFYG3Y2n/eKlxtspU9vdu4q
+DBRgNWAhPSINJVrCRJx6FyhBInIvuR+xqzGrZA/y/ieZNYnwYtMIwhfVbDkSwzk
4ebs/ki4sHpiPGfITFwuhmgSag1UfbyrTkUZ4rrRfTBpH6PO72WCzsIdWNdqY3cN
rI0vgdtr0KJ6/qkImH/G6WnXE8c8VrDeQlrX3fcGu/Prtm3ojh3iOKuXxzbRvRqM
xxi/3X5aVw6O5ORs4FYKeS0MEXMfetFtemUZIuzR5aOBAm1oSQsLrrebxiJAzCfD
AxigO+DtNsiG1sdg5hkSQLh7wNn24u8t9EG3QNxWYj7w8VQJm+q9X19HXl3WaYhQ
RfT1kad1qSKJlSGtFtAEH6q/HQCF0horjLUSe9FSPgMPYZNY+eiDV/qoCaHYRMXu
sadQ7KxUxRrNXcfmOscBVpCg6ji1MGZ8Y3y8T0g10eonTtaHnGTkCUdIAMS1pf5p
9z7qq8XzEUbyeEBqfVqX3mJ3tgT49EPRESdJCkBLoBJwbaX7PZ8gZ+c7PkoEicCK
PKbgrUvyRcAyXUk5etHYF/jBBkoh0hF4bR7ijEg8WHOPaN3vuJ5ITDSQsaXctc4k
akJ4ahQHxgRuXgmqO+GxXBzhsWk1FMzjNwdzW0LciTmKPfiyB7do/Sarw3dk11Zp
ouNIVeBrRxfX/V6vXUIdyJGSeq9rEsQXE0+F2EHSE2HYJ8dYLeABL+nRVEKkTnaE
lJXym5Nc6OekaqnqyoDYnJMcjPvJVVhiqQ+6Jr2cKS2urOwDuQhHisvPExAnBePP
3AlON8WDMf2aBa7FbKUerv+kMFouubp7BbIxFpgkGKs1vGkToL1jwus7YuDBr8g8
SghrXH3+ftN0q479lXrtzS6nLyzZ1/6exNd1nkfYnSM7lgmDCG97GSIgRTilxiZZ
ELQk+K3xjzbywUj54zjAXjxpNWl8z611RVGjbDnKOyAfwCV3oIlR5sGw40L5d1MH
ez2feXfr8kEJANu7CXiwXPVkBb2L/G90iQ3MkfS8RZotinf+ZSZnN7Sf9y4uO/bU
QpPEaiPxKF1TkbzGtGobnZ8PO4jq/rGgS3Y3/AIYfdG+pNobFbXqeqqiaDDnn53q
XG1v8MkdTq0pKyyRHVspc3fe3XwUx7c71gSw11N69m3tR1UmL0U3NAn6UFOnIrDY
01/e/n/QuHogQmz9p8tigb4CBxe3x8Agfi9WhyODy9HR7r7tioUotpqja+D8ys0p
VRfxkZW6d5l/KSqM90Bm/mFGzVWa6B7ul6gs8PW44+qAT+eje0ESFfOAuCPlth9g
NUEeafn3g0JApcJ6eH6eNTIvWMtk4q8AUfP43dE3GaGcfFkJfX+7acvN7vO5pp9W
z2SfbtcfWT/E7BCtBakjAd/2XxfzB3SACDlC3ptJmBI0/xrVgwPGOChmhlIoZzYf
4QK3dr1M007TNxMyOFmu5p9zPqR/wOz+PuK4JItbaNb4M8kAAUtNvV0pV1bQICHx
hbIIHPAD61zogXoBGYdT2PKY+Cga9y3aHxIZX5n9ZVi7w/0jXWOprIsH/8yRwNzI
U6tyhdc9lMvY9chXJBw1JQBVsOZTJDALqoTty/mvbwyHc2TBfF+9DqbGR4890rX2
gCqy9kEIQxvQr8VacuXSJk3bUF3v4GTmcHO8CPHWi9zacCpEUFOdZumIT5ZF34jQ
d8owF3dG6zwA86OzwkKMGelBklytEikKvadbQUewukzau/1OiTUveUGD2JogSp42
QFq+67JxMroIR3Dhu5g+1my8EKSEgXwPac6VSSqhcSP4AND8MYJwJBQ1SX0X3nMg
n5VVkzjynSVAUgyEiNsNdbSe58D2qq98De3UbrJ4cQ3WHSs9PyFHco0ruMU2fvKS
nYIxpDfU4NyNU7JTeDKqttkzlsgDRc2sOIhzyrNo4QIjyQCS35xyzlzVn6j8/TPG
G5BNAlE+AZkWbBSJDVtZhn1s5arxHn179zgPoAZKlfd1OE2pXjnP1YctyaEbK7bf
/8Dfc4k65LcxImSJBmKmFncCSVPus+tZxhm5phesVCRsToZQjscPa1UOBjO3FnwS
ThZDGXKnuzVIlhvrZB1eAF45kze/B9XZ3TsuG7N0dl0ko1xrZqkW13UPvdaQxAoW
uV8MGO1/doyyp3AkDFICQvRq/tXm1XfA9VIgFGNueui1NaIu2d1SwHGsyM5IA4ca
26EKRLAdAFCcbMg9vBvLF52sCLtM4j7phALD6hXKO5Tw03J2Ve4pzSPJG6rUOMoW
LMo/rSjZFDbVt0kDoM2oGf6RFPE2U9t9cnhaWpYxEAZFtKniVRmYd9u1zuaeq0Ed
C5mqXXl5S6QlADK0eG7gBeIN6kPJG/1K90E+PrSJWO8UQtvtogjptbgszbD0Dmwx
PbQ4IF7pTO6NeD9C+1mZ6+EF7yiyQ+IdhvfYY4I1Qq6ZRofPg668dMK+caBp+izV
dXy9AcuHzIUZSrWITYmlgrkzG3AEMIh3hYR3Z8WInCr7RVxtsfWPNBcfM4zSvkET
1AMgi9FKgKM9PB+lCe6XUrRyi28NOWcjsL1X32xE+9GPt9wQsMTcjWVI4avg5dI0
7dPZXcsSA+aUJOqARDSx/dmJ4uGZShKJ/kaEzxTQCMl5UDDcALG9bHsCNjXvu7wr
ahUVONnbtG8GY4keq0NK4G0CkEgQUTW3HScicuU09DgC1AflAG/N0Wik375+WswG
0UYINtH97xbVj9KLEYbKEGd40pYIXBSie35yDDVI0f5SrUG2FAfHlgqjm6QBk2S3
Qn1w7P/XpHSk5Z0ijsQaV+cx+eX4niH6w8UbVKqzN9HHPgxswKyBblDr7LouoDnM
XdTw9UmO+yUcE1iLt8sdNxSS43rklzCBGXJWxaabeypsJ+60wOcRWz8fd8l4eBI8
QaL8/rlSBCkxYPgTKKVz28z9AXuyyd3Z+fk2SWFmqUte0bPm78xSGPPwwsTYlQNu
TqbpVGzYfkiDjsnbTQEgAF+ZtJQXZ0uD8HQGYLgSsQujxE0Dnf3JOBb5P4USmWOG
BkSSzHQUdjzISVGOyC7AMmGD/q5iA/q0/JoZBK91O4wZF/PmW+AAzMJrT0vVaBTz
4PA9kJI6MeReD3A/9SXA5p/sc8faKSv3H96aFAsX5doCH0eofmfBy1yG46VfZGlA
K4kARuRKmY5rpzdgape85LdhgY6pEMcEgf0AkssutszBPUNc0GtG+Ratz2tAcVEv
33SBaEUrRLXvFZW0ySJmqEU83bItUsO7LnBiD/tX9W1Lb70KKDyUNEYtjl3c2SMl
4M27DCn0lCUWSclDawpyxpve7rMWDgTS8ndR/Bgf7eqD3jEhVCd9cS+2CujdvHEB
SzRSNmTJNUqZfU4cFkDY46UPLv5IEHzsLv4zkAdgv/N+huKyeJveDb1VXtE428RE
/NYSIVMLx3eunThCnD1xUHfThDGjkvAFk9DXdqDqxK4dcHPFzanZ0/z7403yTU5e
ih8UgE4HO5va/OEt2ktHZhPZevmc3gaOArE5vtj6pHP8y9QLf7z7o9T1AQaUY4Z1
c1kdQaDgoyf8Ipbn5eRYWMhCVc/AB+3EHquzkwkpDku1Tt5NlA3q92Ny+qst6RXg
BjCYJgH2J/Q8oYo2yV/00EPfuEHVBzd5wHb0JEwYWgG/3D7IXWaOku7UCId5d4iV
cJINaV5iezBaB4ER/5NJsO2m+ycgpETQLbOtQP2RPhLOg95fNMMhq/ojGuRfFi2g
b2f6QDaVX91uOhVs83J8jmUDAgsoyXczisiK2fGA8O7VuiHhVlligEeNgEJ8hehe
qmfYQI6cNmaKXxzTO25pr0WOxXzusptx+dDw+tWbukIAuHXPTMTmLIfGG81LdNde
tuxDYh6WzFkRmF4xbZjgPHNa+AAYyrcAZfWdPfvbjzB6D4txJ4a8ZL3Kq3W2kk00
/wKpzyZn3jW670lL3WlTPBXbmvBnmS14Shvk/jFeQVwFysAOCOVyouVHIKBVd5Wk
A6ecbYVuOk8avah2bbnziDGEJ9feONGU93/WBeDLzSqj4W2zygYGiOgcAuzRhkv/
T6Qs9dGHtxrJ4QMNQRV9E/Tn5MHmQ8jQaBMidaIlVfwgOKNhAvc/BShMmMZOJ8kn
bMIKTiHvZJJgRaUMf6Y3ONebQvrJzJPzTir4Kti7tXIk8LnpQ6kICq9R65Arjch5
t8kb+nxrdhPjH6U/GxXclQoZYLwNC20TnQNS3ADDUrOV8Q/fmFSfreyCfSu6jRWf
tGqfSWkHGZ26ns7sG5LXst9EwR7y+V/CbU1ZmYeD9OixJoijk2/6tIxXVuV45SwB
bnKyZfY+VuOW8P/D62BVQDfiYyZVdwhyoiB4V4uJalb0nKNMrEWMc6uELdDcr09m
BETJiPAhNEmDBT5Dhz43WjQf0n5Q+/iDFWOXNzuA2WIgOAfkx3kv5R8QUgqRwz2A
/ugQSh9L7KTJHxxkmCMCPQ24WPLz+MIjo6N2bCbhv156pdbCHgbiLJfPcaSwltgu
2U2hits5K0ujTuQYqjmv0Kk2Ex/DFQD36sug19jdY4A6B6jwpPDmalz9366Hinne
cfkPtiLpR/390Rsmq8xf0GJejJFfASSUjhpJ6PLs2wqP4ywfL38DC7ysOdZF+aU8
Xqu9t7fuQez10tifLjdMfK31/C/FgvMaN6ILqbansyeI0ZMUEeJ+BxMISjfYViF0
o0HY1uD9iLlhr+9cYEcdgOnZXDl+c0TkdkazNXpRYZn3qitkceHonbIUispW/hXz
IjRh1NfWpWXXL6+LvlRI5MXrNWRzx6AlBu3/GhzBF/IZFUGVmDzWRWiGsAbmLWwL
8OY87X26IA/jR39qL4db6AQlX3K9vjPg9pPFoLd80t1FjrFth6j90Dwpl7nHwnGR
wlGEtbMDBfAsTGE5GQjYiMt1Pvhf9I/Is3F7z/IWl2L9jTOzTo7SW5U/loK+XQQm
IupYDeMncEUzi5WEDw59e2Qm+7xDWJkzkE4mnR4yY3Z6MN+yr+yXMAo72jEP2Tc/
8VHYU+C9NBilARMMTnO36qcakVGpv81D3PIDjKXtQS52H9lwl2xSaOTF8ieQbseE
+qj59w9Sq5tg+IKytfHcACJKf/HMAhM8QF3tiPvCEb5+xZv0Vs1pQv1b3c5xgZLW
vghX+uYJzBQqJy4wmz12wLSiiNV9boSxzzyTt1Ug3RGVd+GhtoDeDgHVfgqPgTG2
ZEsrq4y/oDxU2abVuMbu5FpRjz02h0+6WpQuvtYCEvyOeJUsUtEuKQejoelvYTI9
Alc3STgGaHP9BH9nF/5c4f05sZ00VAPnY3R54JrPlNnKAmH+PpixQmbPfjr4O7lh
M3fieW0pN2cHmFH2SUWKSVaQg64uSw154j8SYgmjH/8vvbHMO3v6KZbu3vI/WCTb
uzN8BwOp0b8hoh95WWcHbBDloN2IwVwSCNaEnFi86ptexj3OSwPVhsIPrshbqTQm
SNRGG24q5ydwPCo3YJHjNE6dNE6evRTSYKXYTbqxJhLBTQm1QZO5OYet9gGiMFI6
YKyK9CLlfVODmEyjzlIB49zrTQek2RXcG8dGIi9xVeVI6g3xiiDfOr6V/p/lO7BG
owTpAR7cY8Kh6r4iXTqmk2pZnF7gr1u92yG0eg3nkzlfjzpg1P8nRzllh1/M1sSC
aSLWNfOsl0ihnoDpI0aZjJGFyTIowqlWWvqpUrNH7Al1CAMKGAZzgjBZVzaiuKy9
7PoIJ3oiV592vNCwyhSJPmKIXgmvP8CPDTNszsOIEx2+tNzpB+xeXKU/SfkF50+3
xsC2mGwGryY4lySraYR6Sq8W1F+wX3o4oIbwEEvyYvlrxJNTicwuodoGithkzgUk
3m36XPh/q6U/fJPdJOfBG6c+LuDyYARU7SK+HT+64P+LGJgkYvxLKvkNpUrgrrE8
/Fyrnel3+ltm++5Kinoqa+yenpfMKEptoBS7WdhunQjNejYJy3LNu13EzB0wXsHU
6JFZoF8PwVcU3258Lniak4m/Apr6SPzkLjSG9rMjcxU0QXHlAiAo9SY5M66AXwZ3
QUZa+aMMRvsyExRr6ybVhuc6bkIrOHuEOYQpIu++kuWZRRIpKusG6Dafk6/Jc6wt
dqXvkyAYPfv0jTp3o4W5u7pMcbqPBT9VPQ5b38wKzNWKrIez4oWTqoh1CoDK5Oh8
z0WlxusEbN73Ia4MMDiZZcjAr7M3yI0AH3/LdABtgfX7Qdz1np/O/TbHNoraQfmw
uPZUNZ/kBqjVPtiuEgzqwSaAZ3tdBJZ3oewHT9e60oNUHGysK3N9ymgOXUksAOLB
lZDM0q7smVyjRVh9NxoIQHzNOJ7M6PvxH+pHk7UKGL/p+t4Tv4/fUmVxKoX/ZcYh
TlzNl3dB5RGvEvDAt4oReyXTx/TRx5Xo0DZmOx+je5DmWAL4yLRD8rTtpCupblAm
JoLqIVWvpM08LygVzEAJ2FfpZQ5F3Rf8yDcyq4yk9nldpmhhG7eEOWFq7G2TEqsN
j9+qzBQHUH1Qep+dv+lYDeR/oosO1qkre6bvg9ERfIu7pv2l91F6wdonZ1H3g7ka
HEFP9vcQ4BdZaRLaAzzrY3wKjNBDyWMd21GIgiRw/XFxYKUrNlNiUM2xXIM//ZLt
3KUJH0pj6wVcp3sioj5/Xls/9yah1jEJPHnjTtzidz1DBrNmvVrSJlDCg9FfQaNl
rP6N/AxcKXMoJrvlPPLI2eH30Sds453ZJ/x8zvOK8AjiE8/RUXqS/RJMXq7oGPhw
/gAmSyN1ppu0aMlmS9uGR8XS53Rtj9JXeaRhC16mGsVZxBAS3UBPMzMy8/lmlI3Z
WJ4U9DgPdiutB4TcZu6biItQYJv8mHstGNjQgbHy3aaiBpxgTukUHo6308nHmSSO
Qnle6zvfKyC8ZFlXMtiajsbdpW6qMwRyRjQoC9pHTjg9OOGdRI+Mr1El4eiEa0/0
79SVUVGhPYSuMUz4sVpYccw7xluwaA7jx+ijMo86OJI7Fba7g/GbmlnE5OaRVyGK
qxClW2R/cer7WK33hTYO+RAxoxFv2FsG6Xfn+6N2XI44vbYcm6Aw+JZ91k8dkpIE
yZ9Lx2r13QRWXg22BBREeAyJrshaUGhnrfNX9Y0Y8kf6yCbH39F2H64+SNCuJJwq
6DJfmDZpKl4idXz+K6vokaSOZfQOQp7AzjEjRs8Yditz8phG7Xhe2JHUe//Mh7ku
/9C88qqbCZ1xnbPdhA9gZQtDpWWpO338iR1/q0ENAqR4ZEJceI20QM938WQjf+Ah
m1UhYjUOVGiDZjZxEVjqTnb3PqS6ZpfumBAbvC89WnBiHuQbeHWEFxCHvlX1sqDt
nVF9AM/jXWwn08+i/YHwHQdx6oH5yYIVtH4zlHPlergjWBGyE6zDrzqI72fClsxO
7ObsFCCfgJKsmWRleCq4S/ae0EKg7feE69576n7eIDOJUvsEfx5qPBv3zPo1IdHW
iU+OF806MCDdaau8Wszf+OPSMlWznECENTt0gUaRWy80auPLuzLT8WBBrbhwG5w6
wYI4zMUG3D6MljA5ZiSkj0i4pUMOkzWRh3NZbofg+mGrgusHjknAwZM/i1NKxNVX
U+JmrbudMUmhyS8SlShIpjU4jXKlcVCOQ2ET0XjSMVghbrArp+8U1/k9J11+MbSD
hCyf26FFEkNrkMWt9BQ6M3QOnI6k6YX26uuWtDpvL75YrRauc5v0k5dgzeCpWopZ
4ZAkaze7Dbtmtg3RljSKy0kgDYtd/FBIIjOsy4aQTb/zaM8B3kZndSWb1xYDJUjP
1YxDwQ4fwncpOJUfroPJapCxZERZMRklK7GfZ7a4CIlKmEXNoaOPfFMXhH4QD4mI
JxiRS8vwYpWKm+O7ELolkK38Mk7pDb18b2RVpnzqvceYnBUdcSAinGlGA2cE8oJB
HnL6Ocn3MwbSp3osF12vClOkIl12hdJjmw1GDXJH9ksazzF/W9MOlAjxYhuvF/lS
sxgts3Q56A8ww0PKifNscNDlwMtmcoe1pkmgacy3Fdg1Kf/rCXrB1PZWde5jkuLI
5JlbrulHAMsEi5akTvkgS/a42FljNkLe8ZkFTsJj5XLpBdFGC2MA/i65c6HjpIU6
sPUNDAi3Uvgjjf8gXpoDEB5f0D9/z49AuHfZCZYIz2WcqFn2Qml/ps94WjWU+py1
1h3b+hghkePcs+YOD4zlWWZ/ypHJIKrZQwzeCPCBU5imAnoBjXls+DfAvgC36Nfv
LlCxRX2204XsVo4A86c6D4E3/AWWemy5lG53uKDG4hRHnD1F45iciTNWv0sZYfVh
TzZwGm0svYbs1iucJ/YTHjCG4EzDGy62B5kPpziFukLpJVPknEoCk5DDRHR5tNWl
jlaH36E/E0RENpj1w5gRP6Vzg1iO0oM42bEbW5YsvLDwk7henQN5GetKmL0Pt0G/
c0X9NvSIQG5/jirVP7nO7XateUxLGXSVroG64WYZtq3zNZyRu6Mk9jbm5IifKKXi
lkYs/I0d8pZBrUnZqfb8m/AwTvmu+Au1/pXxjUOhcCBtp832SUwO7kS18hKMNZEh
QqaafOijDg3bcdrdWHJ0eHsWF5e8710NWyy7hp8QrhcaYpbiE4I8ghMWxaPA/bpH
jqa7ruUcTiR/a4Iv2amIQHo6CgM3GKlPMeXWq0hqAq5wyIG0D/RK0ELw2dH+jwYK
M1cj62oD4ChxvTrLv5iAvk5g8yJWoLnkFEdPo7JavcUkXQIyvMqy7q1aUD7jvjpk
ZKjjB6j8FeGhDL23x2II7cEB5tftgsrKUba1VsJxGqkSE3bY7CBAgRkxNWnJ1XgV
fWHizkxyB30ibzySl/gnyCoyTTBE1vYDVxcBspA0cEocm3uruptv+DPPK4vzxXvf
GimovfsPZRG5oQrrSRxZi1BVJmY9rReDaNHOywP6o/7NFIT9e3nt3+ZD8swOyrx6
QdNsbTmAzC6vIYKkLwH2okDmyvcg4p19NVPypQ2or85JUyUHQ+DhT9Ltw8RxrwlP
Xar9g1RUTAivX2vER7FS9Q7bZocsFc5YOADkZmySOoaEy1Wqe/0K0HDdac7t/scy
CamIQN8QYrE3xZNrYe3v24SS5FsgDr0BOKk40Y+dLw8WkTeNC4f7ofa9m6pNlFKN
BPQkpWJ1Set2QI75iQ7BHsGldgHJPWeejW5bH5mlCJLH1JwucOtXcC2JGfswx6cw
MR+NPjAc3w+5NI8euPrU0duBGgY4Mr9WMQU0NAITqiRh0xxpNk16LV8f4/xqUkZ3
KhiP5ghVwyHztgyaP2gJzFVQW1JI7yAaRm/v5ZcE6d8Am37n+TE3zpScMrYf4SP5
kMOcRNzLEOyaPXkG3vd2FHAa47OK1BQ7IkQ7JgWh9vfjxcBQI7FS7MNLifDxuIP2
m1RptssKrQwtMd6fv9eYdBEIDXSD0Z4Qt73nu16K/Jm4bqNdaSNGAfmD4jW0d8O4
YWVBSJ+b2MHez0utcob1uC2/mUoYTwAc9uDNVyZNdbWDHjsE8POPatNC1AIS67VA
2cLX92Rv8qScsfLeC+y6pREV0XD+EVvOejwcY62QbLQbxJM/GdQSQOBU5Or/ZiSv
Y02nGMUp4YtwYgg7JYk+zwrU8POYTQH9T8qzO3dr1zoBGNF3C9MCLLxIBumr5dPB
eRk2UWPDYkc5ySBHeehQwwxbQ+bnTJdTzOq3L0rrMTqF3WbcDdzWuQM3str1XXvu
HQOvEvloThPI0nuPNlECDtmMTFb/0x7POllXh+/FF+xidJII+8/mHTkM3g93EK32
Dmr7Jb4Tu3sWfvvLK1gtclMALP/OZJ+C2mvIjlS5yxqK/mXz6TmNftJZUG+YvyqN
dd1h06t2h2jboBPCemTgUI+61et/VvnNoSg0CSgtJZnHjTSK23XLS4oUZzCr5IhF
y/TboBBFbGhHsoMucPlsKnOGBW9mtge1ZcCKacVjbhvdgV7ZiWbVaCRu+Gl3N36a
/U6QxExdJeuAmyJsKPxmPxkirjVxI3PpvRQr7Y13E9fuIzspIFgEUY/xeWMPAgnX
xsqi1fgURqlHpAfbmkTv0jxHpqo4wiWyE5XUfprK3sYPK4+dtxWCpLe4SMTtDQKQ
OUfWbLuKD76nxqgSwD2qeDudJ/r6BhMET0uL1LXhMqHjLR+gXzCsLddix8OQtX9n
nO/+GsGgInXhB6BqWVK3Xz7/tmIrO93Acrk0O5MjF7S/x7kg0xDtn4o7gV5l+qTZ
o8q1grkwAyeh8uYa5GAnh8DGXc+YOfjb9b/kc4kYll+hS+kgG9AgZPw30OstsX1h
TjCpD+hsEE0W0yEynmenEBGw2sqPeqt3iJYuuYkE6UW9KQilDwgykfzsUO2wFLvZ
2fXK2frZFDOAulXK8NI55Nzm4rZIOcWLXC+WNqOglY2pZdfzqc5dJss3Ogt9DI2c
SFx1djT4aATN4oNlXYEVTnbw0O4mzNQS0L+eZAP7Dr2vyH9Ktuw6Fo0T5xl4hQKB
fDrxAgo08B0WfB932NYfMNPhwJXw9HPAlGBAfStom0yB80ez5ks3o2WXFKQWutrg
KDKLvVOQrPwpgZIBzxV4al00qzZ+B893LXvQJwMGxB33mCO+sP2052yqFsLbqZuO
tjgxZAVwHB8cFPghT5MUuSR/dGKGZd73kCGg+8+FcQwZMfWjSgNJEzCyyIa0a+D2
c0CTPm6prbBlryNY1vxP1m+OW87aociWi4VTzXg3gA59+gq0m3o2XB08EQrJt1dz
qDq87wAS0bEy0ybW77Sf8xplLJhQc9dTaUMEklZQKNaAe5jpgFCzfKjwpR+my/pV
b3Q2i7Zfzx9De1Ng87b3nul/C2aeGemSaQNZMQ4i/g5m18rcJV2yLPzd2xyqOniB
1/s0TD74rGcS4tAsiRZ+YofkcAvnv9ZuvgnsWoHAuraWcB75BRif90FJvwWbmw33
hU+z0sAF5UAc19X8wgM6+q++jiUJ0jfLc1+U4m4me/NEf7fAtc1W++ndCEqmW88a
rlHtXnfb7atYwCIwT008BvKOMRlgLRsWovyLRjvse1De8QY64rNR5wKF0q0LJOyS
xX/3yDrNArTXhbIjIIbYPKTV90Fu0qInY2krPEy5msJ40e2+L5nuSYAe44sRy+/d
vY7nlQWtmAvgLVe4ZvkE0ej7MgLCLEm6niSJsbsOgSXAKqhmoqyv1N4sU0zcHKxQ
+1Mv9AK1P0f257VyAU83EydgUYMM09na+IL3XPsr44TeEiqf0+LiWBl+HZ9PiprQ
spXhERXXBaFI+BHpLCOrnzQj9sPVFF145RvI7QOvyZwgbeVsWKHdCyywk+doLfLb
YxXAl6qqd2y1tGLBWagqWKxnBQRWgj4XCozgkKsfCIlLgNVAlGR25Rnk3G3+ICnw
QKPTbBkc7o7BnlqtSvTGhmZghz+g52z3ad/3y/cP5tlh6p9hsKD4T/fAGZC5LhmI
IIfJdEw0/nwJ4gVrTPNi67Wl74OuyCX0AR4EcAr3BnV8nMNO+vxrxvKTxzws7vk5
cVmkoNLdvXapTPd7+GURLjom0IjEQfeOiH3Bq4tlA9Cr6/5NZHpmGra88vZhG7aG
oCzLav1dA3NNK/zmFIkMmS2EuAtlXy/jrlQ14mpfZpoRxK5Nh/Q8ZoGONyNLoHH8
qi/Z8lPEmrJjVvfDuFeXoRDJbE8G9UE+1W/4ZS5cm2AS0lCsfg/F7iALeTBERzMN
xywAB3jgXTX9+IWWGqfwpPsDLrcul8AKYcY51kIW86ZCRGhj+6bHOgbMHqO2h6Qj
nXXkiX+qpsUTCjkGWvT1j6WeiDcEh307lPHdrvU8Lmauo9z8CwCLFnid0V7dPe38
IeyHXJclok5S+BGwbRoYRnFT0F9uzI+LMrRA83ETLt4TciACo8yK+A9kH6tgRFdb
US4snJ8/Xhip0YN67yCkvtmSbOBqMmxLxiEgyfjCL0BOLtbD6Al2cEPFIsXwOsSr
lnPSjy3+pZqkg86S/HHxx38q45gU3I2bg5AwEv9hl/JQyDLP5YvU3IVi3UTHwhJ1
WZYcTH3hRqCZlAaHnvF7VMyXYbcar2IFuH1bArXFm4j1Fn2aKHIb0xOI4YkO35kS
zDPiqOSgHVuNG16kok22otxvagDgYGa3YrSH/e153EkQfyA9xLuzBgLmPzOKtqUH
SgjHFmNZhQ8dvyIju8FXZJ4w2leRUuRGtsX28/6b0d8t0VFXvXxXG6YJVAyrWOa+
QLsCzEataYmD0ep04f+Sq6Tc25c5VswXmt9PqOjgXhlutJZoBkxHzMM+sbXHm82J
MQDKRHp+aPNZO1yVrJAfzAlpqAB/qIRvgTKibDDm1WQIs0mN+SMQoOunX9FaD4Qg
W3HsjPTTvhGONVJdz5VECTdPc14V7hZv7nf31s7a3zDde489QT/rR8pWE6gH3Chv
txSwCuk8gasFJrrQGZ+vK+tiv3J+m4fxqlnFv/NKPkN0j49AAOxdhfdH8dUTCzeW
Li9NwYhB3IaouDnRfBZdG1ifA9xtvO0mF1aGSs/EwfiWfsgWyqA2k8g6iiEG5PMK
62Cm6tST1BpfjtQA4gV59szWU9+26uqif0IH5OpCiLgyUeUYyxBl6dGIdlchfqfY
ASKwsbXBtL4VUcCmnv41Su54AeAWILbWwrded9ItVg9xlITshCus8VHIz1sQZPR8
Y9tTvFOdx9u+pbM1WEOKtjuFFFCUeQmX5Ee9JBZd+kGKFcsVfSEmAFJZIvTljq5b
AUHhIYqzfmDCQxdmOHXEJnZu8uHxRLi6QT6jzj5GbU1POgjOHDRYcCz5OCNUuC24
GtkQi7E60Cy9DlIZzZTUhhotowb0K1S/iCV2kw9ybmRKH/gWwm5VB+99qDaieubV
kxTZ/im2UOnHr+GFpWgF8Pj7nJhEGcMrTnM6YXcvBl2rFUdJRuKK0atTyBf5tGLq
Gm3M7wDyIlbORdLDGCyGSxNFzZrimDjQBGXp+4E0KyMpz0yCrOi/raPnMUYlubSw
BVF5nO75gUwBo5eoR0WFJjuE/GBiZ4+NP3e4/b/DNwqN6XUD2Nco8bcBxr+8WYnf
HOHejP+PCY5RaeB2H7geFabA3i0OkiIvVOZsNpDt3dauIbo6qHTQHcZOq37vbhb5
3+JsPlYFlcJGE5ZxwTBSka7bWdP9+uV4GHbf+XEMd0QOEIP9/Nx7zdzRpPgP5mZD
4orCLrh2nlA5LI4OnnjpsH4rqAwUgSVg1YyEUPDs1IqLHh9R5PI0I9JRdQvzvvRE
66bftdjcfYj/YKj+hgJZuFoGk7wrJxRSuqsbE0LIeCD7+0zyxQeSnPqnLS6y+UFV
j9VhufncShwNq9l8edJUp6mMVBCqOiNbTbqgY373vRNLdjJlFGw2CcEZONLgXRfU
rg/XPX9AJZnjEU4ERafnFHMzeJbpjdRR2R+StXc9MiDZ3M4ujpJSz1IxyRbKOBJj
KKY56HJTNyxcAeuGfGlAA0JRXstqE83y8UEK6jVjfN1vuVj5OKuh20j9haIsh22Z
DLuyzsSBPwdxOCHJhdbd0h5CO1OUbrvxFzw4nvKPsrJUNblkry/2gZuOey9YNQGA
rn78fLPAonr4ivqH+fIGGRpmJqeQOkEgINa/rmevK1nsjLF5PxUmyHcxZC87fUVP
WjBwIcVyOvN6PXpzmQ5TS2vb5NogcWg8MZl6v3N8LBnYRe0Hg2V3WOPS4m9kTzq1
TaB8z7WIPsVqY4LURfIwdBTH1vPs4+pwBcc79gEkDQv5B395/l0Iu8cdGKM4XsHw
ThIhRBhAENmUHpw6e3trvUdBSEzHuhWQXgSQoWH8lH1BB2zOCxhLMaVQBRWgUdRW
fC5GIfzxviaouaDw1fSL3EGtCpGOXFLLmKFR6PTSVbCJ0QcgnYg1f3o2Hj1d/EJx
B9ZdSEM090zhDETPBfi5pxF1TCTpCdGx/lb0GC8cT25nkOzl/cqPBAyaYaEHUmvj
GfQiLkKNSczs5tky1nVOg67eUOxLgocATA4ecNCBTw4wuRa6cfTzh0HdJ+eExLfm
5BYC/wb0q9OABZ1xhYh2AFAYPcnXry/v9hp8t3b/dw1JNT0yDB6TyYSf/536QxFh
drERUkhfGrGYToZf213nldLksPHztK8RAA/7P+GAAzXA5sfEUGIn8GTk4kvrFLzU
HvKbmzEXyte1OqIkRzn3ztE3AXoY7+ilwqvLKy9C/s3DTsKuRhlMoTqnwLi9nOXP
4izSAt+3lzDyvWOHXonh654af53iV7DQbPlSuO2F3CnuAT1ZVIuTSZVYD09Mpua8
3U59j2RWLwnZeDPYf1Z6EGTa4wSsjo455vIZ7pjKVqR/dIg4jMgLdIiedzRzDqdg
l6I+TiaK7W9Gfes91acRcydMO/etJJp4b/uuWF+yLeQSL7gb/8MZZmQpzDs6gG38
GCjDHcTbXFK4ay6TxcavduiNz+aPqcG8XmZO+blUWl37E3dGw2wepp3dtJMhw5CO
sqoxELF4uu/MhQwWEyL9f6hoisYQ60DgjXFikkF8C9Glyc0Ha+vIpLITpeaM2hsD
paxxYt6sN29HektDGwYyPOm7/udAipXKQ8yavQ4DWqafVCCPriX4jDd5qCOarB43
2ITBsLyHRhh4Ypku8ClVOBwLEwu3MIvJzj6yET0Y2ECFYD6BkI862TuJqot6aGgM
uuA9MFX6YKR3no/5CG0xFMiWWoJs5GMiBrYyYP7N7iAJ15KOuSmWyTJMdQY0C7JG
yh+SanzOXLlPz4/UDbeSJAX0Xv6HGUPWfkhSRRpOjeYdtp9FcvZni6Q2Ic1AKnrf
6kmGcLWzIQtl4ZPDiuurquFk8+hCEZp9O4pY2BRx2HuwjhX1XSCBi7ozcMtL0yEl
xmcBQcz390DDjyUyTMBw0CdufNndQQVJEkn2YMEP9rW0/igUYGEyiMDnkU2G0ykG
Ir29s8LvA+SF+x5H69SCvPN/gIos+IwVeKVuLe6pDD2TdoFdupcQLztQtDRn18tw
ZzzOP9MYshxcz/osEACQChhRhcTEolXJR54GljjkjtTG4/F3eX2T2J3U5qEH8OOE
QbbJ/S8K1hO+nA+zjMBsP9GF24CuD2VaV8agbs5teZXjCSZEX0ixqlp7k8+lfTT7
uiiDINLzStxcZ3ZjsOKGNbPGrRMEei3107P7WmuHkJNdcFvWUcgB+40PZrluu/0e
1uhHiS06cZYRBqf7K2Ia9Xu6TmenTbzgKw1O/e8/F7QSmHHeo53BUqwK+Ohx408q
hZ36DZ8evtLHamVR1KXEKKDqNwXssLoXYBVh8Ulsj6/0CQjGaHTGxm8flwCLtVow
+JqMUgfaAOp/dtXrnNX+8GUHWt2gwSZn5iXF2wIdX3mpwYb56vPL1wyLMFMbL8gn
EfrkGLs0uv2B3+KFzuC7uBkHuMNw8NdowUbtFzQVBOQDAOQYyJptnxYljZ5sT+Yn
NC62X9TC+L/zf2e3PbkxPgPPYW6vvD7pRxVOmZTWDdOJUgQkaUIKunW2/baPZPNX
geR1T5vjOoyfh7GTxklD5dE2mesOQZM9Kk2CSIS/R/dtvut0sUguNVhgJceM7DC0
Q5/mR7Uhbbsr/g7PMLatJcaMB2XZsQFGqnMwOWH5Pl4rO4su0MsA05UGBA435pZ2
56GCImUFXJNfTmiIzWKQXt8roiMT+fXPSHjgiArvKCk+Jyu2fifFDspcUZqZOrk0
s7D5Z0jQRo0EKaP3euOdNRgxpChcepTAlBqsk5aDVffUbmGv+itlXRF05jiXacaR
Ngl9uEBUZ+S03G/ETIkbk6fH7CrH0t31JjPQAZghvOSxlO2Ct4mxDK9Q8ko/gvef
EenQLuWo3Zw3LUThhACMRzUC7bJORBsD2cdnTNTWHMEpTWJ3DRsynZy7t33PYTu7
Wjvi6B0r5c4Ld4QGtA4I5gB5xCKmks9CplP9kN72DedCXzPMiVQ3uhlZz6l11rrr
Y8zhunppBHlTC7DX21S8xHIWwJ6XhRWS4jSqXXwXi0MDNbaVVE2ECvZLtmvK8jDX
LbKAXrvNNSLoB9Ip/ojL00wZXIWNqVYBW53p7YfJMHifAVhAiiejPMo94+8NfGes
hcpYQpGMafl801SVaEUKawMm7Kq7HLKXmRlts1tmwDSdIFNGX7JdhVWFq6syyHnI
10O7nJUNrfhp1FPUL0ANprW2OsrBXOVmYrEbluLwpHf14HAHW4pitSXqgZZKi1WU
F/jesMkdec0m/09mPFQtINWfHb/unrsL43jZysbzTbsLyoNkGvL/gEXVtcFZ1VLZ
PDtZOh8SdLoRXXIEW3kGhbpxPbPNUrEZ7p3gH9JdYeuBW7CxJ2Zpmk2+G7t0BJmv
F3E5pJveNDgk3dpZq9Z/hc7sf+/K3yFOv5bYsHNi5dDtXvKqgctL85fr0EU/BcYQ
YAD8hDXVymSIZ5vGJKhzFXX6fr74bTguiQ4U9mX2BLWzjg1o5r76k1G/whDikRSL
TbjlfNbQMcBJl6qqD6RuBWq+Yd26NbMhxMjGVpG5kJ0bEBVWmXjKrkVlb/HEfs/v
naVw/4Fto7kzmmijZEazJs0GV6MBoESaF/KkVK+RVB5xQ5515UeThhKQ7nRxUUgW
0Zv2eCjx04uxaKLzheo7rSuSQOgEifW8dLaA1B2vgpwGGMLpsM1n4xdSRmOoUKw4
ByD7uej9AFHVpuCIDBaDZo/0+b0ZiGiqAQEJUsod16+ZcwcUQUEHEegcnxc9zp2G
O6e6X5VxEsiJcTMb4q2uIsGU/v92TJd/bLlEctO0iDhhnPwnTA7RwDpIiZubFVVm
CNjknwO/aFMmESctr56ysck2aj8Jrb70aB6TXyc8zHBQHuJVSm1L2V3BnxKxoEo4
nBuLiCSdbO0B3PE6y+xYdftWCttEMEmptNwf+Yc4x5JBJs4hFb4dLcsuMJ/Wcgv3
z1O8q8jpuiqxVJOAVIqmySzrNnjHiKlqeSb/7IzUbUCfQ8x5iSrhwWwbfOAGH+ej
ZxemmoVNNDBXK8v4HEwqEkyvNLLuLpw2itgPxKIlyPrD/oD33W0TheozdI0lxCIy
pawUGn8PUMWl71ZRsUzyCiNSAlfG0tYr1RNEB5/AhCX+hy8oNkpKRY1Thfb71KAT
FShxqiJf0fziGE1ylivFY/hX4dqiyP79CMQG3yUCP2DusU293yr8U0GG19RG2CFw
dWHEoYQsOu3lkGOTWaL/z1IkstsNdyr6fbbuuOMoZVf5uJOpRbhtmWnwTBqqZdex
aDgj2Li1QOtdoXl5R6aeeHLPHOSIX4SQF5bypHop/8KxKA5Ahkmmbp95sy0R4Txy
9Xzt14gN+T4OiGVc/z/R6lksrSHX/CBOgFJAnw5ufmi8ynf6BJpjTNwq9zJr13Zz
hQFQE1uCkll4Q5IMxEPPf5hom7SluN0xwtKXDzro9fQcwEKOatb+7r15fEF8+5Ft
aDn5hQdujj5jmbsoo9rowWPmoSzOQ+SFWZzdBXd2cyTe1m/TIoOsW8Pao/lcqFcO
nRVuhCZGPofmmzyBiPLwi9VwxWuawiT3+6T1QBh4jf6bycTqurPcaTwAG1/Qj8NU
/eA8fMBaKCmSKe/hNFi9Jg/ppPDAR9nfQ+DJ4qwI389fAWSmJEjnETb31glUIJgk
GaOutvvUIeGJMfiTYtvNObprb/7cJ3GBZYXshvw8pgR7qHs++4hNprNlbMIRdQv3
GWf0NCinLLy/UmWmA0gayu5dFfslYa24HBLQSQi5/AP6LAWH2wa0wJRG/eHGI8To
1E9nQi8RHCaaeilEwckCitpvBUBX8T2+3eO0XrR3VgWEzuqPTw8+sclfD+k9YVCA
f1wbU87mBtPxia5ttzAPWIY32uHqpt97kaDvKUoOOLXeK+06WQRQPiuuJMhw+xau
2jfW60o1ErMD1+/K+rYImuvDJK24AsvnWhulXt1AXZVwSqKzBCwHK6TuYPhE+kzG
3CjgYRElaqmz5bDdQIrHEj1HaaAsO7F5RL9YtpV+FVqOcCucR3IKi2hjtlwf2HoV
e777W5aP8oocxdfFZj1ZxzvpbYPPE4ZaX1lF7Pq5O0FLJAGITCiFcd6kso9EqkxA
Jie03K9rPpU+RBo1Dk0ytPiMaW85JNfNkltMvumvP5cH9eJb+ItKDAqI97XJ7hHy
yANgiwkkYU5S5dUtJGh3duCvHp8q83Qe9n1Y612bgAnd0H6h+I/w1FK7eCF8EEY8
+sK+VaoPIt4Cg+jWmXOyPzthD8FtiQbSjqqscMkfHRxVzS7sXECiO9DIqIdNGimo
XTXdjNLHop3fDCIxrEZkBWjgVMprcZB7qiCpkL1+/virslKZN3bTSJsd69QXzOue
ZgNwHEwdzN+ncpPiTK9DTgb7RmYAm4C6248HP+aAGUdqH8Ur9IUaLnGtMU9swAAB
HKxo0SuvDykK7R74E3tmhcaqzDj1n6T4OLgAsBoF4Ql07Ko4U+CDjPjkkpUW9SqN
7O3yCxwNCGjKXigJILrkubB+CR0K52DVwkoB5UeWBqdmVprpvuPvJ8aQOjBlvJkG
6EmpYl+oHLk5vFimulUpFtjbs/bIOCjjG38+sn+gM3kaaLabaNKrfD9/AnNt4MOk
4+UeTfFmsVP0GomY4bLMcNGeLtWdP1mkiFCNKBvT/5Kq35pOXFauQc47+gY2rzEg
WMA1/ylbMbEz/hNyDxyntV/2a4PTypmrB9NeUkOY2aI8Ekun40AC89sTRK0WYb3q
vqenBF+g2bsTWM4NqQzLPlyrXsW/2/flxxdOSqhAC1R3Jl81C59fVFryaSwFbSxN
zopoNwldETrAnPoC5nx2vdBuA6tvi3uVZpdeQiuFqKQ1NdhZb2RfOPj8MPCycz6F
E6RWyfsKj6mWL87KpwcnalH+tiIKc8sfTMuDjGaU3gTZITFAj8JNN3a1XbNoIRyM
FKEz7j+jJLFNMrCjCQCl8OPH4UX6zezMbmJ+w8sVKqYbLtR1KlFhPT+TqLZSw/R5
jujdZyZHsCf3t8jwYe0xVFymH9Ph+wbZaeyOT/8Z8odXpkE4nlYq3Mo37Bh47pKW
RbqapC/+KL1xhcB0Qy7izGV9Xa/OzmTx3suK3KqCHx4ZCivBzKf70eL4nLj3uxYm
SedQ0oBZouiHVZeSJey/2T4oWMw+0jjKRTp73gETujfebZ7fQx+BVmm/v8Y/6qpy
FnXVNNtbfn7ulMUk9iyXqOk/Z4Vvafl8s0gLNm8P4SOCh9zkfTq2aba5qqJdEF5g
iYKJKpeO1+eKOumpHS+7l+4swb/WfeJL0ti9+6OXj1X74OLqCYee2QvkbKjuO8Ab
oqiE9F0icNYMrWcxlAYC7l6GqQ5RehLXBuhWGpZeo1HMf6xwooDTxMzozwQzrIKI
YjJCOYNQA2LyxLCiyzpCvSQppoA2YlZf2dSZkUqASb+8DdxP9sOLGUww9ysxZyco
G/mBGuA85W1mA/3iuc9q1d571JJwvKMwGCNiFoO5aOyEsjb9cF6hYgfSTcrIi9NT
zfYyQm1I9wWP0y49DrFJBU8ioQaBUrx0DyN7bCPAxRZyRUaJUTJ0acvY7L2kprfc
+dMgjPNWIw85HXGGf2m+QuNHNmryuPtQzDxL/4iIkgGQjeubUlJi1IsbEW7jR/5c
t3hHzQexXAM7rqR1BpdGZklMmgNHSdeoxytT5yRjdZdp6YIfhEsaZ0g4/PohAHkT
hWgR4UK4b0YMqRP37yhLG9lBUWmCZkMecTT842SPw4PPIQHaiPUEedJ218fsIpt0
ovMwO8ZWtwy+1AS0m1KC74NbeMvBYCz0Twu4GzUZUtmuhP28DhyZRMUat5A9Md0k
oA/bHZTa8w0vxHylde3ASmKdXYnQwLGNnZ7UtVrgXWcEwOOBzrnD99jJh0jQBHOT
8bOluR6vUfv6fWdafB7vyhxvNXctfoku+iTPFSas1cJHxi9Gju2wCaW3TY3cJtqv
CpXYmkk+KN3Gp3T/aG6qRVPaxo/VkjW0zOoxihW86V1GOPiP441/vjcibkLJZBC2
6IPAkLn1d+tkmreOcs8Nj6Nh0G/X87WjLOhdca5+RVRq060i4vFpJ4JRo01yooHS
xXbcCblAWui4md+s1P710Cd9M++4MC4rIGi9/LCYefqBiIPWKQLrCfiTqVlq7JcC
OYCMnGNW3iQ4BJLpQZzOdU/VnSH5yBzjfZPdu3bj7fpPcnqmtLXngOU7XfMXQg3V
VzkNSpFOsCucC+mYo2Bu7RCCi3ApdBcq7jyISWn3upgq4a1iGO8uncxeHItGfosn
1/sF7zIO2ehi+9k7mw4wfHbtWtowlf8wbMh5hEkULgjmUmOcWu3E1W4wNt08/+Gq
4c9zTJCJ1ngosq3YeY9eFl95Wn200ThIvpQVZxCoUpd/+SgYJocBaxbqCsFbju8b
oIZDT2c3k9LDWS5D31LAZ7rZQ0rZYC2H0LCMIys6e4o6QJS+Y4lJ0GhLfXw0ZrdC
uiNHqM7YsgwRjrYuDFAWvzu5FspjrqkkdS5M7kCHDlR57bxJ9Y1l2/dEG4dma8tP
IuckAi4PpXfeYbpFcQEdJMs49qUfuv9X5joGhbl01jK+PKrecnQE4OpRzLiji3AK
iaHu2Y/eq3bo5wsa6GAK+X6oSu9OIjnC3GK6IXbfM4D7R53Kb/hnPm2iNfqjoa/Z
V0OYTgbQ0pFI3A8gCdNbmpW8dv4+ilQL/VFFMItKUkty3DdNKF9qZvvEIqA+UR1y
Vqc/g2tVf7TBhpvBXMbYt5GRFEpR/Cu+cgF+fUAxkp1dhkiMdi8iHfrIr2+x3zkE
gB01elf7inEpWxrtCfJzekFVcEHP0T+pavQbIUORBCYZIfy/hKcL/29IfYBUVv+V
FgjbjVSffnfu56eGFrrzuauLi30f/Fss0QOI9mXeoc+PnFFw+qTe1ZkdWJeTORtp
vB7Gu4IhGGlasgdvojrH3AIT8eeJc/I23KPMVZqtCGQD4IQKSbexUk0zWPj3s/ye
2xbdCjByAMJH9Bk88TrPZkhsPoeRub+odVBhjI6tfauIclNZl4eOoNc4eGHuqzpA
sudBHpqSD8xq8ORK5315So/KJzS9HTmcITCXEPDnsupf0R1dcP76sDVHYql2Q53q
fuLIH1GbGWLIMj6EX7N6Oea+mDqddSUUXXr8iYjqVyP7xyC+z5Hc87YBvExEflXk
OIFeaRXtlLGsP1XLj0cl29dQrCRkzoDHCalv8mnATUMOvCefJmRjNwoxKRFH3gMO
kk46g5fj8FoV2+nQj2EUAILwXkCyXntU+jWXHEuLgZ7KxwKyjng9P1dPlJnDRP0r
pNjwTD+ep3UWdYt77lelYO4T+RPzd5lMXA8Kew0Zc+3aCXPODt2BcxpJWtGplwea
SFrkAcWa9GAsngAYFSDyfsq1qdFTNGp+5H3P7/DSdBaguWxy5J+wP0OYuIOEx8rr
LYT9ribgWrK1TaC4p8WR64MzCQ98SjUvasDyi25wLyY98hCQUib4yFkvcES+jiHt
WiN554/tdcdi06iQT2FPgWKx7iux5aYu2nQaXiLrV0sy/uwykoScolLfpuMO4JNH
VuxsX/ZJnZPqLYS8Hz/JivCcROaJmowH0eIH0fH2diQHAZ5cLaam/mxCNspTg6aZ
15bhL9JItb7C0MXHRtDdL++dCeWGj53D468cdtUP6s03/P3i0mdMGHKZ0URWjpab
+6tv4HVVTmjfIEafpweoSZ788CX2aHcGMjEJSUuJUj6ZzGJ9wsJiOtjW5CUFxvlw
b+iHsZ0YyO1n+hR1iMqGFV0Gvnq2gdWemOTG2eXf4rfHY1l2XJwc7HRaRGIOsfzI
ZnGMWkTqiq/cl/YQZas4JMnl/Hmfy1Kqu7aPqCaeCXvxSjk7P7xhvge83DuqwLVP
tMvMgpQ9kDrbWpkWMSpWwg15aYvXo5/F1OgkNHNgTtKlHBTF+9q4xIze2VB2Bw3G
yWtKLdR80HKHX0gLaMXM6Zk8lshE3vJ+SGc5CIABk7zThd98wbAidg/bOvsd/uUo
EDoqgANwVrL1Zv+a7mSDPn4uMGa+CqgjcPFBsjHT5H+oiLQSONuSyuvADt5/OjnH
ryW8wjWdJZC4b2mJJDEMTaaUE9j2jcWcCrilStVTSHDzZ6qzBqj6iDSXmYOzF3rz
Iuu9NpAy6cVgS6CKucQS0m+H8NNkuHIVoheogtXfK7B6S67Ivwkf8OPUB6QnjzUF
PeyXmTBHPHMGF3Dx6JEe2NVtEUssiKKAtzvx+q/87mvXVDXSYIq7cWnWSfkFSTd6
PVjUP9MnOAoP+Mdo5FmX8YW8ZRrpb7ZGVkuITBk1AQ0tAX06RX6TvrXmF+L/pSRo
lBpDQUAWiAAJ7eLfqxEnuhhtf7Gy8ZUOzHRPIlOD5JIcKr+QZD8XaDDRJwAVMXos
0E5wapb1kBRAd9NMmhRuD+Y4Qjd5+76aDYh3EEacAPAEyHIgjm+TzcGwOPX+Qtwi
Qtw0SNsGcNcb/wouBnXQZDlREi9WjDwqr6gcbawaA8nnv1A8ho5Nc32dhiEmRoUM
WganGvTKYi4Wl/r5AfXQtYbas3Ehq5zIkmByaVDKd82LQgCzHV2uCx5rtFjvTRmr
t5ytx3rnglkltUnrCwVISf1iM9OdMzatUpkP8VmvlSZ6qoL+MSceXfGoMXHo/ctn
jtpYrKgr3pgfqzUwIdNmdwSZ/9Jg2VMLfNraCGiFIOqsqBdDe3jG5lx+VTkH8/9j
ioyV73vlhkW9ipV49mTJgLNeJl7fuTLKtyKKAJ4ieIGMzexHZApOjiBfdGLJi74Z
1TQV2BlS6xgXv9kzGVZpyf6lIxKb0XdBXR3YzqVYyRCWyUfW68nouvbhq1fbItgV
qG/m64PLb5Lr4VZ5JyopYD+3U+38XYtwTgYm4reDqtijRvU/znKTrr8vSL1Jd4Nw
GrioYwOgPAlCLY29XB7ppHFICM2gX/BfE4jml0T7iQrGx0IONpEBevGnR/L8/bWg
h+lVDl/Twc2u3m0B92SWDcEx5ugMul4BO+PPGx+7LJGdZbM/2sHgJW/ovqpRDuDE
2P4V2I0zc/vUSw4Yt6gJeVuLD366g431NZ3tHXMHc18uwvPNkpsT8VmopKC6W5kE
PSFUom3gRFLaEsGScxajhomSNvk6OVa+ntuqEBNzrYAo7DOdFRH52uzX4TcWzCyN
Awuiln8iG9hpTkm0HFs6SGNEz/xqAfxvszXvxxmKal/eEezZAxZRuBrvMMrzGvyc
zQH1M1+sZwv2XTQi4cNTJzBYOJd8H2idbDjjOGYYbFPCJbhoH2vJ8WDCtXjkEOei
p3aMUyJYVTKdfEzyLFXbyLosBzaVLNSAgKOhH6OlX3tM3b0EGL/gePv16SHgS/rS
2+Nkepz4sqQHI21FBu/LgADQQ8V1NhvsZTss+xJqd2FJ6kKJkODzGUj98Osny4vl
NPqMidPIAp/qBwuUtXyXFQv0yMK8dc34fsuPkdnPeMDrlHjc1QY72TitShGuoYy1
UClxWfNd3eFGeCuWbml31cuiEqlrmFw7bMxOG3/4VTwi6TSgYZKbEZsKSvnD4p9f
vrgLd5d56IjRzXJPvTL9XddqBU+a6Mgc5UvT8OgWE/+SCXo2/0LC8gQNOaUiiFSh
S1beo4aUVvfDBmztylDQcCVrRE4QYtPLeffDBMmXtOpGJ4ZUV4HPc40F9n3FZB9Z
FfHNLK5eEPIWj+Na+dosz4PoBpNqU+ciAusSYaqcIPnEs//B/BUz5T1Izw2BExti
obFwOKhjphWdK86YRCPbwj16W9OEsh/NIkJHFYR9ePRy/xqB+h8DBsHXv+mBdPr6
XZC26BUaDJD+bj3I2O2Dzpz9MV6LWw5GhxWvPvjZQEgTp/ao9zLBgQdrJJhgBUgK
6IpBUn3nVAW+Hlu/thFBPtMuNGD0cC3KlpxIbTz5Hszn06proXb67RSDlDFksigJ
w7wPdCXPhA0Ibbg2/LNKXtOnz1nVsjZUKDG3qGoDPy+DkDOXN5vB7IrdoL3mYbcb
lUNcSy1T0BKkqFf7Lqtj5aGTsJOYhDJCJo1H2feJIWH1smcu1IaEvaF/O+u9z1DY
GdPiUW983251bTqALEQFTf2Wj82z0TQ+2bLEaEyG6QP73c5PNp0LmPGAXYNDlX3Q
9esTqdgZMTFy/Dh2kFYqePqRC3ogX5oU9j4MzMw3eDuKse0gMulbZaKRVt7MHVsf
2p112vOrWugk4g4NlCDGa7butH9T7EAm83YwjsQ0mMJGWoTSOBcXCq2dZqjvsZ4K
ruR02RoMdvS7sZ10ttgdaYmV+B+wTpg8pAxhkv1qRkiCajL9y9nqt4umHrfP8aP4
rYHb2gME5WZOZ9/mWoFeokDDWLCjYIzUVaGD8CbeFffVbSMXaTNWLfEtAZeq0C59
Qg2OXiTMWLa495FzsC9a/O0ljJk7/Z3rNAGtaQhJFpQsHoGc9AMRPomyvis2ev8q
o79TmpZzF2K8w1in0CJdC1yfY/aD2QmslASKdv6DNk76sTzhC0fkvKr/foYb69yq
UbAzjnPUIlAKN5VunLAlUex59Yixp2H08bjnssRMUNMgc8dBh9zqIzlj6pemcKZb
tXfhz25w15CJmGSdNbIg4B7mUbrRv4dF9REwU25LhSeRYFnSJqGT4R3wCknIL0cm
DLpcz4z5HJXeugrWGP54Zwsx7kO26BjZu3VOvjPJFtfyIG3KGhpEg8yBPIVu/m6O
E5ezTXOG33GAw/79TnGfAzvJ3p+DwH4X654FyNH9CPHBbayZQoBFtk7wn0JCevig
9rG+oqF2CZZXvbKgOlaDEUsRG9oflYAOZP+VyE0Tj0/SD3uPpLcwM/oTTo048zia
Pw8aFG49yjHI22oDcTsubFXljjbHpsNs1UUnT4UnRHqQe/BVUWejybrvMlq8v2SA
AU6mn38Oy98NJCm/KZQ5YDJ3B4i/11sRPICHhcgLdpeRyZHUKg/8KYvBt4oZcLFs
p4afb5VbgqLCnCpdtVrB2yR4eerkatxcEmbkAAKTFdhpWKRXUqZmhiFLGRi0BeOe
hXucCBkvbakwkWxLUO/aURp0GLD4p3qENkt/SLEC/DM/ar4Ip6hEA8xMNq/iu5yU
JWR8DDZrsZnHmZ5V2bINti3tFwiWSjJttMXoLxztlileNJ1v2KnyTX8rBgZ1Iw+W
MoN1sDX7vx1vaZVXXdVcrJdK9j6Gq30Rck2vsH9+OhWoNbmcyra6Jdc/GeMxQ7cZ
A8+CdEC2bEIzAlBHo+Z0BSjJ+KDA3EvXwUnW7xItT4E40o6tiho2csSmkeKNsiKf
bfNs9VPPYGtRpACCYuUrCCxg/LmxuVwH0W6ErX4sD+KjsuPT0vAlZA/Ay9eA21gS
tbA682ghmvEEkA/dyNO3z1oSokAKI/4ofPFfHoOxrqkfaYSlf72Jke9vWeNq3VHd
MqIuDkeBRfXEWeoheILb0Thb2hE6HJ3fSaLyqnnRJbHCxMam7ve49/kggUCaU5DZ
CaJlvCwL+QYSKPAOAe3BP/IE2TDsj+pB5QyhksqA7PKBxSkLD+Y9jE4+8UinAcOh
8H9WiJd8H2hcQNc43cb51Vtaum6F8qcOATfNHkFVLNerxg6t0aSr0KoM8+7GFMfD
cEeIyioLa4kpZ1C9PwH+L05QIVMkjXpj72rrOLqkc5jgQQuTAvZ4fotWKLvHesxL
4ETOsbbbcOXq4c5MxF7Y/Km6Sj0by5JhUfUbiHRpgv+ZQuEVd8y6OoPM4dpAI4ST
bp/XsdjlVjLQM3TF/K2a1nt5Tgfnw8PqMoN7mY93TD/qug1L8vDC/y3K0rWCF/5s
XeDWVctJ31YubcG/QGrbkOzH9Y+ePhCchGmTgFp9IhPpF3v++Pf78KgCQ65H45UM
sfHxfjkNA1cHLghNMg/Q3G9z/LDh2fcr1f2jSclVtJi6zDn05k0jkW7LKN4SFN6Q
Xo/7Xu4g/euUdZk/sTDSMUO6v2wA7yFQBW1g90pHbtFqC6EC+/E/IKLr2uxttM2h
3igJmpiR7sY3ElWNgTMTmqEXZaX62Kepw5gQQ5KNY/m5Q2rBx59va/83uZNztZyM
uid5ywstu2niVyjUXTWIo4mBsDtK7eJB1TAb1SPl+FzK86AIgUPKw/Jd4bpwZqBB
PpC0jh2o6+1hGoDU9cq+dGzIjMWyFNGtv6Dicckuluy6y1Yj+Jtp8u0DXEPIoILw
IqVAMPB5pCJEIxr7SZcQ7/axQWZIH4fOEjzokklWfewhEHDjtlI3HkfbS0UeAdya
+ZljjLLj3bxlCUEyyLkbmktXZ/+LIHjGBO3qX5muCc3KGOdWQSsy/Iev1SsK8n9y
3u/UNVJQWqz825ljrlYpX0vFPbro/+KZJM/UPJ9ecgpsfBmEOA7bE0tzVGqHObR+
x5p+3RH0m1VgO3oBd5dNodgl2Kmb8fE0XwNYKd9cOrwLs2+XaKx8SdYjetk0TROF
nJGl/BHuP01Wv8CS9zMcu2+2KtcEpzDoHzJ66IUZOyBJvI8RzO9zOZmsn3f7WRi6
nJ/MyRZPmIHZCjrxTlNqo6Izo9DHK4e1rCjXOHXGUnCpGAAgUkt2YnB9U+fYBvwi
ApJyXN0n17Yt9x8YZyfwojncF91dsVczGuZu8+vU9+Vp8/ybNbdoHm6JwZVdNmsX
6+qRloqot8GVKKgZbDKXkO24/jg0pVbHdQFf9bM7nHEmDWAsbaH6S0lX8NkxekCr
noB9SiQWOOYNndW9/AftxLswSkjKIwVwTzy7yvxOBkROVz2iK6IgjME4AzBkVnbq
vBA75DdQ1WFu8RaAfDZazCl/fw+4SBMLqCcNdt7fd7fnI1OiYarog3svmLVPRRkt
gH6Xl7r34JfsaMx1p+vXHtVZwFzAb6ftLVX3P2U7COXIgOUTOgw/0vFPJ+VqwPri
m3FEW6ksRZ3gPOf6NOKxEoVBpSLECPETh70v13/qBD+pG+qAgmBUYWGPxdPHNKCn
9x9M6rj5pIgLX7yw63iZUUExR1mqL1R+2YPkiV6S5aBTLCo7wXXue7cilhvCtv7B
ykzbJmSCCmJPZ7MbvM1TxeU+8JOxoVG/fl1i1ANyB4ocpp8wrB3ceOicJ8MTvkYO
p0B12d3RBXhfkB9MQ/4siUdzBajG49jXWRwItQZF6G3oW4bYVJq8kLXln2ZbmlgM
B8DKO3Mrde1qFpagRf4xiucpaOzwDGODr7VshVvIndr0PccJthBn0W3CEU+4tq/F
w/xU8NzksCWp+NbVUQaFZpiuL+0M9NjuAvWPp8/jWsTp85Hd7Ce4NQ3rfIE/J3Tc
hS5UvEERfjLlUgSBQEuZ5Opas1TQOPtPLPQ6Q2O0JFCuDJ6W/EMXq/0NXxDXtE0B
n0RE0uJT4xXQX6tonlm/vw+Yef7wC5uKp4RDGiCNYmYc4/n7SmbH2gYRUMhXxxkE
LXV1YQBILlv6LTD8tdvidtB1gcJkbGpq04K11iz6k5gDRRO0dFVfNsLpKt+OZ3/X
xXmUTYeJ/dwYnfqbdKT0KdeHIedL7jM0pqbZeypff4S/ct40eGL9gqgYVhevV9Nq
AISMgFSU6ZAoOmcsCUKccIkdB7oUitJmw7mzeDnsP5wSpn0TXb1lSdoisPqoYTTi
dDBuUdtlcBw042NX6Oae3ePDUqDFo5JN5C7AMatp5ClIRUNihAchNS9yQNl5M2iq
/z4xQt2t4ME6Z/Z1YxZeEG+scAufL8d0WxLCPC18kQx/TlqmRn8q1rRoM4zwbOle
2i2U+fcOmmHjW2IH1rmLeH9MuVn3XzOH7iUAZvuGcLJ4PjcMc4mvfOQ/e6KGMoGk
fBku1+az8kp7y5swtUECR53/Dkspiiu5FJBSVHhpNr87xnftgzbxcyfdszVpqW5W
WJru1jPiM4Vl0OR2OUk1P3mOMwLBqmI6leHC26z58GSTTURs1UeLrxyFi+l4Cpl6
ZrlvbMsgTKnjiGP4tauo7HU7Y/2u+xGAuWFTYs0jutZMtFOyDUOePL1LLCPJo6tH
2vP2556/XqCdDYdjqpfoyIyimFP4vRKfI+BxKp0jfVYwTWZgpX5+ge9UKfji9HAf
8VwVPgJMEyrZQTqmdnFWg1SjVFPEDKFbNO2+Q67SYGQYbwgInVGA98BNmZrqNhbp
tMDjP9X0TP8Yb82R90LV/JCrTVCzkeZaELIRBWApC0a4RwZ39L4Zke9geM55EPEb
+e8yhQ/ggIdoB4diIwb3aMytJcX9lQe+imz70D9O2cvt+FXrfSuC6PJn7b1fQR/I
lvZ+ooGyILFl3GL597pAVLn9ng5weF+PViWcUDu1UNLW1TNzANEbLHOPYBrm3ia1
qhunvt1HWVeweP2p82Cnc1AdPDUB6DOj1gq7I7Bqp6mZ9VxWwYINV2Fuhlm/bEV1
oYy9TsUxAY+byxelyF6xguhnsaBAqJMbN/88TULcyBiZotFAnpELlBw1eVyVdEY+
2pI5etGqLVISVoKNvcOVc06qHoFlQ5Q4ZlyZf5tigpeXOKDR1oXNppCrOhTU1pyr
yOgdND8CS2ieNiXVRp1DAXJQ8TvkDiwJqq2S9xLB41+K8+hhM6OW6KXME/csk+FW
l2FQYR0E7Vo9VxGyPB8Up0/0KgZTJ34X6u7ZFqUL91SttrouaJParrueIXqGPs5l
HxnGRWPJVfcDPRz/n1zW+TqskNS+oODgnOOf4Nv4ToU+m8waRFjDDgRyj638nj0M
kCglSW2tt5YMt9Heh0wxKXe0dJ9dQ+Y8wTETHjzeKTpzyXKVokY18iTxBnCQxsye
08TPMnTMFslCcNcktaZUzUUYSq/4r9zQPiFXihxFfeIpUCt1K3KOEH6cj1vBl+RD
Its1VkrRmWTsW4euOSzSZxjKegofcsSvav3mCOjxcgN/2PFMDsxaZqoWk+1RlzLH
qkUrJXmNlhe0ebg6ODmy7Hb+WIS5QW6LOD1f7v9xJPUoGDIHnyHsLDiasTlM3FR+
eQJPWzqR16N5KEGTSMlJ/sGDJsD4XyeUmjCfZcxSGkGFCOL2kaEHLEa7Saxhyml4
CRX7pq+uIMK6FCMbZVXAFgRyhkp2tLF7SqFaJ15k/x7aoIA4fiOL1i5HOBJOnEtF
LKB+d9fMJfPAG72pixgEwLrYjVpQLo+UpXpsp6yQq7rVd1sV8ZodfOUiCtEYDnuN
ITPq+CR9Iz0GTryl+GV/4IZI95/eAQNfUk6pmaY4Bmvi9Ft4ev2dFZoxEm3d3oMs
Y9P6NcZC7/mXuULQq8+JsUXH9xdTS5rHBpXYFGPLMwxDTFm6HQUQcxAAa+h+EZE9
fctXgKvQ3DTWo7GoCPVkL8BJRc8+rR+acD/sAuU2VbQLhoBzIbDVNeBjbmzM7mx/
FIdWQ07mL7Db6ET6NB5PqeTo+iphx1N30Gr3DQEtfHf3gPKGcY6KR/bqQulInQYQ
5lVKGVR/z05mJfM/z1E0mMQNZxHrYhK29xJuwFXRMtFY0mX5/3kvbp6++GcBdY/2
ZzGZXf2FtMuUJkmtlttPU9ySMMHtsCxXZRRHtzBtQ/1cCIIPlAgbVjV1zGF/iVJ2
H78M8pL1pFPiIOIrs0aD3wktqDwLUcR3e4p4pzvyc3CWJazqVpM13aH39o09thCN
mvQ6IirQ19rKhNhltju2DUKbd5PC7DrHgM9UcEPzIhFWeDHfIEcHiyMHd2SkgDQq
CaVGNrMKthdG9OAG+9kFGMoTKxR1rkwKY5KCUCVkHDe1wZOMvJl7t1YyghKeZrzG
Vxqz8k0e58B8hWBGdOZ93F6gyOuDmtHEsG2zj3ymquXIfkRujtRhzDt6DmRfhYPP
8ITREJX7Byl15U80ekpttgDr8dMDOTP4yHowN1+QUUfadGeZrBrJzxEkO2BKa+Rm
tQa1ZbE/azEVZOlyqJF9CFTteQTJwOI6+U7s2fQ0fCd1+rvLgl0x9mSiPreGXWDj
HSbu317oZsGRtDs3vILFFMctfcgMouy058VEfC4IONwDNJZHTlF/ueeGgXmOWRm7
9jSAazlyOWL3VTX8/3Nm1SJzUuIJtM9vJSnZcv5Aj9yxK6t+rstz8LNOBZjQW3B9
WN86hdD1MiD/iO136X4nvn9cC72pIkz1p29sS96Jps1TGllSiMHyK2iKlUuCTnJl
N0yIBKZh6sNB7JxMwPjiJGJ6htFVTVOnp/YAUEvHQTaGy52F5mHNRDYJ00C3Q5Dk
XfRblmR6EbTdbcTf2YHy42y5lywLvzFFnfNIZ6oI3JjBsAOHVkBd/XJdLkVIhYSq
qQhfA6QGj4sM5K5y0DU4Idsb92iEfJlApSrvQeKJ3UJ3k060DI5k7oSSSwSzokue
PqozHjFU3stlVDacP+hsgkoVXGvxDm2N7JN1OuIpI2f/9fE+bAiluL+U7TAtaqzj
WbyjiLMJS677/f60dD8j3uiXFZbGOwDYgYjawKIg89fs2UGMGDJaiveLJr88L5xr
g3ygikXIJrcyI6kDCvQGckA0TYi7QgqMmh4FMD0oCi5xpphrC9S9YCS0SUI48svh
Iik28VQq8FVxOAXn6hNWYv3I3PGBhOjtu3Hnh+qoSGa28PRA0MhBy7JbfEpZ3C4L
78ObKyVGAw7TLeZHDIPOG+FYmpsuxifIPZ9LnaFm5advIjpxeRXXSBCD8edyWFmM
0IvjXaB8Du/UH9zfNQB4E8OeCtAFtWHG4RpcPyVCT21I9moRW6Sm6yOtMCWic1kN
QbhJhXKf7igW0/7Hqsp7SQ8bNcVoyPdZrQYwHiEeDkTPgsqS8k3hSQWZ5SdK7TMs
sCqJofEYSfd0JPDHjgppjP5RZKzSv9OFp0yDIBde7JWOGLPMLJu458rCbOmU0mRo
zVOIzdxIiJHb1AjBJsyPPfwpO5WY4T5yywIGEVpmWEOBKvuGiLavAbPRWuzAqamn
wiU4wq4LR8a8iYTzikc8c1/DdsckRdXpvPA51exJYcYP8kpY8slpjXJ0wk+auGBv
4LFcl9RVsXXETxDhsYcwdqbcOtstJGrxSlfgLNEYk9yJlvY4oqaAZoM4VWypifAv
uEwopldfnfB5rUW+/pORbdhyQhefNxO6EXllKYNboGa1b7s3JK9dx5HLv2EhZdBz
vMwW3DkfDHQ017426vuau3PGWzlMCbP0rhlSY3T3AjA/SK28vpiECHBeGfWdOyKh
6Bj68B2lq05osn7yX1kzSpVLuQOqw6835SSaOta2d6/bSwv1sCs65JL01R8QSzIG
yhtAZjXXUXpyJLjqmrxR036BVpfLlx517PNnBGvrS7qfZm9IJO33jRvwWrxJZUIz
R7z/MFzGc2Famo2Eulj3oLGReezNopot5824K5sNI4wkvjrnViJKofu8i50qLaOb
zNDhe8I3Za+6Rhf2kQG+UbHAdcKjl+Xvy2aSu00Mdkrx9bj8xrG5oy1eVQmIRy5t
ljJnMSy7MNVQ0PAmnK2NHMMEoGej2K41opbH4F/UH8JAvNr4SMyfkoXyS5bDb1uK
tqpdfFZXIwqu4yuqMWUeAtYv0Rl7CRQ9l8PoiZV+KGSQrESq1KYQQ1V1N2BVaWTZ
IKfEQ3KQ21wqAsdFXCsew2O1AA2NDuGh4zT7xNwZg9vFPu92hMTJyza0ZD9n8sRJ
CE+YXKZmER3UCzQ7sVrJiQHrBX6XzOH2TvdXaA8hOXFS2PJRNaEIiCqPBlASUmC6
vznsX2xlKO7PQHgqqDvFmlj7/8QD++/Q35LI8Y8tRfjwjTK/5DrFfDOr4hrgvWJs
NF1YZ5TXaeWLh6vt4z2zYU01yZ1MTlfUYZRxTJyQ/+bKPY/+6aVYMT8uRgoNEj5+
R4q0vc5IgipUSZdA/BI8U589fb8ytsitCD5tgpQ7xz2oRM8I9djfme4Bng2kQgk9
p2MyJqFNPwVm/ik6nWznAUGX551tJkmTJ++tR3u77OZKSv+GrrKBGwos1whidcKi
9Hf/7H+8cvA39oXLbKsUeU6YvXPP1rQstuVfClGBuop8q4xG//wRvteI1dyyTc51
YB76L+Fr0rOe5GvwuCsQBmY69/0pT64Rg/UhFCetcC0n+PD30sdXaVT8r6dTzfuk
+yGHZ+KsOFqjYJ4jX3KKC3ewY0btsYhOKZpldOZN71OxxRAG9D7e071mmpAvfhdN
lYKESJmd/i0kmCpTD2ejybIpOZRloyXOBNKC2tzSsJRe/xvcX+gZ+9t+5vzTo+ut
bzQ1e8eXNnrdd4fhkPEUiii+zQ4Pr0ubMtfZJocZXfzzTwOzMUn7BoTJfnhgEakP
/h2X5ZC1xI+5yPZGuwXvVNFjQ9NZk/RBtPSN/egL4Hl1mVw2Kkw1iMcoDe9BRMjB
PLaVwuYixP3PlGlmUFB2dE0QtM8+MbFxwETn5QpIqN7sa0N6NwXfjoZgeqj54GJ2
pEfuM1VhySzPRpF+cqXVEA8BqiDpy6ZNjjOXJaMWrAuLSrx4DIFo3koxLeE2BjE9
2Smzx69cXzpBQfWXYlVEe0QEBPA3hHfci6iiRKQ+vlDTB8seb+IbWaTOq8x/EczH
K8kWlqakW7FMi8k1+dcPsdfxKir0J5ooDGc4PgNrQkv/0WmOX789kdrfKYHgDEI8
6wfMyS8OGetWbXDfIdfYo1AHztk5xAlSSe+Q12dv4jg7qMueTFAmSLkiZgi8uSoO
NBcbSMQh4Ba0faPsq67H8oerJrmlSuOqZas+FmjWXEKZlv4psz+RQ+tvNWoKkMI3
S3D4ynqdUS9TB/u12665ikHvxNkDmYrwK2INLijwYkSkTG8KXckXHcOkNUDBlKkw
fNUqKpxsO0BECfk+QRTyg+pa5Bq8jpoFHbICQEb9uf38kXMoKOJxROeGWruu2Vq1
lzKmM/T3i1egcFFPuoPHVpRg7Ke1nR481TolUNOKP1T31wo8Wdhh5gOGrMEW7/Qe
FSzTiivfEBMWXQrZSzvJOcAv9JNBBYPqzg1RygfVtDG+oxjG2HYwKN4TPUqPRAyx
W+o/OBwLpV8ZiQQ6j1s4oDp4ENK6bT/GfCAEJkSCR0DY71nyLkK0h2/MoP1PLC/0
9uWd2WLvIK4Csp0qoQz7Yllq/v+PKl3pFLQA3PqvGpZGkJVlo2ox/UfWYqni62iA
Hr01Deq4kB3TXL3P7XC4/JZ70SghiqYZ1IGZajaDrTjZkkUrmowsJHAojca9MxQ3
vgHq+SEZvfY8bDxQHBvtG6lCGAAAHK15zzW5EV8d3Wxq2LAhq32kwoCaOqVkm0e2
nYDuDy7ltDKqWV3nuJs6PrXL2CqDLL4WDwa0PuQE3IYXT/L5bNaNjuQDTqal4Nft
qBWpl10jYkvpox04eYehrg3a1k5J09Y4Cjol0ziC1QHVPeXb532zPgXkqL6s74hi
6BDSBPfDYBhC5q/dbfQycII4J6myRgkJ2LWKZBbu82NnTfTrCD86o+th3c76r0tu
S5SuD9t3rQUKHRZ5SDKnEIvc3I3k4ZpVaEsTfeP/dWXbxfF8VMr9Wdn9u1XFbBxj
wB91G/uDM39HmHKkfnyyxMJT2AELVwA4QaNwMacbkyTyaPqlOs1/H226XLMWczUX
vXGlsZUVyVgrI6+PYMBLVjEzAopNPFgd8Dwgx+dkBSW4vLuHLPfm2rXb2EPFx5H+
ZAdI8tnhCWzYm3pQqd1mwwU6a1yaNmfnHILYbTbojh9opm4n3zeXsNQWghOVigAp
fR+OAH/1rkXthYlsIsx2iG9y4hQOCQrt5jYmih60D0yooHi5MqTZ4AxB+TialjCg
mAX2chAjr7w6/221Sj8DtX8srs8AMAMs/Xt/QGC/6QLAtInryLiF1ArQJuZo3u8f
tmY/4j4qER7IFDsLMWbLzlVptaRnLp5I2rUI6cN8UamlKqRKP1tMVTJkm8kBALBx
SMGy/AbdJfX7zBB88wEPIK5WkwLfAExxlxs3SOc8eURMMSLGDY45Lzd08g//mvQj
inD9iCy/bKV89R97MnQ/W1dclZYS/LBxIJnhDwiy8cR6nGYjQg57tRw/VSBzpPMy
E2NL1vM9Lrny6px6/a4aQIwUOuxEqGkjIaguR0oFUQkvWFoUhX3BMqkUYXx6PSvB
IV5Tj3eyPT+SzzD0/jaI7TxS31rcbLAioRalcRb6I3ZElIuE5OLkI8knghz/ddsN
aaGa0R9uIKBEI5W2QYAPfWVroPBEJy4hEOx8seiIahOl9rX2v1woTzdM2wLOW/TQ
S3M8erzX1NlsVMO45sSZ2IIayLjNk7SHCGbTX85VG7z0npxCk8GZHYC2z0zxEobO
1H9pEAxqMAfn+em9S0KYzAlIrFPOLzzgSZRo9fFMHgKtxZORn9aHeAFvpXtD/jIE
J4tFdcrk2IXdma24Y30ivIWvKPKqRlU/Vmbo9NPS5YJiHOq5I2ntpAbm08RPcgC+
bVkrqa3RwUdv1GJo5pmLwTTMuP1UpmQeKKY7Gpx4BP1uTC8xBgV3ntX82dEg/oUr
JT1jD++54Yz9iEhJtO/C6StrQ8mtIsbczD3cOVgFhQx6/fY54uucUFZKBdzOc9Xj
+f3AmLHILKuO2C15YdsUrKvnXT/yvjKatzPyAyr68Kfd/++rdL6h9W04qPbror/4
z5hZmUUSBWaPfgL528h2qWxUGctenocUszwIrvnSDbPJbqspEUIZ/Y8P5WUglibQ
d1TJVgSvtf7bZN0U9RNsONkEOlMtUHhsR/gMabjagxpu84X8BWbkf45PWyNGWONW
K8YhfzMXeGo+qIBF/n4eweSiBgEEQ7MDJG54LmE9cTyP8Cyl0gqyMMn484e4BB8y
aKifU8dwrcd8QCs5GGwFgo1ZAS+UhsEQi7Hr5NYlBd9SGod9ZNiG+dfhxRgpZjhh
srLCwgmoaOE46vg8bYX+kNX+e5Y6NPCU+0m3DRQkiD/gqF6V7c4sEWUZN4PS7uxa
m8N86frcMOqBcaPDP02w/ZaAkiAEnaaq3mfvEMldTQqqXff68zEGvcJaTWytLt27
KGJmM0XxvjohhlAeAr9BNn2uv7IY3k+LooBUwRKxtvWnejhECWU11eN9o2bXLKqs
sFO1B79JEONH7Y/MMfdck6cA1nXgI7CPiyBFsl9UhA6JlqspPzfbZy4xMZQM0/9T
qVbUqbKtnwWR7m+57uQgALoNTOZ/GYbboS+1DU8wYCSfdjJfH8rtBBbnM00u9fWw
YoNJVu4spKvEPKpIl5A1qPFDfMM0Z0NuNH+EcllSQDs41msZq59Mf/5C54IpbQCx
00j9CcKGeTJ5Ijn79PY8XaKsGFLagawtwBYQreX4xZtPNMvkJljzj0gW0f+8lLDO
kS5E+4S7ZNmteo8i5sqxcnw+nREVhQoGliB5d9Lm5mM7npHP5eNzsZOJIPz4qfu1
hpJooR4loh6cr8kkJDvWnJNoQYMB9cKK7Ci4A6iQiHpJCQR85CaabWfGV3MLkfcm
ut8mWPX5t9LYxxL7sqSTkyhlHn4SMTiAFz+MCpW4+bO2bAQBS2jlKltCnyleeU7c
mwYX4jtCps56hfseyREjKh3W/f+G7yELeW7WscnJJHTxLLH9+n0G7Cvrp5rjJmyL
qaoKqF+ohNPlw2v8we44/9rpyOuk5XB07oLyq/2vp3hXcwOyaCREsiMCCgRibtjb
S39+RY9O2LhLRZmzZN2b7tTCiUC2P/uzYQzpcxdPC/1yJEHx7CAWz9qg81/AQUfb
O2bEX7rNPbI4LOa1pJ7lvsOcgwyRGMAczu285AszxPWn+4gxWK3lChmxZGCPrP+s
uo2EZXjQCsgO4HO4q8spgtpVpDazDbVZZa/QV14AE5Sl7Wb5LsK7GXNFL/P1hi4I
bJUilAkllox5GGLtnRmEK2MyexxJ6sZYjev90PHiBlA9fgsQWw//yKtWhSXpXUc0
muf3lbQRTGfiCvaTsiw8EGbFYAbzSbWCb5yoxLQYokyOKCI4FCIC8m9Bt/yMJdOf
7AGYjtFg6jKjBqaG9OeLc4twmT1JhnnAMGh3+Jo8xZ95CHSlq56uwoSYZiP2r9vw
C3ZEpUbJSg5D/6KWoJNEmDb/7E4jxgXvlOzOH6kDLCd09RvZARve5ewZmXIQsDEv
Qs7UeA2XI/rSyDD+bqL6ENiqJOlr4KOGRkkjPuIGhPbRrvX2nd/yTtQnHIga5HEn
W7JHVeuU/hR21ULLUCC4QhPnZAOrZvInmqPQOojO5PFggBbdBom9NUqWKuskbDi/
ZKAfLzho4Q1xg9BVVUXUOAjRMSe4lNlrHcTn54DrtRvNs15Mt1Vb1eDgVVHJB+o3
aKJI86ZJnI/p9c1bhH5zUFh5qPIY8KKaKBPNKVNdgBlfvWYwJqClxJylNvrkxyE5
ksMbTajCtkX6FFf3f6I4b8F9xcNR1ckj50LmfV3uAXYidHfFeuuBpqRqffzGWk5V
AuJ5ZUFV4haoCra0aWe24iF8iISXRgOCooPj7pXHt3lQSej2WMqNU0w41/xovgm+
BcH05IXM6dMPZ6vqlDEnlEXtuUS4uXmBWVQxeTJA3n8ABa/ZHBgeJ9l9Ya89QCr1
yfhqzs4rWLK5fDmArEKAiapdxuGFbfYwpi0rmOR7dE+vHwx0pW/Cv1dqd3Zr7T26
bPKgb1MGRXTArC/0Wofln1pretJAQMRnc7nOYF4Ph/s+ntm7kDxJsDwooq+dpQnv
7cKn5eT8EdEhHc7y3S28YVEDFY28rd+dr0v4F7ILTjYbSXxCOcYlXArxTgguY0ku
pmvQBPDpZWwfmufFCFmUEbrblqziyZM2q58JHGUbCUjLYPR6tmgrjbwHHb1GDWDK
vdA0uDrse6O6hyGz+PLrBvsypkRrLe0gr3/Ryrrvcjp3ZzuLaq59HEJdomdK2END
CQxFES6e6OQuAZNANluh2bGEYmRUj0BVys0XbLe2fgKuTdMRF0q56JIBlpAtupJd
gMGVNvPENsLCSWdBP+Rm7NsfCpuqFpFiKL3//SpvQkS5+VnAzYDB1Xuych37XWI4
gEBr078EgAm5iIa/cADlCffKBGscxkLxZBVSz4uOCUpc764xUZLq96h1Xjdpfi2o
LT8nrIFwadhVLb3bnHAA+QOpp0lhxdaluoRzgC2Z645vZk7VvxD9nAm9pez8U+j1
1XdiNFnDgwCwN6rKuf32CWRIe99ghDGZRn8+PRFx9iIutMAdeonh7bT7UTo+UDov
A2gdGFHk0OdzV5S7/AhAJOXOCU+w8Y76icsouQtWK7kH7N6WPPJ4bQ+JzTGYJgKD
4YMEwYLUx8hUwtkGvqpqaDuf5z0kZJVOwrK7niXRvZww8rWpV/4TRy15cCqf+vcr
l3+GlyiOMBBjNrhtQMoB2C8qMvxsGkSHjGyrroWsVmZ1DdMHlxK3qWvdraYfmPh6
Z8AotJbr8hDcqbnHV2jpgi9i/WJtbTbhHaNIO+RJK9Fq0wyaoHP9qwbPZW8GjveV
oqoYHIrnqa46eXInBGd0elKuuTzXcTgyF1OZmR+LBJNWXlgsRiQYKb6Wl0UT551H
R2rJWk8cmmld1lQ4JCr8jVr0Y7ojUiK4u+8/+XGwYQ+fDF8XK71kziKdw2z+r7AU
kQzcVAhK10QDc/0cZ8T3CrnE7o5twP++fYDUSJmnxFaBu6ax8n8ai1n67bzSJQn7
vHjNw00a8wAVjLwFqfr111S+9pqQWELy0UKHp15BK/LiRPpANZ5CHe9OyCNUPT6i
pppJJni+DdQWXhzU4zpDwy9h7iboTCNIPEYpkErLrZfFZd6IZH+VimGSU1hPJB5z
YYTTQFq40y+VGx028JYiwKccUHl57VJORRI9rgVJi7PQod14nW+POGUukKUlsa29
WTnOQJZsPrWM9qP8v9VALhYwbCLxGOKSLsVgUCk8goPF6SxdF3LOT9ExKoKk13BB
qZzLKI+tqVnFwuiN/jmlQGG5SRuJcpM+87KmqbyDvOLKQifU1SdFv6MK464v/75H
/HiMpW1+150BwqLtX54U71E7gOvBmuj8GnuBr7h+nCc3/oILkCJBfk7Y2Cuk/Gy2
Wfnw5uXgcezadZ/5HDGPmTEFYhK1TT50iuFRrsOkoEofMT77whVGmbrTk39Dp6BL
szZ7N+OqHP7HJLUaRfIWMABtQFHt6ztm8O4fzWvWOQ1MSCIoEU8eSCXz45VBnbrA
VbX+mgcj0sjldUdbpQ6lnfZONde/A5aASs/GvQw86xBjfaXDbWsb9S4XJJ76SeS9
oyLfyaPZm2/WpNCs2z/mCa2/eE3pu+KwTjHSWPXCw+B3DV0Z7tXaj+DkMGmNMHE3
Ii3kcwTNtu26elOmAYZoKo+uzH8fGJ4C00Mi1CvA3bsGDbWf+V8V+X9P+cG6jh7t
W8vKFNPoa1c6L349g8D7zwLbZAdB+nQrZ6brwZkedn3BqM079k9nDHLbGefm+hSR
/N9Xc/gbLrhPs04dMvXLQnveseoGS8VtYJTMYR2AKYtCZ1TswS7ENbYFqdVl4YLy
3ZWAReu0p95mpBZDiaA+Ghm6YbSTr0UL10J9PXKnygPg964YycAB2PSEMAqMlQiX
sSX3gjD1sYWeislijLTV+/11gPWtKlpSEEYxXWjeGe/2THmQ8nCJFmx+UcM3D5xi
RDgWcFVizlDWPsPcggR7Oo8dBOVbKdNrUbOvnEVQWHHYVBcumlhC7oaWlk1DmbCb
FedGf9jsXjDJESlYKG4jqGUk1lK4adeRN8/ptEqtBncQxod5EXx+bmEQoBHcmdw/
gdRtUxtBNhs5kvRfyWNsvEhi7qzqWh3MMWY/Vlze0baBH+6hwNMGI4xNsMmH0gzS
A3Nv8MF9HNQBM26gwDaZjioTcOaeOQbRG8HbzHc/7dQCm4h1pj1V2f9MNK/iZ25o
njSW3xrhMjkuXSOfEiY7zpRNksCnUnJebFqC6FJDSGjl/unpo8swROCEleSUrAxr
2c9j70rpfCvh+vHhSEP4G/clrTrjW6xrwfwynyTRzO2lbRxPhitL89lRVkcv9adw
5uz6pfpu3sStfaFvhHScpSsL1rSlQ3zR6MMSXOHO/Qzf1ovO4y2/NEhhbU0IRJ4d
xy3BQaW11YOMDBMIbNbQeL7TRXMO6Ye7ok0pLT6f+BJTuX6oOdxPscTvUhFJXZC/
WyCLUMpzyCEbGp7FGKrY48SFZT1f6xgCc7JecwhdKoVtpL7k4+UxRvusfE4DDOXD
8TCyXv18lEIqTC6wNflSeNYInkpyRp/CMYj8ivqDDttAAymdbIUTfrpaHqxniVou
3T7GsCBJxux+nN7GIaD2uJTYLYzF8O4uhnaBhZN60ZFFKHy+yz3iI1XyAjhwUCev
vjbnvs8WYTudxTlIuWTvgcogAZsPN7a+pbi60w9AqAaGBgTarEZNajD5F4KtXA3j
WajfsbznkBYTgWFyQr1ANdUEA2hLjhDOnYXLLEcLSL0Cvx5n31IS5bNp7j90DTAK
zxDd9rIANH1O7q9SeiE4vmSJcdGYFlEG8A8U1+Dr1RqLeP7ZF35U9dL8WlYattwm
3+xFujynnSD6SuDVxmU3WPPt9oYCLEaTrCgEIIPKENjccHToEA8OyaRGA4g2q3Y2
KHVVQDBAV30LnVeW5ENlxkLQyx/cNJBIRAr8ICuiO+9BnaZoG8UnykMt+ENSJ06j
xpGKS86gk7muRkNHmpZiE0CnYZTe6JX+BlJBTcsv8V10QVj0/nFw9npQIuwNCsQf
bNVHJdK8q5iDZ35IT+eJ4+IyTpz+tp+RmXalYZB7fKXZQPShNP0oOTGsAPvc7gzz
AnZO37cFqOKrSROrc/LpIrKe2Vwj9eqiLiZqiaq46yVLd3AdFwYDpS9NLV+BeLhV
5kyqmhaSfvXhx3/Fe4FYiAlNzV5S9XxqSWL9qSrKS4p4tDEoJNabTVMWfhzcN3M8
f1L0S8AwQHNEaderEYYhN2OooR4Z4BgWpAsCd9Su/4DVJ9rbT8qpWlJsMQu86CEJ
IlZBVX9WSFK4fh75duUkaE/lX1vJIyJq/9KN0weV/Eaxe177FZsNG62sFc7pj4qZ
SXLcN7H/Sv3KY+465Y6V5zEAwjx3VEqomnqMl1lZS0p3MoY7zqvK2LNUeZqGqkzA
SlrLoS1vx/piypq/OrwFqOw09h77Gw3vQJFaMRwX5hG9g9nXo9cwWPxW3d9j2w9L
Q/lapWAjeMiLjucztW8HpPKeeLy+6vVrXAy3DXpFcs7o3rlOkjJLUMIP2a7iHn/R
yHbM+om+/uN2gKEbemcPub/bJKEjf6imqQ3HugDF1CgTqMP0jN4w5Cc8ZfQHTw//
y4HsZcTxshSx0o/ICwJVZ/Q2rK/tizZ/vePb6mCk7KTMm+hvgl02aonzoj5/Vb6G
d+8SMAioYkeuKpHgyNMu4enzQPXD2vl0cd6t3EcythRoWapMWnLfPND+vcO8P2uc
EBypKRbnS5tXAyr+RBiZAlGiHCpHvTrWy6IfpXHWY57tZHITgDvkMO6z8JebWsbR
NKglftockHVG4yv7oLnZhTSradh6V8BnbHpOZYOERzxeiwol3iBWcCp+OMRupXXF
TmUfNOXq/bwl+V1C8EeUvcWpIcGqNhoy9ZA2nsWXWVO8PFD6OB5V9TR8ToEAxL5F
qfSl1T/AdI8q0nZ3NqLwnIoW2H8zRNC7k1j4OYKeI4jlPsB/HyU6hR2kn+M7vXO8
WRqWbab0d/yFObINix+XJm5x3JnX6MmLeuN+7U50M5WCvkTGotY/Wqdcy5i9oHBr
59RP5EIzRoPjI+bTWDkrs1nnSnB1TH2W3SyGHlSkJ1Ab6hMsbp33sxrnteYHwGif
Xd14n/SoaXzRDP1h1f82ITNGVe9fFbXzd0Vv0drSbH8jdgvB0Mfeja9hRLjaF9lX
sLXtB9pOaAAG1eFbXGnjg3Xwmkbt3UrsEwcCep30CEwbhl8aPXYzCAeAZKM7YY4P
zmuA1UGehOFlrZSAoR5SZugpuiU/pFxtf6PWJkM+5O9sRuYFAwFVscajFAjQ3Fdu
qD41zQ81UQ0DEUcpAnI84wNTfCgY/0BqZFmcjOWlJ9t34zq77765SAh82AiURCKJ
l89hNPf6KVtlpUz5GgFWGaknYPAb/uMTnviQRqkOxL5y14n+O9LPi6w6APXUtmVt
TJooTdM8VhxFSeNbe+gFVn/cq2TrlgtQKLXT9QeOLCJi4ERMU0c1+G4WrNE3sjcX
Qt66bcQxljX4oW5PP9HNYCe6TYD1qvHhokQjnw+ZynnqrhNBpqXirIN6I0x8UKlz
s4Bw73MhCszfOe/wVw5CmbudBwuw5VZxMqxyFsGk4+D4uq/pLdik/IjRIY5zIkrZ
0SYjfLt+WyXQucAKGHKgXLxcNA+55aR+7IMpbPcWlfehk+DBSzw+xEH3gL0aIbgc
GHRxT8VWnyKYwtUgU+SRkFraEopuYY9S5uRiBRu5PmSXmm+1+yZ7jQL8CryQyX3h
wuMdMLC0Bbj39/WRUSqYiGlCxx5+HEHIV9KzloVzGZ43NpFJ9T38EnnqUry3EFYy
sLLyb62LNmRQXALRWfP5wr+P6NFYzX4vGz5r8114CgeN2kNRrrkiFGUmdFiHzr8p
DfnAHpRjUY9Mwsi90InUkugWlsb4j65TjajJ6mLsOXaQuKuWNL2bzOms3RvyCdYD
yfyMIiavhpOCgbmil+wIZ0sihsPtingkypK0Sz5jl/YtGoj2pinnTwWldKICDuwk
V+a/sfVtKa/eXZxz8gKXimT9efo5uZh7PppK/ZBTfZdrTaFM6ZIgxWdr/dQRKZBl
KPhIGQwHZ3cH4n1T+HNb6yzS97Dh7VAoXIBkElb1aJwxhcWbhH8EvUI/Nkv2Gw8W
FP/AFmK1x/gM1vLxDYiZ57ZkQxKYb4k9iKOkPWa66DSAMphwxEdEFY5DTdhqkoOm
6FoVejeTVkGu4vbDuV2jWyFrbG05gTP2Ig9jED3L2Wgvf4PMitWMllpxTRlKgl0u
XphLR4EuyL9alqST0yYB4P+Jk8mTgGDws26GLl9bymqICYXCXBEF5yMAwqc86Kqf
TbYrZfSzeoaES9RnYVzzHbzHJvwwDzZ8vKQF0BkXgCjA3M+cVfnZ4DW7t3212xZ7
DyS58+c3S2I180K8wkvajUw5RDwROXq1I9/w40nXU9/GdEXpoA0EC+/YqN6FLslT
/OPcKq41Mzf2vGTTDRP7A5xmbAYB5p3KhHkBaD1jElYpC/QAcWN30Du9vYEi557q
yD1Y3jlkzLbn17xLTXhHrzU0Z6OJNWFR0iQiIp3xh7yj+DX4or1Mh07ceIyrkeol
+o5M7brK+9p5tD2QkqtJo2uyemB6eVEeQPz6abLNP2D/mcP8YYPkmevkderuiYxc
b4CpfY4E/8CgemuxHRbZ+oypvICcXuz8j1wH7VwxFEpJp2g0+vOaYQcFyqNVakRU
o++SJASfD2EtZP4fn9tF+AGbOV02zMDEe7f+uohGQiSo5tUHC6xi7ztTjwnZfUbY
MhTpu9knB9dCCYWu7qTJ5PnFp14mY+UqiO5NBvg4fcIdlua8wyEAUSBXgTlK/vW7
UffWHsLMWgEiCVw87XvJsjYPygm8Pi5nhUbhLG4fR+03x1i/S5k6TxCfe7DK+6rm
vUhYNL+fLpaLsjlgadGm5jXWE/nhXlcCi4tV0uac3Ir2OfRt5s3HGTGobmcnt6nV
mANXnEbpiqFXT9j034RPCCS8v+8GPUjapz1qqtCfNcpY4Zfhpnm3ykgpDKONu2Gm
Yt54edvKbRK+0+NBQjsCHaADQD9n+jxXA+JYFGD9PHoINCMoHHoARy6HTY1lq0jl
rhis2BVj54y4W4QXZfn1PWmFBYAgDK4w1OJvO1Hkq2q3HF4IPLqKaIhfV7wFsd9x
IkpQ15PNOfcMkUeGD/hwc57XZ3X7azCxZpVG5iGJMGfG41u7XzJVSdRwGmHBaY5q
vA1GxT84+2fz2DlrceORMAXjLRtZF9her8nDkC19MHbnul4/t4fsFJvQs3nfwO93
QYQUDrWXIhLnMw35oZlKNbvv2cwtRt++GH43qNVQCs2VkVZALQbKun2mcxFULOJ7
qEgo+d2fxyLjTg1qFbDGnWX7SwMPXaDe0gZ8Y/C8l+F+Achp0uivMz7A18pmetvb
FwaVopb9Cpxuq79bcNJAt1uMRk5g1OwpDgqTVu8JqfLfN1GwEoNvVzgMuN3dGPMi
Ly6HtwAiejAUwMYue4hZLBrue4DFVdsDzeg3UIf9578NnJ0qabCGmkL99zBuSLr6
8WWrkKaZoEublsaltHySLJISEmRM+aHEomxdg5eN9OMPS8O8K728A2KO+OYZ68LT
RsjZiEsCdhydeY9eObEz1RBrE/0myAWIAC5jSJ//fjlQ3OJQ7ju+1DR11WK80wTE
15z9RelEj3PhJImEejEOJhC5CBCI4OJTydgebLzaE3qoMYDrpYixStDnCbeYfg6j
pTCkrcBmkPrzlZ+swQNBVWTvM7feJT5jHQcPQBgd55wveOQi4O1+6vAodfBKk83W
8qbXmpWU/6Jt5s9DUkuxZgPzspcCZZ6nNImjtMDpmXUV+hDUq+BwWJc8ZLNXNFBn
hLX2zBq+wjqeKUdx3iOZbFetKK60fS2tSKhYOlrwGgTIMbvwlnppS0RRz6HeSdgf
mj9lXg8YDzFKqWo1OG3FlLBfKjrGk+ZnVkWGuFx5rIrArTzGbpZFBai0eZzixo2m
xSKWpQoJrxKDf34RP3rgLu+1aaGtF6X2ufD+ebqeGennjKKJWjLIYM7mJW5UWQ5W
W2GLAXtxZuS9Dvs/yXukxP/1GR17U6z2oDHvOZRUMDjbdGL0NpqsPMPeEfI5NFDj
hijRxrCj9yOd36IVLXNWI9htQhpEwq6F96fjnFMkmnnxtl6cspTVBiGAZYCIjfpZ
Hyf294CI/7uHGV36AvZE4tt0YjQ1XAYFaxb55F0v4u6PGijQcnU1PpVbGXhIBGey
l3iuz7qrJlukkRlEi+xe9M3bb0nlvFHZqLt4jN/Q/m3H+yvF2l98QzZ2XbLYY1uL
qQi40U1PSyZzN3G5/cCNoEjjByXGdfRLMewOrY6avZexctCLETKeg4RTeYIcryYf
wAG3MJNqOprK19AgVo/Kk2n+L580Zfw14wRCJd9mL1kYkrXQnM755ecSUMGA4DBO
QsVRpI0lrH33O+RIPPplz3M4yX16olBk0kbOGNZ+h8XmNNNvcPA6OXa0bfhVWhzL
xxrxguuIKevcgQWrNcznuHc7C59SBeb3Yqs+i76HEgR9nd+2iLaSGEhIfRTfN5l6
Bumz8kp56pvAm4qLEE9jo9HykExF1TlkUoQKZBB6KrU/C07O/CQRVGsH34GMOP1A
6K7P2em7FKdAOYxO3uOof0flthU6gj2rJde9CdlYxsfIG+nLiglzmgyGqlYjsykC
cy3GpUGJ3aSrNE8Lr9R2rWxSR7wQtt1EQzgztOzV2+nyF+sjFnJC3bR0s4RQzVoS
e11rOv+T6B0NhvhgEiBeggwXC34xQ6NI/b/KsOZrd0N6TAxrYIFEXDNSQuYXol2X
NMwv3bEBZc2DB7R74mPJODIolySSzjV4A4sNMZUfUeViShzIlzIpA+zw50YVEVnq
Z6MiIXv3ckPDzsAp8JHOjWEG/nHrlxKQLMtq+hqYJnJiyxeoHtZpR4UpMISbLK4K
r3x6kkkjcLcWt1Pnsc8PUwdNSoqqESgtNoW9UD+uT39ypVEXbzhrZzZIy2zUlpV/
pYBWrvs8JFjm2HGT7qoCtVrh/QzQBRbSaoqhnZ36sbaSLdHgJWv1rD6sH5NlsqKW
SA1DK4nwrTRCS2H6tmWkQtsSp/zcuzz02i/cKvgck5ctItJybGs/8tBWO6JSz8M8
uIGlF9gZ8sri+CPZWYtr0HmyHdGwuLzl0hYvlHe4jVszMDnGqbuJq64hAu6KKETy
1zfPmmgZJCOVBTzQPRfo3eVT2ImplqYUT4Df2vkCS4CfFXDpMTEQp5JHBd8jRPYH
3wnUsCIG0+7lSra9sSFQQO4ml7jJBqaMTWQJXU4ZW9z6vYGrAmIPNsJUaZiY95tG
UKVYh2rc1thFdIVXpbqSnsJfZppWDwvAHAhlp61dFDz+h0wf3tpT1yZg33XqolHl
VUHrRI53G1xbcN7Vm2Janqyqp3ggIa+/6Ef5n9GcTfgI6iSFpBrzszRi1mLSHNXB
uhSKkIeW4jY7P9WbmWYTjjNYG3OQ/AV8JJW1jcdDr2X4lnExaywFrlrsPu4AmPQC
NjHhC3sY3wM/b2UAs7Or4b5gGx9yYAn5PvINBY3f48dNEgJKfqjsjteDOqYMl6WV
dArkJAJCXHK/MJddBYv0FzH0nfi429Q40GajnbvacV/ziU++8PThmCN9PRUBmldc
CaWjDM96z3qgbZgNk+HcEBuZgd63/cP2IRMCWkitJFz63WLS2PJ3P+lacivFsPNr
1zqATpdLpDTMEy7T3YBfPTMVnokXjIwmNXxmZyVyQfmPkSeWPz4U+e8U7DwVOCDJ
XBar3xkuYMH5Yj4XUFcfzaKUWrUmXf/n5SBs0+5wT3msebayC/cCOEX5MgU4gqN6
KHqKVghF8e8cvds14jgCLrh7YAnZ7KhlhNs0kcO7o6+p9CX62zFbIU+i6OFz8kKW
uSEnQJnx3wAG3lciT8pPhTzk4VgvVcxr6cGKBJrFSskYR6VWQFo2pZ7qekDjLzJR
0w196TBZSeRCS++gvsjeVcnTaLr/r6DN0/dUhTZgugP2B/PP9bfokZdOAFunmiMo
3haLxqyFRzmR+OyYEDjgAdoHT+oLWdggU2efzxMoJDcNgXsDp2EO6pgPgHccxOrN
ixM02cOATABOAgvcYDh5aDbxt61I9gqkeLCNqgbFoFwiVVpVuJI82sJu0Y7TL1du
wR6gNyxN5zpzcDcveiaq/w1RYwEOe8mW8VV17ZqPu06sl9qX4HuWdGuq7FpOUS6C
eMhYqGLlq2LylukiMXIHyb3TJjTMdplEbNmTtqw2t9ktaCz2bjBnXnNjI06pYBBk
LZm6Yikh7q1qwNVcbM0RaEgV4sLXRgi79huHb1PNoal3pOaZh9Oo+uKe1+ffbLba
/8ZsJooZo0GG0pVZhzZFKYbQxwgHIqjnzP2S/e8JVxeahjfVtVsRBya8gtte88IO
7rzknhQXHtHRYv7iJ/3geGfehOvbGDPI4z7VJXuhWOUxF+oiNVnxIeKyYfq7mHnV
JcobnVH19g2jJZ9Hnp+Z3gNVJ86YXP4nCPZlxfZvkKiL/EG3At3R/p+Q8cGVpBfF
B9z8Wqqq0Un+l9lwxTh5LcAmDdhdwGkZjTv7n3dKcQ0uObL9p3XMWRbwg8YzwOCK
mXC4ZNRflBO6WQbKtitG1tX6Kf/My9ANXt2ut0M2UXvyzU5zg9RQjZW/7JEAxrAO
2EVNhgRU+omcaw9yuCceoucvUhtZQIcOVxmAjb/SPS43qm/mEFGL5l9uMvCmKrGH
VcSJswQV59HdZNiu8Yowz+f8OWmtA74v+u2t8gl8WVKu30D3065GOg0xI89oVH0r
evhxRp1+1X+1mRW37l+ONP4dBOvRTSZ2MEz5XZ4qC0U+3f6//xSLebLt7QHqE57p
DT2IfWSRlrEFrgcxbA3qLLU8D4aSHHDOIeQiOa8m6JTkxf2N9UwRS8+3pmJ8gGO6
mDxVfPBnXPXAGbFqJGMlP9DNJ052HKKQXWk4RvuwxUQf02oaTfgv8c3t5rdju++H
5uFegVwiiQ1M5i0TSrldW7KEnHT+puLx85K0Cmd93f4EqQZYxfzc8K24oV0TW/qG
5sHFDu9z5udlkPazVOoi1V1v5+rC+hmVqM9DWDaMlrk9dPCNVevHS32ofU4b/mkc
WP7opR0KveODycFU6M1Lr861YM0XKBwIw0uehygdjHSv7mY7E+W5+XUohH2xdUG+
jd8jNhAQNMjps6+dFI9M7Pt+fxJuoN+OPVL/Cz/2xgoIeaE8MVZmSWD5IRcnnxpB
va3qrUq1zUjBEVbG6tRFokka+BrgIpTeDeLqmDwiTIpNBmq934gB8d0xhIv7Du/e
7630NSGZGnPdhE9oVuJJygpXXSpXuVAh0ZpV0VQSen7FNWLdstPN08N72EevOsoz
8hE64dWSbGrspuZRm8mpvWlItb8R1PihW26oHA+lWhX+7U5GmL4FaIyPyf/B4js7
OjEwxsTqJ9bQC1Jl/Dwv3iePes7bELnnHpQCjZFPOGtOtyPOOYbKp3MpVVXCfE0f
PLd56YdiXilv4v8kiN3cmn4Z95EQfLe0hAnopel2M6WNVQ3HMYTcaMyAudtWsPEF
ppUVNOsFYuJfkAm3e3tUmzCg98dthGK8+E/0+vYkVmDhvioSnPx+a73MjvHByAfQ
/ecczz7tfKu1ABJwLlvnmLg58WZIuFHZkw1Xc8+Jmsf+A8n4aNarV+SyzwMJRRWh
52iJmKI8SaSnZGJdNlkGXs0pwthqzpBUPRqzvp40+zrZoiGcdtok+o7QD+QvJBSs
fVMQRyFS0TAx+C7vo+eQ6KB8aibZqbHkqJ9DKkyu/fW/k3725Wri3cyhOEgr+s6r
auVYeJNgKI5/XqnA2bCz/ltpoxkbBIXf+d63QEvP/AqcuT6RsNbmh1xAw+Cdv6aK
zSb7ui3DbAAd9ja1jQkJeFORiZvhK6+P0muTC0zMZCwPO5oIaDbPlSJQyT4GsAFU
pu6qGAEHpmcIkuAMP4wtVuWJXj0C78HAb/hS+ywRob96PC1cdwp3mbRQL1l9Idle
G7g+WgO7jKIjiyreRdzdaFRACW2GSQgTbTXe1h9EiAVB9JH3HPapREzJciVQMriz
nj9XuHhPYqFNjrV+JnrZnBDBSMfrFJ2hXqjajh3wtraKEoEab1L2/+coI67hFWCx
CPPiamPKM5eth9eGxvvQdzo30H58fPjHhKaLIgP7oj21WXpnhgjm03IAoUZ7iMLU
XbJTwtjyQOGrfJR4M7aJFm4roDtQYGoqkEiUDUbjR2DgR2pBsrz9dRYjyvGqf0xf
lwe2XFqb9niOmY2ghCTsTwMElTAiJ07nryvwE7wl36FJ339kG+wSxkXGYMD7qYOJ
qImvdHLOiu50O1vLSuvyDFkNAXx6FVHR0shNIrpZqoi6F0BqCv3sNYIthYV8HlCI
EtIw22E5OaX6FfqP6mEuO66HT0kw61d5wbal7xbilqVZkrnOpA32Z4hfLrhTOZ4a
OVxrYRREwD2yGpc5sedgL65G2I3srdr2cfN6CPb8hHWTHpS/kdkZetDjj7q89tsm
Lw0DmhhbcWm5wIZyFFaEkZde3CU/7FYz7oT9qGhZ7uDyC+8vTIWQO1rgyJO7UFWR
kTaLaGj/EPlnXOm/CkKBSYMN0O5UoBRdOz/h5fjwR2Xheh8SlH9WrtSEQyoy6kCG
AOzIDu0jUyxjJREBh6G8jBrltBlqaGNXju1zFKwdLW4NBw4CBOcDkS+DBYdtEc3T
vpRWTleyKVDGhZ+Vyp/upKHMGdqSSZc07J2ZuYKQc5e3vwlAN1aHrQwLE4yFepkU
lRGBrkrHIgWhZ6MTOVYClduWmP9+EwS7XLeqCKwd0Takk5tiSFs/QeMc0I8gRhXl
famkEGfencv13gWV9+8Io+q9GGi1oPXF13l3di5q95ljf6V6+KAQTANYnf+Db5lT
1vQ126ElT02Nc4pocf0PImT4drtDd9WJEeZYkkJ5nK5L/6/18SIE+kur77OkXGr/
65NelsqjKh1LQfcxxLUtRAmmqk5d94+syFXjfAg14C0ox9vJzPrOV3k9WmiVrzev
YP3mrXo273lRSU4HX+37l5IZWZ2f94k6OsYvehbQEis2b2U9H8cC/SiIcHCcdxPK
LrMNfOCUjtPXLklb6l8Ft+p4VRkQn+kP0kHBvF1DYvsUIK7fCkjTV7FDBN9CnAMO
mBFDLc8qkQdkIQgRkLoQOmmEVUr0YRI8Tae+Jk87/NNKAi/I5IKkGMnPPVFYICsm
Ia5HIM1wXZt+gUVO79QTP7XGTIWh/oYcPg3bph6AvULZSKHp8wv9MZbDTgeezBK0
HcURwFdC0rXidWhJKLFthihjogGZNAu3Z4TTC1wHdCQhk8ERe/gjUyJ/thzdZpSO
F1MJA0x3JWnQjVgM7ccsxz9mQwJQmcVFFJER90MTphBg9rWQZi2ntT/b3pSFCAs3
SQbJB2V5QldHajkYaYDs8MYerV3R2M9M0tKjTgTpQhNlpKG4whI1UHoC5ueSx3uT
ys+kbi5MnHEo96HMGctXmPzt2+VVhludJm2QXqqwUmzvym4/bT/EHPKO49WP7u6M
D0vD1KgM6xPVnWKhQ/dZL/LFvQraS1QtfoSotJMO1lrPBsNOPi1/zEkoyj37wyas
ZyqgMKTS386JgyC+3X5EFvlzCBn6TTCvdnP6tShVekMvFfXV/xmxdu0yKd+G2QEZ
ffYphuBTXnk97L/qfd/2nJrQePhs3JU6JSx3WVkTWOWMHhG5y3NLtoY0vCGXBJgi
dVZ2jdzKPKHWbvvoCt7U75XDpK/a0rzNupKxZlB77bXzvqUi912PkSMECmvmKBHv
K40CAwXELnKU+Di0rTcgWRbAVvAHwjW8KOmq6OKjwaMF7Qrmx/4ivDrmN/H0FWli
5c/2/jPs1zsp7spbmjDPDAM3Y2dScqgW+qYZopOORNfUZM98Dmyp1xscFZdrK2BV
HNQdtToXLLW/yZUeuskg+XUBUnrmVztlnS/1WweNMceZdq9KWIpUfOl1H1GzphGa
q2hspH2vkzohIlW49kx/1uiG+uMPGUq2i4g09pZq95q9SzKgNDxD8qoEoTlxMQ6S
uLhFdhO0nHUJl0I7m7TXCMf1+WaHulAll+grbv0CMgRENebK5hA0qCNE6xr8zlQO
+KRexzRivFWRPoCA2njx8ahnLbxFf3KgS0yJDSZo2s5+DNunrCLfUTXGLWnwlUS9
AdmsQDQbgSe8z7KfXWSix6JeUrpYk+IR8YvJj5N34Jub1vDNAMCppULwWAvKReah
AJiKDRuTuDvO8psZSmrsILJBPlzWt5BUA0w/qp2b5Bf+j46DbCOOpHRQsDE7bG6W
tnMw1N2nSkkwrC+pfN8EGlvGTZxNiCOKk5aGoxvRPz/j6Z1CcAkTH3kh4Ns3am7A
oNliRmXhFsoFlg8pbZMa/4OPt5F91HjJQ0TwTsSl9g2kYoIuCVc5n6BmihlvCx0H
v+aqktfZKruqx9shOg59qTDyLh9Sb6ZsRzosQodXxWDoBI3AbPqfLSyXUTWSxRWh
5sBkl6Im59MYT9kxy9yexR9iAPrRPjTPAC+s56n6/odpy+iWayFJul3eRHYJJKih
zp7dR+YzWPVib8jGlNa+iPE0xXi97OXCcCDhHZW6EIeBGuOlWQ9+Md5i61ewoJve
SutUXlAbQg3c0t7pylSolyw/pXkmTdvbRKjPZ4wl+n+cIDtreO6DAyuMsOcklX9W
lkXPa7ysz8k8IWoJOvFDEqaNaCv4rLr32SVGycfKFem41whQ00PXfrqNS5riuIyl
R+IGAsnHBzL4PwvUjV8JwYh+jI48xxt9mN1TzsS8XRFXq96F9FuCwG+G1/rB0I84
1RQolIKfNv9NUu9X+PBVlHRI1SbOlQ9+7AjeA3FTkhUmTacyqlGyZFE42K8DR/oA
f+FEgzwqmuq5YcZLVV7gD3QwlU9RPFWgDL1A9xU7/bReemYfnyyW6s0l2Mmy6oSx
PW7PaIW20499uBXU0bT1Ins2r7wEyEzUY4kUl81CCsBtonyzUl+IWZxQUHZhzFjA
ZOo1hlBoda4qE9jdseu6GWznUFN5PtZPWANp0NVtei5EBOE+E3jAb5F6VfRqjoyy
jvQUd7ZFIC7iejilcsZxtj4l6MV0rzJra853Coue9U/fxq437A0DejspXosdf3f8
k8HxZkdRWaDGHxxsrKSA68qJuk2j4wZS8n2HKjig+Lso/BoYpylbR8bStnqbLTBN
ySGwEMBlTw9xZWFjAkEfO+/fC8vqZXzgIU2pv+lh5Vjgo4TIVXnT6MlgvyB9gWkt
C4dqB3IdMfPUAoUZ3osZ7msg2NKvCfH63HslpByvfeSBPmNczdPvrwQ7wuIT8bAM
4quAcrbv3H/VLdH9W+qCpoEK39dLZ8YtDxkE+IyW5uPL01fFsdXQrljX7vyEJskK
z5m5abb/3+79jRtHT0EmW/oNcbZxYsrsRED9bzIk1keyKj1Z+s22rAjaaQOon0ov
xT2NRiam+ozjEEFfHXq196tb9gONoEwSYFPDVuq/vV+6m3X8W696iMm3p176m0oH
Dl+i3HR/W0xRBi77aMasb5xOOC8orfs09Jck9/s/RMvtEAfN9CRuQdTXwFfralEN
a2jXn8qA1tbUix7DoKJ5iJatsUqjePlMUcih5CK6Y3izv1uVRYPsOEPicKbVR3Yv
GkjAmytyhxV/l0SgXBSYEEz3HEmsu09I/OsKCaaVZl1X4IgfZr2gSxCehKyNKMZs
hGYWRmGrQykDMMmCUMrMe/A8MZ9N5LAIZfa2GdZGpAUAUawyFk7AZQGbtfg+ihFn
xKYx5E7RO9/ONPiuPhSmp7/JdOT64FMq5NZi6h2wV729Xrc6MCcD+Ujm13qagjUK
5ivL6KCSxCh520MyXZao0lwvo176Sm0BgqQ6WDnr0qnN5yBBeZ9gbINYr9aTaUXz
v5g+ekjZk5IafFpx5/m7acnqqkDC4K98l/vgxqumAsXvhnB25IHqCOabYu/uWxU2
V1cIEcH9EXuHHvimV/j8UZoh3ZhZ8KcQmdZbGSB0blpBqQ0AeN0Hr7pb4gZJqhaT
8XqqWCuJ4OQtZQ36/ddK+qOg80BgM6ztBVITU4L2cZUI0CJf0iEG9U7+xgtc5QML
2O7R3XwQ1EWSEvtFQdkLJ7vob1jOnur+4ZfJHiOoK9+f71EnvNIamhei3wLsATKM
206OBmgS7TJpzRLtP3fS9ev7gdVBrK5wHpoLrvV0MVJHCED/Mpf4nEvWtb/U9Qmf
4QmrVH97p785Bf8z3rCa0jhZ25ENpsF23/VoXoQUrL5Srf/HEMLxTDDpQ6UgsumY
fnDN+HcRjYm45RFJKNzuUA2267TdSXw3BTCUjxrExRdi7wAf9oAksIwtdVrzmLDr
7OjdEnUvdoavZ3TP6sLeC/Pyf4qFkIcvdgaCwzir8YRWEwSJ60pWKqkHdXaqVml2
x2pfYAouJL+aHyO7ldf2mhjYY0pc/Jrov+90MForbXSq0HUNBETOTH27HjhvhUWn
KMLR9KTrwB0cTbDSLDJgpQ+99KD9Ox/uRAdQQc5/ZWtYy4VVWl02XpNFJjQpFe9Z
DU700AuouVmoGIrI3gZpqOdiUKRk4sNQKf9AcRZ6D2UlPTyTUdVBFrHF/hT35SJQ
EcW3wARCWWZoi9PZNyjEZAT96yz2xnM3yrf7K8DQotgVTDrSBdOmT6LwdrVOokJe
+O3SITGkyEr+/0V04OsD6W2Vpn4EMIYO7AoHK1Fwbt+/bLg3lUd+EbSfkJFEwlFG
Q9bpIO9BU3umYSH0b6i0gi9FIns1Dj+o/pVLPxgEg/a5JmXvUKzm2ZS4TBzOpgp1
QjiCFY9Phir3LSsJ7KbfG0jqI2giyCGprMfwDEAQzudYvbKQ6WAEn4j6AsBN3yGl
MKlcZKXHFKYTxfWhjH9iKrwbdNSNQx81hk+dQb0b7ift5mb3J15Izfmdx1GiEZIp
jiTUPPEr7dDsgBh0IXVdjYfZjJxYgBNVUqGXnQ82YjQSPHB5OawOVw5ozstHjCeC
LbgCXs7efO0OZNKRJrsGy7bQNQBLtPg//ZalQwQVes+pZ4r7jeVbNUSbPNyVA+kR
E0lP/8lu4N6fwx+VQamKSnglsd1Y1xNKxUIC9ENk30yQAzo1r3VKgWOkctNewpEE
49J2aR1uiU+SI2GO0lLNWVE8SZ7aMfbOTwM/vgof431tEIESpmcNav6q2s9pFxt/
rNzX9o2oo+MzzpNiwvAD2azTqLbLcWlqr4MXapkLpHZ02KK/6suBUB6M8cpPPf71
P+Oi8Q8bqAbVkX2qpXXlxKgpZ4es/Qlt4xe+274ubH2xuGaFdYn3I458hUF30lJ3
hGDhLLg3xhZ7RHxmcLvaqzlS4KykHKEisWTUSXkrZCUy7PQJJCsAGkxBWnfFtB7s
wuk4tggvZEgAexC82PHfuLJI9yEbcy4Tlf6JKrRN4nJj1Opm2v/hL9EFjGNiyX+Q
foldJ/fJGixb4SWXguC+tBL30K7H3YahHLHUs+BvcIUe/UCbccIFDojPX19DdtQT
e7KS9DHSADB4TNT0Pilki5gydQveqbSpjcu70Gypzp9yes7Lp2PDx2nHTIy3lXns
eAyst90CpWg5zwIZ4+7NQlUUfpneXTtTW9ZeJD6IzhCpsZWhT5FuBjL4aDLw0/UX
llDXlxGWyquIepA7wkEYVuGsg7VwK4XSHTAhmVd160coOSsPq4+aHoFrvoskC9VL
Vl7yLNIJSqiG+EQN0yQQRTiZCYtjYf4eoUS+NwTA/Es/xN5UirqRnk77aauXpAfS
G+6L0V/FZyYPjQGG4CVn8aCPGuMqvaO6Lt/7Tl+GtkLUxm8kn1EfzUmGkCNOYqiB
Ww6QB9G/n2yxUKLlhcbdy7LcmmMsxuxmxUlx7UTkOzewDGjUyIDS0RL+TT6p4UlA
QMN6uHsWH+gBuxjEedgriubOw6pQrP/BXM0LrzCzpLVssdPE0d4QiLytaIKBHsLi
I5cAzLshGb8bDN/pyFJKdBTN5lZWJ1Mw9bGKOnX6mxC+r+Qa6eIhDCGoin+NdWbb
mwxtn1ioxKEkU0FGu5r8i6x+01sJWii5AB5wwMqQOU50muR3pDYK31BqaUYMS7kb
3924hboUZo+BgPfHncwxyd7UKB0xaQ3650YX3ptldGcXXVKClL8/N0zB+yaWEYs5
oXy/es1CJiBIdplTUXfvmVSwM5F7dnQyrdGshorHl7r1iHi2vTHTBKby3zkV69f1
vR19bbcTkqoNz+qmZmL79PJ2+MFIGa4fZ5SJVZd08yPjkZgxQLMMOm9M33C9tf2L
heh79f1KoJBdN6yTCosprBb+t+Q0WXST1nh/kL5df67jw41v+OlQnMlMKaCs7jz1
MuDLsG/KdPD0qlweDFUz3eTvkUcqGiXTKxEHIQTOJ4N3GhDfCLOgOyX54p6fGEUs
f2SsVv1DO6C1wjezmLKcpiw10OSY/3v83sOw1mYH5v6LT5QJdTtg0Uo0FloVRocN
LdAfEyTgMnv9aumUcb7MB2Fy4HnoO8Mg1qv9xMVbqqZwZgLFjbLKH4v/6zQJTTxY
QjvLaLyFq0HTPtCFfE1Og75jRxxScV4GHa+M0KUiHAcT6I8gISU421pFYROtL191
erAtpQ/i1l6UZ7KMmqR7op0sEf6d4vdjXYgPfCVOVd/B3+JUgxjFOaKOb3NAS9Pz
mExfdgo5dz4X4L4neDPv8TsETsbUVR3XCNdRb8Pnn8bJ7tBeBj1CRGpgbgmPy9Ld
pRuPVDhgAvgpzf1ruphWiE7FpvsGqLhtVBmbMK9m6Yir/TOgddNhWo5rqpM573q6
vpy3Cr06QU7f0XqDFYhph4Sqqfa6JQYAWuOQft3d35OhF6rmxoRLwiqiqvxzBWZf
MRSJEAAxnE30Oxz95CAfiISe8bso9RwWWx64t1OJ8iKJlyB8pQhwDpaq/lAvVZ0z
f62rFb3BdfQoZW7SdZr2uk1tkJDKdQm21xXJ5sk+xAp5dST8CuiLtn7LrSZcyhEd
sFChcyLU8ZViRW9BlciG1J5QCv/6YUfZ0R3Qge/3ofWNRcPa4r1PYiUunBc9opMb
DDF+BD1AM6YDmbgH3ZLiWsswjsD68TdqPuGAhXZAXkhpZQzv1fQbAMjMF27AR27t
Jb5r6/HaT+2sKbAlH+5OlKihDjLZnq5VgUL1D2WEA6MhwFkA6a35tXOYyOns7ft+
NBlKzkr/HXZEPLxOVm1I5jpx5/ZU2fNSN1F6uOlAhVA2dr/wrjgt8/t2a22wDF/x
XpHkhN0+M1Il7oWD1s9X6TL07/jrR7BL5umVFipJFQDoECdGcDMStZ/hhxkvt53d
SdDuqdaLyf6JjeJWYUyU3LlYQJgA3KzO/1gP99PHofMx6q6jL8hWPqbB5kbNPlDr
NEie5Jl0QwsxGaSv6MRu9KqE4lYSu/n96a7LpgEz7C90537t0GEqYk9KQkxj0H17
u8lCwJd3KBTjzT1QrB4YbUlw7dgBnu0ad5oc2b3znD9HJTY3Z+T+V3xVEFfMBfXT
5tOd8uRYPGOKCNh1H3e8vrTDy7g8sOOXpoQSH4rI2hcRqapAfO3/YUYy7I+CVBic
CEBeSuYeVXjIlwj7pqJZjOpaAhqh2eAt5E5YJH+pGd3qvWTivjHCwmEg9y9PzmVZ
C+CET/lFyE7DTt32uMdFdeT4xU9cZIdJrNgnnO/SL0Rr9wWfZh+OPDfAVxoPCmTf
WR7nbh2WIIw5DUz+4ac1uyC4ShGhk1rzipIoslM7ZjF/wnZbX1sLZ6N0iVeGfPaA
1b/0gcHDmQt9sb9jansmCYqcGe0IiWZ0VSmLGWiVb31oxT3fAPIb4W8lY2Lr/IRv
xqX3n0EbDh0lzZZSDjEWt7e/MmebHjwADnncyRqLXNVAdudt3FeifEWZq1ps7gGp
BX6CpCSSUBuT7EUuvQlcB8F/mjfQ6N5EZSFOAQ9v9LPAynAG1wKwouwQ9K9wh6qx
MpRajetBYjG+s2arzkC7hf7ECvS4DDF1LAEL0BzBpAn1pfYCgGJPRXMkN9dhYHVV
TegWDNJefaBZPQkrw4tjIhXJH55TGIUOJWRxEx0cFHQpZL+NmADraOcFkyYs9rtQ
4/FA1O9eyGBTUG9r65mJpwubA0Kl+V7RZZv8rFwCYvVx6Iqzk/4vLdoI377/DjlY
6fguiGoM7lr8xPB6IuNhsJpShgW1xsP2O64kFczrhxhkzrp8fjuIgbl3IFnD+vy4
AS8nUlBiIXiqfueemTslzfK9WjZP+rv4hTNn2h5gy9TN+cWttl86vzTYw6KpoOHx
Av4/WJEEEt+rGloJU+rDSfCTCJB5xhlqKjTKv754bmHfQjRTrCGotj7SUpO+eC8R
rPX2XtWEMAK3wMInCmSJIgb702JEPRlQ6XjQCX7kR8tXZIqFmyel6CcKtu+u+Mgi
R4ZcySV/4bDX5cbArF4nDeM2AwblFAXTWncEeuw8bjc7OET7J8mOjhAhKygiVhu3
WbkkkhZ43Ds3LX8iEsCcL/3F5PrR/bxvjVryTkJFKk8NnE09BRCeRK9s0YKDNM/Y
zeg8Jr17IAfzQdBnvl57BA4240hRuecXmJQYpgemK0erl0MnxWBDPMS7W446YvzH
d8xsCClvKgYbMCOE+1CjKlwr6lOozZkuQzhj3M8akVx+adaMLVWEAo/hVi3ELdo4
6XK9qYWjGkMi7j5x1xur1vfd+Kf+o5YK21x45YHnTE/hBWSZfCk72kvja5DA7BKu
3voO+OrRVp1i+RgO0beKcmdHm37uslWk9qroXpfLSyqIKA2f8J3tHpZAQZl8m57G
zZWpnsZDYkLfOLpZzSpklQ4LmjuGn9SiTsPJU8OnM3omnbmwgJYBQW9rSJyKJpn8
BYtozeq6GoUZ7loHbh+GMqtzP8x1OSVnHfIAe1eApKEAub3I7vWnCKD1d7OPkU7Q
rSFaXR1Q9TkTEgCk7oa3B35v5N5HNMSDHJ2F9RGdvAYlxgmp0QF+2L/rhIdW82pi
MFjYbfEnaPCkWnB/uogLATI+RGAVUWRnojKdWr1lxtEjoPLAfEn1X5fjON9Pj2BA
SQZoF3zgqPBoFqOB7tnzVBQ4iUnoD1cOskHeEB28OkweZt9YwznQkNC1wdivs6tH
bpwmkUP8lBimgqWsfvSoKjG3Xty0JY6P53DixuXnxPy689BlJDVl/pvQZSTCAh0X
OCppQan1xXe+nHBXI8oTAMFuvqVz0DYtiH4+KdAC3/YfEH+4gBNm5V3Aqtz8Dk8t
6vE1isL4YSPeLV+N0HobmgB+xssvBKNEcJVHt1LzckE421gImNUXkKwAdiXdJvSG
5hTAqw641DHoGKwvqAyukwwc42RpqSY2FwjpLKQ5vRik4Tf0IbxnAgpDeO0O01D/
Pup3L5P8Vt5zXToEsMvVQ6E8+KJwtBBINpM4ZS/wZXQHmlb2r3aPM+zjHHX1yb4r
FGWBkzRY0F/KpjL6Zv9fYSKqqFaM8kUpjYfZCDHId5bM35sJi0q80T5pd/xIRt0Z
q8vXWe+pW3nlSsC8jBxPzR4SxX/0dgM8hDQaW9Sulrs3CbkbNjD8Cs+Ua+h02K7G
zdp+ihXyOJlKBvSkozEh6mP9EgC2ZgAv/X6En6V8qPb7US0ORtEvoAiLEB83K+4c
nvd8sPjgE53N1RMjyOpNYP8RUzKtl4kU5BreXLGv0lm5gvmp5AUf/FwVkL6DW5FS
bL4lHWGDc3hgKB0dY5hvdDf1lxdI8d0kxCrp9q6edSd279QmgulvW90lkW5jW2hu
CtM1gJMmITsV7Wj0r0vIACkWIjGuJsf627SdYAUPwl3F/xFrRFVKHVLMyG7zh1Ob
yCDWodHdHbpCwhAHj4S9vzG4rXfua4nRxQJZgDf5Zvu8iQkFqVaBvEthT/N4xjmM
7eqCnd+H28WM3K9hlAHPNdzkel+skkGY+jfF5vK7+ooGbiUa98/JOTOhjDLKs7Eq
pA6nDW42Bzwz94TFo9Ytr18HDXI1CIq2iKu9o5xiQvrc/Ca6vRtJKuCyYtnPMAmG
qJsKibRg3gb/FwfEj1adIRdOUsYfAMyNKXZL5Dn4ZaHLrJzwoeOuG8jH9qeCrEzR
7yEqcArSWVOa9KZxbYqFc6i4QWmHBJ0GANdh7oACbYp82UpTS6P1vN/xuG0qBh2J
Y8XxsBGfuHJ9URZNvmXwE2Ksxb0iI/MXfMNrBLk/UpCj0j3JbR6e24LN+U2r82JH
ceskfRFblsRaX/fz3Jzr9zL1JNAJPVzYrkj8HfiW2H3IsOn+yFmoMKQQod5b8JD5
6VACEkgsiLnpMf65Y8hNdrDjpsp7JCE/qDsIyThkq6uAuVY3tjvnCNhA8Z8HdEEU
prc6tr26dHvRk2tFNXll4ru+Fk/ux6XxToEhNnwRqGuIScovd6tJgyTD33zPSK6M
lSBbyoWO36u8oSjIn1Gch0TnmvwpyY4e60pvJbyNF+kFMQIr/Jg0/rEvYtxUgtLT
779wZ4s9hBZx6P6UmMsBy5u5bl0VndSg7ULIzbWhQ56Jnq7D2o8OLWjOIlOy+RNX
/dSiI1EHXXcxZts4JG8DCEuM8DXMU4KbY+Z6V+Q3hsV9pmXuI3aXZsFHhQeV0GYR
/mm05gXA4CAwhgb5aXhPAVCfBZ4i7vk6qCpEGBoh/XrcLHfbkbDV1jvvHTyf0DL1
oEbIISc/E7bjXTJhuvIwUif6J05Sd6+MW3NiQ75/KzLqEsGZyIN3P9FmD1vR1jon
ceA3Q+REELghBptppKXJL1YCLQlh0peIKLsW2Nxu8nIkM82oCHqfVkAxRH65GLiP
lfjI/aZpdH80nXctSyZQfMOZ7qi1AcuMXRo9KOhk9aaGRK0tiXZXJRF7oHf2AH8X
5muG5SQVhpPKGPcnm/f7SWlHNEz68pF/b0RRP0Z/AnLIlEqS0rmtPcuTfo+zjrd9
MGtYtCE/bdSx0MwR4uNbnPCuU5ddsIAP8xa/VVRhe96/rS9g1Ncy5zsgoAmwyS9D
67iCuWlQ1w7i0eHhcMVodQZFPTAhOak8oeJoR4rS4TUqDxUlH4HC8Yot/+VYdCD7
CY+CUfGE63xLO+nERfC6KEFnx8dJ5aZGkwsvxxdMD+EazFhl1BYNSn6ahYpB3C2q
VK5wtVa94qh+J7n41rw3a3QcU5pnfDE5YsUQWK00isNpV0JzRt7BsOmqbQSbFa5a
SSWDXd+3x9yN/oBptMRqQEsZPfOzfXcdFfsZysna5+EEO1iF3NaLk0ztLUDNG84w
q+14zT5NjLoIxCL+bzG2JqEPy+zUOJRGwYGO110laGYGuKF2k3jrJZTsaIuvSEHL
bUkgVKjFPbvDN+22iCfX+K9qNEkJjNWG+UkiyGw32vOGmLQkvKESJPxhTDPPtrFS
Pj1jUmllkoBDOm70bQkqGFFwmQ1z5jInzggFGa6kGjDJ0FsMKFxl6epuZXIzDU+8
eAZZTFDlhXviCzCSdSPofXc3ndncE7Dr28VgF91AvreEeY+FW55Yyfjs8yJR/mQK
EpfsTSzbuYmofFaIhttRIHbMvpruDKxdg7ZcN5eT29cKC2XQoaJ5sAgKYQ+7pb9p
UkUJeIFzuTDqMcWeJrp6NxbJj+4WRoE17IbJIsnCcZv13TjeMAaMaFocC1YxMGbu
rekMlbo9cRec+LUxAZYQgiMhxAJPMQxV92Z9+1b704ukm/zmFH7JqA1mMQ/fdj/3
SSS43Bbh9y4LBUR7nBCiOsvk8LU8F48eq8kB56p0+ke87wX9ELKR417k25BPBnZ6
tFk8HHJtj3Sr+84IxNs582ZfIJQxm5nJCBSSMeH7v8uSiu4U2DTepZ6ZcjwkmT33
LU0kC5xowayeYpLoXNHUTQM45gcjZXBDzEuc9bDplfqQ4Q/Oh/2CBkyZgHpO31Wy
Oqw43y48YcAslR+g8X+VgmJ1zP/0A9u+5ha0wzii1JzinVWctxJ1yxUglb3pYpji
ZEpUWHZb9R8iqgLn/Ntp0Wa4NiynQ1WOLpxOui+cmBJn4GRzEIqQU9sYL4cn8BoN
yLD5+9NZROTFfHKT3SdjEs2/a9YESm+8YA0/pS1noXWXnprhBepAwro+cZOzDkUw
OEs1DzZ7kB5+B+FN0dsfiCzzvqpxLF92SPaxQvEclp1ucCLkyvEMs9qGDxbyyXVZ
vcEjW4czSA1QBi/XYsVPOLbOSDYIxJ79sN/zz7JRUfFsqujDl1cxd32U/jSLxrc9
JNPLidsK06cKAU0dsgMBlYRvCqeNp8+1xCciz3FED3QxOTomcVFrTHr/DhovaQXJ
iMoYSFoIzdVTx47Sttee6IZ0D/bq1yehE30bHIdsyycbPBB77aWnLvpFcfAb8+yb
G64eMlXsuL9OMCM/REUwFxFx0nLsN9MqGkgob4EqtDxOoQYlD482xrDCOlJsWtfl
bPxM4BcSkCSysRePuLVjW9zZVXdsEI5Dp/QgukDhX3QGFWWotfO4yNm34xZFIQJx
vBfjsPLuQLPd5eCRu2FgLZUvXBFnqymrVEbIaVjzcAFvEwuQRA6INgN0FVJzQ8hZ
nhXbJ3rS4Z18jc00CKq98iUWeo9BKkU2EeP+3CNUp5UKfz5MBAvo0feAedDu3GZV
/lNLUWf3daEtkTNoShFQVk66pC1dweSux3j4rlbxT6wKTmbHuW9+154HNirMYuPP
EwQAJ7JYVzVf++0H25He61KdjZEOr029C175TlP2R2V9hmiegPmTpjUUBaOSqgGc
BY4bQwxKTVAQmU2BWwMlHXYG7AXul+uTQXW6uGDyZP0Ao6LCPGEwaSygO+WO8aMD
AqbIhBBnuSvdyQFDjqAefj5avoopMC0XU7wvKlOQYvT4zMizG5TXAcqaldRHTh+e
2xXoroK4uuEI5Hl+5iG5jJ14zlWKlKHwl8ysddc3jOFZ6flvPsj27Fr0lbD8ltCF
oObQUWXxd2CQ1s6ImjvENFzTsjlo86zF3pSs2l7I+u6AN3LoLhTM+Vh/PWRB3PNj
CGL6Clw8F6E9AF9GADiN8gR8CAu8ZxYyVq0KKbqs8na20o7B0LpxH6jvZJzw0AaZ
N+mzynz8bV2jLLAxfQS9r5HbqMF/GOfYCL4d/qvqRNOGEsonQV90gSAKWZUXyHWu
hgsvpgAN9ljHhaWk6UYRtIXKrIeWCS4Md91jFAQXoCG5xq5hu+qlYpPG2y/tVv8N
bqJ0HzbHPW3UzIxYdDQRkxMsk3xFrtzLOhyupP7UX0dgauHZM28CXmBmI7By4lt6
0xgTjPWH3yEMQCXa+5aagl5SQMQms+Kv2ZdOLIJtFhYvPF3fsIvyfiK4N9BJkskZ
gEj7W8c5D8RKtex+5NnTueDcSfv/INyA3ZQFUVv6YxDYVeG47UPtTgKGlMMs1Ckr
KHBVLETXVXIxe/zuYy63E/DxaeAlEoiTvW/OW2bSCWlibmhMqSyeWU2YynmUolQL
jDTbtkkbeEUVnp6pdAPIAa1fCYkSeo05LqLIDKU8M/6AY7tx3VQOGdt1ix1ACY7I
GhxMl6uKa0rhQnBlYgRiyBLWUuEV1SSJPPfp/u0Pta6xqxbvmzmyUDnQgzb4OL7x
hhcd/15lMDj1qfKQi7LuMbVYcXvkPXIbDtGGuRJOgIalzSiMaTqJiGvwmVPLoDmb
Y2C61wfwoT319H/Yci1HKcqsvR5a5j28mP/d5mCIRQKgn57wwwSuiKQRppep/xYS
wAScpCr0XmciCI8UE8vhBXzpA4F1Wrbjtb4AST6EyhFsZAJvJ77mV+tmWUBTGLzJ
uPYzCIMKXFgIi7R8ze6ZPS+w7yesvfRaEzpUeOnV0AVgkwv7GueFiyZxwDuxsk0m
A0SLAmoJOUWYSvgxdAc2cxlVO1jlTnEOEdUELniEDxecLcrR4nF35wFezBtXojoe
PquGKr3D32tr2IzkGIf3lv2TsoZ4miRKArMn3wTVwHcCDNUJe3OYmyHEaijpeJM0
RXCJ1N7pBL22dmQPFkiCrYUYaHH4Lg9LgKGVqdCC3mO678Nm8GifJL06CQJSbhyh
V8irqLPnimkc2E0/3qpHOxBWl16TvUlDAkdFp7gTZZrfHr0ldvJiCjzYwyieAVWr
bs1kjQhmPi4As4NUUr9glZG/aQa0c/dbueG7T48dgNFwpgmYtIb932SpAwbMUCOn
jkNXmF68czUpNXwhG6ExRE8VcYS4McalKe5yptWzXNoz7oSwlh5jG6LfryNdKwFt
vcSbSsgHth2P7SXX0KMtZsxZ9DJbmuYbqLwbwkunVEm6gncfBRg3I9CKgvsb1Vww
zxtg9Gixq6VGQKX60nggjwWyCjFchHrDiDsyYe9zszpghBX+jvnf00AhHPgJzegF
Kdi/wJLmJ//TvnYphd98cty41aNPKCzNFz6NtMOHJLfVsbq76JddaKzZvV3mAoib
+RMnQp0CqOccwQ/Ql6ItvVi6py+JekoxOENitEh6guwig5MhREEvHUEgrM9AWtMs
xIMjbBoiE4Wk05LA37nxgRzMk2g0+mMRAjFhOVshqocpg3ibzqfHHUaBOwaEqyrg
YviQtRRsa//4UtC1T8jIogcmQ0S3xMkLPCh91WvHWWkfEyUW/KiykAwIp0QQWWPa
0uRluP8cMvyJLXp7gLjROUnT1UFQ1jdU8brBN/HXIU9LL1dw3EVr9sw5Yk8KJztm
JO9A+ejrrRNMLBYNXJSqVHzZIMB5zbih+QvU8LFvcPzbXSyJHDRObmrpriWyiGLZ
Hm1rznnaXZTqI+EAaG0fBhIbhw3kTP7QRQOO2PTmHS1KNOV0jecJxpwXN3HaXxTE
Hpax06I8VP5itBaxeAU36M+nvUzmhTB+y7KtbEY8vvlCzOtp1qS+u4UXVCsXJVa7
+C33xyS/0DbmizEJqq5qIZvSqzA9nQNkPIuPAetwchqKOLq0+qRtKRMW5neHEkH5
JGtxRaEbVh+QQXK+LjnD3oKNo2yQnp8mxP8WJ3+NL2XTnQe8J+jgx8Ni2pJ7GIFP
o3NXsZwPo+AFcYC2f9CyO0eU01XRA24du+ZaP7TMGhoOX948rw4z+ENhqphF4bR9
N9ArM4UDDaLO9VFzyhq81PFVM9qXkIPapCWQPs6tAdo3N9LMMjQLu9ALYWUAt36k
Lu15ChlzH/0kBmsmJ026hDWI2mNd1cEtucr50OWGv2HWLBh/qD9oQkD4WkATzYpk
kq8lN1Yhsv8hCpISjjJtOx3t54tTAsdGzOtGyV3szWYxD/QhE27kdopi22HdX+/F
VMqe+17elq8O32akMD+PdS3qZfzXA9A/HTczIpL4FmtW/IEZ2etlj4bRqsgJVuTq
PefkC5PLyWIIo4qRQHYrfTXuv35cuQxdaQpxKU4ZnxKsygxGCMcsgK9yx70AVKM8
/fIWLECrHHHtOA5+Pi+ZuPXhI20UsWrgwm68Ymmz7cJIvgYnqFuNpnZKy/N4ge8P
wzyq68/h3JbSDk0rpEu/yPOjxqkityE3T0nljoq6ACVvFIqaBN7bXQAnb8IZ+pRc
qHlUtCATiw8lNsSrL91OCi0K/QejVpYoumubhvGtt6S0k/09yriJDf4C4EKhFyHb
TkA1H2Bqow96mD+GFR6oh0S928hQehjg6ZA3f1W6O8xeDTkOGlG3WteazSezttxd
2sWZg41OsvrS10Ro4ChCIyyeYcsc9YaVQlarZ0nOwIvXoTkmABfr0MPzO02UB7FM
4c068Pau+z/g8BEFDICeBCWP1cooCZEnDwigG6bNAKgomQs+Dd+R9MRS18fT7dOA
D+yN0f/Q/XclUVnoR4NWMPJwICAbnso/neM/kFq8yOZNF2P2soiPCbZDlzrwXDuy
OVRrANZTC1JpdDp+Jz4B6zoOoQMHrYQ0cHOmUX6QAb0j+F3szCdT73sBYa22io/O
uYQA7Un5nF4NBqkEDLzt4Rg1dq/3hcM5UmD6FDoIyiObOqbhakuuTGBc4KIGAZ+X
MPyxdKpkvzhkSJBf+Kn3DHslMoQlFS7arZDoQzm2Yc4HKqTqHOLxOSSjc9ykksvF
MhOKgE9K55DZL8fs4UnjSrJdSpmE9ZfAF+eYaFc+B9Vl4fjPd90FaMzq8uUzpsdY
CKhWMIcWfs5TtzjEx7OEGTirzsiv8t3IKBverWtk0sMMdgSfiQsHPjQ1545vMZoH
we+u+knRyYz/OVI998aAIgaNPpskhrHp2nCmpop/d0uC6NsnGxHtWwECDIhSBf3m
p+N71bFcdfiU9UtGy2vc9TUe+/e2uBHwAS3NUHrQLKyFFEAKzAIUuTEpkQQ0YG1I
UoacdYstfK/rWgjSAuy8jmqbYLl7/Rc18wcW4fevdLD3aOefaIwtPRaXkd6IFMfU
ldbQIL9oj727pA/Ht+qBwtFzrXnppBRDOV28iCiXQiJUC7tKGo/VJ7is6H9OrkRA
TygsEfVDnLLssFDDXFpbATXyYME0Jay+CVm1cmI8G1EgJ7lIFZFRg99tjSb6sVMS
Y7mZizMF0YolhcDUwgzh3AEmD9iIm7KirjZ7t//Gf8NkEvER8A7CeCojR/uk60oZ
HGh/mDbEfzD20++jzsh1Wm0UXxsHjRt0LW9Eo/fbrSXfom2UCXlUWlz51wYfSLsA
i8GjZJ6DB+1Llj0g0HppRFeFUpz5oDHMATP0L430mRzv99L+lx4acBjwKO6lp9fF
b+GXHOxdRmcpIxYU4NRLoJxKDIwqYbDemRLT9Uqb2wKWjPMYTCf80ynO73gKtCNi
WoBq2LHmeGdy5Q6brYHiOVl5DZDIuQjBJY8aUmzStNkx2D6BxPGnIlU7n4z+J22J
by6t6MH0/iU0abZtuXw8XKRyTcdAkbHsJnXiynZP84s2VVCfI0oY9tiwhditQGjq
3ODrW9v/SssKVjS7aD6xhUUwXjew75X61YOIJO2pG9JSV9Sa/Fm+cQvLAP7K1J68
78TvF/d7jiFB2uMsxsLxynU+citmEuPWr4ycFh/0eKVm+lafGlf9/QfmZ8smM2eU
6q62sEKQwWeEb4NXpejoX27l0QAaQV2oHjTOBlU3RJc2UW/Izpc1deJrGsTAAhks
smb2P1K43iQeYhlkyoNILL3oZiTnI+Ut4BP2JjK37Qlyr2thWTpPGb+B5lfBjBq1
X/tYd6hdl1ThjtnHtEGOaRbZGdc/OPUGOA7lN+BCbIUULtNi6W4yFCjJuXsmTi/u
bNMGAOCFsDCTyvfha1Gq6FpUwRWxcZao02SYYF94Q9jlrNi4+2RmoRfEo4J5NWPd
UtkQX5BCSYfo0eRqZ+3xxWOPg2+usT4S48KT2klfzhf5WSqmsmQCIVLb0YgysWu3
Hj/LcsDrdOLwl14iLt4wJRdUEhjBmexzPU3nqSTjSvfVFqSY2yx+dG0kqKNZfT4l
AVnRWD8HQctJlwuD4a4PHCS7dDzrUv4OMJrRjye8e04m92azma6SyFaTzJ6bYxDA
ejxmaIrNdjB70ojND9Uxo0NA7u0nExZ794W3kJ0EIoHBP8YwN4OgiPLdgz9Ps/U9
SYk4ACY3xA67zkLtqJ5vzZZcjtmlTNiaMD2iZVKILDfqEss3DnjI4xOKRjerd7Sk
gT8SgKkhHXXtv+AN2S+65dTy4VkNZd8SQ5pyLlBKBo1SGGi8nhCg0hwT2L28crE4
ve+2Pd6k8olR/SNmBt0TYW1jVC6Az0BZh6YYmTPby7unKRG8DFr09RXySgB7k/Fe
jralQ1ICBQLLxlqDHetEC1ydT7ZgwWdk4hbqwQHGUZTkdnPz/oAktm2Dq3eS02PN
mgOIns3tMzeUzMP3oeRcOphVLtdbFRDBAcM9kajq9bGDd4x69cHzQcwEbIzZVxDO
/eLDMuLWXrjeOgVw9RGm9Qr/cCL0aGQi8A+4zvmsYoRFMKsx0gemI66M8lSgJ+17
aLzk1be3remgbgwGfkPMzxqmJ9lduvGTTs4nntQPVmRJWYrhDmel/1fViQxo937C
7NOOGijoGsJ6KaPeyuU/4+mMmF4+GZFT1Ec81XBkCaGX5Sp8cplSebNdCbG0mQN7
D6ML10IQw7abVmZ4MluGhGdgZitpL0qheLPBLqjAp+07FalC42pFFZJfMAJrhBvM
VlK5BU60zeCFPKytlmWsqxoDt93rc9LxeFqPJMKzyED/sxbRg7kdt9PcFhzwpwm3
ixaoIZ0Q8jR/4J3cF2RTfpSPFCbWMu2oiclx4uyx8RiVKceO8nfvnEoqlTDxwWlz
lJGo/JBCk14wrJ2yOZmxEMyB2NfEjqPxRREEKFWduLQVTLXd+cD0MflL/yKMPdDL
7GzNsEZ9DzayTp+IGKG+9uMK8vWDxLn9YHkPom9kPKZJpaii1YySp6IdH3oP8KHP
aScIzznEPd/uWBoK7HyVEm21vyXkW5m1LIjqU3g9X5ACFRTB4JLKJFT8mukmAA76
kKy7MYJBFtaCJo3N/jpMpw+7+svtyfXv6uCE+lHq7mIpwNozpdtCjouNV09riWRG
1RT0BfkDYbvkqoBO6evPcm+NGmXg5P4vydSJYU4LMgDB+ULMhbdqiM4BW+ZrtPH8
xtIg8sbWDtEao2pVGOOVAUZHbG+G3vgDn+J+heHkLDqbZboG03EUQRRvEYbU19ZP
HLULHJvwFCNTC7qoa5mn9PgmCSWMuFTTffa0Gr7dX1HaJsdN9ZmzkJb8MKWZst44
F/3qD0Vsb+PHYk+QXzvhdeAZfe5r3ow4W3hLizNNZm4WZ4y9GHsf2CsLebTsV8HI
F7YaIFmOhTOOtHvVnPab/iY1kum8aIFKy4UKMZ/XTDcmgRm3Q/t/9nrLPpgV4tDe
7h4kK7CR+5Jla+sXukrudqGdH3Z8NFC2N6maNG/3ba+8EGqFaDIQa5BXYrMNOkpf
u3S0Wf2y7Ktvl1LUC+mH7MPW13Q/LgRNYKsE5rceq5klZmdt7eQ2I6sOXcEI3YYd
4zzPyzYjeByDhD7fgYRTkFPaRoX8gwumJ3X4j66wOZIAsb71lS7SyRyJULQlzsms
BdvhSujU3duc+tdF7fhypVsK8wqd/EC1gYjxv5VnltRs4DudsvyEfxa+y71yvXb+
IcuReEk0liyB+Ke4X4rDJI1lSEJrcuIpWP0QktfPEn0h9ba9UT62dcJhTSCgK3E7
I1ywjsN2Apxs/wloHm5b/p+gDE+I/OuL4XNtRZSzhxp8km4lR6pvFAhr5ujA8B5+
ypd1abqmQ6RMO5Adml3KTQenQuLwUjuRmzURxItOgJOfUxp39eJCYOTNp6zjd3ya
MTf+kOTQSshyZiERsmRy+5w+lVgZxiZNBXv4g2oFMwBlCmoNs86y9w8B5QozEPDC
i17GFMqMfLgjJctqiUAfNlC3oJDhJAg3Nxbar/tT8pPAZG6xTP2fkfIp9Ybw/iB6
y6k8zTZvaCnAOU2wxzXmkktGFMtHP71X/nmVoS89CR8lf/T/oBcgv/wxH4J+Pgd0
JDevkzyJAZxYayov5yGrw9fTDZO0yyP1kaHZQJT5tfcIZSUlfCUf2tCrgee2K7mz
TR3lY7W4+Xu2DxsvQ1RLym5Qz/p5kdXBXuIS8ZfxaV5E9hMkNnZOzM0h8n0RCs2U
mXBIQUNbmMaslbhysYVo4bOSWpR/RWUp9SzY7cQhvNcxXe4iWs16doL6fK1ipe+j
PpOcgvpi310D2i9s6Z6xGvdnBdB3cpgImg5Cx6bBIhcQAg/KSazpvlcg4RvbrOTi
kaQI5D+QQo4Z7Lx6adr1P3KzpKkj/N7OYj11x1hIXFHxFRgR5urQ2F5YDjQkbOXu
kze5OlEv4fXkq5sXNF8400dpMUx7woCxzQzXvAPcFeYRPAfDB6O6WrZh1aikAUDP
dm2CbLfTGPHE8r3+QCEk+q8wSzhjnWUaTkHFMTdlSUxPhAo/SO2qsZyEFzcHRxrk
G4B/JMh+NmM3BFNd9jK3/iZotQdocpypGYYPHkjmcY0voTzcHGzhQcKw9SAYnAsM
DhNBWkoiS9Os924u/Zk+bBhWoHVFe9fs7txq8lnFUBTvUToCa2fuzG135q1exfO6
WQ0fUnkCW0oBqtdJWH/gdr1KCJVfFhge2JuDBERX5uWQWVtj/B8nl78hYu4hULZU
rOeYboGbrAQiJlqttP9U27RYJiM+SfTLSY24+U6e9+4FJER/52vQJ730Z0GxS8uj
i/wLLaTlZMDJMx9MVQmPOhxsURSKDOdzhVAqL/EzP7XALVGDD8sloF5Tf9COU8Mz
DMr0EnGga8wOrl3inWWrDD4Oi+JOvuR6EquqZ5Gh1REZ519nVoLE5aOf7IPeZzAz
LheCUSzZMMvJMbZnxmQJbditskyQ6bQy9Y0bG6fCK2NSCKtChMDqBpeAwK8FKl+V
N9TyRNnHF+VdwXyNyJWUBGSWsKXXjfocCwtBh2zh9LSq3I2vRXui8QyTxE5rDOSr
kXkHGV2fzbUoj7bsfa0njrmBBJguJIH3+gn02AXJYObvmMgS1ScFIQbfmwF8+sWD
vx+KP52t7FTyO2Y1TGiJtd53LLNHRzP4n3NelGIVVSgcKaYhuTz7lsusu2UflMxy
Ok1cX5bItSOrjV4oCf4HyDf1SXXotmNIG7SDDV8an6XZPKCTGFWQYbCxe3XWbfZZ
gmOcM27I0CBwyGvzNCeOM8N57DUTj2gcbVv1rFSPn1d5rkCviIVRm3siy09OMwRU
2uC1Q8RJjr/OEP2ok7O4nGtNOLq/5KK4gKXosCRYSozOyp8HSLIZME39Lc1OLhmi
Iy+H4M4H3kseXJeMmSup7nU/4LCPQ0rL5RS/cRE+ivgVuINScGKNuWCWrPS1HIZC
ZTcjebZQZB5GN8tf92Z0nfQxH9f/w8Uoy+NUEpmH+DQuoYHt40di8tYh07CxlsGc
Hg++AnLCEZz7O+r/9GV/ig4WlD5D/JPJQkVK1aXxOoZxyXcv4L4PyZTvJKh7iukP
XaArgj2lHYI9OXC4upeAAI6LCxdiEPz7AcaaeZUOThxV0SQdAz1XA0dLhbkjrctD
QC6yrfMzZq8HxaE54+Ot1N00BdWlyPMwsSR40yRumrbDpFHzB4eHFtju0TZQSU5i
6Xftqvp/dsknyRHTmEVHH4rUvWPT5A4G8Vv8s4u9NBwZ+k9/0k/6MyAFQRbNIAJ+
1QdZmLZG+WHEqedpg0gMVnr4/1m/F3KE6AkRamUPjVH6umY0vHZ+TLQZQ760zx3l
q1qTk1weT2oefYZty/aU2kdjYGA8Ch/ZOkVFl41NvkiK1ckQd/lWNOtsF4NZb3Jm
7bCd1sRKYv8HCOYES1hdTHBsYFnMn3EY2W1X3P7V3nkNPQ4KO095nYFgoH0f5bMC
aP6TybjgtJrqOnhjzW5hEDKuMKrChGG7TkPznEXs0bmYHtWrGETNAkbEIjk5B7pu
zy3A1s+bXxtngqmnEJVbVji5U5y59siAiH5dszcQvgqr0luECGnPr7vgJ/YLSGlb
5gzhoiEzGg/ReaCcenti4XJYnCSC2RgPW5XsOI76sGwOAEIvpiR6P1p3OZalKCe0
5YD5F1w8wQxcaUu+OfC/geBLE1m04sJH35b6SSQ2nJdJJ9E+ilAFpaAt3KXcpTay
fWUbgXtjog/CiQw9onUpxaR4kT/srLqSXCQaZrZG+Gx/qdsR4aCAHzfVSWjaOmEw
KVkw/ai5K0nL1W2MNZzPAqAtYII3RDfluSklEgID80OwdhmkLlXz9mmU8kOj1TvK
Vo6+SWpRhKKiJrEvm7fSziNz6leWxDHkya5QglWA5jeeSCGPUqVVrX8K8xsEL1gF
obQ1nHVwzRD90uhJXK+Njn6xbO2IeILXQQvRI6XqUkLqTMkk5Oa4fFNob7ScDEJW
riE0mbJesmkyXAGJW/oDL13JuXiKpvUI899BrANiIEHNXRKsjDpKgYUfrEqP8HiV
eSyo4aDGecNkDo6tImwOX1m8doQhp1IJ+cSIebeENTL7AKAU8Ntfpn/oQoCHQ3kO
Gf1xauOs86hpVObMypSeF+zW0y4tCln2hZaaVp4euIXGHTkBym/gJBw3JgP2J8tO
TTcbTgz0BzKZhpvjuuVDiKgAuS70V6w4HWP8lgTWJcUE7DTIE0E25niXLpW2CRYd
Y15EwYqOfGCIyfA6+FTCITtFWnlAC4Q4cvlyMMFZ5UpzlN9jbyEa4+2V/+kHNwjJ
ZmB+VwOG9mPARx4dwoi+WcwmvmuCv5KUSLtOAaqcqGlUkESIGMo18nXH+AWioZLf
eXAXHA43K8YTk/wGhDhsCPtotnvLhRA5Jj0aJL5HOv5qeUYA/0EsYL8Kr7Zj+CrM
jVu5hoaSyJ2TuaMwymFGTx6nm1BJgFvgPlzSyWiGjjwJW2xFVpn+GxB2vMOM/dnM
NHBjfRivHyyj4SkELtOdSGziwQOVUaShZ928wpaRsATTE4AUNeipqzP2qly5LY7H
kqfv9JQCHPra9x7JeplRzQBpUQGvDtMr6VAAnbVxhhCZtWGH+mVf37ED0YNneH25
meUGpCRmIguQmtfg25o5ENIGaDNASBHluuo4p43lN/pJ8BjJ8hVXgWKxpLxF/7+G
gb29/9SyXOtL8CbcZpPfAqRLRCLfsofwwmnUWbkFvMrFG7Vvj8BVTOOkvzdNvu4K
/V5C6V4GWVpUlY/hiElcUl5XUZrNrXGAQmCh9j3DSEQLkqbfdUOvnrJje4HxjltP
BbDdFbRRVw+Ra3RMTyb1Wo/XlYoWT0Wrmroa8cBMImXayTtaA1HFpV7bNjr0V8vQ
/s71OmQpNoXRdZ1LOnb0OG45uagyzrLAFLTIRd62LqJQ+PkaUEuA/csvPaU4YSI1
6Gm1YYQaUjEItVRgDsANWqUOp1zJTW+jBBmoJ6rfmWtlsSB8Ki7K2PKpc7TsXKiX
CwVd9PYTsmOFn73TDZuZY/rb5k43+BOP4uB/E9KFOUkWER3bOEnlg232xaVjDgBd
51I1st2dLeEe9eSBEjgNkQQjonnmZ2V99kfPgbuhZNsg5jO4qGZDVzfn2EcbCXVd
LIZMxZSprW/A4jHo3/IDLKkxfMXK2T3EMQXTR04yGYfUS49ImfftJ4FwV/SWIwHT
n9foyB8R9d8u0wyTibKOYIEta84Ybx6NE1sFKTaZo98/aP7nFgNyBTA8/6H5rg23
d+QQnTEe8kf6VUX5iaXxq3v+RivtgLM1g/meiWl/hhnVhTZB2PhFH9kT8H1JZ5CJ
rIVwpJdMosdcANOQy0mJ0oN5Q24jz2c+B+m2SYSxqFwg4ZZmnE3yyTr2BvSFjiDX
dROLbBP1FRQUtk6wigPY2gNB41/kr7cPBbCeVFrxTR1Te8FGTm8eONYs3mb6BPgr
xmYTo5N15GHSxZ9Oit1c33rCTFn60D36+zeuvnLJhoY52zcXg35MRf+xIQJTYY1g
TOUpqbITRrdgs9y9li+++uSBo7WlpC59yZ/e163McdW1kER8j7ECHuJejVr99eQV
2yoerEy9OGhukI37apwtmDXWpPGpr80oW4QM/Iva7UMHGUuwbwredALbF035jetJ
Ys2otMbF8OXK1V+YrU43MBzzw6jxvJjVltZXUtifImtXMbj/PwoMGEFhoek9CWaa
+CCSQjI8Q6Wtdqj3dDOvRrLAMyf6zfEjBbz41/3kkJRxhPq2Wp629ZKMmeCN/W1X
PBM1gzCRCHZWGNfVbWoQ5sOSDwz6gKdf0dA88l9cJWxNAEXHYcHQn4xU06t5x46Q
3RVqjOlnB/RxpGRTnHs1PmoD50AjKztsr1XSYXYBKh8VGG+x7NB3fd25lb2CARf4
DY42o66edmDYWjkph5lNCEv9yCUNIWQ0Gw2sY7m2Il9eBA0U+zkQkZ8V0pX9xpB0
QJvjd79Nlkc5SyHVbtuUqMX0aRoWiqw2tDhYU82YYy++2DWIAwv/BYQyOTlB6dnF
o4in+ZBpJ9Q2VHv7S8qNwMaV1jNcNQX3r1I9KgEBG6WiT/mPDUN3cqQ/xN1ZqqnC
CkqP2sA6cj3mrKSQtgjAVEdQ2bu4aM2VZRL/tOXNkIOCpu72WdrGVzYygBEmxB5c
gPNXXR5k1vWgLyJHu/veEMn3nGIcp8kvSX+z1ihlwoH4yJzU6FFYCYx7zeloRIW+
9fzqdfa7D4mm34fbnESzkL8hz9jUT2POfNSBLeGqHtl2a+Q2vL6IPy77h1lsQDgI
xpeqA7oc3BlDlTvvOIf0H27seCNNQMzLIbxPm0WEhEp84JEUoEklfFvxtjqvffkj
Ro5NDKdfNctUxlohAR4MHmhZMIa9XUoHscBVFXzEKYZ3lYjw2Oi5Nb3bYLf0GwwD
nchAQa7o+qM+6LhuQfI1btqKOYozJpuAVBAmZeZ36kgiuq1zyRDNIvgmvq12CeHI
GGEmS0q9sgijCtYXIg4DcWcM76Tkc2Xx/E8qY7Dgy20gya1KLOBbxT8fo+CZhu+J
jInhJ/0Pwa3oOo8WAggEGC4TLRGC2ul2JmTwB/eTvR1CGrAryhwKotljn9R0OTBS
vdkVGtoDLNeYKjDITZR7XQAmNwQZAeK/vE3hC4DSwIqAg2SedNmQb3roPsrDXbJP
GYb8XXv9c56HqKFCKxZiwIcNNbhdFokhnVAWb6Ig2L2VLJp/iQJH1GocB+00b2GC
23SogcUyFblgrs31ATMTGizh81ptdYgyoROrPnnAVXAVnhx7O1K/NOMkvQJddSQ3
cPb1Gh9m95ZDTB30DzVnRxgFqgxGqZKux8sYpNjE6O0KDcSZGDLhh+/+FWCTZ7wZ
p9FOcUE4fYRA0LX6dALwwiPScpqRBDmRizJdf2LeYIEEMh9U5dFfrSbp3sjLzjoa
vLV2oBiSg63oB94f5YJkPESyrzzvBXZml1YMRDNCqZEcQ7xmKIKnuPoi5vhWD6ZZ
BdapGbGkkWqq1VyQwQNq4BmP+7AKY6b/QIgkjoiwa+Cqzj6eMvzn7N8oybaTEP1Z
ycDhIwcazhVxB2OgbuEnqNp6uFBpEGMPT+l2qewUcQTt/ieaBH28324uGrfWh05q
aFzIeV0Q/97F6PU+uxl4gqny3lIgbILWdqpqQ5bmoth8NNNguEX4q6C/4hmc9PMM
Ki0zD//jAo0HEhyOnSiuY5PY7p7Ei1+FtTwzgyVIUBezPIFwBXF1ai9ES96HGITS
KUZxhhCu00a4Mall7BNCTAmc9UCBNbCoBdvfujFSRUXhCS3VyzhElqxK4lxBDzzK
1T+JsANLVe0N6SBmUFx5CJAiVKZAGCzfhYkmENNwz0gAP70MApPPPK9JA4dsgxs6
bEQRG/0wTsT5dHs9zvXQeK7j8cdgEzEFUGYBI0sZ5lYGtTinheYLSr4Jx7xNFD63
fPSfWa66HyaIW3kLjpWkm+CEwEPv/oIEAcmT3fcq8fzL/TyGeV5MhIq/fmmcfwCN
G1mHi14ZWMObzD5mzY5psjXs3UAWpb4fByV1eT7a3QUR+iU5mQk48JkhZFJidtXt
MAWKbEvnxP/H110YzPoPV8HkZacTtmlgJ+yfP+h6eMtRN/dS/4ghIJGr3pP15aEj
iD5Bw+iKTf29lDyuqUsxMj8KthojINPlyC0w7NclnZtSRGqqYcm2cp6/7MrP1yLd
22Vs48CRXCvFj07ueYTC8PZb5541uxHNh4E463IRE9v0h7kl9TaEnywgHKOoVigV
uS8+I+M2XBkOrtb7hWr7In5N9VcUcIEu9k+3Pra+sJ4xKBPNGXoP0CSsxsHDQX9I
bV3PZWCs/PKtrwZpJeWZhjkbHOTzxRK1Xf/Vf2G8aFiVSLA5/EMErS7VQ35Yn5E8
CnbPQOmw1nQAT+ECc2nG1J6dyXCNMDD5/41gGqDp+ZNp7xlWUkklspHYu4pe/RdO
Kkg1ZhXTcM8pU9lx2/F8A9CndE520YDGJch5ts3CDbhTsVWhzyhG+r3voElMndSd
H2TvWYaNLq/trJ57KLfsNBVgJqetPkPA71sHMOHMSdnecCD8zX5s4oRRfL9jtFIl
OlvgD6u651/HrI1uVvqEU2NP55nfB+GlOKnpRRtrO4vYZuxKLtoVTwqypbPYaSgr
sgprxsuQOu2bwmYbcJIcDDZJd2d1tDFA+rDEV+RGLVzhaGzTMfozttVwv5Nc/FMk
wKXlj2K/lrWtdt6BhSyIMys7FrdGklcq9FgskHXr7sT27xxxjcw6i4E8DczY/+RD
hlhPokCJ4276oOJMIgMpFxAxHQlykHJglF2wvI+dBmTDuBdwvbricLXVsVTWRKmS
5FIVlDDDG1rkJ+vR4rYlxeHQJCanqnXv2WBc5xzzD8+AT63bmXgbo4AYyYABRK4w
Yzbko25Qd1AXCBckkinHPHTTSV6svKLUWkxrgwiS8HPwxjyxma3rUDJm8yynu+FK
V5P0ytvwByXNZ9foWBYiHMmKYgegClZQhkIQItC9qSKaGZPkvy3lfx7uKNNP7uBD
fY7duByo/LdPh0eXsxD0nVjPzeWMp3HVE5x4qBfqBUYoCF/IT219JhG5wdc6Fo6G
7c064V0jLeJ3h8YitnCzmpqbAPgJHaDQMjLHTUxwTL7AUv5leIqiy1rugwEK0cX7
N0ObnKEhI7LuuFtvUy9bvsOqG704QNeQsYBnFvy/b5DSETBWnKmVL8AIJCHZx7If
sraJ8ul0yw76y8P4nBAnjWrJOt3+ZBTQNB2C5FdPcpR3GGPEi4SRuwEvVNakWQfU
95reyMfRF0ew52rD5BNGNQYo/o4cQJtZYdHBnohXc8AcC548Ft5Xt5g8EX3HeHfi
84pFcmJOlxl12AzGNrEJj24y4GWCs4vKiAJ4/S/q5bfn29oaxuSt1WSR6I3lAOFd
dA0MDCeMGJfKBIJqxN/78VGSPcPxIgJ4lRxtyavt/Px7cjWAJx0MZclL9CcemfNd
mOWye2XheDNZ5+TMFCTP+D0f92KB4GawVtfYY5RGb0noWv1cuJFO3vBJS3z0VO6P
Oc/11Co58znm8krQKxWUlOWY6JOPoNqsILbnZzn1VB+6GFXPV53tZLO0C7BIJq6m
Z9tzQThNaEb8Zf0rGVXhMpEBMj3HF3rJaVS4lG9jZb3Vg0PaD3VemIyBdYrtG+ws
FItCmT2O2V2nhAs2dnR+0IX9jN9vIpNopNJXa+NQqkZ7VCXtTo6BmellnxhYplQd
Vw+zA0APbUwVKpn3YOaOaoePjL1uVXNJcv/s4UiDOKR9FN14nSXA42eV08GDxFdB
4hW67w41AmVw3R8zjQx38wl2Up5pvYiuQsCg9ZsmQA5AAb6XLyQR8z1/gskb74q0
5n2Fi73CbegQ4/fnynqMZ0dSCVMMZ8xvjNPnFdFJ8EluNNzolaGEp/5ucc1zn+Yo
GTadey4lj7a8kcAc0YT6ohlhWaSipNbmPUd791D3xz4GEMm1Joty1muWC9OINPBi
oCWtGUU9felIh1KKpxUamBspkkK3WN5tLiCUFezLQY7uq/3Su39SRFtgzMzL+P+r
D7IMq7O32RPIIwxOa06ITHADTWVD2gpS2DUIbAHgmqS41eIRnmnOT0jG2f7F/rPX
cMvf5KgMlmzLfYIwrUk7hfkjFZGBx+urqP2bJzjVgRFu1JJq5dfjldl+QhrvlxUA
9x+ypjrklmpbEQGhBsMRikw4iQjFBpef+sU431Q42I8dt7rN7BuWg+4TmOghazW7
NL9Xj9YEDXEL/fxeXrh8gYr8lRbgDVYWPcbUJpNA9sgWqw3eRiAjCNK9V8IRDVJd
c89jijejxcjN9T3hlBOxjsQTinWpJNTW1ar5oLn7duZ/5HiwpZ8HKWUOlUpRrb6C
lzWHri3nv1pxMO0ZGX+0/DC5HcLmLKVcJv2h14ePUQoVnmDrcKFPCw5lmTAbzkmh
EScjZjsBnhsA5akS+rRAJWlqR0fXGXqOBQ6NR61lKe5dz5ovrSQF6oE0C1CeazLA
hznVeNxYr3Af+ZC/EeT05pYhq4Kmvf0McMnLhHJgXeqPOWX18zRwMBAEBQtO6otl
DrPrZD6wnANRf7lprO19+0xCG5b2UBzVnHHZqtSbSZMQviNT87SM5EwH1LQs45Nv
saRYmnG0AomiAq0FMa+olQ5sMR9dh9ZK7d59oQc1jeaZct0YeTwrJqWNy54CFUdH
jY4ql4x1XFNEq1+kcDYOHh80SFzaBeP5IHFawy2dDVhUAdSOOFIefJobpJVSNpoe
+Jy1Q3PEi8Fos3l79naNC7WVgmx1gyfSL6ox5btAHlmyuVvHMxSAUOPze2MU22lb
vFLnN+XaKgGP3NEcnzH0wAR3gk2Bo3TbslPoST64K8z+QEShxyalG4xcbt/AzQ7A
TJC6W2fZuLTb6e2AhiYhWeh9GDXmSZow95jnYG+HT3OtziS27A6Ew1SDmUlVf9vP
QUVnvkY9fWPLpoLRls0mDBzKY8+WxiqaSzQK4WTAUvn/ref95a2S67nxVbkIZ0Gl
i7g3WJgo/YlOoTRQnbrddvmM2W5++Thko3xS6EdmoqMuVGuYqmX3oHKbx86mTaEG
T9DGec+SjvOJAFSAFUzjMcmK2MWrkOSgxHl6L9jakqAlVkdWZ5p8Blw6A6P4m8oV
V6i8cwH3cXaFBbUsgyKDXa5i4f4d+z7qCXTU0SJlMPR/cHOzWPfmXkXqCpt+635m
TsBG7yZe/ie6zvTGLdfstWFNVKNfUQSGEK4UvST3DVksPQFmkfGEkA7J9UphM4nF
jQZfZS34uWCwPuYTOqks6y1KEVy8eLq4i5vKd/tMZ/AZ6Cfy7qFUMD2owV7y8arZ
DtQ06lcYdK5ZU1vdVrGiZX3HF9U0vvCduY8+IwJnZrZb3FBFhJRq1VhxWPNADHPd
VxmpoRBHv9TQQD1bU2uk9C26dDwVHtSy11MJ7osq2whfBr+gDWPJ/8pajp5BbBCY
Qlu4Ql0Kqp+I7yHn9KsaqxHhs++RIKzj3g1oMKm5RHZA4XMPovF3wReA1+6dijEZ
e2lxTWkE2um70HpT/DE8nzrNlrDZNeSjybdErTmTR9EEypYKmrvgmPZKArlbxZ1V
dF8Y5z4OSWiKNtOUg8BqD8sUcWiGOtKmV8k23SHXM86S0g4/Cx4m2IUntlNVaVsA
EALedQhA2ANOXI9mGzt1baalvZ5WMpjSs6/K8zSFeZlyskCSb8c0U3aFX/nNunDw
w0K3e/UkVIqI+VsBxwyX2AEXYzf0r9z14Mz8yzTfCSrzVYSvpqB+hHE/QsM7tgTZ
UPUBvbKOgc4EffS+FHKT6oWrUFHFhIjWVE5+0NeY/W+ySgOi5qY96EtZyY6B9bZt
rJATmEW+7y9cvYtf9jmBgrDRMR/f5nuF8cQ4qLQcOpOb9SakVy0i0T4x8kxc0g83
lVWngYsBCGqE5tg75/m4lwtX5aAcR77/B6ht50KyVqyWtf38/z6Wv1t30wDPazTN
dQZoLaAqFsd8wrpQ2vaejpfiVOdLWJMhhfixeV0MlKnoYuTNcGEuFSKAGsow3vHg
9kfbwZzEALmqtp3THoxGwevLhLwKqU1b85UvBXpsLA2t2flNPFZEVt+m+QdO7UVA
df7+eciRJ7X+ZqgO06whEGZ1xihUoukZvh6ipvv0QcaTtMjIvvgsbAfE3/ja4Bx0
SrJeMwCUvOw2ahS86ch9/6grA9rPmeTD8BVQnCjBuL482SJBRAVMP4os1GSnnPBm
384TcyQ8MRC3hkXSzLg71QTRVtOld3Im38A7OBp3hEgIYY4aiHBhPuNZc+LajORb
LpHEResqNzSDjFIC3HVsP8eVukAw/2jeLu3rAgvRPYjIvriDyMSSH45qtx6xd1zf
1qXymAfKyVrX0/YUFXWOqqDy1qeYVY9IEYyGhLaqdW5EGGHYWtYT/1VcvJqcBnUh
D8smrcsiEsQzPqy6rIDzLPDSqNiLB87T+iMVmB0Vn0NtPS7QAG7R9d0v85v1cZYb
fsh6UBzOpzdKfb5LBfTqOZm9ntM+fWQwjSiR/8hCu05QOTEuUGEb8Y9cCwGttqSI
YE7nQiRYWZ/HzEIqHIJ5HhIMmMu6dbbX4OLlzLpfvzkrJiDbNrvuQgIUSKFoTMxw
5GEdAHtOHtSALMlVCmNLdT7QGv3qMt55f1E5SyVsV5q1KVDMnR6PTWopB7F1htHi
hjTDDFdsTlMzJYsaW2tw2XS46UGzpXXBlQvVzrlKpVq+wsO2PSOmKQydyyrt/xSM
g4+WDM4G6wBjyEZeEViNyHt7Xg0aLWWnPhr/TH2Ghn9dqaIUiW1d9cqDbDAGOsLA
EKlUiDsCuTcGo9iMDGuYGds9ql7eso6GiXDMyBq8L1r6YIXIvJQK8xdZVlPMW8pO
6UAuNacn0/uW7g84gl/8iFKYnuoA1ewbDyz1RkNZrZ99wO0HR6LNC6O968DAPwC4
iHyuMptpAmmjxrcrzxwPOTmF/ob597w0vzVtcDMjwc1pqs+lVGIHkxoBDgsg4ORh
1a2/WXc+dBtbV9vrIX9ku+0gDX9+IjoDh6yUaeD+wCetRQs1vjjj6adCa1M0zKP9
41B1nQxIt5chehwi6SQ/e7vmBYREHJmk1l8lLfUa/PyGS+0xB9JnRHxiVyxp82xB
qFOJksngFDa2cmt0c8tk30E5N1oRPUPKudKZMM3E1g5TRh4snHYFrv3o6BcarRO3
ndUQtle+Yqt+n/4O0nBoOcXJAAKeJLkk8y27fEBbKz8wDfqNt7eQ5zdIXxWD0tnL
iMuzZoj+Uj09mMw9RWuL2qZWIHcwaqEMkYzKENqj2PhVIu+up6lrpi3pBkOlTChK
Ke4d70fw60LYTuNq50sDndOJ2+pKYKapf7fdnig3pjTpuEYaYL1mWYRfVzS4hdJf
oG4DBYuxIeavlxooFIblhlu+VzWdicHWy9Q//Dj69r3X6dzDdzA9GZOIEADYOykY
zCjVEvp7OBs/kvRk2MEZPcJPfdwJ7DnkFF/eLQ0aPG9QxSwQv4qDEQJyDFRfjQ74
IIZHDnk36ggw8BTd+TSmt4gxPjTcsOhSE9Hc2cgPrcCuvwP1r1smT8IpT5mxcCCW
KXY5z/ZhmEDBsMIJF0LJWx2hnykgXt8iIzOqTne990ahltiOjgA9RNHF8yGUuv3o
vLl1rw84khW+Zj2AU3RFPQF33R2QugIyQ88G8H2KwwG2Rg7ZKC04eNRzMbwPiw5z
FhmAFlwPLhUw2oAXl5zUOmrFjNh+JhNpx+w1dUbV2+ebh6snCtChca1ORQ9ewhc2
acGcf3WJVLH9QlZaz7GnLzYatZ5sLMLzwpn/KyNUuMJgIuWzH4UfmheLCu/E8hXE
XbbmwgryGNFRyPrKc5Aj6/QSspK9F8orBRJlmQYpN39TPoCfyxBRq6aTOZpAYF3J
PFL0e3xeMBkpbyip3g3A7hnx3pkhzVP4xLe3fPpwZDrKa9QF2k3tFHhfKEvKB8Wj
9+U3FoJKQc2gn47vwT/Acc10uZQNR+Fc9K96k/22uMzHFspzVag9SMGSqODyBI1X
b4Wgtfjzn9ssrMbZtlv+rybebtyygtSnpl9oLXIR0q4OqTK1aYqiQNsEfR0JOkx3
zhzgFR4IBk9va5slT2jR9Rxz7PVUcnNqnIgG4ydU4DGg28VlW8P8LrwjJ1HjmZqj
+2ABD7xthk7yiO0aKK+sBY1UUG3IqkuStHRFaglVGM/amdjl6kxj4CeeciL5iAPC
6bdfc0rIlcY13PKlwEVldWaBraqKu6fFl8ij8i2XcK2uBGcVptUD6/xWU/GwDqCw
jKfWsoBcDginnzTrq/lp7chpP+VN/THtOVI30tYCshkI6pShJztnBRxdWAhVf4tz
poeUxxWMywd3CB7FLj1W6kQ7FqbAWdU0G8hw2ptXlbyzdGVeH4O/c6YHcG52o2/u
oXuNAEtgw+UhIWP8Bo0cnRKKPT03ofbSyTkijzdtjeL2i66xWxyOg5FhqtVbwX0p
vLPTQN+fQs8LnCwN8PrM7dVb8Zp9m/+AhzE1j3Vpl+JrgCh821wgCZPLCYakY7ht
nGlisviSEjxk3GTjTgRFJkLKORxtQSah2ZEk/TiDjFaEHowUzL3EVtYYQuGc95CT
WIIYPSekDvP/pGWqwMlcTqXBQ8sKlzHw7Q749XO+8G6PKKnESE4n39dwQEAvc1BM
8PhAVF9CHp4W97s5Dd9u6d/YvdRjh39xZX+d1aoXYVyWg6i5xRNywCleD+sMS6I/
LS1ZFgCXhdOGjBAteAd/0ACDHev/9KSZdMFj7goMrQJfz74pTG0WZR1UUbYm8FA1
OrVcLDIml6k8DI831VQo3traYSonR6qkEOZcz61ynAcjFm58FlCOFbQeP9+P69mo
nQMzCZFMccXYLGBoVyb7yg+UvSyKwkacRau+F69Mx/BtZb/SCl19+lUFNH7WOF7a
Ci3SSQOU7fdFpFc8Oi9H7JdndmuyZ1aszmhflvREmA/sJeokwGffI3j4bQNVVg/j
7ld3tfq/g972OtvehgGYPEN7TO5WP37fJGIkAeU+AN7zjG1gEtycl6g0VWOgwmq3
P5I3k4p0fjOUJBpKZ5ZPNUTW3hevuaK4KdLNrnSgVmI7xWzndk3cQVpF8coq3Aff
iaBYjc2o1L9PV5NDE0ZE6rrZZIedB3cNFQevGBNc7IoFGzAZungkB90z2+T3tFJX
XDC68B36XprO0n36eq/HpSmaNLcEy+ZnI2N1z6OWAaCDBk5c7N41Yy/aVHN0d83d
RhcLe3fe1nRk82arXR2YzNlzGP5W4W27ARYJRiPf0Sgrr5oOEROT0e2aNqhyruO8
LUvU3kYNYHp6CadFvELvBpHUT/dQ78fJXa6CMyf7XXNsLZ+R7/Hs2XheCXnHuf10
FrHnVuyeFwlgl1KVs0rHXDYOEBlHG3eNsUsedq6xjaiwFi4Hd0Ba1gciB0LYAqGm
dJul1aKWRKljCOFJ1zrZIUUPPRjNFn7HphdgDmZjiiNkdNQZ6mEfyka+8fzhnnBo
x+iHvPyw3ZwJ00jtB2XnTLQL1awoW31MhGWEmL9uju+y40b/OQiHBV7rEtpZgfPS
yYJHUcHv1iQ6wEPayM/RWzYxON8vPWoSbkw0oygMXNa6KzISSjpFFV5uTZ0KauF/
1CSuZkhzF7brEcjXyrtozsdWb1yVW4caOm8R0noCMCil0rYUfxun2uuvRilKxxXp
XpUE/jJOI6QBNl9263Eg2GPfoYmM8uvFeW8XGc0Muw60IFtCh0Tb3tksfQhsOQ4p
69FPZxV3VlB8gDZ0DUtc1pWuTlzV47tS6SQw4u7U4d3MKCil1Y2TnWYxvvVfp2BS
HZ4fsbEbzyHmg90lnhnrvWzr4LZiJDQxdkpxTHa/8n59SrUWgOVyu3Tz2XCdlSNg
QYWq7N4pgqjh5fOn1Ze3EONCwYCJXGb/Ch+AqWayjR1X13fGDe1pE0ureo4DOZ0s
dx2u9ovHub83UBWyhqjm2dOBNBzm15JRm3WkFTQkZWJXRkSbJkJHkWrYmI4a8bCO
WuPZnjgZM1hJl4Q5tYRw3TxQN4ybfE2h4z/vGYZ+c7SrNMoeCpTdD0VxFXgtYH9A
VsY8RfAgb3jHM9zyXEqBaz8OJanOpWOShX1bAcuRvtAhnuKaSPim7hItscUmsnsp
/BQQ2cNhFSKcDBnU+uTgWPaZxgE3UuzSDhlWhwSXIF/dFCgGqpeAZNwsBiLs/q3k
jxIY8bST6caEkCegZC0fgp7epc/uHpJdycgWEh9uqTB9S7wN27zl8qSJlzOR4hai
6NVSkjrQxEKfPQOFUFt7v+ryzEURRI/xU1AsIndR/XkNzbxdTjg2gaUgCaLenh7R
y/IdbiIpg+FKN0GfAmxmBsew0GNQ88CZppn+MQtoiTRGFcCtj7cduTR7EYuitiN5
wbQFGaid3+xPzmqkuWbcaNpfIyZD6B5jNMOloiq6NkU6fHk07Pn7tE5YePSQWo0C
4XueWRqUumN73JxNLWB4kF5tXWU5J6xOC7O69DYQ1XCQjunUUUj0dSydWA+EJ9bE
Uu/xPFy++ilGDKHZyI4vX0KQ9W2fXMBxA30L00yBov1KQQRK9U5OhKbOO2ab15aK
m1/7g3FqMN1n0xsFVc7KkqIeWfIW6mkHiFHfTiPLNYL1DiL6XRIRvNkUz378OddW
4FnbfH6Y7Z5cBAAM+OhXNpNO1Obqf5I5wDU0tRlS0DmQzeQQi70qEM2lckztK3sr
xI0FCxZRku234rnxz5d2XBRuRh1aQ1BYZzynma9Ue2qgpRV1llN0n1yDXyTcMv6H
BqySZhHGMvZqPQQcE1mwIxxLtAm6mDmxNIAgSKTsp1LUSdPdgJ3qLPyteZvSmyo+
yFf6Xtg3TVp9E7pnX53kb4xXNhDmpbO+l79JZx2Kt6nmL8g50OQF6JRmsg/r1535
wX7NhFbyEkGwB40WEZEs1musBfkI4v19QSDUnHr64aj8nlOqDCjJae5U9tAo55ir
HJNKG+oF6uMhhgJJp/PU345wAZ65cY7IbJ6YxBmx0d1rcfO/rdLZvBGty+AQ98yh
Zk5fEKF9F2+FniKp84kQXFTjdVz7poMqGnHo9gjzixsJXYcg9a2pHa5x07s3DM41
hP9h1rlno5lrZa0Z1ePrcPKDauivECfHsOXAdDwYROQMIDk/3tnzNP7m6mmYJIsG
RaHQ9bNc0eelOxwo4HGhHelE7aHbuVqo4UmpDPULSdmzk/+ENz4Kr8wqCAyWgavS
alkNsnmfS3kC0BsW5goHilvles/TmcRt3z/zFPIClOEMO+04lpzOkwZlvr1iaMgs
8rZE3Kv4XclOvfvtbBdqY1PVCMDCQIfAyRyq9xvr1QQ7E7SrGSUfw9hiNbKiqlLW
jhrKRhay6l5ei4EpVCw+Sx4vqNArv474zkHaOfQnigrh0bo084Wb/IAEGrcz8/Xg
iAiTh3YYfWaodNGLZznHcB1S/aSDm/7Tp43/TEGQU3KVzPsGCr81gt5uZmS9dk87
0T+b+vq7DBXPHN/W558f/KuRDpmBx+WbkdYa9xL/gAsvBFpZr6IFYuRyIHmAJmSj
zSFiU27SgE5TDuXmxa5TRSa1Qe4kcDoKFScswcBYHQyDf0vPUDe7UEWeR8txDcSH
oW6xOmJOTIWcRSAeAW2/WP5tMWV+qfv5PbWioi2RvdWKiSECHMUez8d2/CtRRqBT
hLDC3YdIfGhlkdp5yTjF3yLhp0r2IxLWpReFjptQNhwb0SunwLiD3h7Dd3pYc8Ys
eHEQHdYjktu9F0kJyTHyD8ubpIjZAIfoC2UrOLVZ//gpKrCGbAsXq60HGwvHN7gR
Ax8KdZHjuEtKboqRvRUAgskt1IuyXrPcamYIWFmwfGk/94g2c/BjokWVFkNPsG8g
JOhAqjuOSmYiz7bDh9rx7Gg1zdvXDDJRe2FtJR1qerVRKAZrO/M5cxRAntRmWJFB
CjrFVKiukku00uJ+VH0t0HktC89PBQr2Mo40uXXL01v+dbQx6x7tUkpPokcvnC+y
GlCECvlkGNulKb5nlcP1dUk/UdJJbU2nYK/E4bsvPAN3VRWlTZOArgJ8dpdnYxYm
uvWTT72KlRv+9Wr8Un5c7zu6RbjADlQIzAqOpA97O4G3IIUzhvEcwljkcvo37dUN
slxRpC73HBMMzD0nPNVg1eUPIYxjqE8sCrjvpX84pOnmOKKRG+ZLfaylX4V64IIZ
Hr05ZHs0ejqLt9XWa/6ufE7kpBT8wKV04ei/vIufpp+g00ClDvsJ8QrlcSjt4GnA
6fX5GhuxyVUMFyrATh21hBtAIX+qyDVHIJ+i+Lc1xHtOx4QI0viNMOh6EPQVa+pr
p3bZqarAYiBYmEJr8zZFWAfZBy2SCAyP26y1CxZkUyZc//c7A0xhY+PfXmMkU/vJ
78iEf4eeLn95Ai5S17iNeTb+38rF41dgDxdV/BL+P+T75QLTvSqxuTwDGUH4RLhF
96cgayhosJ/WV405HmT9FuXvdZ3FLpa2mqf6bm43IdzxBuzxCvNIzqjeXSm5MMXr
q1YF1LyMUvgcdk7GM9NEIfaZBqgrZ5uZfbfkbrVG+9OckJvNUL53TrNhEaG4lDrj
OfI6dMqVYpORQgHxaF9Psk4j0O6pSe43JxbhDOvFoPUzjpBs82xhG2TjGiGecP8b
Z94tloG7P9+IRF4hg0XCsRCyth0TiA8NHi/1COCfkJxMrvDxik9x0lmhbv9ukzZ3
bfxwSaMPDPkWczb7j8Kaulq9gK5XCdiPykgbIU5tJ5caVtJ+Ww39yai85U/COwpx
vaZMpk/v/PspPY0WtFIkWCyUzSSjbSd/jNdULQN7QeaONKa8ygHT6+7Qlf64oD8/
pJtuzUbmPpF987heCmVXixJji0NLVJ0IFFToqUdMjyvjVBE8Dk+t6Gh1UHNaKla9
G5Hlc+1g0Llp20XBnfEICMBmls23+oC28+Q7OMZ3C+WfH1T+TeA78pyWHyh1XXt5
NjAtDokDVcxji9ZjSQ6QijGp2tOAzJvZq2gpPdlWtFVjedIUTWW+/tFs1ViKtzHW
WDdqy+J68iE/uE8JRvFGlXtYe0fyb0wGarL3aH3wwTh1G8+VtAxZuNcY5w5M6YRx
gO025fJ5iNtnTkIURYQaHRCi/fOYclggJQdYwnA+54oZy/HwvuUHrCsUE2KMntop
MQQGb5IYKVtt9+7LdLM5Ety34/QRVOst0ssQjGcvf+ri/qg6Ud5kOYGlxXjJMHCl
aoqkMO59m1MdtlH8XepCCDXSlVLAX/UAjUbgAW7x+3jDX7/2NFb3Z4wirfzI/uz4
Y8n+zgkmW8HvNipaygX2ZSI0VMN4+CzgL08TzVOuukaknseV7DIJf0fBJYZLVwg9
Op0ScHCta99vFaUOX7Et9s8QrKjdldpW0u7y1WbKSJRL8LD/N/DoSP9ddn6Qm3ye
oZM3zUr7RL46bZT4857WxDF7zmgMudeKHUClnzvDbKhK7gzpEyntREdy/JXvGCPe
7Cv8p2NNUoTbD+v7sH7zi1TXd5v3Bpcygr+qNblzWfTUKyBaiBD04xHkm7zpo4KN
qairAZosWMJGNoyPjGP9mtvGy8AiRCEtVQFDqi8ctXfyOYRHA7Z8N+cVkBlhkhBJ
/UxwIj8/UFSKIwUFGAWUZ3M8IJ5pTRblEUpozUNKrk6ZIcQwoo9o0DhzoNBz8NOh
do2wuy5ApaXd9Yihi5g/cTN42oXAW5T1sDrD9kEcbNFPlYt0ILNvT9rG3Ro7K3Lt
7S7FEfWYPj5y2tiv64xO7V0sTga8Qzxm/eSw/+y0O5YQXjwIYNBwbH7fWgdcQrxt
on0OEgWmVxIvodEVcJw5P+kNb5tM0UuKCdsg3be1K+exsTEnu4vf5ozM711YJff4
uL3tpV2Pm/T1K2oHe2o3ZQvYmcp/95voxwi0+7rsUwgxnNU/WF2fmB/pB+XPS9R8
tDHCnOgUkXPKuYJmhF3hq61hZcmdNmv1kMWxQx5GXfSrbn//Nhk5hsoqOxL4ckqb
JMAx/xSOnPrUMex+Wstok1wd08KV6agkkHJTrqwV43yT+e+JPQdFikJBe6Uas4VP
wBK4J6mNd3pt5RRlglj5rtnK71UvA4yyuN3MRYJIvECdK9UNFl1hw/5bHZgAN5Nz
umS0h/qyFbmF9R1xVaPzdgS+NP24oCD6Q/tCiOO2WVP+2aYL69io+2fQNcATLz3l
meNrSRSmaQdspjDk/fLzRSHG/RQwLeneNYEkUM/+pUqq8ekeA+cEs509jJd9SIOs
F77p+BgkYU/7SwmLCgYuYk4SzYqVfghGPZkl83aP0LW8GVAjP2pFmOGDi5MHSUlK
pFeIWsm7dclqALU+vmiuhxUKWTEcr4C+AjDf2TxnNzTL3F2tVNUiN6FxZk8y1yrM
ghX3gUCDt0ghQ+I265WPnF0qO1hFNCiFodqPKiFdv9nRTNmfjDoFkuAe6/BlOPXn
ZIR8lmagh2Oe2Pvd/7Gr+t2LNuFMfm1sq3Lh2TFGYO4NPM2QeRwL6dYxCi13HlPv
YngZ6IhBDyLzM/s5+snAEc9otmfItMbJucV2kM/Njgc/VDuz/zu9Ccmia8jqsAD4
WmQQBG+99xNWKLUDsscXT16sA4yVspTQYP0wZQe2T4m7gkv6bx+79k+T9vAgveXS
ZaccrdQXSJEJnipmJ8vQiwr4PYT7zhSwNeoiw9hCXuW21VTPeTuY5DxdRvlp2dFa
XxdMAoorA+5XVS7bvMf4LHPKaxKLjKpALB+yfbXHKahSesQ3hPCwnkdISwgMAuKp
g5t2JIKylcxc7raABZahMA4rtvIYfMUSYZAhJEY1nplhMRLLyZy0xR9LMEpgBqFE
J6Z8Nn13urHxHSZO+3142hZLeOGbGeAg1I9XUPXMRsD7Fj+uix1n/qUsZa23eCHz
kBUfmJx7BvNYEZCOJKDbOMFp96v4iSOtrOayv+w7JFbq8jMoEZ2W5s4VPK8z/sdz
60+LeCdnG/kgFPh/eLYPdKJyRFWN1Z4eo89ZAD07+9Ruqh2N3rmzA9ubz2GYDeiN
Tr6T1uA4HjBNRVQYornuyi0NkPJqYcpdTvPkyhhJNhrz92Glk5qjCZh7+BQ+78JQ
bpibQUfgXdPE56Z+TjAKb/uwmYn42gB+Vzgqi+loO3MGxmbNbMxOELTWfkqwAUbN
5P+wV5o/VTp8JXmhtK8sMW3qsAT9DPJgAURUZkVbfRRXjT71xi1HyW2MOnL25ORF
6jmVVazOGJITscZDDDWDhtXXzeJRk7zgsnyPJJjhrdpmIPpdO/LQ0SEv+IJszrct
ktJl94juozlKFBUQu8N1TAQx+9CKKEOvnQNxs3tkHdiySdofs0ypwY1ajaFnkKy/
tkc7kWRp1rtzV5ubpC8hc0ZWEdhZG9JAGJErykQ1yugaQJ2OnDqfqJ9I3RBD4rCg
LG6Bdq+jWwhRkHgSG7cHvWtcj0jxJ5azQIDRd/l+ymAl2sY152j4d+o2FghwfU4J
x/4+73F4Vo+nOTRDZwQtcCTJNxk8hpO4zh/807LsV952PayAXJFc/TJSQZeIfLdV
7W/1XOvmFkppIgElaZKIzIjphMaLcPXJRtYQtaLPXOptL4HuzgTKpyeEwKM1uBPZ
lAinKd6LMnRCbBYGbyj1Hag2UFoqeBIRyZwf+ft2GM8yeLUeoFyWIxonkKJ5BFKv
1VKZogSIEpSYGuYi7bLWdddc/rTJ1ftK7KE4nuXli3hMRM5onx41ozN8pufXyBWs
W3u96jewS+OxHPVz7qyS8anM/bbu1iuvFloZpGF7l0dA2/bUywhVSTO+fRriCapx
fGNb1CkPGB2GowB3qQhY5ZcnpBhT4LW60CYA3wZ4QqG6dvaTTUodIAfU1JyFgWJ7
FMB5eJXcEb5/mcRyRcVkt9jTmBM+FxNdyWZtJd1j9bPy/8bONC3GaNM9Zhq+4QeZ
Gh9T8V2pwmXV0DcFWBk4kWK7kgiwZkNbqlFV93KHLjk/m8TPL+710spTd6ujS8T+
K6OGx14xqzNz2MowlEh6xYSWPiAk/x9C9xL6c7ij+SJ+lPF2MLABcq8SoNVb58AS
HRRRy/m0oiDMCsH2ttbX0XmHGPwU3DwtbqEUrPZNgdbNFAWtOKa5Lks6Ut6HBfng
YTp9qiM5F3j8bBy9L5S8iqJch1sDreQ7pa3qxxJ3w+CrtC96TvfCEfIiar3H+107
TsxeftPBBnhHuLx96k8FPgHHLhUY5X5DUSi2A7knrlx99VZL2wZZhJHR/PWC5ghf
ZOC2vRCvQnLqJ/Mp6/WdJgBO+0phE3QIRmHi/8bvcU4qhvWPvE7Xi6m/oOAAT0bK
qYdV4/IX5KumkiZftznB8bZ/CKwtmJur7iiRng6aoF8vscBhkwFGiIxoFHIGsbw/
TWbKvsgJUiFxw3gQ8Gj/TeMDJNh+/ix9du7/L4bfDTrwzjt5pufzMwwxunizGQi0
VHmmfpsKSsF1wN/NNofM1G+hmmt5ITpfut7rDGPmcY3UJlLhEd3NYpQ1tLw3ZonZ
gadZh3gJunKeXb3aYQ4lonUIcIl/FBgsxeh18BAdSYxyVP9dzUfSx5uGy1//Y9UG
jvQO9PWdHPl/NmCh9Zcd65ba1/Mu76egheBx1U+oWuGysA2X+lTTQkvakXnmM3TN
j98FRXqByZmHHXNYE1FVJ6BTWhkYFFD+RlM0CAJtGb8r17W9OUDSi8zidW17Ctho
cE2XhL1PZ/a5QPY4TdSPBiiNxpd+8F8Q4wJFygT1mm7C4o50wJMoOnU41eoL78v1
fQsyskxjsF4I9ciY7uTBU9qFLwPzFhpWubg3/y3yt+P17xD2GvXy5XILXAbGxeS3
K3H+YdnT2Vk12p6UA0EynnyNPKrcdGbphWB2C0yHJZwCBOXh8321RIlozwFsucHY
augtmKjJ0BKPtnINxTMj3fK2u04QXZwwhF3csoM0MuYNkFUgK0gZchpWIV4RoZ9q
OMgkJCLoQybjgeiejOdWEWcM1wXaM/gfd5g2+0t1kt4ENQYJeIckq0sj7bmZfbfX
GjBKFNMNxNusrxfsgyugO4qvGGazmJl/VVFmurY0N166UPDNaAlYnFxNO99+rwLa
lm10zCaC5OAPL/PbdWQm9rFDscDPpg89nTBtfsiA0cF7sFAh2VcfutWO2lMfENnj
WiBpRm3ZJVp5l+BUwygMjiWSJtudHJPdVH3HwOTFkfK8pZtwPlNuAQ+Oy1oblnk8
l2DIjxucL5dpX9+QqiEixwClrQ5pMfGKCaCvvHgmdTpNF4mQgvAZjTIzzFL94/qp
+vbyRBkqXIXLyeC5xK4pg2U4fa4DrNcMAOhY12La8n+09LawVMxDneJQaqT4VpMZ
npVmmW4iV7sZFwtzP0ouOrNg0UGHN+sj3xw8xDPOFqDbYmCFz9LyKvZ5Nmf4bQu/
1fqbCMq9snivwvvxt09VLaJ2qVw6FOnRta/9rT0Bvw7l9PFDd4Ai4cUXXjjry78J
9qmHzOqO1fb2JxI+9tk0ieyJFK9+YtMowcx2sQ2Z+rcY/PHljG6gpgLRqrdc3Aq1
tSHcG6/n81iV9a1JpZj67jpvqOm+qy4cq/sjg1WmUGi7j9qiAN4ak3u1GS8E9wze
l9I052XJuvT/CHTFiMLtMHWVJ/Z+PzvZUkUKzKoKZJwekJ2cnYmuAkKCSma2YImk
ke/4FUypfnoU0I4lgkYgCXFKYA4/DgC04oPYzqtXJSSdreBeuUee5siXfy/0DrZ2
bMuvED8J+Im2cx6XltVNqRcjDluHy7OgNcx4AxqxYtoT135If9qfZnMbikt52ygn
moYq7fhveMh1ot5IRz1FwhiAzWOtNM49hTjeXPlRtKxqOjTTXGvXbE86GpSpWJdP
LZ+592Q7E2tPa+IG7znhdwU6DeV5O99B/J5dZNzKL5d6L52zELTRSqs3ZJZnW7Zz
JaLHgWJGZ8eQ1m9QMQx2FXbR1DAUlW21lZISGjXoeo0HzM5HG0YZn/coqUEoXidm
NnweGOPjHXyNTQ5sBCOL7yCcPVj6eLVpINmm80Nc6da05HtHRiCw1vVB30bPyNoe
DmySUSJdU6lVMbQM9pRm1z1hOaBY1t8eIgbQQyOLh5BVpyK+GTZahXQiPHpuNIp/
XU7XPJqgsRshbe17FkhcYwcBzquzl3aqXC8QLFXNOtUVaCQfNiYPrNkc0mY4ANIK
T8xF0K8IBj9o2MQecc7pjGWlJDRgh+UpxxRgg47ve7VZ/I++50Y9UQzFdYdsP1kF
IQLFnUiuSZNZHDftkH6k6XYT9zYIb/+ByEsSq+jb8vla4hoX8e5wcYZJ+t95CMPz
yMG5eFbDllfzJGloKagKVz5oBQ6S8ApSGsa5Q9HgwRgs7h2nOYIY5dCfBmxSgtDm
IWIYiQgjpelxVwwANSbWXgPKcYyODGm+ayC6Z9IiSugcb/A7a7VBxnafRJ0vCKI0
F3ypTBwH58HUW8TGENpk5r6vIbcPh5MxJQnK+xr9AHvp5vk9AKcom7aL2ZLQnO5g
s0B/+4yMjQvFD+lK9Ua24ZzYEab/veHTdUiEiZ52E1RST9GPOppyWWPCKBUnJ/3j
olrZDRS1xDHWhr6k0tyeCdTUfC5CeMsXvan382CDpoHDF21cvbeOFpY3PAd5hXdA
oreo9X7WxOKhV3B6kw166VZ0eF+RjnhOVy+RoDUdYJJ94AN8ih/njLOHqWqrpPDD
XxM64suJIliVIiVrjSI/LgQaaK3iQ2knsan30r+3YUY4OVUjQ5a7E/F2sl50EQA9
BNTjtEBZSX5XBs15YXwv1Jii57861QE9XP1YXkH1De3a3HOr35gwL+Cwz7Bjm9bL
Kbk0jByFrCc6fIpIbJSwmlz7KBKAsu/kMHwnelbUoaIjr3NHswxPifereu3gcRQs
L9//57JzBlMpjvl27nf8c16QNMvB9BnSdytthnhRPj3DKBv2xjKuR9wzjn1Hub/J
XkSiewZnX1tnqQQCSMyOF66V1BO4vIBZ+C/6UNMQP+5YMiapMAW0yiAkdUd4YFU/
sTRtHpQmHyN0cQznyE/YWZvG3ygKO8oohuGDMh5uAxN3aKHYScSMCUfTSZopqgZi
1DDcuKYJObK8kPJLjnN02OrUV608YTeG39HFPrjRgR2J4GCyi3yL7nJ/7o0YILC+
z+w5ZWI7lpyh31xKj1/bwXJ6co8Sx2HSkO8Zs+eut7JgnJbjGXvaLOIXIJgNwWjO
ucKNrOnjsdR+FHraaejyYDp/mzxMZeUhE2HfPPw18Vn4y9cwxCcySwaE/CbCwWMc
c1fTNqKAMIiVBEPcBMt8+KOwLK24gyJK31fzE6Kvl2tSJjv2ESeH52R6j4PnD55f
NSczniHPapMzKrcH3qyA5H1K16ifC7KCSidBI0+QX9/QsAoTB3xCOav73ZXa0iUC
RAVtBH5070JufOsCdVFiErm4Ka1FtZVKQh4NSR3V+LJDpTMGyiY/Xyi40mQMqb0R
MIELQfypaRxccGMesT4dx9xq+OxH3IxfndhcJEOBMiM/Ebb9Ln5ux+5DEJN3D/rE
LfaW/VtSWoVKm5MUHmzPD8bGe4E8g56X6tWOcOkp3nKD1kO5VsXM9+Y8KBLG0fsZ
Q8HK3dFATIb6eBdAOHozROxRzbzVpz5wOQUS2cMfrhX57sXOWtM05DR5mmISuTe4
miprJfn9uIhxyVEXPmYUIeH0o/f7cZNLIE0LINJTzT0V4xavqdumj8/Q+zEQg2IO
6x/LrygT90xnFaPfWQ05EflAMePsgUbmGSkbwBHKam/h8c9GuhbZZldyt9XaiirE
Gx/x+FdmYHorJQeRbGOwPW3oD4T+xw1qCj0UZK8B4Od2WPOENz4rKpK1KNEgiipl
nbMqdm1uv0WqZENyVyIcBzfd+kpVILikQNTom5jh7BQsXkhA88vfRE/1tnyT9/6k
UyAjZKrF/E2A6LkJ1vMq9IlTIxtu4Lf0xj0bP8HCAQ980S30MfK00FvkSUfhk0W/
i/EAvj8AhA02pLXHKSgoJV94EQCELZbAQ37XHmVZzVfJgKq61qg+2IDeZeee7YIB
VTD8kXXn/ZKNmMMee4iortbsVkRr99cgX4KxIROh1AFa413NGp1TDwWF5q+yMRK/
YNw4nmeB++8lZesxZc8QwKSxa0QyJ4+RCdrhXQIjbvR/8uO8l3OqvjdPhCIQNOLB
OKs2ZR0uDJ8KLZy4Q6Tuio1aj7NiSfjKx8usYe770JuiUcotUjicjNbkuGxK0lT7
m5FHiUQC0GhGBjm25y45ClJnkfFou2Cw3JSIoluuJRYcpzLRNcPc/ycQ9mqsARzF
WnkkVjllagSFfOWk3jzeN6bp5NdvR/H65s+C1wYGuatv7UzRxb/pyJQL7CdypMA3
oPM3OZJIf4AVIfWClSwfFRZAq71F9LpxREbJWUzBA+1DcrmoERS0xWuzMNNmPOqx
wBREUEMSvf2PCn4WlsU16Py2vQhtrqkx9moWVjWJt7RAKRTJkfIcmY0PgDxI5IJR
hIpWzmfgfe4DMIuAFZultGeZA05ddiOH7liQJK5b3ddUcqw79brjI8Z15NCZjuLP
0G4eoiRifQmdbfS+AJYdzpqebpufiW6QIiiKgc6nR7VaR8wJt7iJY3URp+rEUcCy
M8RgQ8MZTsdWzMSPJg7fUE2cCvHCZrc9WQrbFHfNcL2+AqdqchA52qYi7UrGezk9
99smONtjHQgyaUO0JtPZH5yzbJ/LJy1lpaKYebWRNvaBB08jz31w51PHFv7ByEvm
5VOaf9YqzdHcAP6TLPxsaQbWN4+ItR8V1uCSGpJiend70l3LyX0m1HvevADHI83A
9bkgkHKRxVL0Z4Md77quVLu+jXBUeR3TqOS6sXo2Pj3KFXeyc8qm1vKnfNYxrLbg
lTEYCJ3f1VRG3jEk+LF03KTWTnNT1HVsLERaU4RXyYlcwt4Z3NOYZ94i2+ZmZqbq
CdqjOFE2jiTuxa9i1G4QPooGo+khEYpr+vsw5f3mlJrpaGcP6qcNpJ3Bz/p4wHov
CtUaVAJu/9ylam4DoD7XIJvro0kJFzBwLSAbLakXp8/OhoZ4TrCD30kVUSGCzLEI
GjOuRJ56l82HAzWjNwCySCiNIwBkf7dfE9gKipRHgGvrsgmUEnB8Gmi75Cyyd6du
U4di9GbcK/2khnDD2OAHd9knQmpq2/Y/3NomlOvgYlEaaDFehXn9X8QEijfM7VnC
7v3EnCARTY//eubnj1IZbvstyYakihzlUqx0MyEkOIjqJI926XeYGDt3iBhW2m69
4fCdGN0wwZCFuyIhxeDu0TpFiE429kMfkkxz7kJkkoFk/QwHkM+czK1gYPnNcJFW
DBAE3kAZG01Ww5pIlWQLpSIqsrXdopJp80tEXHE4wfLjFYD1hBqqdSW9jbt9nePl
zBxAPuTb8llbRGHzCEVgrEtHPE/7FCbUbDhaiDr5ZLEVEVDwJMqbi/bMOtDljaGR
wptMpSemeyRujMUP/pnYo5EqvL4dYsKnB8LQPoykb+W96Vkz8i/c8ks3pbHUSNpi
ZxS98DstW+7swTd5efL+ebQ2vk73GgMeaHmZz+/YwOj1TpILpY3vuKyIMGT9/daq
0EudFRXhVIWXrFjutZojK93lNU73QzjPOM24PD4bY+Ev98SLaVSLf9U8hA5hJp3t
qse90qdFGz6E/iNDP6xAsoex+pUYpr64i1QUwMPjH72JINzqhIDO+2ub90+yx7Nl
O895M7MlG4qJwGUj3mMpN8Kx4Bcil9tbJU0/EK0vZH18KBkFS2VXJrcR+yJa+qng
3blCOI/lrclwvBJ/Qo9ZSOTgp/Gbtm0rUWduIaPhqfTM5gBDuTKBnww5NyegysBQ
9AWBe/8jbDzR0ZQmp8KHWdtq1UB7SgI42Uo4xpR5Y39d6nzNmCb8km5JZtpKb3y8
QaV0JFdP0F4zedic5i7G2caJSK0dbH9MunlS8trIQ42A9D07SBTWRTV7bT6WY01i
s21wCTTe2gz+0FP5QDjdOpQ0eYT/SxsiSBXzkaKADTZw1g2qwaIPPfOZgyWHycVv
xIjm3snA4dDcPtsrzgVKDD/JqzYRao21qZs9m68LoWcZ/YnjGnTF2tqdWFn/AcuA
uSQUwbpg/aur7Kz9wRLTMmodHv5SRiLo7bB2r4zkQMnKt+KfxU0QWgZ4VQvfPHI0
lGVFZ7Emg9E2PbKO6c4konZpa16b4oUZ8YDn9Ccz+LSw3vW4355DWDcI0zsuEOaI
KofNQRTkQrOwRSw8vurOL3dSsrdkf+pg2fYc2x86dUkkCxQRGXMBnbYWy8SxtSAl
HSt9T3ouRlH8qCfKKJcM1S5W5ThBY/gM0ccUAblmW9AjXh9xKEH6vBe4hUH7fbuc
nl+6y3K94otbiTPsTTKQeHL1V73zwWeyLvw6WjAscRKkN5K+uG/pBnnUjbaUG5WC
79ppcT6Z9XBWzmIGfVXu+OoUJl1VbubowXxGUiFMFiiq4D79DUp/9F7ZhhFshZMX
oBhqJlVx6x1IWz0z0EuS2h9zMaWGLLYHsJSen2MBP5dJjlCoWZbd8ItQV7wQssVQ
14fyKLSEoecwj45OWJ+o+ebeGOi3tKgLlb5PzAf8tDX5kq22Z0ftBAD8izp82LJG
upoIlgvSEiuwVStq/QeBclnaBLT3kmKxZtGtQFJWEztiBGUF1DPNOkl7S4k9enaw
9XIYKo7f4QNmife+YoQRRpsaGk/UkTJHElgslcJnjJ2KWekEOqDcht1DPtuDtLc7
TMp6vLIyCIqnNLbKthelv1scl6kC7dUujdbNIXVKoNuSQApbFNbHnJJeiBcM5IiT
Zo6KecHzZ++xZA0+PzkyH625C7UPE+aB/IPA8DDpkQie1uBNdGXCFRc69LAskJQY
bBFJLF6QB2ZGN44sEMbmzm1NA0DdZ3Hu7ckxnO7amtAuQhvrjdNLiXq3NpxIBYSU
i3H2KwzEKsYD0k5v18ZXfnJvPGYORhFJdlUb7TNTBqKcJ1QXXt/gnmQLtCnZ+QYk
otXf5wr9R8MlcwRMDEazfPjX0D4bEAJzC4LCd5Z84rMjt+RZpRJ11fVeCuNR9UDz
ukR1CExwwx2YRO/ekwV9FdEZ4zAp4Yxd2+6/61o/wkeVOOjHLOwjL0q2q4g18h6y
BNNExGZxFoyoLP/f4a5Tl/EF63fwT7NhYdvcziXwpR4+LZysqN5Q8rU+WHTXd3Vb
UmNZJERorUars4uUoT+mEyN5QhQISjqvfIkVHecTFTaiPctCK+1cdTcT2JQRndq7
CcGTKLbN4Ho5+ZOmuu2qAKtyzd2eBdBfoBLMUB3QBZQ/eVKc3RLCg2wtRAbS3JoH
Tl2usBkBJzQHZmG5jdDWJ/GjWzBcyRowyUN3juM4z3HapGzM4sM/oCG90ZqxeTVU
xZvFyxU0ImUZV/E5nrUBb0tGk6whjPTzQ33zSa/dAlkqLSiIXcFa/ySMcNYbI/eK
3ml4nRbGopYcK3AJFoBr9AeGV4m9+Ovz8fQ47LNQgAW2IIZHhAf3Fvttt0rX7JRc
wneBA+X7BD73osULPBXZEYIY7L/BH14TEgo7TMGyVdUsVzeFIWumErwPqdZS/4nu
m6kP5KzX3C6jb+HOy8tKtSpEv6rOrbAONtV9eaJqjaWvLPOoNPE/6KN17NTbmphC
9J341y7jsoTC0LkFKFvkyd3BXOgGVwiKNAnVq/GDInnuyulR5jwi4fPCGAyab/sL
uPIC2jsUdBJRULQ25P4FMT5YYcU7QvfiJ0HKp6dZFriAWLK+MLMSVj0TspwEXQy2
ZEVZF33JFVehlfmaWe3tj9c/24gDr2ImOl4LXynih2YiH5TC4GDE5qgwV8PCMKyA
2rhIVu1Dsp60HSAQDmQSXXxKzpsBjxoo4X3chFipjrki4yOtcdzvAFOGEIAN/Y5m
qIxmNfVlY+I2N3Jiv7oTEbGfjp2NCdMqHzg5kRLAwhq2Sgd6KIz4jjNLn+fVwSxi
Zi8NqiSt0/BuMDB2/SS8ygJV9P5hnjD4/N7n7apCK8YcLRx2hw05vB43B2C+OC6b
hp4iotVHzzycn4flWhDmrlgYeGT2DJZWaxOhYGoc0IPsYgALDhGkDKbOupmbQnyg
QMccspmqOA2F5NaJmJOZBlKNgA3oes4vNR/AXhnR1w84ZhDsE/agiqLsvcWiOLtj
BoW9WYpcDi+VESlsTRiWTUTmfwYg7fM0YQ69FNp05dzJUkdB5nImPRvNlyfhZ0G0
uIbZtBmZMyUpjOC30LtnJhQsrwj1FeKTlMsEDYkddvTm+MLx7u3nzgedc1jmE0el
1qTFbCy20RL1ecZ5U9P3am/OYstlfcfxb0HQ7A+W+eMwvC/kiGRCZQs/uPictm4o
AcDovtzSt3CmOcVmFEu/8S3VnXn2F8IhyL7I1riXFuqsn4Htu893yDnwyG1elGjc
tQV/kJqlFTHGCAeJcDFSpRXs9w8nWLTWRUBghsYjW1/yCerfOKs4ZxHZlEP6CrWh
2fj/iiMU8xZU3c2W1b99a3B0X2T/8tBRcL6UPI0ROK0wlGOBUHK1JxyWQ0yYy8/U
EcBHlAWIkexXMwjsN+nAKUBC0JTINHK5N3Sb6k9RZVWHoQBQQY5JSzVJcq7hrenO
jAZ7NRf7/0uBZe8hYBxICvD6TdqnzlsIkZ8CYwM37wJ4Fg3f0LSieJ2r0OFTE7aX
kVo302JwwXrLNwplTQn5Zs7NVdvoQzxcIFKcL9IbpPBqcki/ncXZ2d7OIs1sgcn/
IYbGJ8t0eAWcjKsMAi2Xi64SDpDBtrQ+i3mVUImg1JpPmRA9FAzdx8apUVzpiZI1
YPtCxNiTv6tCTppg8XlgWiJGlkAD7evf/pjbRD/wcOz8bbafYcpAjRLH0j29yNZG
8fOGIuOVB0mK1Uqh9/WetJIfSNr/7Y1qQBh0dh2cI+l0Qgcn3E8lbFnwN8rRGmZ5
ABaNcTUPr66Hkj85l+5YTR+GhwXjBitDs4SvQ68CDgW0Dir8cqFcoS/ElClSGtyv
cd4p5M+6bZZsdq8cmna5k8SHJlwEjfhNyuJ7Z4IScjSQwqqIZ1AC4o2wyiaiFbhG
nnurGZKn9ymM60EfKzs4qXr/KqqQcwLG+AeoFj/p1a+Qj1JgfRPqOxKXJQsSW0FN
JY7BjCli2qbbOlzBPAAFKvGhTfLF7E2BBStlUSD51CwOwacjtMi8mH0NFX3D+O2K
upzjMmIjzscKqwW5xmPSvfggTJ4gei2tISQMORfUHme698bRsZCwQIc7zEImA/da
9o7aFXojgkjtzqpV5t9Ig+d4/aUQbD1S6dgHNO7NyU4+rzFi2E5M7ybSRYWuHzt3
qdA3KLSy0SUu6Ls0FfWBM+SkPRWMDR3KkuIf4RZFBruCRUoQR+SVpDB5CCjSSKQ3
HyhJHF+wCfTQ3bUpciOOEu+eGcjF6eYGx8nvLHqEcGTfmQrOHGRw2Teckr9WceO4
PzLvX4yLPvNUKCTTy1UAy0dZPSv0eCHlh+g07Rj9PjlEvetQjj6P468HpGWKtY+R
MhGFX/Zaxo2uB20RaAGkxEiwG5d07uFbSO/rzimfs6r9yGA+DnbG3HQrGmGUS4WP
hPHo/vyI8/YwprC2DCgFjgTnGpRjSomqTtfEOqDedTohW2l8irTlpmgv4/isalPM
QC2JsNq3caun7SoQeJN7ywuDExT5zxJipphXylq1Sy4r4n+Hh6LyzxkUlycXMYyy
inAv7sHpuKbiuMusocx9fmEbYKnSQ2jF0VOoWClsvkDd86N9ULBEqqLJ67wcGu+p
HfjQP5lmf4mGbR2BvnNpwVAgepDD9yiFLEfbTEoUi82PdVcmLZTM8yYDwmOvxgN6
MYNa9DLZbVJQ5qfeyuE44aGKv66PoHYIwV1UbwChSY2DAFj2ojHc5TaQA358sLhU
Y8R23JWnd5QgH2BimYSv6fVSWar2hRHoxowZyXjOeKy7fWgqhcs/nF5AL+4hU6MO
piyWwPSXD2ljn63FcaUGdZywecZQWmXd25Ok0/sN3IjQifJ1vHLuGVWRHitJlv7e
psCawI7y+jnSC7fMirIce8unL1/J7Xc8jZymtInJKoSFVCqOT7Ch6pbbJQs2tF2J
dO6j7a1E9f+VihRr2DESY83vfeJC1MSNjy0stxK2x8pCqcE/uNIu1QIWHzGeR796
p43TuGchqTrRet2LGiTevNF1F7u92+BaT2zGzaMAQaArgNR9AgDeZBCMgmuz1eWz
EV/0eQP4euQnr0WmR/tpd78Blqaj51hm1Yp18bA6n95b4+aksCd0af9GWWpSXWJ7
5wZLvYWydkQuQxH+imD4snshu+yHLb07f9XJseJuoQpcT0qT1VsW/8MwCcJ5zZMF
hpZ8iZiAhUUxAq3B2S3dZoc9cuPRUcEov8Wy4crzVjWmublZPaUJF1TKM0MEbHZ+
uCfaAgOG8ObwdDofs9oVEekyggl7dxNyRjPX/oLAxxd105ZI4YnY9yT2CDIcQsAD
t4WJMGHXSkGCj9G8Ea84FZxXYV5c2fl1abucemzxaxUcu0xndI0mb6MUkJD0ltE2
KYYYsuE2tlCbSKCRPf+TPkK3mX7Mf8Jvokn7vZUwkq2E2ov3LB1NgLv5djNn49fD
zvPF+0AZTM2ePb5A3IhrMKaaSp5Nwg2mZQGGFmwApWh+S9us+oLodzWkm0QRuJBB
CVPqHdwJO5QqJqrG3ZNBhzlwZCzHY8RYZ6hvN91peKlyTC52G2J91383/WUIZMLp
CW05gAv0KAY74cSsMdto+tlt2Mz0rh0yU+EV8MmxmfRiGEkOHrdLBUQzLe4sawOa
vmYnWKfRnKQXCktGK+ZAyLd47+GoyEsc/lI4fvb6/SMZajqpXXOpra1KM3iQlD/I
KlJZMB7Q+PssYtmFXn9IUagkNbd6FhLpwVl01BEPdxR4wG+2q807pvBdRIy0O1GB
rZvZK0O8VSVMk7kGcGA77GJ6I2Fxqp2XqISwDHjUJfdJp8Q1BGb/8ZChgXjL/izF
YsYy21qFEEiW51345U/JZ0jP2YX54dtY49INjpv0d8VjSu73npuQ56ZrHIzaBwoR
AhRKF5CNKszcyFFPXjg5ho9vb8mYBG8SemkPH5CNMeIh8ZvEyuctckSSPGVYmgF1
q5ViTnj4hK3KDc0TUpaupbPxKkp1+13QjNLiAQqpXBpjIoQy9FGSFNisUnRnnB7O
JX21JIYn8CZ997TyUBJiz4tn7b+8pp9zrJDAkGFv5qII5PIdw4T+0dIZKRBKinoS
0h9g2U6R753Q38td2cNyIbRJR8yWZnKzA1ZhzXSp8/N2ekFr6EH2HrFAO9A5hRUO
aAyskn579kEgBxL+e69wMye0WozUoOm/G3hXHsOq5dbfp2UGsLThtD08xZTFcS5c
P2abLOQT640l+Sqm47PxJI1fqkPokuLKsGwBZRSpS3akwEf33vqX/mgRsioz1doA
VOJ4cyBn2i8oJEqxIcEVEuH2VCekVlHwmKXir1wz1w7VrMJYv5+KpBRxUn9nHutp
POjS/aKXwFQJuGLLJL6Oz+10oHl5xgIQr0WtUz1mrefVdfflgJN7mbTOQX0v0jHQ
cJU5M4GmaJYIkGG7lvlMvw+c03qNnpHm5SNjwhlZaF+VLzAQiZlruYAbmLnEYhKU
MsT6EQZFoTIsgKUhEWS9EFZJQBSzni/xBZFYTn5V50Wfw8iDvcFJcwOUbTGo5Ni4
z/lAzo7ZnfW6Ib14vbrA1FdOE/4bUS6BqXqbv33O+XG4ZDPBv6z7+ggWSA4mp3dt
dbCQacTfwFTmKCm6Ex4BPX5gXVFdCn6WmrC1SPvVS6e4xzS4aPi7JqmAFe1tNF8/
grRiJFCaYZHwPdnZK04+/VdeQO2J9oXakDBDzXW5VK3mGl+++kJ9Nc9IXFuxbEUb
ORAEG9zu7FoPWF1OUqMh2q2aL9P0WsB1q/YgNhJJWbos4a9aLDOUHyNNP0YIlMuW
Cjkzsa0/GuYmG4v3+1osjyqkFNVxbpZWwv3WFiXn8oFWVM6KITas2Mw390Pps7pG
FKBnPrKinPctk6u6EK5OqEt3Zb29LOWW2GEDS0fo44UHJs7Z1g2/KoMCJteHgBSW
+p6y6uV8muDpQg84ITnElz4HKuvUgBihOnCnb5M9pAv9siKdAJ4N7wQQk5XRqWZl
xzCh88m5f8i0WT6Rtu/4eGZOd311lHekrnl37+ib5yhpH9QZa8PORuNDch4VArH3
5LL7VdbVlLTILwCJXAzoLSHnvK1JomaMh5FjpkJiU4Zt3VVcWL8kyTuhit4x+5PS
C6lQDn+DOk7RuWOYv2Q/dIi1FuVQShF7W5xonUlDNjWCo0R4PUGBLPwRnTEctR+V
rnsGnNNTwl7V07XtU6gWGrX9eWLcAn6oKw9vodZ3awXitF2uvbSqeq2i68CtS9Gb
1TKmpjsjtVnX1TT7He3dNV/H98aGmCRP/YyRnAiOZEvGRH1dd8eAeJpJsyfMxtBD
uTeBEP4IANjgCrl7mgQkmWCh03n+/TTpxFo286WoqfVi8P1PSmNx9MR45060VS89
66RA8DWCxnEfs2BhGRPhcpXJNe5GVpF2h52PzTUQXb0R+GbrQc9ZPVXqQUowm4JO
Mel1EO/qtpOWcYc8XJKOAs4XM9FZX1nHr1vkDGNN8TB92mjIVO+aklIl8wH0mP4m
mEogz41LY6A0OVkxzZpmvSKEOhQLeSMp2wlz7UBiLJzLCjdOSl3XqtHdE4WsL0KX
y1mBd+jCwo4FMIeJH7VYKU5twIrtPd6U4IYZht1l6+c8hBBYgHAkeBf8+G9n+dN8
VmXr+fe9eo7ia3ce+33cSh3Xl+WJW5ZcjPJumjBOsSwtAx/c+UIgnbLFLCTvjP5r
I+Baof7EB1XMta9DU7I1HvHmAGu3pyuU+85V5VId62EPaapXEVAW4X3Cu3JA4H4j
MlEdwYtw2MgElVo5O2coiSY4BXLANSyKp3BofCtpodPGSwaKWRZPIZ1aJWsxrC/m
hNKZQfYffv2sAxs0ai4odJ0MzmMPhPHFaCc07kgD3/SfcmqiqWmYHNBEtNOBbj93
udB6dm82kauDbZLMrXR+pouCRhtl+Urea+tHgTZ3Xm1Ar5GZAT89DbTkv/xCxlq3
8+tRk3Izyq4O3IxI3lQ0R8SwP90bMnL9amMge6gHU6IXiZ+oKQFxALh241cGD8k+
a5NqHJ02LYjS5bORwYXh+sIRBJ1uJYPQv3Y0S6gVURRzFBesqLrwUkv9Pjy4SDLi
ZhQ4WcdqzjYXGA1zmiK6ApoMnTON+m0LwolUuwDs+ppm4m1mY5WiceZW2HzWvr3y
cUQEL/tbWnDFBSGCvUl4FlU0PT3lzneUN34gBlCmKr6q2U/Gsxn1s3zxHE5d7i0Q
bGJbtx1aTzAP7j+UX3E4In2fPOvrk60dE+oG/CVKNRYybX07AmiBKoIEIRfWkAnJ
WJKVmfR3nRzzEV/hdF3Dzs7j4kfEdGOMKexUBSSu767XrXnAZgo/aNmuhjLlyCjI
T+GEjERcM5laIUtuCv9kykms6WikhcTg/1tjFoFoX+8G2zj16TNZ82kmkU5qg3Es
LedxfxrJc6vZbjh1A72IagcxAR4tOeTWo2mazx6baKf919fqtd3OqauVwSehaGgS
MFdrqbb3z3DNJR2pMYZCPKy6XrAqaPB33V1LRa9QQGDQOAQUPrnEc8p6wAp4E+MM
SadPGjLAGqvGqcbYAi/nK8cnGDWlyOEaoHVUToyJVbCg91HUbzcGFXPlmj/wKvGY
qPk+psZLa2s+ys092F1ja/UP2Y2RE6qdnK+ak9HXa54OFmzkPCLBVrq1XWDgH+dk
ELaBLnycHaO13UxRdkAa79v96Cp1g8z37nO+2KWbkwNBwU9fd8aTQZl+QV5zsn/p
ioB/FfX97X1V9AtZ4jNjT2cqCKIFvRHQ6ceuETP/Tjt0M5eq6yZhjgBZy98kXBOE
0AiGcSVfHh2OnKfsI3Tch8Si62I+uN+1wAtFArAQ0f/dXC3C9q9QQ0lXUzbDpCwF
4NqeXORJFWvnfvBUyyqGFx1y/bDWcfu3E2KdpoO185kWrnKlsFWe85iPkDumfREV
1s2QlDF/k2s/La7iY/wnk4mpLxdMrIhqcE+kayi8OUb5QUzXkgLXue4bvcjxYOxr
PK2re20/ebdExPXm+B/AqBjeYzaNhc1nWa49Y0nTCBUVaY7Dqkab63zqDA0bjvPH
wf3igBJIakqSemS1B9zjby5OK9FbU/HPvS5bGFovvasza77HytRURWxZj/WPlh1E
gWac555oRuD3zduhLfs1uFN9NgC+m5BVOdjsrcWeIsbCUDDPCgy301PKXOGYmHoI
5yGws8cTfiW4G1DPmgaZDmaNe29W28IxGHvuw43vkTDDbH7l8OL1iLJbJL2suYpH
8bsIVg3IArY4VE2xN+vkfSRLt2n8PAq6ZHin5exAq5I5Faml6Q9T9m553uh+FEat
K3+OJNi1pDDTw4LqojOJMcLjZS/zlT1I15jNDt66JTFugCRhIhznNf1BDSxeqy3p
FjGzLJ+3fJySEIOZHleslAiIFPC0caDP4pgzj+sAk4XbtJWN7zncDuA2IjmPYvar
2boes32BeXw9+B0SyZ2BA7ukqs8iapBieADRCok1Fg4YuJw5UWGPVJCz0d0kZweb
cGMa0XyVxzo58pBqEkTMGj4vgBC2dOTBead7qc4zmACQw/YnKeQlCQwdtfMi4Iyh
blm4EoUWY0LmwsKsgbqRemAqE7BcBbejp0cH/jQSIRVHrJvD2xCpN8m9MB88UuLH
kzSk8FNW9gKeEK8qctn0DGNt99ENSUBl6qCm/mlmSqMsjIc+dAQtBC3vOH9DP670
6DAchCbcdyAUOYu84pnLvHeXaZTUO7Oo44aJ0x2I3600LDAd5KCFFybKwNyMNGmB
vNvwqSv+NXhPQCahYceckoQNU20b3bDSY2nU5RcS1Cy0BDXpoZLroAf4JlhEANTi
RGBCtCJpueBNo49HsejtlSlrUOv3mmKptdkurcjEZTUaWyZh4PHZkVyMzI/BgKfH
8cbNQf6EhDIHCGKA5aVOpxKrMw2+D6DC5xQw4vJ0T5xh/twwVe1Z2NmULYPP5+Ll
niFfpUmwXEye6NAiNQ+HigasKhwwRuFG2/FQPEFN8t5S8aAlGI0ebS/NDhDaBA9m
2s4LTBwPv0EFthE7TAMyVMlkxkypatnrCtJp/i2dyAkn0KUKkNOTl0jNpgJOBaYo
T8EI9csZy4PnGucUTnlsFIG9eCLn5A1tuG1WfkZt2BJv9AOhc32sS46pBZA9R+0A
YYO8mW2ELLhdWHiqMnF3NxVVemOwuo0hInpyK8e8nfnjYwxf/qzGWNfnoFgrTAKF
15WrlSPmnSwC0D/bTMLcifQinfxFhZyBUj534oGMvWGX1BYV+s3KR2jhwj2edPhk
+7PegDZ8WA4FrgUISS2Ai68vGKHH93KRrh9nJt2uJ6XQnVq36E5RgjUfCZGkYzLt
UMxhAKNUj895/CSItQW3BFQ6s4VeGarB7pnghqwWhDuO3kaAp4A8pBLM84JwoERH
ywfC9xLTnbYsNBZqPaYte7pNjnoGwhJyOxzwnccJ7uAhGaGCilU9vcNz9a6Uy3Oi
sjnt0uchFevb9SwMnazLFyq0UU8wNsRrp5L3bxsRYkkx1BHKFtMawc/dnFlTM5FS
XFj807bVuQR5QSOG70taeS6RIxP9Zt4E0O5mU44+jAlA9SDBap+o+wh5jEqxPeBD
DDm+0SpwOaIB1vY3eBpX1ZLI5a+8aNVXKCgs4UHymDw4OkpeOZkW287KyA7thOYn
wAXNisLcindnNUb0XPtlO2rUjYnMXwK67oqgMhu8340h2OaymlNEOBMa41OXISOe
cGviGLE7fqwhkFIoVpnf4btmSpI/fgPfcOUdxXPwEeZotzfbnBBNIFCo2krpCic0
fyyREbEPTLQhFbMpftW1mhlezS9xhfZEYpFKhcfra5CQvlp8/nyPrXzjrD5KfTOz
0mtIJ28pzqLzRY1wlKRdbYWr3rEecrABNwG820u91j2CFVTe+hZaI13sK5NGjXf5
PXWW8uDAN1KFYi6SzLLV1e8O5jVHSyBi2welJrU2MI+9g71D9g6zjfJR25ew8dUJ
AF2jOC1kpSgS6k3m/PoxGV4OtxyPVYFga+nNXd3hxQDJ5gni+EtmEC/Z86n35yzW
IE6474RdnU7PjUzL6kFmxTkpHqR213SedU5PiVJgQS7W0bq/+n/S8a/tR1UVCpgr
uXUZ6wq0CcICErxRNVFbDqBBSBF3WhADFzbmZhGFBN3tMGwBX8hZi3MEXPlPSidE
b1EfJYe3aRoXvEYZM4GQ3xFqWGAbK2mzPBxqxfhBmRlkM5zoe0a5XVf4x+dwUcUM
9hmNHxvrRUPq/IO2SV3UnvCvRAlcpEQp/G/UsIXQTJxUBiCey+7506z4UEJb4CzB
UyTb/UPxhawUw+c0nrUI2A6IJm0FEGJbuk/V8jCC8RLdpBTYHdGasakgcOohyT34
OgQGgtXxNOosu5Y8U9Z83H1JEvV9Ql3izHxgVFst7T0d/jAufFKvKRNbTQ8Jtcfe
UdUcRxx3piai8E4iUCUmFNo6LRhPf5pvm6U4Z1Oia9W8lylDUBeASWsZu05OQxL/
kbRbzq2TrrUfV+2dkrT/t/q0f+JVftvCRNUqHTKMtdH4a3duXqyjq/umNK0SAgYU
10x+y2fYpNIT7XJv7Vr4MwR6wZu8P92eGMUEwpCYmodkhdKksLUOV2dpymWm0YVG
pbyD7g52IxQ3rScJUvKXC/lR9HYhhrt6VVvd3D6K4/nPvlWTEbWhje9KZNmWQIr3
+Ce1wJNp2DiomZXqVwtylNxupQNzDkTmqgxZADl2It6K9u57+KjSmj5mhv5U1G+F
1QR9F+yhhCL4eGO4gRFD1v9RIp7EBC+y/AjWYIQbgnELOc62BP35OqKWxH57vAGk
eBGIPWF4NooePihFe02EfxM/GZ3rBlmOCabS7Y9BHgGmkXrZZSs2Zx5BN7vbvUdy
JvQR9hvAT0sAzcemp4ABqHNScOxx8iPCZ+F53wdLp6Mks9DoqhmSG7ki1AjyzoXp
NLlNasbFHDiWUG1O7sXY5meL8tG2iYnR4x3NsHvJ1j45G2C7P4L0TAbbHoWV8GB8
HoK2SMQoGUgwk6VuBaPQ6SNfbYGL2UvIZmXkc0w+4uqyhEgOfVIC06q6RQtGyz+E
89VOcCH4jkidApCHMGqOzsGx/GQK2D29x+/MEPp/LNb2HkzWicy2peJZXA7Gs/Tv
j8bfcy9jImzzwZHdP+bEpG1sQz8DwQX30x0iT+omcrm8TiF2KRupX+RlzMcJ+Vum
4yQM3wBENKkAJkH2EbOpQBIi8Pw7rb3fFMEcfoXFOBLgciyaSNag+AtGX2kdkFUl
cU3y+UoqlR6ZUx2w+NmVHrbs1xiNjF505TCg0ZcAwazp9uxyXHASQM8Qd9Nmm2fq
5u87NJ46YFkGtSDhuPtPnFlOciUQCbj6Ssbd7RZ31rLoTh6EPqlg5926B+BpHNZv
+uXLlOMq1XiMAloYwz2lWPbV49CGl2529KoCwUwJgP8hrhBGlbJ9hnfd5kdLEIPV
ZnhfFdDq70E/PCX4N7uBqbEZu1+S1cdora3wliHCgZbVdh+lleLX8qoJ2uRWY/El
Gs8Lwqv/3UKJpN4uUEaKGNjoLmX4IYAjtiAY0juWPhkoueStqkOnwh6t5jbAINGX
gfuuOZvWYeKMw2dU7QZlHPWrAMPVHO0ipdW+62ckPdGeofKWiEmYgVC9dKvJk2fj
emVAq/B3Bg7NsdgwdJssXjrbgiogBtz23VPeHHaCWuOVW4WoxZtH5CcOlCekxIof
JC4epnX5srMHMHP3r3vM3HLffYc/40RT0HRmk8WOwi7bozNYGCof316+FNgteoXZ
/Ng83bwu8XL8mCjoebkdnmbJqkahwZb+Mg942V0Bi0d6YdpwfTclYoNxuujHGz4U
QP7nUqU3+zStCmX9ziINoLfMn5MUWTDuLneN8Zm6388fKFD499/9flQCJGJCfKW0
ixd69Q6mUkSBmBOrBL+FkJi7UNKhRo4S+lxVLAT2bqIjXz4+78zNlspfLbAzEbQQ
hTQf9gvoXZ1NnHag9NO4wK3ev7roxQYQBCTDSxTEjPdmaFFGDcFTEQx/JLzh61yc
61FHN9yoxlcSQShWZreQJm4Qi8WhroW1Gs3YP8HWY3CvFsw7wcMDqS3YIKoNXy/R
CIXWZPbxP8iSd4J3gCrQH/vrj/hLVqcxoQMfb8cwn7RmZqGzZvaSyiZ8n6aePKdv
iKl7RpstWKNi1BwO0HokopXRJPAqHouAAkyShTn0y30gsMXmWcPOrajCLGU+TzLU
x4ln19F7dYj7/Ip9yEoJ3Nad5NxZ3hW+4yH0RT9Yj1a/rK01khhVIoyoPmSw9KVW
//p9ywrGko7R1gRo5CLe4c9N0zgoSCX7kSF7O5syMW4CIanjueBbwz3sVCUU6mNf
3JXcYvQ06c5J1yCPyqGlUHmEeYXq4INoxIt2mPNI3Mp0VICvjCNKd5ETg9jXHzoz
I35dT/hWiDDeUds8CzjKELPoAUnyGk3wj+Tr0mYPQdpOicrBtmvbESnE/Anm0EQN
xRhyuMj5ATor85KZlkcNYpGH7ISVv7SntGrQo9QToXSpx/AwDwE8gmCFmvpoI5tx
u2cTc/IsSJTKv5P9mn0/4gW8b30x4sHauTSLQVgCe56FIL2nxxG4Pz+s0kSLDsqs
r26e5KU1uK2QWdOmiA+HVLtjir4r2+ldOtlnsd98l9HUbVv539OR7Xln1A6Gm2hs
qN+8pzOSOmNkoyAUeedWD8EoJiKV2YllsvXCYa6dm05SWOtk9eoxF5zBNzs2W0jm
qTRjoiKxZcoDBdX2KmOU1M+x84MkEk9S25pSxZX+YuvPUcAfEvkkFD91jfZ9lhas
9BFUna+uaEIvCt7BN7cZGfVKAjFg27vIKm1jaLmuqcNbpgSFmtWW5EtMDCTlW9rK
q9USe4QQZTYpkmJv8Kbbe/L43kem57WzHo97Rd0xQlv/YQKa1SirD3qaPXZuwhA7
P1kcMUqj8E8uj/W6Z2X8wsk0H6v6nwwwgTDWSaLnOSt6XQ7AZMGmsCejnepkupEk
6oPthybfRZHkJqo6Y1vWIqcZ7Wyq3UKI5p0kom1jfUckrs0zq82dmtu/MqzvqyJC
zxpoX7Y2I4Gbr+ykV8hpgP6OmkZKAw+suz+y4/lSVdsFdUp4v011kCoPVyi0Ey82
e7M5OMdJJhOWiXKxH4kTeyN5RiqWOiZgx9VJsfIRrQ1elEfwC+i3GIMqFuH7f/Ik
tfFnq/JNWVsVfsS9F1Wyk6XNhO5WcwbldcPgPYYVC1u1uFbm7kfRN7daDib9BgH7
Arjr9LdPfNCVZxvB8hYeo64S6Si5QwqsneOrqWUwsjihzaUN14Fg3qiBygavV84A
8igLzZ9/aaL7B+/LehNpO9xfWoECu4csgqLwheiAHaUw+emBtsJbh9APTIYumRKD
/aiQ2m9gtaFybqw2aK9C6E4iXhkCZlA02RClhwwRO0fC4SR/qkW7rXyDfc3t7jZc
s3ZDNttD+CaWtDY4sgTRHE0HGNnDqMcyKT2RJ7WiDeUQ9p+X5idfZC130SGpWE3q
TOa4+hRsBWrkCqWWGR7DvNv8Qc52RaHIYGoTatf9ZL9t1qx/WGdDAHrGneiE/dhB
NZG4WNrjblR8ZiASjVJPtEJ53M1FZrju4DM/bjeMbcg583DXQQ6UtazNCSugI9aw
C3bUpxiyqhIaKb+p/2E1nZUBW+8glXbNt4542yAPxdQjciW0iImyS5pFRHIFP7CB
M0eCyoefnCtEMWGh9069ZRiaQnzsaPoyhc4ZZ9cNQqQxf+JavYZLQDJ5v7n0sItZ
HqCuldp+fG3iEHVOjsAHQK4oZWzsK30Ylg4asWFyL/Jml58q1pt0IVXHDhWMVxuZ
NO3dw0qY08OnpgwBxXNS2aKvzzC5AFgCfnVpnT4uqP9mgzMvFlQHREtO15LraAW7
eIQOwKqRKTyJ0ZpGZg5fqMeR1W38rKvr6ocTCYEnbCOVByq21MaBgn3uV1WGGa6y
vt/1atjEbBLKEto6e+mO39lg7J3QqAKc1ZCRXAJfvllBzcYmDjLoLjhtDQZXYZY0
GVONSqtSNUsZjD03zvjipC5zfvIUl5uPo4zeMedWKBi7pYauTWv+pLRAcfYLL21q
+oJxEMY9lykBlNLKqhG6by8knTfeaYFqaYzSHXkY/t0p8lyztTN6famMVcvdPtUv
L7tyDvSrNJLUInm1TDwzykikHSFWj40F+fe6Q2R0nMJ5GYw6DRUclT9TPpjbfFLy
HJcjeCMbLwZHGFSS8odDW7QPhFssxQXvs3qXmBnzEMtWWOm7GtMD5Q+DVcFc5MsA
uWM9Yo+z8ds17Wc+wzzzWKn9KaV0NWVbX70cg5ixFk6Iw3HbX3eqe5b7d1ajCcwe
bWQx74kJVdM7sQVi/BRWiqqyMy7H1TWLO/oNe6N/fwR7XSuMuiXSitQ4OiFzvk7k
7dc+migaXIO3an+vwZ8u9MkjpAxIp328dXfuTet5x6bN5GgvfiKqLh9Eadd/+L1T
L6LDgQphTYaknsL1Wawh1bpEL2QIngsWB1Z+HYG92GC8Jxv51CfcvhZ9wKPR41dR
h3jyth8xPy8b2vcSoPKup6q3VknCbsU1pCLm9rmiETEWufBnU6zQIxkWC3jRDzkw
6DmMICSn0xN3OLiQ1AuS53RT1rIb9QQJLYkqOVhHH+CxCSVWWylJHsCMz6ymYs7m
O9PJzoN5kqgqWZgC9Q4e44IVB0+dmWhgEl41SKbB9aw9jSul0UqIyzdKVHBi9o6L
5kWC2G9EAUKFkmxKp/vWD9edL+EqcydxX0dQN8iEyiqWNKLHVtK8Ri1/58pvoBMK
XzM9oHgBcPX3hFpGVIeUl+wjIAZK1FiE0KIvEkk2EHV7Jyy4Pyd83BE13KtSwuiI
t7RJ2X4cV4ns514Iz/szSTXHgfsb6X1NNdJNCkZrE0AVrXlUkg2vWB5CcmFMylO/
bdZHIv91K4AU4GIoKo2Hcm6GOhuDq02a4LIl4gYXVA2pqoi16AMy/lkVVHmO/vR2
oyzqH91LDdjBBQyW7f6+a8JSvrGPD2vyhDmOrXu/7QQDqE/tU11bdTwP5nHZ9P+Y
55ZekejdEoXOx0kDeWQm2pwczi13aOkqZ10E2WZdNbXOZK0Buc9voLSIMGRnRE4A
IqEfgmdPCW33fyrl/LthQQluMXT/GsrZBEZRsXIlIrIL/8avT3QWpJeNUWV6hFxO
TKBFTCxYiWNIywOlb3OxA0Zsk0B2FM4syRz6XEqW63ktL5f1Vz72vmJHsgLaeVlv
8B3ruSBpGaewcB4evRphSovTBeOFDwZ7sJcMnyHK3ADX7jSKXLHFvRIZK6r5a0SQ
vpYsS5rz0YmP9hE5LI8yJPekUTS1N4a/e7LvDyAIHe9k4Qo/MstTqFO+cQubCG81
DH1ltGYnp8yJAlYrJote4h9i1tHLKQxcchEMKw9frucNRVFZKSW8XbPkYkH5d94e
stnup9bAdzmRrt0bfa9KTY35b2QA67DgHSH2qutDVOQQ5eT58nwwS6P0KsRVRbbo
t+BVRd/c1E3L3qtdwR1XwlgfOaUw0+37lJwM2GJZWmVw5x4yIqzd516DkBYQN3Yn
4824732Y9xqRMrW8RInRW9tR2bOoLqrT+jhysEM9jt40jca37oi5Q+FSgxUEpSsP
E0s0RfDYSYSNd6CbnrY1Tut8s4ONr2zYSJJdmi0izEWsnyHteAWVgUaaw7EtauiA
uwybC+3SPcGKsBVhJ4ar5/0WPjlKCPLDo2U+BSbnHNIXn+r4vzpVbni8jItb5EWc
GL8xSg1kaXOWA6phAfCd7LxLfsKpBcNZY1brPHw+2c0tkGKBsWChFH8Lu0dUeg7o
5aHjZyfpLlbhamwRZoMdgOIN5Z0wM5etQaTBk1FYblgfVMUA/FuZta9k0nL9oxuS
B9sDHtJbqbuY1jqH4M2zujfqLnEKFDKpJqP6CiySI+RLwF7fL8eVxGkodySCHNk6
uL1Y7HoarROBOKRoE5ShN0txWH3AuVIFQX2iHpTibWji/XokE+KNktmx+1UmvDhi
V9sQBQQsD4252N4JMJ+1NFbnW6XxohDmqa04mHmrELPjwlp+PFEJvWL8Y+T6A0Ii
mbtiMA2lhf/ZIdhH4k1CFFqK/prO0YUeCSAJCwzya6dB5wyjlEWsrIbntwgTA5RZ
aSsIzh6E1oKwz47P4Cjh13kgq9NW0n4tHdl2vayvnbD5I6sCld1HBqD05QKr3BAx
RJ95tb194dkFVeFAOi43INsFAEVBbdNyDIc29cfvNYbuZ0MACugFxUEkQAoo60rq
G9y3vaJhS2Im7FICpqk4bL7nwaGxyCdjj4ppbNORK1kVlYBPgR931JHroDg06E1T
pMi7SOYmM20q1PVrNRHe3gAWOEK7v3BM7SM35S7ciVXZU5EbIR1tEzIn8arAeUj6
eXrEyVyMWu2pXKZlh46zFMr3AZZH/jrb3ztucONSM7LlAaZZ/aKpOyFiuu8HQIl7
38rjHcf+F9CNHA4cUmPMUK+eleiQqymQtqoZdGWwismzRvNqUmCH+IDE84MJYPSC
Cf8Xot0xGa2gX1dkJ8r6ImZHXbP4YD3AOkf9HdivVgkwlXuFUTzoYUFkywkG66H+
EW3fTEjkE9cEW2YrCfHSNnZmyLo0eaoYPR9At7qfi0L6fgCJeWYpN8XIlXxsNoJ9
KkgPFgbCmBraoRnnKnUuwjjTb2I2wHQHLM4UHF4T/OqrM+jPl0tMbWqzvUIobsdb
0nPQfAz4/bT0a4JJwTSZoku1MjFeqe6tp/QGVOmDD3wH8jSyJIfkAFMNjEvQmRsQ
/YEXVh8+8jdpAvdDl/I0DEA4rtGmo4xv5PUe2c4njxZ96MB1LFavL/277jxiYclU
rAKgdC0u4Kb0QiN8TVfgRHCJdzHJ+JTQMMUM0z/4zGSKXJl2dO1KxHDY0zwRvRwW
JmOpDKnWErAaP1IQ/MwVJHrKbcu0rqJOg73SjFcEcXi8J4c5SDVs6jqwW/83sMb6
CPliv6zGgsf1dVke16dcWV8Q+s6V1wNLExOrhFgmTcRm64LQOoXpgeAYRBjty+EJ
r8yosHNDC3W/cukVIUnGkXhx3NUJpvYjoAmpYObMyR70yOqX6Qvg6O9DsO2iOm1A
ph0cb2hOrKsAbB2L0eHdO9rehX8c9s2SX44mdhVi64NwxSSblMv4i2B7j8OydYBX
Akizq2G+x59a2TOVp3G+qwYrO+T1n8PRJI1ANlwDKWM5iQSXPZmjyiDsqTFpAF+Y
qpoczV6oFQfgZ2C6ZDiAGk8aC/OcyPkgAsUPeqRZQrX4gKajQQWNdXsuvFCv7eb4
OEAHLwWRu06uDO6QAy78pO2NhSWZOCSMOcnzsffk0ewtx4P3bItDHzcRVa92z3+k
FrmJhycxhTjQ9awevxjFk7EfYTRvUd/YEZtJK2uDHo2UVLomMMpY9Z6hX+jKXspq
EJ+as95LdGwHMwfJNTrLpO5+eDq6vUgIniJXLG10U4Qv9m533c/6KtmlK577AAMM
QmnFJfEgEzOSyY1yru1rCTOnxfYzQvUxH2A8m4sgkJZngeeqwUSWAzT8JBKuR9hb
QOlv+z7x3cqrWigeImgTlfW/CaLej0Jw9/P5AL2FvKWuHj4kxHuxxLTulg0z7FtA
jh/8Ec0CRCvz4/MlrEbe+6Hy1UGXZNQnQI/PN8L9763rGKW336+kzdqY8cE+tAb0
fsYzTYEK2dukqFzz3nrfDiDgb8f2VWaDF1Zk9VOXDt2NOe1V75pGIpZ0zJan89Mt
z7EfoiGJKgd8MvaDIBdDDvf6XATcEQyYtEXjbc082yn22vhh+gVC7s4iYNUV9aXA
JCAPXNA4HhHeu4Dsoy2mEXIn/ly0Zy3/jWpW33ZcIJ4xqiQt9PNzadju5KyF5j11
+c+UC9Nm0VZV7Zb9mJYMcjZs/Eg0llJ4pdtw31Glh1VWpXZ7ji5n0nKHOqDD5Tq1
btZC4/x/ubzgKKMSWOb4uTbcDVHyfnSlOV83xZiIJ7RNnyFWFBFaFtiqmav/YPe/
HJZStftl9znisrj4rVjsc0li19kat6agoTlFX3NpWdH4B/SEsnKXv9C7SLjziUol
clD02d+JvnfGVdokGwxUZE0t5qwFo0+M/msnBKqhU77ga/+clkxhyk0dD96ME5K9
WzGnHBrfFVdvP8J+2KdfbzGeCSRI5kfHcbIc+PlIwy7EoTEm7PP0nD9tDA+MQkEk
uGkL0o1ZDvRXymInf5l/UYuhE6mZYT74xHD2k/mjkRXXC7huDQesUXJEMNrkyZcd
wBjpHhMud996J9zcP3lQuKguPAHWFAXDH2zJZElcu23QipVFlj/21eGbs/mijM57
yPpGf4U/TGS4sxwjXtifreutOb56AMB8SBo1lBCDh6lltfiT7/PVh7M6ju2PLyj4
x0n1twWTKmBHx00WrsQD4Sx/ONkuIYeZq1ssKDm4zTKwWH9JKxojUsexFYX4oiWk
eGIYKWbNSkyow0Lt3nbmI0h+Dh3Hf5/YtcdYROzfl1ZY71Z2rjoeV/kn+xmery4a
fG7NFs8JWc4u99GzKkldhi/QxP4nBLJ2nWQIIPUcLoBowWaU1dCNZeFfIKCHEAKj
1SX0fK2scQl8n7eOwTKZuYLFm85es85rv6Mv1uVgCC+U9G0fCjXA2Qi2vwbKQD/z
WyjI9eNG/jfs1dKRMjLXdop1ChIfFwAaC2jFZrV5V+pJewuzM2v/VdTpE+cER37Y
6df5YT8d7nLhRxhg5PiWnbg/ZAHQaWp6TMEaldq9wSg3Lq3CWcIQ5jRkFWcjKShv
FSq13MP30B77Hvm+jR9Sdq4MKAheB52EOm7fp9dYjU0F2W0t1pfzj6NQKU7nVF7P
C9+wrTlTdCOFRsfXnaMciJFL3gAWtvQj2rqr4VANV98LyITHW3xXgy2ZTzlJbq6n
rvbTZc0Gawx7bZkcXWY3mvIZinK6nY7xj98en3W8g3lpsF9YmgoAbNRhSCvImhQ5
mxfoYBhzGcffS01oNZagIXiu1Z4IJ5BV0b5qonXK5TZP0tAPws5DB19eF19hrWej
du1pXVQggIrp2QQjTHfRGjPv37s6r5cupJ6Cy/e3UF2DDQTq9X4Ai9NgnmMV1JEL
tb6ilq3sCYzDwoMEnV35jjBJwEMAoBiQyUBJuKA01IVTeYsWaD9SEcP3u81gfwf6
i15kA+p3kWji+6KgAhPGeNf7eTilCqhHkNYQPqHEaR2ThzO+nhWm3qBKtee5gLPO
5De+Y/dyV5jAhMfweuGXlYBFJMZ3voPzG0tPsaVrtcs1iYBHAUHsvz1CwYZPqtDF
64kWTyZ0fna9bX4UyMVPqjXeUjBhmjd2zRph5YsMfKJ1/qj7jJqneq4LgwRjkIV5
JAAknBUC/+rZh6WpGhyU5gTMzf/58ulLt+nuvxpQrUjBWB6w+5WEF6azmgO+J6Pt
xj1ZPWP9HqiH55n1uR70YYawN3LLfTqkDOkWZBhm3nTahQfMlIS2ffzoNblK4e/m
MxWy48kxBCdnOFtQ0UC0McipLbuxqzFAap6VpFa+VQzGKhGzwHUL8/jpEKABEZlf
A5bPtcPEScDC5b+ysKvklt2Ouhl+St771PMTWpAJb4X7X93oLUJnrJIXZNiOSxkP
xWvzid4ptMomBVxOSp2F0+2iwYQ8R8hskHBCbYkSu4v0zRX/gBG7fqxvqFxlYWLz
C0yq7h9JGNE6qYQVSyP9s6/yOU/pFtt6wXchEAUZ+0X+8cqFEE1yMAfWIS8XeSMH
SBQt2Z20YXWwO4sXJTN4FiINM9N+JlKctEdyOYQz5ym4xkazjKhh1SvlrvQG1GZh
CcNH1mV+7eBtamhGMXbYX9j7IWWlmc7KUJELGcPvkXTefZYDQViTAVq+3wCIvZSY
TP3UbH5S/W+aP1UgVLYvBd87EvIvUhq748ep9NlPhHAMNZw0umlJsBZBuP3A6c40
khK4yiXC6FT+VyG70x4R3nvfr+ntjdKyw07Lydu77OhWvoQaWApjs748cwS0czqs
+qp5INbRrkN20k26QQSdDscWL7VlDMcFHPIGXWy1G7IvmykxrPtTtcICkVav6UxB
dmuhWbZfZ3O+EFhZYjeZVFxOa81PfzM2VLY+FHez4wHrvwSLY1OiGlVG1WXy+Jff
k20PuhFB+9SN89/kF7APrXjx1F77kXi2SaM9FGgYOxDDD5+p26XU1a7RJbclDgWS
Ymn3dCHNpW/0hekmD4h7kSvGsdMyCbao2wFeDA7ECRQkYDooWwWbEZP3wRrsVYuz
IE6PIttOU19MslqznmcgP9JujEqvMHuS/c2i+O6xmWjAvAavJ/doU+GY9bTZR4WZ
5Rt33uZHqKscktyujuWk9vLhHykXbONhkSlHRYaxFAsDUugSldK3Umil8Xt7D4eY
Si6gMapz2BnnlH7oY0KOPKqIALcikQyp2BHFJa5+0JDpYszZ7nsxIfCyye6BWhR3
etQ8C48P93d5xhA3wT2Yc2s3nzc0+B8k8vsfzL2zEZi54oXaXHCnXQtedRELPseZ
0x4zMzPVjErql8Xh9YjlacQzHTlXNfYhlggKEKMsxUPjr45+Kn/E3mqubVB0gibF
P7J/dKVuHZporEy2GioD8MSuPRvM05aW/zxn0LMk4w1G/GwVuPmCCkgdfax0+njg
sjyzsXnsObtTOZuo2akGVzr+66sNJ7C2Ci/LBZidJeDbDh5etmNf131MZFx7XGX2
HAStxBO1EobO5uqaPwdKgciJmVMBUUeikecBoKbck+jk+danTBB8v27JSdrCz8eE
vX8lJzFeTNbuUGuBjf4+Oo6GTZoIj7CoQuM1GKn/ME3P2m5OnA/2arYSNoYGAWIf
DhCRRhD2eV+IY2Og3BSKmnRnCAE799QiKD/nChHmP1WbrOP+S2Gj3685d2fFKmzr
8g5hcaQWEHJhTDmm7QtxR3b4yuTC24DoxeWuJcE8Ra0e2C0jhsLKcXBilutaCSzW
hskQjBkM+3ShAPgNF2LVyYukjBif5Sn59n7sqlDZSE3Rv/vnyRLt0U4Va62ZIB09
Khcmj8nFqe2HRI7812yVWRPJVrkoZjhTxpD94gBIhTTQ//myE0BuTTpRdXD6300Z
6akpbtLJYSBdo2/5gAI71fe5D0B3oQQguoE8JREpju++HFRvsJ6SOocCug3xhFsN
SzXeun5iId2pyu1nkBxb9Km22afxigjZn1vyiZDIqOjsdRmozX74onMgal7XOK2V
siL/R3VY1COqnLFzHlVndDvWvY69rhINVPXJsPWaCgVDGbwtrABSj8MKfpydTa75
spk1tziCfzuYEW64xmhfksM0nJQ3/mud2WpI/5aRX2k0MfAMPSyNHZc9hCDTMfH7
53OxokwF9AN5Z256oBqMLxN9TWthjLVjpSurNwm1Fz3UMDiOOyQioZEAmD7+sqfe
ZdLXfAVZiTuuzWo+KoxPfQjd/mZxbRkEN5YRSyL8wMOWffChL+pKBES3pKjoQLPw
OX3Zflg5DzIbaS2y7z2lqwqOosps/j9Z24/fTAWJ6+FyxVAHtno7FAGhAIJcbcp6
id3UVHR2CLPozBCev9UpQSlKJHhL3srhDaLBo422PA11mBi9awvlDhiOoDtIKvaK
BGzk7bXDWWOoLI2QRgatDSPqU0IVn0eJ4EwHsH3UgB99PZ8YTXyTRg4vYUPM/Uc5
IS2hU4LfjecHh5GAy/eXH+oRG/X+5+NaVf9gh9vYxs/n5uzOZnnBppV//dkLlBmj
nLubCrVZSfYxoz7qyr3KFPZPkAwTWiNseTrEkXqhwDbnqJ9gpcCNqaE7rJ40zV9C
sZhCXmAmaTXQN3gprU7Xwcu1tHp4fPwBO0r2xaj62JN0UJYCqlMPjpWf1yNNlwSC
irHyz1J4i7Sm2gl1aoHLbnilqWDT8Mc27Ag7bKLwrz9ifq4SQvwejcDvYfqptvhC
uD2PgEmLls6PT+XDAgTgpfnFDJSFXxR4cOYpXmu2rEilGJmDJoH0m4s9tTRBMKYi
KnYBXztCJCQ45faTqBJiZXOZBj6QGxYbGkx2RdKJjy5TuOmiVZ33KFVXIA7udP5L
Ker9MkAHEGckR6ctcbH85EgTM8dW6xCa4xevAXxOoXOcxZyitiRqE3F1AfF/702y
wKc7kAQ8wnoF+JyNa7UuWYKShvD91IMo3YaTD1MjCRjlo9fvkD9ebPN5mUA51C8Q
qMsjAL4kNWqunmDqihNrnDv8KwW95wjg9xXn9UeuGHd9dTd42u3L/bq7WOVVXJGN
+7JPtxwhktEzrTcbkZhWJ0PaHAnj9PojcTamptFryu6EqnzlZlj1kHxi0c/2I2EX
pclUmh4XLPIv/5O4UbHuExPccsLT8jbFCGUSGPSYpj7nu1fbTePzTGIyygaItlVx
CMr+7oD72MKwiia8ZmFnDoqL2KLqsfkA/Jdc2v3APYezc2fm6NBnUtfIx/wTv27H
v2E9fRRgORWG0CH5e5IZ/CtvRGGtcyoTJDzdOmJ1vXq5NXwuAYmqsxc9j1MHABGK
3YULMR8V6TfNP4ixsqQ+6YYCxxuaauQkRcFnn+/3Xjc/d+Oe5Mjb/F0uZZ7Yvhr5
QWcKrFV5TLDNxrbDqB/pi+o26DvkBxp6/8FD/grYOkNbVSKmrXPoN3yUk3648kVp
ZgwYoYwkuEC1qWpGxn28Gka5cI2ak0ogoE+h6bfaMwVdGz2tTdlxRmi7FKyDGhUz
0NIMmtO6jZQ7z7/G3weDQp7PflMNYd2Mx54kdzzAtrF/JNlZKAG6NosF3PHCdx4a
8C0MNc+zEwsQIxqZR90bVfsGgOI02Qg77AfncnzDO7svtouXcQ2M4muwp04k6X/M
smMG4xOTiGMwC3MoEE60aeYJjtY+HMgFE7Aw0KzsHfJAbR7Nc58Cf2Qx5rEbSBLJ
wG7J0oitWksb58Dd3ahmR47HzODOFtuDJjnMyJqwaITtwGU8NiInl7kXbJJP8yx3
HA8kxL1dezMVm0O5PodBaIcSlc+EwgWn1mAEh0d+rAK6pWFnpRcfufML9qZHba/V
G2CMgK9i/P2K/RT4wMAEVuKhPwW6QHw+/ToJWKwfCYgL/PFlUGUGsbP14h/Jdj8L
nCTa3ddfdr3Vnd17lvE5gOIsfir5bAGF/guECWKYkBdZwTqopyMsIUXdDcX6hJFb
EEpXyb+ELXUXfj/zHjmOMgS60zP8yMFM8pwj6trfWuWOGiSQLNNylKfWJnQz0+9a
i8nDfGvhsT/VNDYnXlFbImQfznMk5lySe4qPaB0Ps7j0P8/cTUeITJQ46S3Sj4uB
YfEIsC+E5LkrTZbjCyFaMN72w9t6pB/MsuTTQNOhhf7Ott9sd7WNeSs+R+vADo5X
yCpbA/HlTaZaTTHLWLjGg9d8YpfLiPUSjPOUGBDjSkYNQlhdnEuQfwmlF6A7TB8i
A9EGihwB24YCFRCrqdtlVJp6IoWhaz/DFpMjBFrX7Va1ZDfkcDieQECElVGAMPZ3
koaHQkOvg7VfpnHwcrn0O7cRd+DQZSRoW9Ml/5DTvv32eByEhxizsIXOFNtgw/iZ
Se4x31qJA227UsgOJYLyxvV4M/P+/nL4+cwCx4fJAzbuPUKk7UTec9ZxCW9k81nl
fhO1MaIOyGM40j2RDbm/Nz6sgOyei+MErbrDKIB8tMCwcT0xRZQkfAUhPEAS7KnP
0JLsIqIA8nI/n1whM+q540KUXXkqRHMxtsU0odbnBKf1qvHb43Jefa1P9hFgVivH
/CA5qOlrcbW1phkQ8dS2d1xKKbcNSTmSabgzPSIQI4ucu+JXk/TWZEmQbfy01bzV
vJZd/XYDzxwmbZh6/rHYMTOGuMersr3b2M/reWu4dE4qgPBd2SlbFNCfmEtEcJrp
Ve3ZoPhM4UHziSgukfDpQffRMDuoyzEvuJgfBrHosdGK28y5AATz0Br4we/NYeyV
m4lMZJAwoS+T+5VkKsoAvQqtwwmEcDPdj+lGDQr3vzydN+TZPghBflPouydWXYH/
VruVfq3ySiwLcoR2+9sKB3Crku1YmYtAEouv9/15lfKbF2UG2wYrQugqhJnJteg8
YbO2uVpD1TcBQdLCp1HgJbpQCjm+vasGrTIZMgMRE9C+3l6lMSFtpG3QDzEMXIYA
R2HKrgUUwrItkN9ainX0pY8QbDGTeF21GLf4mg7FCJKjMVqFaY0Pamz5e0qbqUcF
1Kl5qOuzBmsE5aHazBcBD5QAd5G075iaH69qcKPuTm1E/ugwCzK+ErBgP/L9i974
6HI+jLloE8/Un/p0Nx3Z7dJ5/JfWXKuqJG1yArkHsCx9wtf+8ROvGKsBeK+Dp/Sc
E0VPUGfqtkRcJ74rlCfVC9ZwE9fx7swQVlh2Vyl+QI2j7zE/sIr2OopLaQ3n67r/
yMbdyS2DOZ+SNuGj23KTz3Ek2tesmRqdFfZF2VLtj2Cn4pHWOjJ+s3HqLGtyd6LH
5LFUvSEY1S0qJZvDl6HbKR9kiq3TqEFewgkVSYluJgPLAIK7LsLBY5XFyeSXxOIv
b5SM7DzuD94OIPJ/rOeBoztYO7tMzvQWPzhzxT2LXgZSUCsz5a8Xp1Gvg16iPPU5
tFvvfycikcSRVZwayWsFvnud2W1OMy+o/Ly9I/LR2BXozpbhYvgMXtzFs9QC0FQr
vpaNai+PI2I1rzR6cd6Uuj+aBQ5aJ3SEdW+0aOMUhSE6CYQ/eZzNov/s/ZwHDvuV
i0xi+0jMxL18OP7UOHi5m1Ykoc9zimvOiuXn+7CX1xkVPyPHlxEFHf002WTWE9qw
ZvHJ4kLGSTR+pUpA+m79MPJV4nB9qAjIoW1Sas51Ci5mXUASWqzv/mcD3DuP+vqj
6WcSwESnV/5PIK80mDqQKlwNby6+rhVjHaPC1gIZmFYzP+ORhLCr7v4yruTz+AXD
+HOOptVvF2yZJpVUeyP47DyUyRtnJS+2AoZk3KUY0d9ER99AdPVjynN5MsFgZ5cu
IUzbTRKWadffwssgmZtnUG5161H+Oj3MmA+k80lgo5A1dLtYaB+Sg5DJcc8ZXlOx
eHyV4NLDDc+Sfl1u6sFruXi0v1BC/2Az7hv5u+g6E5naHUxyAqY5MnUss9M+8Ttb
04vqs/qHwyErZf9THw+CdHo8UCUkNPc+kE2cYloB/mfF/4ft507oKijVWB9976Gq
Gok3bqGOfOZHIaeBFzm7TNIYA6d+lVlTs2ICnkdEH/gmRuPrELiMX95Awdc4IaRb
M36NX8ws9MMdi8dgMYn+2JGAHFkoZtuqKKlCVF8JHwpEx+lJF5dstWhACZbXttnA
S7KcMrKhcrDXtaU9/wh2xS3vK7uojIisduaQTe90fJxM/zJ/m69vtjCy6+t2S8aA
uF6s5z9tXbrXRl6EUfsMcYvixC/KMYPUPP/Xxw1dL+fVP7hGENrswtkYgH24qHI/
b3hHKihxICCVpLogLp1TWukkkobynyBB6+BSCiyq2b4AsA2chvmKgwepl9WYn3B2
k+opgnNNRnLWWUy5RebS5QhM9lnXeQnH4AeRIWezi0Bi5lLRjwAWpkioBf58NhTx
ejrVo696u+be6dpDeS2DgXBTsQN+5lA2gjQfwib3Fv0dIn8fMGc3FgkUl9O97L0s
0d/50XgsZCtNIWTvWsqTCihA3jCklVizxOHlFpAmgzKZf/hP7Y84LFEg/SVQ300+
U8cLTqNP+MQ2d29FClxJOykUxe6OjnLqsDDaCMikaUFIt7Crojfpluhzzyx4dCPK
u8+b1ZevadPzvHZM9Oh/Npc0tghVvLEc52PKMp2SKn8PdXhvzsPxCjpZRrt3gYw1
EX+qrhndea3uaCkKJv507BEmuobvZNsScAqZhX008Gt+XjqCv+yjaqhit+2zSwl4
gD5jsDAjF8/9Am/Bwwq4ZqFo1Uha+AYH2k/YKXZ8TMDAmYe6r6X7j2soHoalY+Di
a2gj0J4CS2RtfY9DCXOg5KF3xXxHbtlafZUMM6d4l/oA8s3DXed2j/bhgsy29B/N
Qax0ec0A2SC+I5aGfY/oVQlhgQp6ODtREn+ej+rW42szcaCnOX5PJ0z4QjMHH1b5
W0OW4s1jL6VuxXrbpKEHukHVrMsrwL9fMeDw4ZJ7l8ZOnP+Xo6n/RK+VxymqwX37
9FuJqMNzIWTZuXwm1luQofOz31tPJTLntBdAle/AEkUe+as7GR6H3jNw9Pk+yaMP
ReHBraMFWSSFcPPcEZmslHinVOjfjs9jSA1vqEifknsnB1iV4qpOyqdEQ99tNQt0
JvO5jJUy4r+8JKn3qGleNctcep2x2Y+QWmpO9JhlP1Kf1n6ZCccRvcaHTvE3t3hb
XqB+OQkYgi2xTzWol82LDPKQAYjAvYYXblc5LsUl7wPhBEIBnUEHOu93PkfS2E2+
uEAwuxahb9LQmpbWAQmPXexwfYJRO5HJyDETgQSgbYm025wOq1TlsnVBj2fPXcsX
T5RaScTALODdZgmhQZ2tXBi/Jg1t42kmkL1HVoODsU0oHxE1vhGk9bhuvfLAL7VF
vRwF451FU976Mod+fM4GwjLsQm+2IqAFzW22rAspYGa+x/FnUSRf11MNBw0YmEQg
gnxcDLLEagzNu3dBq6NCJiFvFcKEICE5kYPCzNK5akYI5rkrAvIZTOVLOcm+taDq
vk4PG8uMLX4QwK8l4NPqyp7BdtV6hsMrNDINPPdWvLe+HIjfYtDLzaSZt3xDV9tN
RF0lSNRF4awQuNVcpcOG6A49GLQbqVU2bzFLrCUvmACgYsH2ugHiTdQylS9uEheS
zcAQuYqz5oLq4k+beqTYUtSSq/BXazahjaGdcZd38GLjtp9XiZSTwN2sI5Y9C1RR
1MfC++D5goX97EQPCoLT5oWruCOW+RoJkc6UqNGyF4W4DI22bKALMKTeS3b0kRdO
EtpH0djmFGAzH10H1nPmN8TLj0FkImgB0rmDCvac3ioXA5rmLFV4Nx5nzKtlapje
4U4d01e3eKgj+eoebRSzL+rwwEsc5PTwZOgMa9XDIMJgKLZ1mWitW+8agSedQv29
1OdhfRiInOvvn0OC7Jyjh3Dj6shlvgk3ZcUfzrecWGdbqSs8FTFZu82a66cn9GI3
vOVpC5QqMMNegkeQXlz3e3XFS475kVkE5wNMtBj7RWSdp8fF5NCZLRdUjCEfl8y4
jPMIWXJ8jIyQAKPkLfbzKMDA7ismXG6SHaM2u+4xCRQewb/0JoBwssQZtSl6nYvS
AZqmpoW0kb895oHmi03BDHKu0g3sq8Z89DY7quS2hH2gvRFSqy5ijnLX9mXebXuN
6o10+bnoaQsyHmJdAcF/Q/ed6/SRohxmkqnBkJ9oBU+S/I31aGHjDdluKrc+o8vN
8dWyaz/SHNcUX2Mh3Tsj+r9CrLAv0YrcEVpmLV+3DWUQqbRLIfd6f59DbNH0Ilz0
f/qmIjh01HyeTXmL4wVV+zmxLbRknxi0/kZay63UjOzVoW8ZVC8lQ9+OkHaZ1+oY
QkyhuMZoM+vZLwxPbF6oOLqMMqNI5kJgY3rEXxetfvNUCMnuOwL13zmBZv5txQ+T
QmItA7x/iM7nswvHj0rZzAXk3z+n5hrr2bIa5mdaDEllP+erFRKzKh+E9D1IkUUJ
TmgpUNAwJw4lvvAj5U8xkKadIrAYJRhtZiGEuLZ/b3pmUueFg96G1HqLJVAGfGxb
+XeEsxUSlh77ssEAdKTR4Xx4gHkDWnk8q6RNyTxrk7pXZbKDAzvOR0OdleEmcBVt
tjpeXp7XrnON2NPwiDYjImCvSosYTjAHFmx8Lo3OuoBok8FH0qMsq+RZ6rSDpSP1
sV/SaStu9qImOHoPEUsdsyzwzzyy5hixOw2xsT23V0MkCVdV5heaAoqWxr0xnK8c
IUAkxBPnpAUPwojPNxwpWytKm2rsO0nZWGmX4JbzQB1EE7EHYFDStTkrcYI5sGaU
oJS45jj2TyXyxl2OnhRFi4WQ6dHO5D9omgrFU6Dz94U5xp//2pL2hkIvc+UijiO2
Mv7zVYO9YESUVBOHQcCiUH9gIWXplV0SVL5icBpEnh9/zLJhGc4YqEsrgnOKZm8l
5dqJWudMzOOE+2zeBqwAA21dTIatsmdQg1uEkAMxau64UqJACOd3+xzd6yTEI40r
F63pvjYHKS/dk3CmpIcqyceR1Qq4GyYkhHA9zXw/DFg2L+YuonNoA/jNB8WOacEd
Sgm1iVPXpzK7y6zcRp+9ZRiXcqP/eoKi3WeOEMub8eatOxy6hmzJZJOhl+n0reYt
3KHx+lWTSC+erB+QBSdxklz717K/5ourdU+IeYA03BWVthm2KOTveEd4KUMsAc3b
gaptoBosuN0oCRy+TfERbOV4AybKbea3kyIjnY249ug+gt6LaTX6S1AciC9lh8vl
NTja6yYMFdToyHnxFrbXcJ+80Ugqn84ED4UrauHOuTs83LrdhE2weXIIOrYUctsc
gZxwVCZomQzn3bno2BYWVXV1e7KyeGYF36VLVErLZb+q1Pz+fKWKuBkybnf0+X+w
C/S0oNSc3y6PIfC6JBpzDXk59CA9CoSz5hvvhnkt0mx4D89lESzchk1dt43SAOM+
kfnfxH+Vx0KqhE7GMXaTs0CwfdBVC8p2yNvkZ+rQWB/WAcRkWvPpxrQSUckjV3gT
UIRt+/a1+nBDalaB5Bxc9jZDRzauCbxmyqdnIr/NEOPRpqaWPYOoKJU6hcFXvmXs
0BKpyLi3pXkyGJd2iL0IbMnneyBq2YIHLwXiqfVDE/rESbXVWecZnHhnK9Rcx6Re
724V+1MiI8fTrACrHF1xgNQJXO5wzo6k68RmpOdD0HOgPUM5mIk9K1FbM1ZzxnaC
CxKJcFMmU/sLV+1hhhezBh6qBRB6CdVcw0QDYxqKQQ41b2JrqMBVHwBFPaxzf0EX
n3Ey7YNHzB94HInA1YGx36ftKhhC3kdoN3xPEr/YcNsNQmCYPZcAN0z/bU6kHd2e
qOolD8nxMlwe2fGGqPg/y2cGphLpeHLUEHksaN9tTUrUM6V8c+HbZBGnBX+cwBwl
QkbNuoOho2kP0d/TGlRwZV37iqecEH2CMkhn3AyxjC/zPQ6Lifb4fxYbLAMD4czP
tr2AmzJwb5pHipvR3hfPKJHS0V84tNDozyP56RBq7nwlr1aC2YVgvvPRKlsCTZrg
40bpvQgsUAJ0E39VFoJ4e8QDNIsMRMzY3piiUlSrw4K7PtQrI75K8P1vTgV5vkhk
dmkuSZNt7TMyBJyfudjzKrDbV9z4ac//pjqTQURFO00/+yJQpnhulAZo8jv4GrFA
BECwsq/xjlOqNvw/FxuHQpql+eTTGCxKEYVLBs9ZAuxUCwIFMk89EZbEoPC2XOxN
1pF2seH3d0cfZtROJBf4mhrrRCplv5zH7srgbQKFNOpSjPbY6cuxVUfEB3hn9paW
4Ry1ismhP4fJeCvlbnJ/6z/CZaUB0GvuQW1tx2uidKX/EFWo9DCs32BbyIHfDeQ4
PGohqCxz4+tV1tP2mhv0qPCrSB0PX+rttyKHJXnmCne9PCABCVMOFmbSb9qigIh3
N0j2p7uRE4cpQHwIQqggefwt5RFYJCHWGjPkN3qbTSajD9W+xa45XkXQOHJWGjmv
h1/1xOq2gTC6roplJUD2DWuASnDJOzr9EsyOzTxTpK5sIRgeTasZGgsrltSyZyXl
YqOWPrV49tojSl6z8RuNGir/+c2WKuS3nCvCwB2KlpBqDVc6IctG2Pqr5i+fdJXl
nBvQ4rDiPQRd06yi6KZoq1zgb9pgAqUoLEY6LwMxi4QE3SWWXoFveyuZy7rMeL4E
03/fivdFCf6Qaw3T2rlQJWjgRD6u2hO09xxk5PO4QG+Ipcz30f+KE3Xyvymifgk8
h2Ase4/0vyHjPaIRKl1OsiWJBv45HuCsVmtdJVaxH9wHsT2EBdI4YLnoN26iV19D
yJh8Msf7utwIna6iiZ22uC1UkeS3yg3ALbbPHdAsbKG+5/50wouSbsw5OO+S9VkA
WhJl855osyCd1gSEQBlFtBxjctszdX5uh8dOpHwg6Kt3BWeEmPRTqM296BCgjP1v
xFldpqFXS/RbiHtn911s4KcDZsO+4EGCnDkCAWEhj3fcZnoxTx4e1OS12hNdPqWE
eQOhMoEq9iSuvPnKcujD4+JOUZyh3x3rL0f0KpvikNekZsMWYOrdvGl22217oudz
pbira2taGRcjgI3kYgbl2SByhrJGTcFEPmaojdBo+TrMrMv+/kJKmWlO/sNDwHgM
311lqnuk6BX0kym5o4Vpn1A8XJUu6zWTVTUWVa6/JiiWr5w9GExOQ74queCzJzSH
JOEK6ylwGTWYm69C7OA39yfIXaM5QYBuoHMGP4anpRrhzZLBYHhMxnr0BcreVqyk
EirDxN2q9M/ShSB/LHL3ZyKxyeyAoDw1DIlwCyRwUmeCLDbzyVxB9BG3bxTgqlhh
4TrzoOeQk39bfb90Djs73a5KASVmwphFu3bjR0b+uVCAI/3ahcCxC51ybgrOy5NT
RWKfe7e7dWn8HxTn/Kq2LuIsgDP3quPmz0/QSfGPAUOhX2IILdnqq9y6GsNWSZ6L
zJggT6MJQY5qMac1OjhaXlfhCpaSf4Kbkvpp4iD2twdKH6AlYaJiJHojPoxVSd2q
jcBKjzUv7GCAM03eo4pZyHlZosckNb7JUs5Eia82rHOC/kJtRz82rtOCiVo/on9C
/tk/FWFAtB7xmrvyN0HaU/ZRQ0u8NZcPKBKwGrcRTqQL27dBkaCQ3FwSXaMzCdUy
VLM9o7Blpf7aLvQrNgx3AcRizHzHjU262TgTDbtOyP9ao/LH75NiezMjBPGUrvRJ
YuFruXvgpL+GBqgSsy6N/DoVX2KF5CsVKa5YtcUSTg2+LgigqnB9b8a9/ScDxsYa
ykMs4Dc3tANs0wIQrnVm4VkjW73d07QtaGe3diCtG2YAbJ+nu4ioE8TkR8HqpFBv
2sjP74nf3H3PUSlONsMx0GmSBmj5sHPUawDmDJ0Y+PTWAFQmi9GrI9Klwqd1dIMn
BV/6gSY4+kYkNLKwdCD8T6RkepxxVjUBav6eof64yjeTNnA/q0CXs8lgGQCHGSpQ
0yhBl2MZIeAysfWh5ELIxs0rpIhqnY3aw6fLna+3CH1t4aW9qLj+8z/xb938od8X
iWR0n0d1Pz8tVn2aT0ALtSLuWNeEJw6rpooWDmLbBQ9s1Jicjd/MLVYP74ybCChs
3awpKvYoh5SnUKH8kMmjXKZ80fpzQGp0CUSuAaydU4h45eOT2AJDAZrc1XDppS/r
US1uCrJJ6n4cWMGpgHgXi65DVaovlrCwP5GVwNzmpxbSp/rrSoPsZVWSk/VdR1oL
yExrxI05DmOxJrj8Q/IVg5qXs6adRt6oUepPKlHtx6P2X0YMhYo2oDAAgSwXBxT1
80tJnGukdtSBEoLyYuA3oKcmtNh+/k9/HlB1qguNzd3pXMoedzKdu+Xb+yTjUMCY
Nqst9ihWr06yQBfXlSPF/qdpu7pkGH/XENYnnKRs15GN4Vwkmtgx0/m+Nj3IKd8t
89ksZ5dr5ASlF2TBjhTyZW04uziKLYSKdU/JTc9+zAKD1g+iaGu+TmqRnnA8ZAEo
UKDCTLpzDr8Ime9NIqSFjWFujULMBCfNLEL1E96AHw0i3/c+6L3y3k64e6JOn3oo
2biD39IrkIcpLFwqJgAQtqMKB9UMB/EG/C6boBRxl+jYCRqsq0KWG7FixIzz+Xxw
nMJW4jt4zq6EwbydlwDJIJ1GToYDJGwI20nHCIuVLyELvJOZJT/GMcaiwQRdU7YX
1F0PG67tK3HAyG4aSjKO6hCYo2Zf/sDK8IFgI/ea3OPiBurlqW/NeEuWWKgZ5aCM
ucZhAcJRMzLyaFYX8PSQIAxFEwN94GtXVtXnZl2roPW5zlSsZlcZ8fUxaLCGGrib
X8hk6QTbVVZx77M/Fh7MIncLV2e4zq1/eTC1pBng3xGw4WXxn57XyrYTpLg5g+Zr
m6zERIofzgLi+XQWMRfYfw+PaUVfIrQQH7+U+O9JgcMlzfTRdcyhV+IZVi0oe/ns
Hl8Grf3xWjWHryJskKLzHEdlUF8mzLTjHRi4GdfwtY4GymD0mPeqjtwmuBcJswXn
6BK2BaUm1aIJlu1OjcmQRANBy+jp2hy7oPyqQBRbsJNZudQNYi+87ftkB+CjZQ4M
FgcMko8ViQMCbWoO7tr7ZnXgFOirwBAWfBXqMzHrafUxck3AgPyv1/b8qNh2zNUT
0hqk9PPvvY1TJ33+lSbgKfb/4IjYrZf1YW+CazMfoi5Q9IbFUX//nX3L1dq1arlZ
kY7gqdOKAnVCIKaG7LlU0LMU7xgK3MXfC2wna1vjl4lN70QPY2p5MoV8IUR3YZ82
PxhguM2Ydax6lBZ89oAyrCHNI0tosgMHv9ai1eHbsAF9sPJiXpFNiBOj+Wm6bKTr
p52D6i3gjG+5y7OU1G/2lMO2QjvP2muEXR/0fX2RDxOgTigNY6QwBjgmwm45i6uc
r33bwugRRq+zayxvNGYr+0uATk5YFsdilE3tcC2W4Nlu6Dd9sR9+Uanbf2dvAtAU
Uubpxeke7BaeJn4Q1ZIeaz46L6o1cqvHWTDTcw5RozweTp7to2lXqZNNym87XTLn
dih9/kNz0AbjVxcI6KQQ1Lp1TZ94CGDJQ6mP2UEhxSbQ8TgyGUEv1u110QmX6d83
O5HgTb+qXWmx5gZc7CzXsrjAUKL8peK8RP3im27u/CTEsZrpQXAYh7Y8EAvpGXhl
5gsYZ+2SA7OXLRE8G5e2pl+E8tgqeyxzpjFJRbJb9el7+yZWFu+cN0YawAF7qdTP
c1wAn7iGPW5ud1PEHtwBbHfEdoS4g4DcMUfn5xlEmQ10tjHQj9MCMlzE3F0QrhXN
HZ/8Z+0UCmf5MRIqGZevquDjwpewX5n8kkmRtqkU65rEMTA29FHjU8n/Vm8az6FQ
3QSt1enwSUgz/4ERFA9i2NvLph+lnWJgXppHgR9pRTi0OE0GpwVKOFvWHzvx0BIg
5D4vckT2HJlQMf07/O65j7uHAcVbp8s75M0zaeurfYXWWUHPCtSlgXcPrfOXXJ9W
kovaSHwD6YAl8I4YuIgCz3f9K8ZcbP5WBY2tguwAZhahlMUG4Q1KOo3dYssfqwVV
vRO8YciwAWvkIVNp7Bz7T6noeIKxDD1NWiHPDRffqZsdp/8WxZusbS1zmTQapOvQ
/Ea6JzF/jcNmmhAj08nyFKfWNdAdSJMrEKLIGMQyXzFsjgh2FYuoEfnFMK/6UbzT
vBROXtMYEfGrMvtzJfAtIF8AJ0mfio8qT4Rv3cqfTflZLtoUClM1rKDz6LDg240D
vqAGGWSjmukFayaM5DxWPkzb0iSusL3aAuYgDmXcnD1XR29snNFmHJhBph/pU/gC
9kzI0TJ16cstzGIWnlrjkxegK4Ng9KEzyTAUewqkUqxTCzxMHwPewHCLhkkjRrqc
c/oKZF315FHeYyV39YttZhoQWD65eWSVS1w92ilGu4i2L2CbH5npqLcqwt/vI44N
c5PIFdGPA/74yMDO/Zb5YIkQB9pSkiIXLiRak0BmaX+PSoko2JFtPOog3xSvHpsM
WaXdpXcRwrC4CHcNboiv4P1Sg56utrJ7W7+JpwvElQGdb7L8nj01htmi0e4i8qBN
LKoNVuKWGyLPFoUvdkptK5xPPl4GXZpBxPm8XgV1rkH/B3pRqC0SNbiXbHFM9L63
OkQNOcdDR4LzSlh3xqVFMg/10SCpjSvTMSBLpcFQIdtO+bacZYF5/YQjQeN0NMlj
CUIkrMMHxMfiBaIhFC+jrNq6AGujEi1j5/P6YZOzyxKABTK8oaJAaGklNkV9j/P5
bzZJlaV3B7JdY02yIWNIbA9iA0PAKiqpMHzIvsw2+k48VHhrHtl7YqFuav7nQ+nZ
oyrK+SXdx0u9Apfm16aVfY7O1BDM8C3R8Wpq12Z58lMfBNnwYQx+pfeJ8g9puLaw
PRdD3hA8zzNI5DyGhQlrMUtNg3nJKjfhptBtZRMwr728HRQrDMtIDFbF3xPXBC07
YCq8ZZA4nlUL8+eoI5RjukuBYXzGG+6eD7VF1NSeXlXDxZz4GNm1EeOnNMgWnRmG
FzUKItu4211JmJockaEri0QC7LKrwVNButbQ0kCTGXIW86wGFi0OorRfnOuHP7KX
/PL8grRwnpPV6lhBBodDPi1oDAUabGT02T0AcXcuMY3hZDhxNJdrJPbLAlonMYgA
P4F5m7QfzMiZ46lErhOAAurqKEtY7oBRUPCGkX/mnk0aTQopCCywNzpOIla3ph5i
Yj1TaXV/y5f883NKYVBguUpA5EXe38T+Mn7Id81KYSBKUGs8BUscLIrs1rPnhgdA
RuJmXTtjKNDzVwPqy4uPY/opwuEb0PPl3XpDAFReDrljSqIMD1rlcIJhPWo12Jwm
eMpuoK0yIhizXm19OvCUOmtvJ+KN+YkPqWltv08DPyhcaT4nfMHSdTfrVD1Gn2OY
ZInB6cLsspJ3tE8QQBqdkDx1sACWVGh1dAW9ZD1bQ9vCkHWjtdUaa1yJaRG8rMo3
2a3xD2xPNTYfNLxZSTBz8H+qyVtSHwES0rOgEoFe/uI7ybJZoYidTsTBvIgv6ZIs
Slz2GxyoQ67We3HMhK8uth7zWO2xPeP66UsgIy+gSBbZY0XvgPPhLelEGsyFUe8u
0RcfhM5rNocCr37bUzCTWcKe7d/0lyRQ1kE7l/+p8eFRGmFbnykLMEhRCeO8UZaq
SGZXzW8cDfLmQQw72jSG8lgKSiwyA54pVBPyQfUB8yX9IDQ0bUBuSHFy6c0Pzzty
9YYPuIgoghEm/ssPnxnkIq2gRCwqrDODETOnm+JT3netVaULTGwsQr0O/t/aZVb3
67UU5lnxHcQzCqN1M37GfJFCDkLOFI7bAvh2plU0/BFvJCSKS2ZlwaoD2p+FSRGU
U7CC9Fgezv/TPKky7/hPU6y+IFwPOrKA1Ig0V8S6fO8cWutiRZ/pWaCJ+L0xTW47
WXA+VLx54bq+Tw540wEP/Yd0XyLQY7TowbEWLv2A9hU8RQJBH7n0ytfxds35y4Be
AJyiMQzL34cckuConY0yb2tfUd/b/W5y8q738JGwvxLIpN2pT56v3IVU1cvDj1Wt
ZWsPs5NtTnfPcPYUo6d7CoMTbIGlWY8Ea5KpTVBloVJHmnk+sdmTp9BPMEEWoIw9
7EMpaopeAUc7o64v9VjqKPBgAogYez4mBeGp2iMAfBMHtanSCAhcgod/D3w1ZCw0
pc4Wxc6opwrm9ffntfMBWokUfriRNxSDsvRRBMq9Wrz/tZZUItAZpP8+aIFnrW5/
NvYhFk1SS2SRMXBnD/YhoqAGfQZHbo5QMyLjzxG+fM+2FQ1BmhOq84U8bkiV4V3P
l5vYJTRCAbuGMcZTW85tzWLz1ga/RgXyYJwZ1ilQacL3mqlDTjFJAAkL6pmkktT8
R1FIkysj+1ZY+2O+3BfBRG5gpUIWUx5weV5LRVme2jKuFHdFHP/FGSRcAeKkUQGQ
Aow/JrCTbfdv7pu4ZXHw5zzRpZZM+696D6LFSoypjl3zeDxZ+Kgivo2OW9UAulRj
+B+E2mFKIQ516Zr0RCaPA0pAWs5VdfqY+IXDy3HXZhh0wbBkERvnrW+T3bTqqo4N
rOwl57k+PlDXdYIv94UZLn3+ZskEpkNkNEy+FShhVihBun4CnVILVheNcBqngQ53
tXHbentZPkOBWQcuHVDzs3ZW6NTCbOnucH16QMX1ebOfu0PTcH2dw+UytPmKgEuu
b82Aw45hciG1r0AgYkBvOutLrJZXGkvZukaCtGTvcckN47ZMLXfT79aBRPpvuYPK
w4H8LekFsuHEPlr1JUXlsuxoZfVKCh6xQy65QPYL/LYdF5i49eJ9qmf+1NYTHVYH
OkSVmqQAz7THFYgWq6t7ji2MpkT9liPCqsUbDVFkx61aPyE3ciS/yZ8uy/QTs23O
V0pF8zyPJH+cTRPsD/G5xVTfWWaF4q15wJ3wG2uFYWJfRby8TbdcSw6j3tcWDWzm
mxbYd570Fe6tZ0Fb7RkaccpVI0wndm6eU1CUyJ3eW9q42wiGmb9xeJAAtWm/htP4
+kdivGBoxw8v45k8t/qc7XoNzA8ItIaPwLFNwFx0pwVhBK41x3oc+U5HKoEiKOoo
5Tu+EEEWp55/QuadoRv9CHZnd3GW6J7M2CHzqne0PdeRW0Y7Wi4IJbwxQ/GVyL6l
XeK28Zj4ZNytz43xK3Ua2x3PkEFsG3IZk5Y+6ALj0K9Kcw3ECMEUs6RZ8r6bd3Fc
abh1AuqfVvtq5fUeMngVzVR3hVj2kbZBryn9/oB2gStJCXWvTbL0OQSrcnKsizKK
LEwY07Plhwypw9//hhLdVlNgsH61Hwo+xZnssZ74H3hyhNS0ZUMqMUcCI4AU+9nl
FJT8QUQXmkXPAw43ZUr1jYTliL10g0EzkRsw3opF4SxrWRjl553nwnY6sGspYk81
1nTimHGNTQtncl1SLIJBMWfH/fW4nOjXx9wK7Vk+MOA+ODgowlkFBSH0GWjhbFaL
YOY2B78oLn73Qor2G09UmpdyBa3cE531DDR/fgf9C3+s2ZQKJmr+jHeAK0hVRhwC
xd5TELcEFORVZ4RLSD+cZdyXSQFUQRNW2XkGTavfFekDx6XiNclqE+b8TVKcBeJq
a2wogWsP9DZpJNeAOQtj5tFiT/w5+eGVSIk176LxLMyeq74ceJGF5iNCBs+w1kb9
zjVKB50rrnzOqdRaVw2c7DXXP6qVXWCcMSDq9ZLxGxxCO+HaLrAi/06kQ+XkCPGR
VkkyLIEBC+nHZnILBaqR1K/VhbExlliVMxVTKPw1S3ZU+iIJpR2JqrHfm7xFPdHP
EgXHle/dcXbBeA3HUAJ8v/2JBRgZ/miZ6KEVi92QGL8YtRPGaunt1EimxfxHAky9
iw1BfRgayv+KLmOJQls3PsLTGwcbFzcJA+1/luOM9xgYCjDuObLwELMwmmH2P4AR
n1hpW+bS2v2cZzfd5YNR072NgTBVAy4uuAf1RLvlcZy5Z2kM76BNonT7weBUxc5G
YIYvrquFPJodPwExdlPHVsygjorttkovUlkKLQGHeriiDN1ZBZhLkkTWxigBIjrT
7DDTAmXesXzxGmykRqwUWJFoxSTA9sSX6mrVyUjKAn3EXzl4thyfi7naPyVEhytj
G/F0VPvak3O/yBQ2dBR97iv0c/JHnxJZMhiLFIoxcT7L0K68Qvnw6wx+5CkzWmZ6
HAxUnjXhfMxwYjrmaMQgO6wIfchFFr6sB5ZFIl19xVybml39cMaGFoWn2Y8bcRUr
IoOdWN1tdlOYOcG04MjNzU6NdDXKPbKVsX07YGazsAnwdXRHjo+p3tvBiN2zUX45
mMvgtfjDBvyI7DbUKGutkO1AKh9NYdjj7mqlsDzIrRSLdrs9onDWZyo+D5fG2WWa
8NSo2++CgHKt9bqCFrHwzpukfjNPP0w+sOAtx7dWPUlzoZVX+3Pp8uvRMe49kjJ9
CbaKZUt2DzfSyKTyTs1PnhfIJImWX/lhSsCsanJbfG+SKreHBUyX2s5WEBL7noLM
E+41tfZQczccsrc5RKTwLupLK17q77bsnVShLrFz3jtp9z+tT35qfU2hd/ibm6rI
gKnw7UQzKbyEPO09K8xWSXeq//6gmxQM021vjEnFU7lXQzvAeqUYQ2W1wqaA+tv/
NOCbfAPjDLzgiPP+DRzyhDajXex9Ziyxl5WBB/D1AP0k9cxLDQW91vn3NPZb2ygM
OX62RejITCdVyjMrPWdACEFJpkmWQfFNROBpiSp34gdhF0lyhYCQMQyASOJEq4wa
7fFjIXZL18CelQ5D8CToEdER90pqJJX1N+mi9m7ZFk0Q2cJHciAOyoqq/H/zSFdS
dip0o7Xh6YcCPSXUy38v1yPigbbErLr6GpLIt3Mv45F8/L9lkixjjZKn769mL+lN
RSJx4Xw3rSPYXhQzTH2QCaHsWic2t//Ae1Fj+wDQbFnZU79HZ0V2kDBHJCgB5pVj
nA3zA+PTX32IGE5TryOeQt9jwCYd+KrV9jkW9SlavegIYfc+IO0QMHhhtAuvgaDt
5UGNC5o40DzEX+yrOhOiP9FHXpJ4j8zT4sShIxGlynh7uYhn/rEW4uM6/BAFbi0F
o3sKnk5wJMduwIFQtKIp5Yf+XBjC39S8S8CekqpseDI3VZwLpAfK67hmox88E93/
xDQ/aZFhXBArfijXLLwF9kUcddwl1Z8HPwWLM2Qo9iSsnaUElDVYDMpQVFep1mWD
s2uaoXZxsFVoQvvaWnICKUjmMnB6LbjZhQGLvt851Mw1UrT0iKI3HVFYj4yBVVXv
XvWPqHqfB9qGNTewLR6p/v98Qn64gKO/diCS9bdmLkJNIhTPrN8vJy2UZEt3Q04e
9X2p2WsWQJfENB7Fu7cKDYcZf51vzeHQE7uzwMaM/swTzTM6rzsAozIYfzOiY8O8
DoABFXvTPhzM9p82JJU6q2gtIQ/Kf2PR5OXIAiQoOKCJelkM+SSVWi6rfzXnyQdr
f/TvEqv8vo4op2OjH3ZcTHvdD34F/DgbwH/AhSJ+YAZ/HL0HJ6jcCO26TYFyCABp
4JoZ23556MDLQHdk3hupOyNWOUb3ja1zaqXImK7KQ6dyprs04UORn7JGnYMeGTbG
8dJLyP4Ks5cYM2KOE/XDzxeVnSRybbZ/h9xOoUAUhoNg4xpNfH/gwwqOQB8lkTGA
uNxgbw4Q0lnHQN2qtymvzWg3SZw+5K7L8iJNJUyZnkSpmTKtmrmE/piBq+/zwpb1
Z2yrlQ3L4Xt/FpIMcUyRnMFWCdes+cHdlkEvqRjmAiUeCKRxrjWF6gcHXAMQ/1m/
Fj1LaEdSHdtMwQdLTKKE4gFF/4xFq3WfSiwkGPstC81kLeWWG8orn8bPnpn4/+cM
U+AK4DF+dYWdhvEwYEH2Zcs8GW1hRXgFqrd2PhQ5LThw7hWXwkhpyHqXg1ltl/fo
ZPKLoFG+7yWUPNBpHiabruMBNKdOXXju0fxQClZ876iRbkzyiywvkCrgVgT68cfA
CxsAunpXv3O+jt6JApixJkglQNwycCi+rxS31PXKV005F5WUHHFlSjuyKUzjEfuf
gYYCIG8CcRmFn6M7TIUpQlTJCflI7GxRcBATwmooSnN2b6VTCmINN6E17+l3AnZM
pOm/OwPU0JyL9hCsoyaSRqBy3+vqeHP/cnh7QZ1hePw63kVhOqx2LUxbsfsNFBp4
NUn6vdQShD3uK2wVdlO3bWCtN9KwZbxNmuW1d4dJy75mYn7xKDynU+KVSkf+r/tQ
Jrnz7fkWmgYA5rgzZvzu2Ejfxzii6jj0NMPzTsszsH3NDCb+whTt3GTPSAxUJvHm
FsJiK5lvb/YC01Wrw5BGZmu/7z7U2Gjpjj8ESBfyHLaX2GHgNfvErUe6RXq8IXbd
CNccRFE6H9cww2PVYQmAebyz9I/Poej+9s8PBXUI1Nn6NtoFCCnOYFeyZkStR0TY
nNXS4jgOmRVgAK9JDnSwFojsY1iI5Lk3TAnUGbhb3GgLjG5JIOodcezki2j8CC91
jkpKfUpkq6eXLNssVARuuEEWC2iNlmxarg8/YkUT/BVHRaMKPe7aL2izCqTRGaTL
gqYr7PDu5FO6Gm0fVPFg9oN4D5zXA8JXbKeq/0nOgyOCT4Rc/j3xclD9FqiI1K19
/9sVUgl68D5WX2DjgpG6NwMA+W+FSrMqZkO2u+nWMycuAiRZMCTzjr+0ruTudXFy
o13qY2B13NS27EwT4OzR/oKYDofBNMyhEnkOcBO7CUynaCArtHQOkRLEcbWTABr5
pBesi7YmAFyxtGnIabhlXdXDEPGXgZc9pbW2POyeISSMaua1cHTCNyn4VMkTyIWg
NJvN8xODkZhh3XDLSbCEq308JrAGj2HBYRJlzUNVWyHrabOh09ggJbWf6zPqq273
WZWFqyNCznMoy9P+1n/by+kBz5/s9ElU1KkSztirk39G++MsjvTEsOkE1gB6kEEZ
xWCsjZqKN38rh9t547t2ukpBBqcKLs5HW0oi4paAOEQwKLLkWXDA+4qeCSmGqL5M
pBlUpLTWOQXpNCW6uRlKATaC5WOxKYzFN6ABVBFjXSJ8c/eFYooefLSzdXGqxHIs
E6Cf0g9gGB1FFPx6t25RgdV46qzSVOi6F0kE/GGNpocc7/DaSHeO7WWWw20g9tjW
3SgU+EnihbdFz+S/Wf9Za7GRbkv0yaLcf4tqh+FlkyX7o8XY25UEb1kzNoq07+v3
L073lHEJH9Ls1ul0Xxtmvs7roYuHAayzAB6FJ1SE4hTqS5HXsrH3Aw+DmO/wJ+An
imWCy4Gne7/VvHVjZyKknZzQ65TAMs2BqZ4tTXGy464SuV6EbQ1t0r6ohoSLjIqi
HBX6rF7e61JVdiY8+yOIrb6gHk18+4sPq8Lh7/NGO8mB/+AgHeAC0oLBFw93fVtw
mVNIo3Dz12cE1vRj4oNse5hSLj4OE0Vf+SCbHONkyUzAXRaQ3ZMnr95J5hFNSdPW
Tx21XVu+jENqOnrvFOcmbxtFsOwg2ObO2V+CZAz9dsvy+fbJsK2SJQwL7K7IKBxU
ZsmbIfCaB85RYC6030YVpyMLnQc/6nVw4u+HaaGoa6cH9tua4f1q6/Q2z1pYOb7k
PWNauJ8hCtsEr56mPdZdRTWwwqmhV+RICXX4zVEMQdq/Yofc0HCSm5PYJXd2TvUz
2U23Z403SGn7dys/6hexxUMqPCDb6yl3oS2fVjzW3cyHS+4l0XEYAdihkFMCq+5t
q6kzkEi0NdP4ye9t80SwXOPAhxagTtjK8hktL5rs+NSeMl07TMKbjA/dUd+yw61s
132hn94by1ObFe5Nsg3auBLMmZES1mk8dySHhm50R8Z1xhp4xVzTVDlZSDLlWgwY
wEFNK0r7RWJBndH7ylk9yO5YV5UaGEg+N3m2IhS3UKaX4z6dASUgutqD0zsW3DbS
cuHxEP3+eVnF6O7AyPq07x/VYzvFaEoRueskiSIZpwlWv/QRbr0TuC6cf3HeGclv
jTJb28Y6PoKsj8HdxkXwCoQnPDHAIc1w0oMtvWYVtL+wamAnrvtEI0+Jqnmx6eZN
jDS9fHs4q2+gTesE/FDBwGAUvAJsEOoB7iVp3Q6UTkfLqI/ZAMwmRvKwfYAxynRg
Oe2rBJZibHjFgBM5kj8STuqGMdHi9/k9MjXKtD8b9KFBxONg+DSmKH+xupVwSdec
UszPa7pgSXafJ509W5G7eXRmEccPy/qbrBdYCwiZU61wVQFt8BAPO6tUOd6fS9Yr
2sb2+cRMHjVQUWAb8sjtasDzQILjvinzUCvpO3Sadbe5s9yjv+71ZMVaXIYydGNh
rDJSrlpCsSxaBfmoJfFAy3hc+RYEbNBPgRAihxyW1TBr1skuGUJRnQsuy5E9QInz
xqnEEWwXianNUjAOcPXszpR/y1e7wF146VBfLMHRaG78TCRrk0P1R5q4qcOsXof8
khWdNdtOHa5fOoXQpu4slFejsRlWrnrrycAZbLdvsGOflJQJzppEIkr555MTYWtS
cytVWuCr72GzMD50SNxg3gpKyWTw3iWNu0xw9RhDdsDSwqCgMKNkQR85dDcDgI1B
I032wWfts6mBSSNr7SZUdAjk6RfT8E3dvb0PpgHwA1Su7aOssDerNtpIgOMfCs8j
xaLsMUa5CADJuKibO5N9O+K6AJ/0sTJq/Y8YQkSTl199F1vDPkArAfxGuWuOZwIG
UqAqpmuZWXMhcyJhWpS9icKe+MfP6HE2UZqVmR7d1m3N2m6C5gQhBh0b+V0Emt4J
g7beVzRKEUwJV5iSFBsUGAvpx08GjOLJTJmYFBGlkQQjet62xuC24VGXawFuZgA9
9wRYCvJa+e0Rn70FmoEWVEqdgo+hkxHg2IkVMrFadWn8FvscRGmKTQMJcFT2lnki
65MWHEsSOav2tD9kUrLty5dbzUWT476KWzHgKnGXVeJaH/W9djWi97j2PKWTnUxK
jB9d8+Uxo1Rwxz9QfMLJCVCA8OL6uKkzNFsjgSkhQfh7gUKyK7wqAUvWcDBihFZA
DUgKBsb6LOqVk7CABakvA9cTAjgsoed+rV+ro4Q70/ZWnG6X9T/99KpYsX+un9lw
hNIHLoAlxTqwLCYaf7wS0VUmtZWo8TzppuTJN4B7PGa5aMNRE+8wzvvzcYbrJH0v
RTGJ5xT+K9fkB02mpM17cx/t5hNWyPfOvPGTdLYVdvNegoA797Di6Ql5V2trOkUO
e9O2DpnJ2jHZc0BtQ4Dutyy5BTg/N2N8cSaeLc4qOKd+VUA8VIAa3pa+OK3Cx9iD
+Bz8SAkDuxGF82k2ygHsH1GGSc5cLtPdUWgOYbPeyAPYVDoFDMfi4UzbwOMgdGxo
zcMz489ow2gO/8blKRQi51m33o0XrdswjshpSMvdXoy1kEbehfhpxxQOzKlN0ZvO
YY8UZP3gmkcsH0H+Q1FPxTIpx/BPiXuQP4OEZjPmPABbp8y1KQEiBv9a/vh/LWwD
BmY9AF9bnCLIwrvaLCIvJ+AOpuIoEoxIJYfn/1lmtoj6njVHAafunzZ0WAK0AwKb
ieM33lKVP1i0DxCxtE+ROC5stvnQ3EXhtboF/ckycdEAw7siR2LwoYUdk/bOmID3
OT3LV15jHkt6Z0EaOfef8dfUK9UxuXMH2qsUnuraXjJRi4piFo7MRAc5Ux60xdC8
Z9nLlp0joyix8Mg9MFGEAXhDK4z9eiI4YHzurvOryHqgq6e65Dfi8qQcRHREWPrk
mmNlYouYtgRBlk41BAAYq5D958Bzdgk4FUe24S6siy7XJK3iaJd9sx/e3Np4g1Ni
I6d1mIRjdPmLIdzvjhlYql7YgOt1W29TmXmNZ/Hqndztdfj4paHxv/2PEkF7sYrI
yfQh9yoz8pEflPtszGvazUgkdLP4SN44r92/Uc+kpyYjigt2/+Z5HSjXn53UfYXB
x+M0gZlaWgq/bhLHMMqAArDEThrvhzwl6poYjQ2qlS3cj9qHdMXcn7YM2roMzdw8
4b00PqBZtQyHwzzEJKcJS4XwYR6xF8c4YxnnwHUBnsJeFubTni3inGm8GHyVvchq
aJQ4kbrKy6wxKKNv9qVTpkCaZB1zy/lFsr9zlpTAGxU3Fhl6b5fknZ8FXLAR5Pk3
L9HtfRWXPRe0Im4whRhhi6U1SaWmKHWys2IVjEetKm53fI3kIqA7Sp5OEhu9D0Q1
37FbcH7zJymcBfmpc/7xm8QrMwwyntw6df8NmK8L/iLYm2gVOwr+Nqzoq2Nlv3Zf
X/JW/f9aAC88UXfuHQ9Sop42RwDUNKczQC+Z75v8kNiQi/AEJkjOBoDGmwF/sCHU
35rMIXGmrhBrHmPr7BGMkC0dgrngtgXf7jC32gMHpAU8fRke3/lvmnLs+0t23Qt5
m9tmuFwFMIcap13F49hE/OpHaByVs27IqJO0iY4INGDLNtTHSjsl9QaLnY3dMCBL
ZQIWaKVQCI7zrmyv0Gw5tefnJMCEU7pv+lADw6b4UTEqirn8cb1DjNWQrzrDl/aL
XPelji7Ll5ln1t6ArRU7a8FGsl9oYqcMakYd3/is1itUDjYmf56cJzGzby978s+8
sv3FVkGKIFcPPM8vPsDb5H9W2yfEVRuCEmV0FxE0XeOyP5CxvE7HGuocbNCW4m8E
+XmlSpWFl3HZZfALdw/gnLchI3XfMg5n6lLOI0Xffv0E3KE6GZUFzTk/+sPc6XrV
c/CT14bSl1zZpXvInMUDz88QMjGb9dL7hkJT9NqTkXPZ7dUJx1OqAJRrgEUalbBW
eik+ccL3u0SdLAfDWAUBDjUQdrJ6p2oSzYutOZr/fQVGeEEYTcUu5eKnI5R3y9B7
t7N4sdIseztyzRz2/LreClPB1h+2G7l2+QC6DuiJcS7Dpcv1D2w0i4Bp0VtW2vFz
8GJIYroBpB8REs605xNGW5/PzcExJn8zLjXRx5DZHX5XhIFlPpk93WuupIStMKCK
xQRa0+miHyi6YfNINNN6q8JtuCY7kVHZJcOrlgPH2lFWcmpvTDw390C0nYSeqzn+
bjFBD2Y4cPhidj+rNcpowHIl6VPcoAUkL9xQ34nXtUrfq4UFMvd80c/qqR6QbVI2
/EKAnfuUTPCr9bunL5e6PHEaGGGciGMmqxpTDpx0c3N3FRfX6yBmzT/aHaNuo6y7
k+Ucs4ELrNcZ4xyLCnFd0bn5w4otSD3HxR6gue3VMY0hjZJ0OE9XMTn/kE3qpswC
3NPUaoSEnwSi/jmp2q0q12xz9+nETyhqup5MM+9SkAzCHdr8eiEyYyf+00rFLRaD
FvlJsmN0Qn/JmRvshhqQ8nYQDbOYIHnrmYgO8lMpsPWZ1ulunoublAke+GYYjdbr
vA9Vhq1v3V3F71ch9Sp8qnUIxzZk7rOMKs49FIykjvpKlQ0zON1G1pZDAvG4R9DV
/pSZ8u9XBd1l+7TMtMORX3BmnrFqD6zPlZrNvnL4JACYZ1IxqxTwippL+P90YqYm
7KrRQJfbbXYp7ISPuHRCbKANsJbPsQN0evyVjg3nsyNK1lA9keYJK41QhzFWK8Aa
4RtRHnpU4qQyZOQMoUmTAIqlw62ioiG35vSOqTBD/NxCfU+PxtKpQHwe+hgJ+fpx
RV9W25yC3PtqSX/AMbSXqb6Sr//zfku1TBGFXO+VEo1F1DE0mWQ/Q9qhIUYYfOfI
lvDtbnI/Rnhb2AHPceiJec+ugj1OEJxOuIlDS0kyv6D99iqlYWXwrxDuHmFeX03K
xvJJTY0AXEwMEbPU2ngTu7C3b5LpD8Ty6D7vgxlguDXsnopFhkF/HyzQgBmdV5b2
Z2QOsACreVuFtLuEI6iGZJQ8u4Qw0OdEOhA0RQ3b8krmWZ0Ldc5CWOsBaWZ5a/Jq
XIVH45I1fjnPKbp9SPMJM6hxxyjfVwoLcpdnRufnBosMNOPmx9NVDWnWogAprLbq
5GCoKd8oO2T81qucY4r+T5wrUUgJPSK81T12SeeYQ0InnoDegM3XvT+y8RR783lF
xxJ7771ITTgJUZ9txZyqWhS5gFUvbdh47uiBLgwZkIEpXL/c23RaYqnoxhJyl+Q2
BCE/WiGfROdBsv6a8hp3n9zfiSYeBeJyJBEF3biYK4FBVP+rgYiCDmj9osAnRe0G
3c0FM0ZSTfqdjJTPS5nW8QqUUCZEDEg3fGVEKEfO0DKfzoDHbpcl9qd0CXkeSSpc
NpzzFcZ5AEU0zF4USM4mVCOMpaGz3Hxfs4eMvRUu1Jq2c4tDPP3U4ofHSX5vO02l
YcSId7gVE3hgI1sQRxvFeG40Dr6SIwWxPvHSnJbPD9mZE3CQD7NPOTXzqCLZ/RuR
VunzYSD+HQnLEGo+T6jub660z2OWjAZGvrv/LdUx8g1m5enU1SOUgJAjUl5U2iN8
SyU3D9XErelCqSdsEccH/DLoSTR8I2kGvv3Zo5QytW/kjuf6DTK4RCPc9z+NquTZ
b0YioddQSd5cSN5hGythGZGaIGMZBzgUk8x7VrpFUjb3rWOFw1OuxMWcqI69EGTl
quYlXlaL4gSwUaGUjmDE1hZNvmoKYoPs/fyVx2ndrlBP+QL4U7+1mGQWERG0ZTAm
CsLheXJW8IxQx7NI8prnGTVD+nizOb/Bx1KVyB+ZRK1VPraQEbaWSx1wK2jXpj94
gR+9cSYQc5Zan/iis+T+gst8CAJDtuqChdg3AQZdLhJpmp3R6SoT1+gIP7rSAZ2O
ZJZ4YfdpeshOmX0dY7GrZsZXRLNfQtLOpXL5t8OfDkmtQwUtcH+6EtbZWxdXMobt
BFmQllK1BaYU/trBhA5Uxsmw+U6gw1qsyw2wFZXTvWTKa0sPxG1SVrO5wq4lr7Qg
746GAw63fD7udKp+9zK77sAXebkiEjQnYprKyidoxoxOlyUzAJf+DMXiJx0QxGDY
64pcZXoGi7KN1SK1HaVwS6/H0H0XSIFJPW8DcLQpFeIpqq4NW7bDt4XPgHEV4vtO
VQQRNfE/hsiQzKk05bwMqUhSIaA7qpaAfSx+tYosh+181YGDlEqhOooTVbteAQGP
drxWLqh1bT+SkhSXpDXOfyyu7EJfCUWuhnEh+nKQ8sim3/nLXrvHEbrddwC8A5Di
/IVIVGnBKEFeH3L4+L5TuBSuo8Fxo5QTpcYKuAm4t0EHI+v5HwtfD0UHI6i+Qm+B
NqVnxZVS3oHFPOl8lUHJkAP1n7uvmdscCZwNua7lz7iFE7FMFWSsQs/RYogzuaZe
X+lSWBbjxsYcEx24k4/0EPvM5KnNwmjrjQD7iIAQL1dcxFR4XhydVNz4ylE2IRBJ
GUdBBmdM5gTkIWWpvVodPHBSr7PptSDhOk7AoT206xEmC3SQVBHBYZoGf1tCPAom
tt99c+Qojy9yL6+dWWgvBgQkP0gfJv+tX3dWCT82jJ8CM5hznfrzE5smt5q5LFoA
tGEHKa83BYo0WQpeHwX6/3FjvrCx9CJCFvRXKtImkRq6CoPs1rWiv2+nqIqcoTQD
eJld3sUg6gvPHYGH50Cv4hTmoZI+YQr2jMo0ESO0YJsxLzZU5Qm/mPtv4Sd/iXZr
JBz/jDKfA7nrKoAUyzFElz5O4FyxWVVD1gfj4ITx7BBfTs1+nL1u6k0gzBBfB0Q1
GWCwbN7q99uBUf+dRCRwG2voOOzZbVkAILasZKDUAQypspgSgfL6YZawUt3mfZTg
dddIHV9Wx1NgZ3uVLyktXdq/gKlxdRhhOCjNWikka+ej/IVEnY0M+yHETdsdv03S
13ENTPPvxCjgV2u+AKRMMa77YdXmHouwjriRP78zGnR83F0FKicWU30opwQF/534
rJ/Vh3GDwkH++EopayWOADQimNSx4vMd2Y99xuzBlUOVpIpsHAyGrHGF4PrJTZ4/
PqhI4e2X6eCtbSzbzGbwPQHWRUG8Ysulpxw1CJ8M+upB1uUf4uYuO3LCDNaSk/8b
fwKWUn61vx5dipHa5zNIRdBeNMB0+GmSo05Lto8YVcnzsgHfiYepn4IT6dsbbDYi
wr6rJgZuaUYwC9cw7cEoi2FJwSam4QtQFrDy0NfuZj615Nvg3j6494r1zBEFVjRt
vPniGPU9+8LNDrpQwcj0Fgy6lREwtsQKN4sRPoLwwFH7falWiwrGuA3V2X8wVSRp
uua54WAdCIblctrvtK6wMQsqNGKbejyWHUtEHjsPkGL7x6LAr/4o2pCQCU71wk7m
4UrvS6ryNhmLPJOjOR3zYbgNwormTXhsWbSPD/mDsC8zyk30BmHBzM8HIoKcB+dW
UChpXe+4hCBNui2emsS3KntE+QTMfNAGV/muiH67M8aIELvxVQ8qI/LAfYB8stsW
EmnmVuupbGsWUkQUVGt/nKQHkl6r6qt71NQ+DnGHiEJx8HvOLQ+7rfNOg+uzsd7k
e4pQWCv/YVRQo0hxyzvSuGSVNxfJewvMrZJnFqkmGF/QmyjW+C9MPAQsY2hjjlb1
6ACTXpEid0mMWFjQdlXO1j6XgrxEQpqgarJaQufbVeSj0+H2dbD/c54UySEBIWIo
llvrPEIPf7BpDE6p5mD02857zdvcs71JweFuLoljqrzVaohhy8SWwb3Wt41wHNW/
4a9Sxbxg/Mzr4M/+NVOkKXDBRPsB6Q3euHFzPKzvUuwtH2oK5O0QkSvvE2/Z1iX9
ox6VDsvQpd2ZbHNxBlueojAk3pzoTufMshnz+udUB9kS+yewjrdx5npTEJOXSJvy
yotQPEUziLa/IvtC3oPkCaL+nCD8vS3M9TPzjsM/Y6ypIjbPM69objG80IwOrESS
M600S6nYuGVH7EK0mrjwWUYqa3W4DzO1QzK1nrj2MTfB8gGipiF9C1roN2IQLOBk
kuQIr3ug/aVTuqGYvx7Znd1TV/vBwGd4C2/6ativw78AkJh7AkjoiNfn7DwEe5r0
2dod5q+rGyMUt/0u3kBrbyXVtSi5jz/k/s0BUUPhDb0j2rvrfR35P+8ifWzyGSrv
5bBfqWzJDHcBV5D8C+KGSmOUnYvktMZv03kWf3PxRMpayWsIK79jijBiN5p9t5yX
Y1ro/mR2T5E0DAZ/XaGJoq/NJY+Y0ywN1rLGR4O18YWvJfAHetlULE+YflO39Mio
WNLxTXz64TSod+8O0qeTbUeMmV3xSxEN5Hlnbdp1wVDWwA3aKm+3DWMWnpVwctmn
xOipQKRLs1kxmx+rLxCwbEyElGvJQyoWBdafMl8X0qsVhEhG+c13tTCW7IURStty
Py4KncPs5qut0WFJhY1Y6Muka4FIBP9giPw0/dUVXYAPb3V6v6qg4+A/m2Ii7zVY
IAJaro2JvupWev9OR7ddWNXcVgCNBtxumBJXyQm/EQMY64LoqcBDRJ9J8jbv7sGE
j6MVjeazPR35NcAzBb6srSSv7XNLSgl6xz7YxFE7D02tQanpWrFL/UTC97qr+ruh
y+3/gKQ7I8UL9dq1SOLoID4iEcvHJjl12UPl1f9TiI4mfisCkxjA5fJ6f6xhwgEE
0C03LM/QjVBDisiTvFp2Z64Kjt5fcRHVrQ663Y/JmUZXYYLbl+tBYQPPi9LLLX5B
m5AzrUpgVXr7MNrt0aVU4OZ88xwrNmD7/9HapMXwKDUQO48FGGfZacnHaB+xUACU
7YBqtFTjSoznVjvRuhOLw0VMc5r2OcsII3WwkO7y65kOE3IlJJdb2cLr7elgI4/Q
dsOv5S/frOZVy1VlHieU69AV1HZG/nGVwKthJ35lG+NTkgr06Jnwmq+m5nNFzq6J
x0jJy7msrzudk0352zQpFNYnUqefSw6jFFflMsYU6CNQ5v0QOcSQz6snYrc4EXnl
FPrcHZHLD+9+X8b/qPCYoRkdFWWsQWeesBYcV6YTAJqIWBpygfmLu6nabphqMjgm
Ur0ku7q7AMxXGzDztvUorqWcW9QxQj+iVCOka6MQJzG0cwQmnEzn1y37T86oKavu
ncWXSbDZPq9KE/SXGPEnW6F6p7ulSPnDh4GJXw/xWYigqE34j9BdQi28I/+dIQpl
jBi1StKHK8JtNik9gBtZqqfyazfyZGN8Vi1+DUTXHkzt17UAK+swAKierAkHGBFU
BuGb/lYm98lL/kMdBe9rnkuPzZ1zxYCiB0Z9QITBkZJKI0mrTAAmeoaU+Uv5xXg6
scDTllpNHZZwj0dy+aLdxGP41R6VOjmjEfWLAku+2L8KobG+nGIzIozrnVId3tNK
KZbVUQD51vjshrZ9DwK/rtOyks75FnLcBbKmkaNb5tCIgaNLAK4wG4iRQ55QvhEE
aHkIuitwSAr67Bgj2su2EZEQsjPEL6NOlg9nScbZdPbyO9LBGjhQvEFmMyR2DyY7
rFkyMlMJekBf/T54JitXqMvsL70ypd6TpMQur2pRT7E5+VtEf81EpUjR6ALdkxHh
G8iQIO4GjGlrSsU15Aiggq4o/t9Bq2dN4Puk36K4fQMCIu7tYXYtZdvYUxSeehPq
2JNxsMf39B92Gy8sjVB5Ui3dPbMxvrEbrfGQ4IGYUu9iPkV7TSyKn9Mwxyc8sq4j
ey1o3VciRZhyYLWU67AlLVtwM7y9+0S+FWYsMUNrjcS9kiBPqwot1Stm1PuXCpW5
B1cNrqh9Clnc6zJG2lAldC6Tluptb7smp4ARSc7J8lQdEugiiuTZW52t5jdZLFjL
vZUtR8aASpil4rnbNIc5+b1sC9zosoZONA8NuULyePL3gAUkRhKu3/hMYu4728lS
aF4FZV8g/PviT8wQ4vUp93CJBlvXoNoejZB3uS3XoVcnp8LVcdzE038Cdsc6p6oZ
TLeAMC9A/KiQLLgrCs17oI+jso8WFcbtCLCWOFRiMuO0lq4zi93ayig3NZfHTCjb
40GQWQTuWbBOQPRhkyIl6Kcq6T7Js2Wd31BPt4pDzbbKSY8ty6ocpQ5PSW35iRhm
q7/wZyoF3UFfw6x/5zh2O1s+xNhxOUtLT5EaBP6EGktcm8+kTb2kZxh57XEQNd3f
JeTxl3PFJ9zxWV48ER8k7H4JSBhFqVAPnue4tvPdrnkj/RMsABopBzgvkWKDjb5O
X9lgSQfdHJPcBrNAmLxFjTgVXfo8BK/ff3dgvogG6quJRKx9Vt2BSibrc+KOXLe2
vVgDrwzoix7AOQVFfX76htvC42IqPDrfoUu2OTnIgHjw8WKwelAfHiPh28Miry5P
/a/9mZhdlKawSQXS5qN0C36hTrMyo6UFJedSbgDnxTIlJ2Z1H1WvcNFjjtiDpVS7
7blZS+tuCWnUITjn0gdMZfP2O0Ofe+LI8LTci89k+JW7Roa9qiaMgpjgOn+HuFAu
oCZDstzELD1i4KIH3EPPlBuh6Yuvju92NdZDuQF+BuMB2AGfyPXcnsR0RmlxgNqJ
aSjzyhhznzV1wqDaK4oNsuVrCw5NIUfJDmxaYCvphUNxfXHtcBrq3a4Gc2wku9b3
9ImzUDPGTbpms4q5ftspV5RZ+xzuub2VdWcIu2bwyq5oDoJX6n+sjLJYq6V0jKSf
JkSfRDLyeqri5cHD6LntXt2pwku888KpPGMVsCxwyYGVPPr2hEj7tgAXebp4AGGk
UG+7aXVfVZW1233cxE53P2e6AfcaBhHyUBHTU3CEJykPlCc9RXHlXPrpL7wPDZMi
T/4ofkVd03zhkJJR3K3SnlYWsS3vHYHvM74dSUHHqdF0CaQ4H6P3+VQ2jCfNxufX
GJeP75s8NMZH/fQSVX6e6v4lqg+wWqWCxLI3AwE/gIlBnsRGYuUH/XWufY9jeQI7
l/HI+goldHL8b/BVVYOKMcI567m5GLX7rVWJyCbta1OkrWnAgLUZfT5swrxLxmni
EsbceaMBFpNW2n4XwtBbB1AAeu1JpjgNLCwWkCiKfNdeK2DZ5D1a4dL/99inGg3i
IcuKOqPt2QsifEmASoSFwCOnDSjhnQQSaifBwSVfbYPVP3b/1CmLcpb8ah5s9p+C
JfXreAIq5V/4ao34uKj4EVlOw69+EWwydj2JHNNcjhEjS6kBTf4GkydG1sRrlb3D
jWYlvHuSzQzXqG0ATDlCpUmvgGXm+RDa15w46nKnr5EOgz1hnUQC05j7oGILG3vG
eqbysK/YuUryvolvLeF76XSz6PIQdCMN4LuqR4ZHsuZEsJ6pph/sAABBh/W75+9g
HOiyIeD2KuyftdWIgQAIJiHHtfqsj1G5V3s4doXEl0/kIIRQ3iiAsUYDWvmuDGqA
cw7sN5y441a66ihIlVg41dtffkXWENebI9qJUThrc9wYW8vj625YCdsEwSW4oRps
inJLebsmk32/1XOgAjzwT/Eq/Tbnko35DDfsplz/7LMd2x9MmJf0JkN79GuvAOBd
AVr8UyOwcf+FQrVvu3aEYcp1HOaMKrEf29vK8t4XIe6feMiBgKLmTOfM2eizSv6n
KGnPsvYgGgZPppr33a5Ab36iSd30lw82KP6kaNDjGjlVXeAcvbFWsGz0LbOVEt7s
bsSwXfBVI6WBAne4V4jPR41H17QbUlLoieHC5gteDoQUkuXpT8tj/gpx2ORbseQT
bH8p9+bjtLNFEFvDfp1/9r3lTDf3g7gJoMAJ8im6QAapG743c/jnTxBEijPbyC3h
2GeSxnHWSvtidHOiw9W6Roo/5HKBPKdHGhpJmc6M2NC57eIof0OdkFU8H6gOYLnK
boi7IjRIYiB+oAl1eaCt16uLLKi6q1PrQpe6xnw/uJVNK8WLSp+1m9mS+YTCg0ci
iHNsNbsOeZB70UdY5s6ypyLkI0GuGiWN8xd7XF4DfiDHC6V6EZB/tKv40Sh8vk+l
joNDu5ONZPYE6ByagTrFBZD4+ULPJ/GeY9ODi3K43sP2MWCXzQIWDhm7a3ieZZzc
4ZOgwtx0/l0d7vrt4+t8XoADnMTAmx5c0FSgcjU1it9IxE2TUjBB4stSelGQtRbo
XIqzTcjiqV3ralTgUS2Qf9se1qf8s1kR9rTQKe7LBEopZkwQfRMUGIJs4xB0EY74
z7frsBO/reUfZszxeg6NIcp5LBUQeMOJkOba05O6J83LAB2G3n3dNZwS/cdxHnBJ
4hVMW3YLUwje6b4e0tKuKe3OS82dOYkk5dOrFPsWWhK2bMvkgBn9HCKBOJ8L3y02
GovIJ6EmXEeMtonx8qzJ2z8ql3RBWfds4WlfmlbTA9bUPJwDOXZU3CPbKlLVn1Mo
k06VGC6HNqm8sNJpik9Jn8n8dY/XoVVq+Z1Q8aDZzzRaYFECJvJAh8z2E/4KKTzq
4X2mvb4X/yCGbxh+VFKTVeVfsoNGAW+KtdCnxheenhKzr8OCPp0GGjpRkyuG/FT0
orgWZnbb6QYhKM7ybcymRcqaGtVdyh1njkVIsCVENmhcYgEN/qNTpCLiLA4gpy14
IbqQ/z3/+xyGwYEsIdtHgFcbytdGnf+ry49A99vuW2o1V2NL6692rru9JtvI1cBx
2nuofq5Pb0oPROMgchDIf9N2QT1rVPz85j+d46uaCjVqGMGinmis0v3pDm8O+FT9
af8zaq13epvO5TSbq5HZ7nzli7ef6BJbeiMtAoe2ge3OqAaAAKzd+Sm2yk80toP2
MKqmKUQS6hvocBm8ctW/0fDDFWlRPsKHEhbI+G5jsJCP4P5cqHLvJzVBf97OR82Y
neNdbHtuAP7OI3ppEuMrN4SaHX52/Rr/9QDAwcl3JQM47g3Sl3VR3jG8GNRY5lqF
LtzV72plKO+/mkSjZ1qU/ubJXu6Tltbh/vuj8RxNaZqGVH/WeDN7fKCwINfUrie0
FfKU2uhdK7ShVCTg5vttfIjoPe+8XOsT5wm1UtMkPqxp3BtE2BYrlj1ArbUaULvn
/MkpYRwYPdXOt2NRJlb6gvO086HDMb+yUlD9FEOy/i0YdfdxtpjF5zM98i93KSMG
upRrHOsFk4vJpsI+Axdl7pNS5tqS/TLw7/QS59/d7qOzxcP4SV69t2DaFoTU9xv8
G1Jg9sjU8xB4tNERsAQUxCE0b2bqZgmxtzKmDLKlerk+yyo5z/ABzYZtDnZdjvbk
2tsM/EQL7x/cZTmAnaqENIIxNUgXGCFeTEYztJIfBfBd+e4W1ZpslSQr6FLgfXZd
QxyiAOXb9s9d0lqiYGuSdnjx6A/YgURuwjmWCqK5YYSZD3F+R57UMqA5hL8vkH04
+SN3sq8B31Od8vkNb2QbYVxWKUFDQXv3F+6TPz+s5lRJ9nLoHtlN1/S95eF38wHC
6TJfXi1Eyh2c+XdvnaaraT4TzeD8k+Og0eUv3zUkoYo9qsStSaWozJSjXWxWB0Eb
CcQp3a+464r8PJfdrPTwPeNnxnP+BR0057TAgSry1Nlz7BAVxozcSZuBuZeAhXdN
fkLSEN10FdmU0zo7eL8BwE43toTcgp1LAsqnwwPoD+OT0mv1vZ5KuNuLGVf6JI4J
imwlAFnR7yB9BM351kYCQzN8SOGlYCz5n/Mr0Wqn0zBJ8MBBPQ0dbwk+zL8OpmaW
WAxsFqVkXcApSuF5qHJ4msFKXq4y0JjyqeZ7O1FL+VT0JcpTiJ4yYtrsP1KSXtv6
mF5HD9fgEtVBfkU6EZ8FokFktzn5dmQEuCVNc//yL/6sRScgCxFgc/nIgRTI5nCP
ebKZny9FEV7I4/zVzDRaGnsnQzI6JDoZzn9+9Cdp+AB8lbctCOjQbRCcCQjIw6GF
N0mwbuFn6YeFpSswwysGh8cwqVsSen42HVO7Ub6msQq3Tb8EoX4hjsO1TRzgm57B
pUghZpv5OkEfR0eBQis+YlAI2D8y3tDT8Eq/ezpzmjEJR00xYS+Pla/K6K2DTl65
v4NcgSZkWkvQl/SyreVPAnmPjTpQBlZVb/HJgQafW1yKbgZv121DqZrXjcf+w4Qc
yFKcx2zXWRWSNTXkejbUW7D7ArYxhZq1t9RtMcyxl8+RzW8fxeutTOzNGVlh52cF
IJxv+IRW76wwPSsQ0xZzzJPrjvsveqxeQm06HOeD8xOVFiXDMS+oJaiHtDkJGM9p
2wOpnMGn1baT05PrrW/t4ZBhASRW8/1jWuDfLNpbY3Da27/p6l4Ua3npCZDqUQme
ZezGzhKGNIwluB+GLDAbOZejQCzVgQKyKHl44DB7+D8tEb5GtBg8E+OsHU7e83JQ
cYVSoikQNDKBg2NS2DIcfZAVUETbWEG8o8UWHmzrkOz/9CyZ3MrhaUfNiGalVY/K
IpVVNolN4kVsBONrbZAORmZEvLf7th02JWsj5NXoo/wlELzORvEjaXVGu/9KIqFz
qch95F1Xi3aVf4VysOxppaC8Zy5K6SEh6xlvW5MFnhrmJGaSy4gug9pbv5BW99p/
mZXoxgRlxfeyXcA0NYu7J1bpT8VqW1yr/rIqYd7AZ4k0+IKSTq06VqAQexvPB8CN
Akg4eYSvcJlrft69jXAmY2j4ihRwI4+7ICWaDwnPOI8TduCOk98u3qDDmIZkkNQh
RHEZGyNg2olRRZ32U9xVPOcSfe4jX5nfIV/0QKm0r0v4s0SWv6YdzN31CK9khSex
sfua2nW/Wz9t775FDOQnkbzCzzmH/sZwAGh8c7iQ/PWrk6F2Z/vR5doI+tN6zB94
4xUqtPIvrLNPpDE8nqPH9s2HD8/Z4QrdkuJXPM8TxnprAowWr7x086dOcnc0rUzE
nz7+48QeInFIrOYcOx6KrFCob4+bsGvo/EQaggNeGhp38ELrXx5vaDdJOW/mycxa
OyEqmyF+lXGR1rYd8HSoW+K6k9bQyNrC/LUHTfZ4U9tYoXnE4H0/ijK8rdaeYkTW
HBTuZ6eC1n390gzNBSwsQg2JcXJEdajlwcAGopCqA5oIttuebaXPG0ipzNzGxxZD
oaMzKV9bhdh4nNQsK64IbrRDXrRBroVziv/7TselASd5hENHc+7K4RNO+E/GDk39
a1d072M/cnjcCFG/wP7zQKaYO7mfl861foZ4rZcmWA9HETpqaOIS4eXGijVYejGS
Ki+ehzkQdv9kJmY1an9kCQcwWVjt2N+AAUv8neHDPgMvCCS2D/GnL5/nL+1wPwxZ
CmASEgxvsoNFAZzXms0jWbVb8IvN726ilCaTbe56FW6O1JK7f7D4QV+44y/V1rs3
R7OtzaWv2S0caLNSUKUMdmRybpm+mAQiWe/GDSLyzGES2A2+PAAHD0epcFqfJMl5
j0xa/zjCtSS9YyNqHSxfD1gCsWEHRsb7+R/7mw3/kwNyCcygYm6jW5/4N1HUnHUM
E4JwsAUadlz6yZ2sTKS8qUA8QUKejzFX9HwIHrKbdu+IloDf4b16OxvhHXjkk9yg
EZNWSwZC+m0BohqLUjJrm01iG/EljbgqGCTmhCqVNFu1BMPaa7z0zMLM/KU0Wst6
p924fWcbdZNJs2iZMcaebql9QXqMJvXvDxl1DYZr/U3Tkk935W7JrmvTs+mhPxnf
nPHrfCz9zxvoc72zqOQi/waRo/PQisOK0n7696yrtKRKhzrEG4nYzMGfh2b1k79S
z2AJohPEJ3GAuPy+iNq4JbLGf+UOZp/PfMpe1HkUeQarUPkxQwysP+LJ+qTa/xJG
wRck0ZTDlm9YYQqAoHD5loy0kWWmh0laGZN7bwJk/aTgPAPY3l4KBGmiKd2gp/Fd
Ls7OvU7y7jeSb2bapiiKVXHHQmizM1IhMsyrxbH7511urIcPrURXm7pCOrdKWua5
RGuFSNOOu+HrmFmBqMI41BdyrurTkFK1Z8NHXde2JpKFc0gb5tx9jMVFyffjcWr1
j6AlL3/Fb8OtuCmCWD/UJbSTkVmadeYmauPynkWE6svbC3udS+Vzh/D+Jx2PESWY
uN6SqOHlAHVkwJYiDsGFY6+augj9nxRPEB0BKtsZaFC2qQzdEy0tA0CBAF6q7J4R
DcOyIVTc5wWIAQUFUTHxbCzZ+g2ugr+nL40bz+U49tVFcqUbYjXmbraAh+breTX8
vXHZREFqKZmXDgSFDl7MHDFoUb5COCzPUo2hCA72V7vXvtYbSza9UVYDqqtxZTgN
3Czwn/J0R/Si1cnSINdxhTtMCwf2flAz5o+DEdnivLmd+2UqUNm9oMoTS18EtBOo
+DhPpSDEEFtrXffv1nkTgz+ntyRmpJNGBrlE7OBg5mbc0uIFN3wKpWIJdzHLsgm/
1wVcFLrYXlcLh14NpR90cHZcJCjLEiT8AKaTA3zNlr13WApjguizP8AVX/DlerIo
dJb9u/qwmDQSp3w+Fn51SZygTGkVTxt88b0gQTL8R7Yd0Q6DC67u8lDp5wIp6ZUe
hdd9cpaayWJ2E605YaMiL0O8fxJ3eew/rTtCbg68tgtJ2wXCHRdkMqg+K3jlYoFn
pjJFO8UhqTKDg7G2/fdLuy0JDilD90e8hapsbhhmMsUjUJVgOjoWyNYB4ffnGDD9
TPzDerg1Ko/Tz96eIZFqUqp4Uu1yGaevvfUuCa1AFVe8vgGsMAK8S2lKRrRBv5Lx
ddKGM+1Ffn3/38o+UJ0KNto4AD30Ycxmx2s24Jby8x0tjVmFmZnQCIsi6+iIvj1a
wrVekD+GNnWgcYRVpuRCDkG0AQNa2OZchjO+7iTsNi1aa2aCfQEFimPWqsLo15r0
f+K+TBZGyCHuQbA0mRt6ahe2xojXnvqW/rW9QBN0W00GZ3ihkJsa0ghk+oDSP444
HD3B8yN+YuL6rOiXo9KGQil74PnAPQUg2FkqYneT6bmPKVf4FhVqTzz5ucuIlPtP
X+BvIlQK90CLes/musHMfp7AJm4Fuy7GiqrjlRnOEkCgWY8YgEQsUkND9XF/minY
zHmv/FdGl62xnXsBktPSZAQqA0+gmv7e4M6b7uQ5pFQggdWJl0z/P52/dUv/5awz
tOEP20tnR9E2599Up0Wu83DRIJ0R6jN+vJQikPFglxP4JubbQGHtUQDr4d0Foe2G
MmxGJM+8PAm1K2BKKh0/+RXSKVH7o0RxL6ngmMgErk0FzCHgQDWgNRdBlCqoh5it
YzBcFOmmeMrHve8/aMTB5YFKd3U8iD/2rzf58zV9hcN7ZlckGYqsdESZEhCWZEy4
tdMfSTpbpkepdlxbeTdJyrlYnnEpIYX6vQk9mBdZW+RFM5ofZPxQRlcph4riAeR5
6FY2k2J+AmiMzQTU0LB2SLvGSW3LjhacJ7CxuWzSiYCx70yYfLwbo5DwcGcB1Kbs
qOV6unSAIDaY8C/SXeHvouR7cK+XFE0fRj7C008UFbL/xUVweYxWD6jvIijEVPJw
K09suT6CvvMxaCsWzaMIsIou3PHZNkOUhkTkUkx8B85sOsM6ICeb6sAvPE5yuVWU
V9D7FRpuyJoUbaQ3p/iXRJBGhiTwVSAB0JhekT+bTDFp6HmP/UNpCIS8UninU9as
pJ1i91j/CbJkxj5LJ6QkhTSTnfO103DUn9s7/nj36g9BgJGW/d1En//wVDLQc5FA
8FmSfQJxT8G0yvNoUOMyG5ftgszUr9kPG4VlT/yslYDpGFkPdGJXYZTDpFb5nriP
l0RKAyAGB41KAv9oKdkODMnxGU/GYAwE/ASzIh6m5VN7F+/utnLpqsMgBdiAtEoT
+Za333xZc3+/qsSoyauVhQVXEFfHa0uX8JkDSSd9DQ1FKIFW2SG5YYMphOk1irEU
0J8dTY28YMyvH6Q6HSdpXVDScyUC/2bpDuBkxuJoadH5Ly8Ri1vmk5Ni9Nm6aRIU
ueG2uRXNXiiTUSXw7tU7+b80TsRKgK9tuwD2M2B2gL+bRXLJASZhif3mxctoOXay
zohpMRVy8AgWiWV5lIWGlZgNAL17zOoLi7nRGUJOWIl3i1Znq0AAszes4QFWX5pP
MmxJILCSxdniCymdpQJsKfLCfR3NtNSqk4OqWgd1gi8uQtlelCE366ioHqlFiemh
RK18lfQlnXvl42fVsNqggxZ87+mPlr2ArkHIC4iysEOH+bkTogJ25ajMtj73nxh3
5rOlWsmzw+SizInjwsgD47U8Bs1NZa6HSQeNdQzDP2DHv7lJSdvvf8czAfoNhBwQ
brOQt4DcBGprT69nzqTWDynd0nfMAjmx5DSJaH1dq15j1YQRaTMz/pGuB95yD2S3
y0nDsP1KxakxvdUItv4RCp3zVkcelogRR8jCMBFfS/gG153KHbjmwGnrFv0OOPgA
FUw6Sf/ExjjGrHNn1xd0eBNnM3RgJC6BO2el3isZNdDfxtVUl2egfM36lbiis4vW
7WuKzTKVyjWd7ljvFzX/yn13AJuvsmRFNRKLrz+6EuQlG6PB+WqJ2xkOP/wvF39Q
orQki7MusFVTb1sjSEXEJqV5y74Rd6Z/dMA40hOXcpxIMXx0OtTe67dpxacs3E/h
8NE+2wP+j+SDjTu9MbrRWnEOADk/pLHkjsvm/cAiWHYKnzQXcKqNPEelaia0tvZ8
Eo8/1yHMYQCTDdJ27tlt+IwcBAJ6WUienyI/lJztDjQCZBgLwGZDYslZfXtorE4i
xIbviguOzT74rZVYLJodQG9kHbgesoH7H2oslrMCfnG5cF/U8K45yoIGOEzSwjPI
238hRbTMbTlVlT+8X3dmixMKnajwsLCLta/3p7G8CZeB+VdMf9hpyPia9AH2aoNm
ZYIn6J2uA2fPwN54akk1TWBi8zia6HOuyKALKRpwevhip/3t2QABr8gsPVBgw53K
GzFpd6qq+HIz+pMOSsRliEkX3SIB6A0M75GAFj1wP8gIujfi1HCxf5YZJf5aFwU/
SbSQRjZtnYH9h/naTUzcOesAp6k/oLja5/L6/ufMhSdEal42G+S7osbpFho06wob
GPCUfMoW1ffQDLBbfE2fwUNTQ7cpuRTK9K55lHwqWA4uzMz1awLHe08X+D7BvMgq
QDX/25joFFCK3ybuFMIm/TgIg6FRsdO5NEnACkyY3duVBjQVlpy71SRQC/T+Se8V
c8Cs3cMBA23pBN8w8HRu6hOydCVy9UTU9m+SuPibI9gDAReqAHD9YM2B6e//GiOG
06NsAatize5bB+vNMBcmtjGrshuxRjjR3h3CJ74hdWhqluyPCiYWA5xg5Zz/byMe
B9jrsGFxqhS+ETiOxAbWtGgfk0WL5D0xQGZq3+3LSOzgfKf2RW7sCHbswOPyOfN1
miGdPiwGX9sOMRnNv6BbDkwRHHOYsMtHthy99R4S6pFWwqjTlxqrKTZiVgq6Lsp1
Qt7PmdVIQvVmO3rZbhnDwZKVnjO5q/Z5irGpdcymB7QIgKb2QJlzsv2TlwKigYRK
KxHlfl7dKDUWRaqOUlhro6O0qTDifaKAdpC20dtNfJxvUyajywUGu4w+jnz3Fdsi
tITPhMgrmI/XjMOLwf3Wz3NpxMXYx2HZSK1zXb4kkfukPMOpzM5jzMhQW2cEh9ys
tp9xl3j4uFuK7cQF90jopVgL234XH4p44YrM3VgtQCFejxSPe3CxLd1pUfbXxDoq
SLBp2g3T0cODZ5IGclIrlIlwtdY9P/mvbt8Rbe7ea8ImccSQ+9X8x9nwzWSLhvJh
3KPZ+O/EiG/hsG0nGb/sr7eFxphcDgXzICccYzAeS1YtxGuK/ioho/Q0m7XtHVh/
ov0H8iNxjxisXulnFGIFKuPxvSARI5xYcP04VHKAZOQIXFgXSEHh2anJSUwddwrv
zETO2iW6iA1mKugZH75AU+v6sLco3RkEMObLDFydFPVKf80HmINtHcWeU4Gh5Ghy
ejuGcii+i7bGqkDy1QvYng+U0QGOGwejlUAOC7Cky709bAyxSRTnFN9pugnhoLhC
1AeFYxOTs25E2JRETL9vYufTZ1BI1fhpKBT05KczUYhmp/K8Bx8IlsSMDVd+LFgL
7LnuXRkpvpAUbzm/aDYpmNnxBVpYzJB0Tx7FszeUSdiulYbf/jknFjV7InPp9F4h
xsCdAd2N0FpMAT+rX4nCvDbhcAVBz0pwFfb0ArytX1nPMqLr8zBffi/6kRsDNs4W
vHAkSQdSjnLZc01lKVxqrbKkbf2wBxD4r40VQtXHkQYZziEQ7pYvq0SKZ652bsDa
QOPUYK+P136Y3rCv1NiS0iOL3nFLjtlU4T+a4nrAMnzn/L2ynWSy7Nquat12i1oT
3QSfJVgsyPl5mDzKbgjVn1Q8fp4JG006cWrWBnnXh64DZVLrWRcI5RaDeSqgUlFg
s+Vx7qYXxgy40LV8aAx94lEHQ42brbasoQOaKCmRrVVfojXtQ7Ob9vFrf+xEQY/c
2tmJbYR8v+nX2pmg18xavAVeiVvHVIWQSxwdOx+jw6mCz4Rp2mYI1wg65sRpRkMK
M4S02bdgp6s6ObjOBvZgapoiM4SXF9EZBFDBDjaP7rmF7jVs9K2+2pny7cXAwIWF
7cpX4a9p5kPnwFfItYyGbz9kXnDE1DP0834pVGwKN0hf/CmZyOAvyv4gEEfIweAu
fSDwv7i+ZEwpKVgd9Ho4z3tQ6BvuXBVdZvI9U7QO4CseA3dARBVTG1DuKGwOL8Cv
WPWm5XVgzEAjWzZtfW484dh+fE6/hY63xFc15UM/jA15V7/czIKrfcklnmdKbYzm
evMFQENxPT2+B3/4+oAOV0ucOT/TB+fxST337UTNFaUGFEiChB3mDDohhHTVvBX9
xy0yeBlWXHvfeEE/a3wCdy3t7j94469QCIJmgWHh+1lXYxY6ZuSuhW3CKkJpWeGu
O1EGA3x2+jioNi/1t4nQ3Dwl045EhOF6JDvACBR8sjIYXD2uzttT22H/Q+exoy8e
DaCnYv48rZ8MtQhpYxC3wiDY8jmLlaAx2jRM4bQAFQYL7XNZGkons7QjlHVCXSIq
BYnFz7XHek/g7Fe1Rw8Me0/ka9PsCUuzfhqJ7AEa4j9VPtJAojZG7XhzI+lhuSpo
3xglGUIzF5Tb2VrUodaQk9g8J5FeYNlQFeaGMpBUBLCbz4tXcPGrhdjeYdjOnvsx
vhIxwUvkDF4REm0K/DvbwgXJVHYkeDKuwOQyL8BbjoEXlbXYiDzfqlJ5H8T4E8aO
NZJgbnJqMwiU17rbrqBALaNRScfqKR81nAj7DHKeAfhU/TWb6hVYphsDPjRCGH8/
0d/rXu3DAEwk6clgNi5tBssmeejCSxOtZ88xP3L3bbsUzG8r5P+afa2ULUV3ug3B
6SA9H6A2rLcHRhJimsF+Wr6syCbIzNJguvW0QASTmr39Iaa7vQsuAlkZvU6Abud2
fcxr9TQmM2yK30ytyk+p8zrjar/0v6k+eFMKl4ETdnmODXc8C+RPU8a3SlbNHdTs
ifRTLNaPwAaETutB5DzH8QjY9Qlpj83aqqL60djOEOlilyc59VTRkisdNQvS7nJQ
p/lxwGj4X5Gi5FuQbwcEO9tZEfOPMF/u5oEyjiZbH7xn7+YYwWQaGJoJ+z7njn2j
HOGkavUipd0ycwLQHoTPbIKL59/ZCM5rTi80zBxB2pp9ADaWzK9EW1qgbkD/OuiP
1oGIGL9NpqkQhB2I+ubJurNTvK+D12uP5usAzGUHcnMqpMbzYJmgmAdi9OejclCq
LlleTO2rgfg+jtUUMAKuhKQC2Qt8eU4YCm0qdJq43rka2PWNPeAJa9clXQUl0TXR
wlhrmtL5kh1PtU2/H+Bp0XRdy1/8iBeSi7ubdKMqlcba2DIacW1U4HchJTZI2t0C
OsHm/0ANU456h1BHyRNxFTX9trxHiONLvVWYv/sH2OPpJKy2p3heR17wLZ8x1Ypr
ZGE0pSXZM+FZdi8fujRkw3mEOZykCXbwcVPfNn5OzEqkgnnqDhKwMJHBz/wNLdHq
v3n/a/yDYOigXzoD/3sVsEZmqMPP297MQoYc/WnS5o3tPrLjXscUpNpb0ZB0EOF/
815XQmMBquHft9UqdkKbs0cLmU4APHw/0l86vVOzYylQFNTOMCLUFljD2vG8iMdq
Nxx41TZ8ZUBeQoTnBlpSlUinoaR4LAGMb1ae7+CFCS0kYJMHKb5sIuWGSp/iE9gQ
Sc2VtHRbQhOMYRbbNvinq3kQBHScH8tVpMvawanE+B4CYwJAvziSh+0kbReWq5Eh
5RWXT6ZzbJIw/Uqh+TzbfuFsrivR1UYlXjuZc2KDtY5aIrxRElY6aemIiyGUsxQ1
2xNrokm2BcOxVdnPGESkKUCUrg60r9J/MSQ3G3TD4d9g9WfrgdUyxY2RWBIcadq8
eW0f3FzU6xI0nG52qusS5i3tXM+8XYZutTk9B7Sn7Ct9Ksd+H5+wH7z2FujVFUHa
VF3r0Hae7DrmUo+7KGdW26BJ6AJwO6igNXWO5wl+osWGWk76WIgNCxlpxst5Ftz+
OpZmWayU6Nyt3v0aZpVdgNStTTGHZ6Z6JAqGooREmczwrYoOswIIUV+Y+TA/I99F
b+GjgYrJm818oTz2DtI5aVm62H4u+QPMCNf6MqnYEwwVSdH5RwGJ5aIAId1IqPYS
PXHQzPW+Q41KfQEc4wpP02usTzu5k4XTPNE4d85bcW36iivk51CJFG0VCdc0lI+8
O1MmPLRcRXXhoUEni7cm80x3QoRhv+ycNlqLurX+F7/KOn3iWNIuYrxWxC6N9G9g
83eA6CtBzNwxVDPpATP0xg8Xhk8m46Aqi2uv/ArtJdOkLF6CCnXjjrACHa2vr/u4
mb8rxEA07xnMiswiupVkPe36r4PMlkt4UZYYLGpuAEe9cuFOIrt9q9Y0go7qFsa8
orqUrT+t+ZLLrGOacXGpQw0yIgvtxQbR0JSCJiFFbJo5yV5OUsyGvJSeScdled3M
FX6nxsIQmp/9fGk4ydVgbVK+xCwQylGtA1Ml2RGRHEruBj8WTaU+6OFqMQSMxyE4
1XXHnQZi/gKNiTbhKvZnFdz5meuSIZPEKKA9p1EZDOgnppd2BdAR4SmorAc7x0tl
Ve1B5nB0TFQ/xNtuVbyu8PRaIhE7jKBM4tCfCbgcpXoAfy8l3URl2yehztD0Q2rN
IIT220DRDJvvBzVdVfQBtawKbLRe5NA1RBl6kGE8LwioeLnvzxlcJorh7y5D4Ka5
3p1s8VejvGk5p8s+SDC+IkO9O3Pj+8Qy0SZN9M94VFgDyM8qR2eCusc/tvVphlST
nZIddtls6pZWXgdg/Vbql6CJfCfWUptv73FZHI7bXUsoiEF17ySlozPeHJCTuVLk
edxm1XjfX2q5m6jGKdVJHLu3FX+fUPdLt252r7AKVy9nxNM1e6msTeU5eB9XTw/R
wWkCUS6/YDsBvoltLv2SV8R/UYRpr5R61iTQjPqn1HXzKX+1Ysp2AUVpDSICiAQB
ovXdXscaW3QPfBVcxLcjeKaWTvG/ixL3co52mVrApeYMEK/s48agUsnAMYMN41Ro
sZgtEUSdcrk4r8oZIXFjNCgdlMx0z4QAfT625vqz8HiZxaeGZ4gfqPWJUYgzzFS7
Abr/bvJ2H80zqARiQju3tdMZ0FvKGHfKc/60fHKe9ZfgKYc7McNq5euTaSiiE+MG
bUNGFjXVZwVuBLZbBRSj9pmAMwtheuBF7aYoqQw9N6S0l9U+i1TvMbu5JstHoc28
i49T7WJ/rSm2qEevLxsoNb7/DpUfX9CfpGWmtDSKHAAs55oDkzPDZw1pfgqR6B+u
Zl5uJvuPfAEPs/irub6FFEIikFlydySoBvQn7oe+NRM6bpKrTVxZFuWcHrsxLxbv
+ohNkxbYF4lOMSanrq9tTM5+Bv6cM0t9DFjku9Bdxodn0OKzWux7H/ieEkuTQ0U5
B1GIxywLhFRnkISmD78GFYVUDT/gnYXMsOW5XNiu9HE90bkAi/Sd0vN7QrR7ksWJ
I1vjAlHE4BRcOdQftf2hPmBPEirlQkAYwD+RlUZDUdg0DTcqQAZ+9TrON3A+QztN
wAkX0OaZJwP6xNACVR+KLPly1/u/8A9JXFiHjuyZvOpd1GYeK3IAbiCCgzteCyN7
hHtibBu8dtnE27Ppe6A0qnDaFALoqhQeFnRDONiPNIVY2eFQWjMt0Hl8HYIpuaYc
eON/HIcR/TN6PycihpwsrLFUTriNnV5CU4ICYCZ79PLH+wiF9kyDMbbrJnz9fuM0
pRZwCjcZYmauDLjf6BVwX+2wyUBovG8dBbD3mXWFzCXuyYwO+N+ZBROkfjwu9lv4
fc0Xmf/ZQ03QHowD9myWa5lDFXHiMHtSL+S8m0PrXAFZ/sMw89O7lvKdC7kz0kzH
oluPQ+xx/hj9AIinKGej5BRb+fLzBiopD0SLZA/vMBayeksv6tGvOHvVPzEE4jJM
zy58s/0nMUODCHPfqzyFvpgQHgl6g3L4n5rcKFnNlJuzUAenAetT1F0CbcUr9DbE
ePv422LfLW0FVtbVMmMdoypPomjdOtk2VpdF4pv5n5IEmMHT9erL62foyHE5Bbld
l++6Byn/7b3RyrmhD7Gu1mxEFUdmtWwX7TeZvOl23Rm91ymlv7K2Wh5Sg3PwuXTz
MCy4LPRwpB6bD9ZvHV3gjiI7wSP3DOs8OSOYsqOqKMqLw174VowqKzf/XRfaYa0Q
gbckWsCWqgglxLhN3+gayxrMbmeDo7DfqNQz1CD3d+vQxGfJPmrCLDipsozE8H7s
dUjP5gGRORj3kkY4//TOBpOKiGtKwrw+Q8DtnhL13Ls/9y5F+Q89fECAVgPjvPI+
nS6sqQUtFYxEZ0Yq3B0XfEBqsv0rleq07mbF1SWYs4r48sHWb9UkKTfKNjgMpkCj
FRnR+ygKZ6uJt2VpZ2M0PnxXIS0yaDyhCooH05+clMxF2kahKUMXwXH/7kxFBWjE
zX5QuENvmaRBp/xu7nlOG1qY+Z4zsow2WDJA6yCo2cbVfdQe6a4soLzUfYoxQhfl
kq9tpyqOlBpOuXokhm6RGlyeAkc83ieJpuSfmlti9rnEih1yO1yiBbZKd0oUQiDW
XDYb0Or98VB8P9nU1odAhG5wn7mDNWCWf2D4pisgE+HGRxS2Yz4hFtMUX7oJ7U3t
UiuoyrfwZiOMDGOipiEW1jm97U9Df2NSSe3+TDFG4XnnE+a0NIXzgeFkeyFib5j1
fumgfadaMrKyWboTtdvxutriLfCTNqLF2oeAby2PWmCb7J+bqBpgopFN+F6icWwD
5Y5UirpvnJh1FNT9m9JFxB8aera9L1kttD13YBzU01NVDRt50dS9TckndbV9Apdo
v1dUf2zIw//nbEelCYrN4DUWuymnxts+9Uh7Z8eGBqbYDDNb/pl5hIlHktL0spjh
UG83bgztg7GNGuofFUv5b6f8mQ12E3QmDRAt9J6U24SNKteHjE+q6apSGm7csvpy
u5GfwyhN4OzdWYBC3Igz7A/gIlSVjXviXjI0mVn+CO9+KJyzk+y6qpE+CzHJh5Ti
1ByEDFk5X9u84eoRPgGkp7Cbek0MTJNgLkxyzgsJaKelnpw+ccySXH5e9qtzyxYR
mhgYy70XKFqatd/9r/xQXJqS3/6zXqYFmlVA11A8NHUobJZs+Oj3mvOUyAesLi9Y
FtspGVLGL5VCU+USfRjYcbNoxjH0uepCLnRcObaG7abETv7/yvxD1WU1XVxt8xWO
FqebBJG/oMImr3VLIvzKFlpl3Ly53QcBhWItrIYufh4eb5GmECDnCh2E0pADJKGC
FzuI+pX2zLIB1bLbtMprKa6Vj+5LT0uB6GDQLYMctSmtt3jShgaUyaJ5GLcHwiUs
+Ppt5k6ycCbQb3OuI2gqLENz7C6hlgNLMgFSzzazKacUo1XMo6Sxf0JCzs3mvy4A
MvBjNepx29Qj99zS55MXHzZxlbAvg/ovhwEFzEdMX57RaLom9MHtihMI0ZEa5Ah7
VJ/JEd+sHxzLAkdPzgR6TNkcxNjMIR++0l0xHcmmQAMg1kHOKT2OHOd6vzjti+sg
a7l1JGnTcN15+kuavXPacIRO9alfo2YvbV/rafcdgZA289rjA3a5NftpYQJ/NOK6
`protect END_PROTECTED
