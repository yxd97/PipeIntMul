`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sKUIJucW0jY/2TePyfR5ToYn6mtQA9s2WBvmv9XjT+W47s6roAZ8rTlXj2VA9QDi
oivss19vIgDMlxARKYRijN48TqjcLN0v+LN/Gjdl80aII1qnKjCVKkPKh25rXx/+
KlxbaDVVhDnF3MD5ntbNHAL+MA75efahi6QxMovhqodwOk4a6x3VhdPPZaD8Avia
BacZbqtkDhWa/gOtmnpTJ8OwMEG76GkwBtdGSLKmFJt94qb8XIcTJZFpRVI7+kPG
t/R4R0wwOpIsOb2/YQ7i3pSejbi78a0JPWg3mP5Tt3/6lBGyUUCfyWbuzHujggOn
ZR/gwvXVv6+lpghwcdzdWw==
`protect END_PROTECTED
