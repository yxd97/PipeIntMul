`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gY9Pcad1UhZi4jGTpHfTo1EoPAq9BtkIWCqWNMzqxDM5MEpDAu/AWaJdd11nv9Vx
5dCvQ7YTm+aBWbBd9gKOT9ln2a2MqpijfBoH+OkfWbPiglRlc/aVDQH6tmTsM8Vo
9rNrfBprMVjgtGywcMI4zCMwmfBjGADPlOlDDPuvgh40YFCTbG6EfpcjOIlHcfnO
ovrO8F2d3FTlvcRfTTUbmP2dsfI05nQEuY73Mxr6sBUpKpQ/k0GosPGFnwD6lOP3
KiskaWOQaHVZNB2PWG4sdI/Iw/TId4SNV6XFvNc978By0ba1DlKJEvio6QXPPias
FuzKucl8QBLjDY+Kx5XewpxebtdCYkYtZwbHZrXE+eIYXcUjKYkARrQja1ASWPWV
VKZFkrRn5FQkeh4GqnV2K80RKB9mHzGS8yfTNSqOAvOsLagV8gksPOoz/TwZOLa7
0oD7uxns4CJkUYw7I2r2Ag==
`protect END_PROTECTED
