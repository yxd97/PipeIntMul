`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jUg9Q7GBEiIpFr3LvxoX3uj7jo3xttg8gGE0SFWZ8Rz1yICuV29lUk8nTK1BA62t
BxyOmavfHAomWiLjijWO4kcm2z/721P8OPliiooL30/OX1m24ey/sN+lM2Be6ePE
b17kyWq3m1lGM5YrI9wG6xDxhEvKIDaRf/nYni9+SL0rpZKCzVuhIOwaa1/0eNTs
VFa/vpfUB9XACQOphwiwr2bKTXjO2830LSMIlXAw17aYPetdR9JCMYue1iHs6oBv
8VTC2Rtg2XcsccNKHxxbsq4Agxsbkxs+CsRfLBy0Vgo=
`protect END_PROTECTED
