`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTDJ8fNnZCtZc3fRYnRJTrlvkS7EbDD9OPR/9nmAwqFN1TluidxH0CLvBT4jzrrB
bWipvzxsL0EpDSNHxA3QpshY4kPhlKZZSbm5pJQFr7iDHP51sj/XkDi+zXyUJiIG
XJOFbYOao9lj9G6bL5UUp6SHg29NrRAn0brqjqn0phykwOW1Jr2OJ+6Ju/QQLHj2
nIiOHFnLmJqtb2aRnd4Gi8cjENsBj+6373gGfVIgdaUP/nQAUtbwcc9Rbpw71bm9
3xN25FRxuJn8RLsmhETRCLK3xMza7FPs4zwBxt3AYdhiAK6YQZ5f3+XrjsAz7xQo
tFVwStMBIXHDFxsumFgBZ+PHS5PvzOAXruovkpx3robVfGJyp2t8NJyhO0Hfcnjf
/BhrLMNaDPWTiHYDbbNRbQcafwW3Lhlwj0Y1v4ABIM3qQacLDYyN5tf4HNc3VaMA
ONNLQkXmD4qpYcxvYzl6yc4kg6wSviku06JphiGpwi0nK4mswCwa8rdt5YwsnPJW
`protect END_PROTECTED
