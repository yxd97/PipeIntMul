`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JHyLAJ8X6jfy5MXma2b8i0mWMJ4RnhEX7DLUX4Lv0upkf0kRBaI92whWmYv+66K9
R2VhZaykcwaKMEP3yyo4Sct8/YO6CXtxtTtjrLnyqA9QPcWxMuF2Vb9LsgjW5Xxl
WnJa8qz5mdEG/Jpr3/IwNyHUGS+VqApFOZL9ZThTd58hv8mUDLpCh13j0R9earxF
i+AuaE1D4YwPua5nfWd9xuBimixmtHLrhCyUcIzkyIGGhpotva5qZ1mKGyQ+sNj9
j214dN1x0kZ5CD16c6EYKQ4vwYQRQjo+f9hPB5vf0Ka1U+LqczL7HoJIKilEAi9L
xyHMHPhIwCmGHHAbjrnz04iHhtDQRg7W0ZECE86JBd+3EG6SpDKHm+uDerYAc+LK
S2RJOXKO5h+yD3VuYfz3TzhHtQ99uyy0cjO5q7zbyoA4lUqqVug3LgQLik+zV1rz
8+vaFMRWGr9SGF5/kvlamjER2dL/9r/ud7dPIk4CLiCUSROLUqhhigSKV+ZoGIrO
lB0cMLxLIeZGCGdVH8O0+CxQfBz0BdVdhKuC8uRxpmvdycxoKjrUo4tldfnS6TlW
`protect END_PROTECTED
