`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZaanU8CQGbAssN7VQdD09J6mgOyOKhjT2CX7R4AQ9VfdzAwpTb/XtNedSCKNbng8
dn26hQVb2rQxY1QdyYYFkOaDVjdXWfIbOgKuNEPJAxSwPg6GctS1+k42xsDAL1NB
TkMlEXaBHmz5XBroIbyIENX87kedozpWVumG5lFlgok6OELJwMc49Ls9mU21uFWA
NqWBV4LvLXAy5x3cXWme/63h1xNffAPawGcwTGjBQP1qRU5w+pImxzWAilkFaGMd
DX/BE0hC8TSrnezZ591hWoTxGJ1K0+Df+wUUwbb34++bi+3K/RlUhENK8xC0Mrv1
Rv3lCsW9JznJLh3DL8AO5CwLMTSpgL80va/wOZEt8tZCNpadUYH6U4oAmI/Nh7tv
slPSkZDKNl0URcP0R7vdrGiaqT25cVUR4VeZBbeoWfgcNzj3yvAGsIONkt242EiH
9deyKvInA6IFLoEjlZF9wHS3X2d20eqwvrhaJKYDcou2GD3P2e2RDNcsxNqxwBeZ
CV71lmOcZucMcmXMbkt/tlY7P/n7xuSjIHY63uETIW+KSs3MSPUG0Z/70koKp334
7t0nBH21/s5U1XQSob2mhdXj4u3KefCXWtDPK6sC8Ym2bHkcovmtLF95U+bsQaTZ
pbnMefcQQZn/2cpftQUORg==
`protect END_PROTECTED
