`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fk+MXrUfQ8l0txEsRAwoxQpnXC4/nzyYOgC3rxJW02DfwpsyAoX079fNZJfe+0ts
HCHS6DgEMwfK/G/gFvBHFSGCoAKvyygkdwHtc118/+rL7u9GDqRDe4nYiCtis514
Y5pn9/P1NNQYT9gKOE4sV0N0gf6KfrlHypR0XYu3YplsWP+JVS6wuUfZ9TjdQQ//
COwZfL6dwP3t5xvK465oXt2mGOe6P1g13hAxfmX/XsDK/idAHim5R532YvEJpzS3
fo/P1evAaXqxFcKp+SZ9wQgzJeeMbef+4b7IJkxw74wsrFINE4RGzRuSbLjV70dY
rOY1KmSG38UziBcrOKGvxz1Yq2d1r1892LVDCdv/IkGIk4mAh/2I9IroAdVqJGXM
IYuYDu6wIYgefVRCQ79RfRWqjnZC5Ti/BmF87eS3jQ/Xlb+gpi8cXR5tfIe0Xyp3
v0DcJxeyna0n9eMXzai4rdNzDcSF15r2S9/g0LJCppyudIp+xU6jQhIQxtbgolaB
MAHQw3o+vABO8jLsWdwhIeYq6WDNnJMX5G0WM08yeCUeaWrIMnNx3vv9RK2Cj2D5
`protect END_PROTECTED
