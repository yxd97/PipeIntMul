`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSlwxMdUpz6TiG6Mop2gQ3KBKX5REMzdPtCmwEh99zewSPZo/ZlZwLGGT0lxkYGZ
7hkXIw+dw7jXzb2DWrPkH1xdjMQDYB7C70P3BxDAV6kK2819KnHp/M9FXzufZe17
srzakZ204UwLYOOjTv+IYQYmTArpsOO3R4WrPTt8M2PCxNSjHpRk/h6jcNjNYE/p
2B2udTNqcozCSKaJaEM15NG9Qh2yrf0dYgLyg4F/SwAovIiScwpXoxLsqIhrWsI8
yPPJXEKTWQBxdIbzSEBkQ6vjOwzI5vXNSP4fIJPBNAIcJeYBF957tLn2fENBd03f
siasADSg5jA2G6jvDyGpiNMq6whWUjnwxH/Pwg7LR1HKJppsPGVXDw4zmJHizz12
PYqREpcsIfGnyHikNO8aqdL/YniWfOXpu6GqqfGRhNg=
`protect END_PROTECTED
