`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9VLeJB0FGn+IqrO8Mo7fNxPBcfiJ3PEzgJ7FzYE+VWzwvOkGUDyJHU5KOsliXPTB
CdIdFQfpqIFoao7XoOyfwyuX6gyG4mt/d93YOu0e0j1nFDYdpI7b+ByxcgOxftVS
PK/56tjGYfkEunY+Zm52kkqP8+6slo79HaEtuDYpR+64a8M596UgnL1ewihB2jDB
Z+CLR1+EMgGngWVsofgKa5i31ssdl43QCMWUgLlXMILVI0Lp84PxQOSf52K13Qsc
Iml+z5nIbQeLDK1T6CTIpXep1wYXAqVWPHvULdwQq9HUSP8aso8yMgUNnEvmFZQb
nbmOq5jyE2I0hHiIF0D3Tppp3ManUbk+ZeWwNSkWXCF3XFAJjhBA37i9QyDHjqWk
OYXY8Wy6wllTLBrzjxWph1uRhcde8z0JLeLYL6tmwBSHarArXV/7K5+00cJDZNiO
+kXl6N5y/Aqx+cAGiKhz/M4nIY+TFVAJPNwmMSA/OLwMyqgJOUOuVZ1oMcJ/EB/l
fMuudy3uKknhLCPfMf6S4I/r1YX3zO5PkNcT1r++F6buTnUhiWKF3BOhU4+VMGaM
8245uKoT4zUlwr3knKQG0TG4wEb2zLeU2aQ41c7oLgzupFgS803mEQzWR2oufVW7
`protect END_PROTECTED
