`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P7lFwQKCztazkJZOCF8BMBcO7uobinFxDkxBzNK83oSVdpUmMHbmX0CjIjSp5cBK
nJF1tOM7szOShmklafXofAy0cxXV6IoQd8HMn/UZhJVzpTNfKchbRRmeC+L8mL7D
dReZV4LRfge/GOmRE5VvTxBHJmg2TL9Sa1zBOc+hieNUVf4mjO0M/K9w9E5T6LwM
sjf6x2h7H0RSD8RAInCw/4ZgLs5AIRcBey63Fep+1PfF7Pqlg+Py79LgpNCUtNqx
j5EGX2NYzdBAX+Dx3b/0mVlvzGREZOBwkH3QVbYNERSfZNaAexuAh3dOqjlroZRc
z0p/8EQQnG5QxTOgLDFzkTQzGBFa7CkbOpg+7DaE3ACLaD6Gckd05wB8q38hyvAU
1HFf05qqrfSN4qm3AvfIZBIljxZwFRPnr9Qwi6RrcqtQgaANTu+KlLQGYdracMQy
iNLXyQVVGTw4gDvp5ZWDo0HaKlHv0iVHPg1h7N+EW6heorAturTmQRHmbzL1siHu
W8hKnl9XZB/ePAc98QHHgnlOhEdNiY/SE/Zzg6joZjKkHtvDUHfukCP+BICBVplG
cBxR6MLjSi0dcCGVhyTLLFIGeC7hU2CgXFP8YLeOJEl9QVqKSBeeGuLfoXIZPyXg
/UVCHRNqDh8tBgd0DByDA7U7JSh39/vqVAJtDPuNQgVgZ2IHZUDIQZmiBFQiclir
eAmGaxvAeHGpUgnNaqnl4nrTr3A9EpjYOxUQAgdftNbaKO5RRlGX+v5XkwPfBsUV
tnlwuvf2qHlnhnTkE0JVm7/aQh7xi2BNlZ6u03BKH6kmnsox3GFZff33jiH7skJO
IZLrYZoa2F9dmznzvsuhp+1HX0F2Nxh5BTxt2nhniVZAOBg7RbrfOSCSnLwQ9JZW
OMoFbHlMyXM1puKI+7U/XS2hu5/kUROEPhYd5P+obrE+825VWrWkZKTqFS96+E2e
0riSe0uh514Ac1tOqCdaZ4vd69lgiZFk/Hx8ldyugGToj02w/Fj37H1UvXGtY81f
tyEyl9VQYVBJ+QXG+iSf941ehVFbefgOL2RxQfrSWbhbHHQd+UU3a6h4dZFdfYWB
V3esMn6/xf7Dj07bGbAB1oxkw1zNa3+NNSl6bAnHerH15EPlTiFQ4kc5veqPx/3J
l0XexsXkF6dPjjRa8bxOxz//8gfYrxd5qWn4kRuc5sH2SeYrWAVdNh2huYl9Y/oI
iJeiomQ1nKappdTb9bnTNKY8G286quREZpafp6eFHl/J/KSP0IsNJOaTqzgF1Tw8
w8Z3sFUuFDRYWDtMKzr4bZ1Xcpu9M9dPdwwYQyBYvkw1RhYjtnIUs0yi5rGnvP9Q
B44I98cPxKj6uDte8cVfAnmL8sXcGVVnjJ1IeUL1ilDXbQrzOLDPEmi3L5cFCtmz
wpsQbR0O/8KioXpvesudVOk+X+yhdq4nHkBRoRZnkDj9uoRg16YlD9X3I4kxD58R
lsOPsabImLG3h61jB3i5c4tFBa8Yq3hbe1uyYANKPbtnsc8LQsHej1wM+kc+MMoO
/2YxoT2Cgmrkc1eTf9YqYvKCURx2EhYACWA2Hen5AGWSW9FMWvIT2TTE1hnpFt9+
4vBdnkAmKpinPvjaFBI6/QFbZL6HJVmG6QD9jMLMCefshNNF51GvVrZU2uIpD5Yi
fzf12hge+W82Xz+JU1rOzzThaEOIekFYA8EDwO3PrFveKGUqDDH4zRt0POF9sPpG
Axf7+C02TqXy5NMLXPy8TjdLARKdcJJN+4rBMnViGEjtlW3oD0kOHx7f1+EHav4a
mA1qSktov+7B7RaCaeygSp6Rr8/J42yJvI1OjXzoYNfHazywBmTMVFJv4FCDeVDf
khChFlkZGWJHm4xnHmv97OM7QKCF4aV6xvjRGVzZijPxSrFbA+OwWour+mx71eSn
GMtWJFVN9l0+U/f1svcOuxE8wA1y3557LCsCEL5PTCxgKgpLmhE4AGW0QrARYZ5I
+8kp1fCkKI2cnSWZ7NTE3OLoFobMys/okeUPABXkVnZRu4E+7bk33Ym7lU4/J2UB
7fYDsgcMSbg33w7Gh5pXMOwvxNu30Ymsmy1TyTZ8UaTmWGi8wAFIKCMHpLeCPrGt
0kbgvwQnXqRXqit7T5B5Rzx03/sLsHoOdGkqi33tmeVWsjpRaQAU1+jTY+epfVMs
k9u2DMvGWfJJINZpDmYLDnEifi4vNn8A8H6V+buuf+Prkusyj0RaKxANDLdYVYWx
Ffu0A+gZY1WQxN6tfkhsY1BTalzzYUG+TW90L1si3lCMzQjRXYPShS5p6xMnch1H
vWEmSqAvyYmREUl34so4GCGFstbqNVV64cGT/tpzK3u5uqRWZX3KFViDIjnn3+0+
L4vwggaHFjAToJe4xngniZm6wu72Iomw90A9nvQfEKBQGfTiUM872YnibsO/ispn
RkSxhw1hJ8JglaLeziZex5BwWw8lmTC7fYNtDGaO+UgVaIrM0bufEBUS3zzFd6ay
WEyKDkPUWr7kj4Y3bjczSu/HOhkU9yoV1DtfMtAz6OAMBhWILdQLjzsT4ikumx4k
qDVVoTrEMHHnxpgomkR5bWRNNBZ5Nv92XBX6ivkgfOEsPggNQw1BUEAfa2ik06fX
t3e1dNZMF7K+Xa8dFVZP5C52+dwVuRk6v6/L0H0WA2GcuOBogWwDH/EN9/EycF7s
8UjfDCXvmFYJu4eEN4ogU3PgUjPNFBIdSD39UT/UbaDNci+JuiUcIfDp3XK729LX
vNojsIp2LlUHHBI021Tkhk1XtHIWpM3y7VtQjkf9McbswFdQpojiAHnXpg6sFDBV
GJ3vWOc5vTMSugxCLiRWMz/pLHnLbVeRrqpJEp+kovcxE2zyeCAkQPAoBCq/XtbF
PSuZ7p3R12gL7MjWmHYNaVsEslPejjYLLI2RSt3tSgMmrhdrlJX8ejdF2ZhwSIUz
ik+1YKmNlegf6Q2Aj0CKU0yKExEYPcZCbs4utGHWkFr+S+gQCOmUhxfX11NoXNJY
XKl4YhvXU0Y1e+3wqrgsbWwhTjvVrVzxhbh+hTgp3Wb4DOi1t76S22K5F+nVJMQI
ZErxFufqkwMsZkwzNkN3nvOB436q+m3auYhII1/1aTulwYKZjpQPiyz9WExqxyUQ
IwzHocyf3faKy7uzIM1X1EYsIbtHrhnYbSXcqU9copPWu4EmVEJQXeWPyDSsI1Tu
ikK0y+7l9k2ImKjaCxtBawldcwYxjQK/egZU84r4UIuuM77IVjmzSBj8m6V9//ZU
eMSUEezIwT8T0gWrjin7IZzVSPzRWkaWd3cflCtYXVn+Trf2AJQABdH1lLfI+O86
c9u4DCdoTGpwdgRlX32B02zLD40DFHuYLFGxc+EBW2xdM2F2ZAgzV/Zg6E6ikGcJ
esep+EIL1jCHciUWx4yFGG4dEdrrqKs7yqu2KEbG9HwtR3ZPE2PjKNdGVe1UuH5S
uyIPIXaLiN6pZX7qVkpZBxlUiwoZmU3Dbz24f352oLuI7AMROhCtjNwGylfWX4HJ
ICySzPjoltPK0I/DOw/Ys1X/AWuGoF3AxI8zBz7QVR5+0N413PsYtJKxTPDmo25O
jXy6CLqUvWtVdZPmOJ0hRjgxdVgGew/XmUAs9uWgPRLzZDp25qR8n+y4TiclID12
KXNfVo28cOwoar7XEQWKfJrQelBEi3c7NMFmH6gIGXl1tUHbwDDsoq4EH21Hsgmb
EBzjmH79nC6yU18aHNeN+hUl6b9XXGG3PfYiXVWRr9Lxi8QdHP31b0OIMaE7a4Po
cK86DgjMzO/eM6MHaSFPQ+WHjesCvbZpMPUGd3j4wwUv12x1OD1StaocR0BASdDu
Pzu+taP7Z6ZqiwJKR0t6KbJ5KD/siCctI1V6tiK22vsJZnT9srRmSY1kojsFOAUZ
O7QMuQMCL2hHH2zOy9QDVrxpudK/kKvxqyXIfPxapOY6CRKKiogg7ZnhjBDIDncG
JYev0x7KdCA8n9hN1IwkPf25AK4nC+B8rA7WsCABM8guGJBQ7tpSkJDQH0rAOiKU
mMUmRLH4gMn9T+ZgcPe06Q/eOmrUyaTBvDUym9FGP8mZhiYa/IfUXXjK1OGutG2f
TCuW5Q4dHXuCGA3b5jRALOd2TkeFst6Sf/3moD39U+MivAqQUHNNUKseElnxlulR
`protect END_PROTECTED
