`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wlTXMK7dBYrNvJ/XF5TdNmWdGOLz9DXBb4fiNKimnQhd626SwWlLt4wAPZ3ERd5V
bhx7cbj89aWWA6otltLU2GEupsvqO7frx5GOhwxPNcibMBvX8xgL/CsH2T83yo1p
AZ8kvQPkP1+afHbPCBSxUfAr8tfwDai5SiN4zy9gM4jpTc6pF+UFUYTHLE+fbxG7
oWfwRjIgX7c16KBYRLFHsDX8WOKuS2RvXgsQl6VsI6u9rQIwQTaMy2mba4YSBxLE
RfrHpdouxOz/CH6gAIPrGyZFyWZdWhwVDeHBapyrljLs1nPu+mCSAMHxReV77MJN
tqlleM/OKY+gldNzTj5x4OFXNvfwvQFhn9lUrDh4eKM01tBM6IRu0tjHh0OuyJAy
/vO4sdODmWd+plYmKwIIIg==
`protect END_PROTECTED
