`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
60XMQbjipopLin+DcqLmcg+A3PfUd+yy3TJzwXV9fyR3gsQnEXTdIhPximkQ36hH
HDTBYd17kXsUNTzVfTCzT1HtFG5Pz/r+9g3LIHWhFli5XoW/XuGP5FFvceS2T7Qr
/1DbXzZ1gbW4wCTmabfJCjuhFl4cUw2I5BSy1nrxhDcWDdz9XyfpRBq5AuP4bKsP
ryjYua0sQ/r4yjFQrB2cuhUnscfVF5atwn/e0cRgQD54rt+5JsmmCPReJxQJdPEW
aen2DDrTvib9Kl0tkZpvplbhw82c2inzh39SJgXhHZpqQnP0UWAbS9Flii1JNi1c
pRbHCvKa+7c936YsH4fJyAy92vixRKwgzqYrtO6C+mmfU835QvpIfImnldlOHeq6
00jYpEgIXNDh8nf89mSrkUJJEBN65rFuqrMtgaYI3gLeJPw9BhHPT/xggyb76FzE
bq5N5h6wS4I9lkZxvhco4D+tv2xCVvJnvEAtGdWP4mhSGnqpSG6a74+B6qdhYEIu
`protect END_PROTECTED
