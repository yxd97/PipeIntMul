`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gADBAVv3TGVt3tW+7tIFfaI3uJaMjDQ8LVSwvzyjwI4w+SKyEhX4SfUlI8TVxw5f
Ly4Q4PO56SPrvOKMDPh92cEcrGo9f63ROtegExRcraPxYa7i8PPC6CfW5aR283Rd
NoZ2fwezN5EF49AD69os4gQR3UaJ/D0GuI/5si1G7kin3lPLNEF2cxrkDzgyJ1dw
TlRK+xSL251F4h6Gz0XKDnHTMQgLRLyLre+DiJQcXNCIqfiFQvwwr6y5ZKNpAqBV
gKj58+fp1neA36SEbVkJYfWX67Lw7lgNPDaAyk5mxBi9S03ig6aGRd39RA3+XohL
9SWdrbSKZtr92hMv6TYHW/3tnQxqVU1F37PDUEtZWhnAtiAsc1GvsdnmmFGSlYFn
W1UalJPFJ0EZ0uINMr0E+IgSQ6sx/S9aOg2GU5/IuEGzwA90ApK22C0ljDXOLDqT
yhY8JkB2fL/5LImhT7o9dM3CkTioccSa7rt/ROOmoOYdmihkWpULNDW/UfLt7EJu
9y9fpwL5UZS7CMcjVSiBjQ==
`protect END_PROTECTED
