`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mGp7Lf8BjP32h8ykg9EUjl+ruCO2/eb+N+JqkvJpxJSusbKjTKF1NFxrcxnDaXYW
VuHUZlkPJ1v5N0pRcjjRl+9fWxH31Oz07Z9/XK5K2HMqFbeE3uRRAYvlpojNAx7Y
CLrIhAEFax+8Tp6qtdg0+tBUWA8zG3fJE5ragmRxfDIAlQaqozMjoXnGqWUtm6eH
PSD4yj4+krrWUHlOnLlnvdRUQGeetZv/R92s3DEjlbM=
`protect END_PROTECTED
