`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qvty8tiSK961jJZZUAWPbeKmYyvYMPDkg1QzcOo7x73Dq2l3Qov0V8sqEAafojIy
edm/x991RiplO+0VRCqz4htrNHn/aqJ+NVSR+N+afBOKB80vMauSCA26YCgWtP8u
x51VsTgQrOi/h+gPldVUNTfj9d9SRh1MyffgBwKg/J5PsIAM/RQf5NHGnny7XRYk
zJHj2nVg5ZLnOitTSGstNSIzLuY/EsfhNMmYgjFzHY9zO/ipP3AQaIwCbXyuUEUQ
tg9MG1MsR3lFgYHKNOBjH/7miESkQLS7iIWaFz+LwbW0jyZhtREBgHJDskfY4aQx
K88VgJsV0VH6KXPMBqIL/hodooPM3QXHn4PYTkayRydBOgGa1Oct9RW7xrdemEFh
asbDvkYJToRFsE6b2mV2rrx1mLzf6uKAGrApURwaQNBwxXZG1BTdLGU4psYU342g
SW/ISjKHUjj+RJBBVZ3L/WRGOiphlGdJ+52wsNfJSpkoabsAl0ahxp/3Ommnd3DX
89TRdQFhlIhRizsHyebO3pU4SdOh+4DLZGaXbvsSJ5C60p0IfNHKb7810VCprntD
WktlPSzqUN0E67dmi3Q7fJypMSHgNTa7eOAtwjuuhRD0yBK4s0f2/bu2GoBcjUXV
uRmox8Dht8izNUchZzIw0eG3PRDyjMkrYB5jc/+DRKLhuCjPK5zbiTyrzNbiaqJr
B47TnbCQaDFyJEfNABwjUrk19RuW8LnQ+ugDG6DHxknTtaTvpj55FYplCQoHA2rJ
4fgHT6jGQwXNvZxGlrYxmripgXDekCqMvfvphBnQBMtrcCSMJgZXlRMf3oGTagSE
kOE14hhd9NYKt6F0UIhnPw==
`protect END_PROTECTED
