`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IesAymzweWnjXJgQrQGTcNpQ7yRJWHN5e/YRE5eigaz37Y8FDY578kZIBjghDV+u
uHpfv2RYOP3grUNKDk6Qj2v4/vY/TtW9E6KwTOHCE01x1poysWs+7AFSBAYZuCa8
AQE+ejw1YrlscwSFksPjGGBnAveReoUw1prhFY8TnVvq4MaC8zdChb/mDW6Dn69o
M92zjnlbAHeCzeRHMvp69GU8BQtst8QJvarpnFQjWcqp+onJGWX4e6HOIZVTID+r
md2w+iSogcilqHkWQ/Sc7XK3oakncXfF4vDRFEsEVmn94iNkppdOh7863KqVLxqD
2C93ZhSRiagfTFx9ggg/y2wfoYaJi70QN0BbI/pLpcaWJ0fTXONkYbOc3Vu/9j5i
rRPJHI63Q6SI1kMCfgDtKt7yKFPBh4nZ4P0L6ua0/TNgiKUaMmdUKomeKj8quVD/
fK5wYioA3CdjYVQ/RVa5Gw==
`protect END_PROTECTED
