`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOSxEY4FdX/WIw3xEf1fdJhq/7dIu63aZMaFeEzD1XcwkdaXccq0iA+Q6klAP+ko
ll9JWMGarZcGJtWQl4iDZQQFp3Bk7ZdOW8K30L1ZIg/T4C6CKsZYx15DuXp440d6
YSYIkUq1rAYRj4Lv/O4b9QqWEib6pDmWCeYxJAM3UeqtjTMfexWRoVgyLcKDrqKn
d32Hoy8OY4J8FlcB21FAIiaJVEJK9Z6+6M/ztEkq8xwgx4jh+Xs5fqLZQKFvbuSY
vOzdVjoeFr2qQqs7RqhxUukXBCAGc3h4icNPNHl2i81G5yoKnufghkeEFD37bvjF
LA8Qdi1SDOltWAF38J5ZotP1MeOdVSWhyuImF8gARNkzQiOOIS0h3//guWbIvGU/
pq298CMwk5eHs7Q06tZKfg==
`protect END_PROTECTED
