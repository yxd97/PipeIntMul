`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PfBl5R+KLLtxMPoVdvKqzwcJ/zyLp1Mje7W6aisVZzA7IctxuxDV3h48x/DAdSTS
zGf21QJE08c6YK/KeygrSiUvPvuPgNyXQCR7e2NKz0R87mEM0LRsFKU+Bd9NAfM0
h6u62+RHJqYY6YBxffAbINQqO4VOSiMvAUpu/hWa23/jOIhv7SfxxgqAlXxqQPr3
Yblsan4lV/YEj0xqx8ll43TegVAf6kcIFn+BNx/GlQSpP9hx1PpLoL/wTwdAyzgT
ec/JEUk4Qn+HFaZcpwHAkg==
`protect END_PROTECTED
