`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LcFRrrxMsvfIyGixkjpyL5zk9h1yXcCXX8aaGsvZyd2E0T3jxtrYICA2WOipnnBc
LTENFyuMfEtqbeMNkH3c3n1f26Kh+avxoo0odb2h2BeAHRgtDYluIrPr6utNU+Ey
czoI/NHC5fXYkggJ7E7J/KweQAZqt0Z5lU7rETL13m/bzp/mo9n6t9usiMUr7FEU
cDIjQw0CmJempTBE/ulgKTnIma59GRdfI6kkFyHekhSTS0pk0vtNVKEY8cOWuT+k
M5g2VFXMQ6MN8G3WVCT+Z3kcX1gyJVTou4DY1khk2CRzhSZvjgd2LZ7jMZNhaLE6
v+EXBUJGPdSmKo3SK3SSEMBzo9qumHjyCyGqRzFxwKdMtzkPupEUDhBFRT2av2+s
HqsgCZhgsIny0qNvmkSfSt7m7W9D3Ey2f225dnVRB11fMCNI385Q5StBpB5i0suL
DbNTMoZbksEQJdVkXInHonTtXDa3AQDVJDrcHUbdMUc2Bua8h+JYhTIuTSIc77Ss
mz2Cz0RSGqcaSIQ5HJYaniSlx2tApcu4wbjJWjYkmDI+pFpTPH8+H+mcYCjT1z94
iBSqmbhXayXg0ufksa6qjw==
`protect END_PROTECTED
