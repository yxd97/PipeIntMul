`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59/KYVFjGmPOPUNyNtkZpO8dbKZxbTy9T2ULxWiHBW9i+kfQJWBVj1DqRxEZxIgK
jCUQ6OQHtTnkkpJDyciD3fbmsMIYGznwttK8TVJcWL2yazy7DUOZgaCniD+Ev2pE
xfijnN3PGTmRC70dHNmplZWWSHH61YsbOr3fJ+nmADh3xkO5QQn9ljps7Hmcn/8+
rIQ9vRCxm5D9XHQmLy1Cu+FTAiNzH9O2TfY+jHhfetovjACl+SKKO2AbHTAn6BuW
n4N//jHVtrTk0xiPdY7eflP+8MqRy/ZlYpvnK4cSYQlJsMFey6rVk6jcGxLOKATQ
Msd1V8gaTUGfWzigLZTxeKakfZPDr3SIbe4Fj3tEUMjyPbjwdpB8PIRKf58JqU8R
+/chEPN5HPPgn6kQG4n4dQGvzL1lAuv9ten2z0NI4fc8qk7aWv7CNqXudEooS0Z+
`protect END_PROTECTED
