`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/ZFWTcLEx9mAvC1w6vulRLPP1HibQaCJXl+bUqTuna5rdzpGkDL470N/YoljLm7
Z+T5tJc1I26Sz+crMxmuLMpFyRNqjyGmc6JSvHUPIjEPNMBfTvCrnr9yFVMT75oC
9xKPHcjvx7M4j1BLaCsoEVpjmzgNqqjIBkOw/ROubtH4aQdq96zHtqvRwgf+pgTZ
IrAibiDWULq0dGfoVnlB8W2nDihTjsKfX2mYJ7DPyomaMvgcDjtae11+X4k9IMw1
9sZxx/tZRtqNQqxvtf+cRYnhncA0BB+RuKMBFCKKeeoYFOQW5Kzft3kGG3R0l0LW
xSoqNsv5qgv8JAIYt9DVa4EA1Qf6aWt7A/td3b7kIvxCR1v6QZPQak3JoGr3MofF
AaK+M/Vr2D2sjtEDCzIUlrE2xcV3IntG06G9ggpgmHPxtImQKFmrB1YrJ0aoLL5g
Gl8nfCAZg2AUE3qGRVq+UQrSscB53qAKtvRtOmFSjzNQuqw1ysMeiGyWSkML2GRc
yTWcwaHnoFnm1SnZLSsdUNSd/iuT7YAhIOYuMKVkPknSAZWFkkAZxMI57NqIlZj0
I6aMVUjSbcBFbJddar/T4EqgqcqgJLLR8ydDnVAK7wxet9ZQtqtsEwKoCU+qbF6L
ahcMuaIXaz5pDLfSk3HlOw==
`protect END_PROTECTED
