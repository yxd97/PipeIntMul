`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qaInRdVKUCR+2iAF53g043fBcwCkyss7IX1p7OVK8CD5ipKpnEGJFvW/fgWh5fuN
mc1hxPpzX87IoI/5cnBWaCDwxjAzEkWS19O+oC6PQ9iyDeBnjU3PTMOPm8GGXx9+
ydGgvUfl093H/XBRHzHisysU9E6ReMdKfNKsWXZhif1oNySZ2wfp+fkZZ6uJGUTm
3otF/HcCGefM99RUJexWmCuXO35HsC2+ljbpsa2TqFpgyZHKiEK0PWPOh9O5i2gi
Fl2DRazDHVqwK1BrIGT9rKnYne+C4FpOqg6Wb9hoyTWydop2LRX7yHuwqwDPAGmo
TfcsY0m2x/G3XLbMzz66+RDzZE7HMZeGLWSOcUY48YkONp86IA9JWvS0aT5lGMg3
SfA8Srfhzi3AId62b2tCT2NhINplI72qdpqe0MK9Yp1MDVl16wTtmqTJLDC1b3/H
VV5nJDPslKKiroX+BGyOU9AnGoz7ippVSErZAA6b1rjCIyWw6mqFR9cJOTLSgVuj
4VJThEhR4yvfTAdP9C8IibtGKCzYBj2f46kouHL4wCuje7bkrIiRqsY9gHbt3sLC
gGgCdZKyGGKsVohPdZNOpFAcEkn2sMNwGUw5fh/y/NgZ5iZnWPZfslg7Z0B8Ar3W
0YBtniEvgQytzFUhg/QYgwf0pID6D60YTMHAB/kuO66CMFPGusmEn/ofGmvchhGO
2FcykcCE386bxvxvgIcg+68mmhxKt5q5AtwbeJQypKril3UtrBEtZBp59s8gZU99
`protect END_PROTECTED
