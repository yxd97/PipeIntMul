`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDjvPmQEsJ7i0QPUWlwJ79TdItBS5YoBA7tARVM3boXRs0sMvPl/mBUpdIAAQqTQ
jTNBH3D7nI1JytSnTkDC4hJ3fma+JKRm+VcV8AONnj66qtTKfABzDMZOfJEMyXsq
TgTnzsYcq8AKdcJI/+S3GLCeD5Z9cf1Mw07dcUPtzeo46xGgYWUW7nqLoVN+azY2
aCqQW8UCnbhieDsnlubAeS5DGS94mUklt1+syOJgKHMF2mKxaozYRKXGOQSZTdAU
MsESzo2X5wxGbxpLGFYDrLDEvNkMW8ea57AhEyDyo4ur38ugYwGvOMBMBLEdFSXa
LllFzyak3z+CikhO/27gjTk3/CEOv3qBIHUrzSsgZoLovvgSUppK/pHnrx1k7ly5
bfi/Ii7UNicm/sjz1BQxrPTTXc3jE/il7faKyjWMSys=
`protect END_PROTECTED
