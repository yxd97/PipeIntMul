`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UTELz1AQnxthHsQ11kuSQ/LXbqRADIcWDm5P3dLwXkLWHpPasV2fIFkE5Sli2mET
EeJZOLksDpmVHlDxhokR19AmsidQqzf3qe5wqnn2ULpM5uu5YGvWIC0bJ4+5GjVj
I3YBg/YQQSCDbzZVP+uNPMSbwER+Y8RQkH2uiwy/vANMeHdPIc4Mj3b23wJBU1fW
VEVPQ8uxEc1ozqzd4kKPAbOifmQG8AmhjtGcdsstTPS9glaCmvyzwNbGq7d8BJzc
pUUw+KL25RCQNXg3Q2MOADlyFjpiCFx6ohEOxYp+IKC+03NmyZZHhTC4U/xcQGOs
smyx2k5A+YtHkzKC3az8GWD6kFP1JY9h431m2om8nY8/klLe0G+0rIb9vwY0aL+u
Y6XjDm/mrXAQklhpayAp80kb7iGGWEdmJknzT5WXOW7WIXRD6a9SWEqtNLXtOFf5
`protect END_PROTECTED
