`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VE68msxbdtwPPdYJkmYeajEdkPTi6Jz8EnqOVRngIJCzfeEPa7KaURHv12Mm3jGp
jg0o/FtoDEQVZtNUvEK7FidU21YOEEKCWG5YKkHi9TpYZnYWpr+zLujOhaVEP0Fk
j4V+CSRE9QBYPjEn1ObbDXz/PhsVGe+osAs3jM3eLYmWEvVZCNguwEUbTQ/LS9Wp
LuFcybrJI4azblucauuqtWUSdJT6AEIvi30HayNBPesli4AhaEs5ENqoQhR3hv7N
p2wBXMJagZ7QaXeoNOPzU4ofeJkcQiQTbGSrk7bSvluz3cLdjef7eXxqDBgX+tmK
7sB2WxGN4XBmSU5sHR4PTlNzsog28VvA2fNCKXQS0OTL3QC7YXLqPN76XPZdZTJk
AZeByXM8bJqioryBgfdpYrKmt3RCIVRAaVWDeGn+rZ0495M9WlETzfACxIpRdfhD
e1TNbUXZeCp9hMhIusyoAmKbYOgJBMS9EMRVfEmjnbJjrbiXR7NbCSWoqTWZMN1+
br9UdOHsSVVFOdcI/YrLnKVzY6sEVjDolavSrGT18vthUL75jPCZOJjt8HROaHv1
SigtM5bh7trDaDqOMYiRYcG8SW4piJ8mHpewGNGYt2I3KFr3Z5zEpSOrfckALue6
uH+73GEMH9dXZKf9dpdYn7+I3KEM88h8+F3S+maSQC1sMEgTn1frfsDWLBAbM134
YIfUMvNshyNS86MuT0A8wqKt0xe6Dfy2mu2oipphb3QELfsVIq5XCJTH9VJzeW1J
wnnJ4V36uhTQAJ2UvLPuRUXTy6VscDGq7bg5FrUTaGswzRLuyaRDTb0RXVpetBZO
IpAV/rkeJaKr3zU9DmwDIymgxQzXtkGFs9o8/JEvuOTr/Q0FpoQKHR+lHK2KZNww
MbjRVCyirovKnf2gWRzTl3yW+VyDo7l9mDAtJgtILbi/nLAYhzjHc1Bq/ULl8AMK
wdV7KWO1sOZ9zrxGKkOLpwjH+4Tve00eu6pBotF4RpbUkuL+nKG9rMyJTIVIbVr2
MiVaczMv7b0iXii1sfWahv1BMhOhfHdqlwsVSYEQ1GDl6Lh/52boDlapxJeprqdZ
PTijtMw1SB2oTadCTNbqlbrSs4W1vbFYa1P5ZRPNu3GQyPfuFfwVyc3/81R66qah
G2wF9z2/m8ONrQE4ZY1TmZvHbVuyWHKpzLw/YX/FmNtnSYLlbWEf0NhH89UnWH84
4Q1H3JS7NPrejgIIb5+Yvh+ot9azBP86gYzbvmQ6WF/trOl6MHEWWag0n/oSpK4I
JMM+usMGf9qurdRoc+Ohh8B04f4DhGsBWuLnZUlNtaiQJyA8KE19Nl5IPWiNeRIS
8FuN/3ryiyFKnySX6lFLlRMUhTMDJPdCbM2l0MzAdKzLCdyttY0g4/vrtZrS/Uh1
nkbZzFSP1+S1DnoeJ3WfZw==
`protect END_PROTECTED
