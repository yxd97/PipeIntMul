`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B8JBBM9TgBbONoN7kIqMMF2MBpns9OH+n6REZ0pc5I20S1xCaJ+ZYjHZ7gJft4Op
2qKruFgP8ikFgFgrBIf7HvZrBsqykNk2ZB0vA1N07kdOx1pmqeiXjDepXVyX1Q4L
m7aNSyo5+FeGZyl1zZELx3sOn9I+awVdKeLQPZdpQpXCMe+Qrc810yQ3OwVrgjhE
0ZKUD/NtyqmGDd6emTLl22iEpLCjyE4Gf0XEuC+BNrknltvBlUiREMLM3Sm67cI6
EQbatHS0fgfX09W+SGDXOrr55o10IRNRykyDxlcRW80Xi7Q2+kIRslX80WLVCCF4
XMSgrI72hxxCuEXk5hJGeQSPlHVf8oTWsZ8o97UOLt8epIYyxCJ0tew/b7VSENIY
yln5v9O9NxcesMAF48nw2mtQvvazPr8ASqBaZD9xCYmYgrjzIV2OPAUfWluKeuaZ
X7mbSNWqsFobpEihUoBc+w+1xkDJ53FH3ZD98hPBIawl7AXvTpA30V4IwMA0wV5Z
YoAFEZblAPFZZ30Q/57WXkVmYVQEMkrTpwLqTZNpNYJ5nRGSrw9rbnqXXSTBC8nK
`protect END_PROTECTED
