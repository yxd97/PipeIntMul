`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uuRufZJRwzpb07zVmDQmdNQ4ynedyDAyTexFXIfJE1aYX2jo9kaPVo/xHxH5paw
CpdGchZd1jfhEUJFX1PrVgPwuFEREWJhiDE9qUehnImMrh93ravYF/G1eGaP7R+A
CGCoh1Jc9w8lf3I+AW2m5N0cxnYYoJPOQzciIKtY7k2D9yoOAqezh6TRh+ool8kB
lT1w2r+bghU2AiVos8y/WrDj3K16jnslsW30W2xICIPMK4yDbCsJ8398S+iTNV3G
NRAwajdMQdUr8Iq7ZqAOyeoMRzCoh01MUAZcoqZD9rcwF/ZP3T/6gxGLbikU5Qj+
WjEJbTp+I+wcy4TawyTBmQ==
`protect END_PROTECTED
