`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QzgJLS1N99RnznKaopuy/ViuujEg4PfN34mPtboey0c7rKU82JUXzNVtpgY4ITwD
ffp/cURkQmHEIK5lXq09Q2CzB24mQBc2fW+8Jj8rXCOf+Ya8X39+LzRHBYRK0dGI
R7i74zdaQNSs1dAe5VER85SnPnBLao9yMWoCk0yhU4Yj+Mo2e7zx+g+qWp7xdTCi
ssGBiXV9geQhv/VH6eIYgoJIE2fqa99uYFPn39g1Ga2XujSGRMD5JnfnUnCV7r0B
PUKdzAfK295quLLQMSVOtWPV4sgqVHoFO82qNXlxDfFEdM3WMxsKvZqmyuCow24k
9AqW8YCHWlJAzA0vaZ4Qmu6R96+Serlp563HwgZBawur9r1QXI2fp45CtaWNIZYV
10ud0klH8GLC0m1nu/OQbPNwOu7r4Sbob0lakF91Xjo=
`protect END_PROTECTED
