`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZULFA91TNcau6DKu4CH2DjY1kvUYvIlWRKSDEDxo21Oyo9IBhR9ENmIFUOq0s+u
OI6CLyGtt2r0RSgXGiY9fVGDjZVIFGVG2JkoIcRgMOEmxlZ+DbwwV0AicbDaHssc
sl5tWnDHQkuJh1+c0tIWIvO4l7kvSBglZmx05PrXVrMaioiLP8aiJqkR9kUVzv1l
0YnMRkuO4W+EQolN7DrsVD0lrIj7N1SEaPQOv+JXiLDUoQbRULXvgIawYaE98Ohg
5EJ7qcDGqbLScitYiHTF6YvrbAeB9qranJOilL28DoCJ+MrUlhLiWAEgcfEgTTKe
Kgbv8uOQ17GKBqndw5uaZMFdDNRlIp3hO5Tjv9ueH+mB1SDKpnuigQdm2VR42+9d
08FCiJUscZQr+89UNT/SJ8nhCAz9Gc7n/1NAEln4zCTb11fZ/kNAcbsD6iCAsBm9
s7GqxuwrrneY9vzL0qllhZE3h5C67W0bTUEgkKYf/GyUR3ZEGPLjXw0Wa8B3r4rc
AIaquJ07iZnE6m2VCn9jp15rpKkiCGJtOmFdQFpP5KsXPTh7lBIHX8cpd2D2r87u
pEu6xUQq65U9M5VAnphBpmjmkj40dMHa94X6mgQmM6x6IGfp27kRYP5kPlfL5FGe
2oHzsDzsVgEVf686S4VwZ5cdSFobKWW3dwFV8HWVc5a1PTpT0r5+s5dpnV1ir3vi
XHwbKPp+CHuGhH2gP1/bjeuOqq3kLO/FAHwTM486gR5DgzCn00uW7WWvKnsGV/64
+eTWgqx3XBatk8S1/O/P46s8tH73V8VNyh/OOpM+AbMMau5dHQZ9WhEb29+dNyeu
+WMiktxQncyKnwltavOGpb7jxi2z4mAjfnbbaet269Mc/MiONj7DYifV5frcfSYF
yMMWDGdE6ivY8xtX4zGkdRLJOwjNp8OkcmsCnyyfE5Fwp4n1zJuJ0WUmx3aOk4Hc
3LGX+6n7iq+BW1RJUetMPPKTFUfUZy7I5Dfto+2yAUuCaAJIEof0LQZkWilgph/Q
1gnimQLJBkzmrmeBi7PfHlRTrpRJHgmt0UaF2TttQ4/EJkLT+rrVsbV5EiY+UYeS
MXLVp6abp+Unwt9HGy3q/do/TeH/i54uAovKIDRDntSEms6Ulg3j/th4By4hIALT
`protect END_PROTECTED
