`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2P2AYqudyWzpLE0pvWZMsrExZfv+Aglv9vKqj047PEj5WktYZ1gnK8BzHKDL2u1z
bB3OxqEzxIgTxBd3efJ1AAMPgncp+k2xGBu1uw4Wa199y/ZXk7hiEji1UljFvrC1
fX1jcENdCh3oE9JxbREY4hmM78YbXOD+OvCT7Yk3luyV1SyiYTj0vQfKKX00yCAD
nsOm/lVWgnWyRRwM+xC9rq2gzcvvtnIUF2b6pCpWWRU6OvWgp1jUuSqPhEpDrQGq
fsXTROsHC5g9zd7AxpqR65abc4MtuxOUz3NuR4ivO+CXaBbGGUaSb5W2VDTP8Lpd
AUQfWqeTQURritQq/03m34jTkLnZj2vAtAydP+5u+b0MDwYK7pfgFHURO5BfRMmp
Dcw5AkwOoUD2PNC0qF072pFPDnLFBshzeS1f0UWMebc=
`protect END_PROTECTED
