`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eQy0/XlwV5FCrJ+H+2rbtZNUlRR/IzkMgaFGcVpU/n76hxVVNUHH5qB7I7jrUiyv
gYv2zl/a+G829Np78j0S3yDzxRQNNfaIsjvzCfQ/btCUyS2LJKS3bj5slYlw3YEe
mxWtM11U4CIRJDQLX30sQIB0GGkdI6USyEa/vOvxVJ9/ifNBkGdOuhSxCTe9ISPj
I3DYbNNQO8rofxeaD9141LK7UkKJmgwRO3057poTIy8/FPiHiMyaHrAMKhOP/NVM
sFqC5/dInUv6613RDxgbuW2MPJyMMZVFZXC5OkDJAI4RD4X4hxOrzmN1+s9k2MgV
Jkl8QclcB/nZj7Qltxq4Kg==
`protect END_PROTECTED
