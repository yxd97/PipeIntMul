`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJrlpunUCfMd+WKRMLKHo/2wSmV6HFvObUbEH+fDAhxEys5WMCIAcPtN2pekpZms
kzruefQsPdsmCyf3hvBimktBI38KXqid3VhBHqdioskAD9CQ8pcHzlxqHIm7+xlP
tRZDXXl8EdDvpCXmuAVLV3XQzJMZ9/Wn8PxVtg0bi4Lo6aa/n6jQoqopFrGY8xb/
cGCmuDeAa3rDwNR8VVUMeNzdhWqvpjQgDZ1QKOjsrUL0CTY8UnqOKKCMJZEy7m9t
WdkZeFOyNNWIhWisE+GWgzLQKzqU+HuZUZWosOmnvEIw5pDkChsbisXQf3EKtCp2
F62VgT+f8UysW0CCXZ96KTcwF2So2PkKHJxcQclnVI+qEd2zy3iubWtzvSzt3/00
LbRNREunKNqDTOnSDkm/leaqO+D7aY8tNffCdW9L1eXrsuAPIzwm8ToX9Wx/INt6
0dTzaprL1M+QHvmdZzIZ2PYHEUzD3DtAfDTdQmiHPvOGf57mAQlGlH0/ZJr1db9+
0HEw729chfM3djiN+BI1mt8Wx6e/sZIHDVxN8RDoN5QATj48Y1IGGPL32ZvCuG5e
6ViuufrH5gP+oldjvRWPYomVnP0u8zBG3dxegwIXNMT8497EBl7pgsqsDPVgUmlP
g+TdnZrMtw9vCvSKx/nK6JFBeSyflCYyBrMtPfxwXl02757fB7s/ZoYS+D3XDhmE
nmVv5fiKUslWvu2sLXMohHxnv47S1BLaCXqqKFAprRbQjJEYDd/LLZ28+gh+10Wx
h3NnXtpOKftL6//jF+lu+HiHWSwrbh3cZ9w8SrZbB+LaoS2wtuF6j3se8/woV43b
WmaPSK3p6wshQZ+wp7z82v6TsDFZJVV68F9xJLT3q/OplDojnkH8uNXRDb70/9xZ
6dbVpbNSWM3CgZ7X+DKkVvD61J40fUV5SMiJ8q35bNbyjA4mqng0WrYUjpGSlh/j
1xrz2fDvzdNYKQLNgjqyxmzPWhEgvllLkBCmIFVPVDJy/Q/F1AtQeRzmwDQb1MuF
kyAYJLv6UmjrV9OfJR6/4aEwSJQh61PysjpgWjitu5yrq9mAW+t759G6EG5j7Hra
m9TyfyuOtUDtzRHigs4Vb25CeE9/R53etpG5ab1etkXeS/Q0WNg8dRTO0nQAeaqq
DJgDS0tXReKc94F6O465PCwnArfagJgKjBqaRT0Gr65wuUt0hZSaSP0/gGUOY7sX
wNLTEOb884yQzI1VGHHchV+ohuMYUrg7Vbw9x/1hyoP8i6eV9gHMWp29N+1i9DEy
5QZCXLQLuXnk+l7WeL+kIEeDfU1TzMbrx4yAS8o/nMxgXCfQ84TrWA8z3VMG1vMU
ebFPbSKqz/RZkmBrUIHw4i3n3dmSl/CVCH4A0BORNfgkS4WtrtiZ1ZNmYArxkN/b
B/Hx4ji+QkZqV+SdCkOFfCu4qBOKSdXaE8PyDnr8cEteWfc7v2DeQOoD+Sp/mzBI
tkSwq9mpe3ZbKf9b88Cj+YEYrFT53XU04PLOhyqyz+8uTSZtrmAbqeN40/cEmUVH
NWDRflKVRt1bmbQDPWpDmAeUbYJ9KmACs3+4V/6PY2UXs69HulylvE0nF80javJP
Nl9/tnJYAH4t/llhqyv3azGqMePGpmf5j9i7I6IlrnSmIJvLFwrLajdfpyrtLbSM
S5iYIbj/myJw7slpFokfeFao5dTeGvywspzVtmc+vO6ON7WxNF6KJ36U4uqsJr06
4ZkEjxYQIXSCyJ4efeJzxNNipfi72+VP46T2kVzqbCLXbbJnFZrLAehGyz6eh/Ez
bUZ3Zqk4C6/a5TCzVa76E8O4nf2q2Nsh2Yh7RsQb92heLV9jtKAe+vGpvPdPao86
PTTm+21UlPboX9qXd+NF2Z+MY8T7P22C7h0fVdE4+x+B0jH61iJ6YbIccYN51P7o
yUJPw7g6zzi3HzylgCL/feI7zXkgpEhNqs1TRFE3A/sP2Vv1lCfDg3ubEmpf0E5c
GEKWbgfQurjr5a7fWxVvJCyftwud8f/lDh4eUGgYqGw5xYzc/aSCIrCbH/O2h5LD
EQPd/tnbjzMWD6ZEVoVCxEEjYxxsCwTUM5bABb59jEF1jhdbQbXbeR/hmyhFdU9m
YJFLYSfUwxFYNKaMVjPHu2DxQTv5dtBjC25Txpy4kjWefztEmSBRsdJecdHnorWw
P3h4Rnkm0Ib0tuAipIagzS24HBpIfmwaE9Km1aj9WjFip5BdrnS9WKDNzNTXmR3D
Jv2Fd2tO0f4DvLJHocdAx62HXtvkNicdbEoiglaAvrVnaxHmeLvXfTKUfyIFFxjm
zpuRovrr8hRYgkkNjuC0AEB+47+R9b+8zpeZQQimTfJKeWwKcHhAGKYS2cXbXIKo
JcpL2ms4ZCn5zbKSnf56ci4rv2nJjBubsCKOnzrMyeoTB/15o2TuJ+GU7DxbvFoV
vIGhJLNHdARH/zFpu695V9XrNLC1B5vMZrycjc7J+DTnV3lkdBr9QkZ4OWHdpfaT
zNtZiFzwtupVGCHV5j0r5fopwGKu5QZvhYhXPUPXYqcrQ34Z5OGHdLzebd1TjRGz
aJIdhtkree+XjakdaLpSggLBlj2MTtumbvaxv6oxA9Zvuh7aBWf7ASfd9CqiwFoI
pfjCP0WaaENme3HGnsjl+4g4dyy9kPtAU+FKOAc6wwbGVAwuNWLThGKCCY4fPLok
JPIq/A7Tww5zRLc3T8aYDmUv78EzM5S25y+HLgb4gCor5L7n14dNYgM2gZgcRamt
TT44pBk6bVxZlZ+CJW5PQ6h22SuguUmZR4Ura78AM+3GptIAKlMo7T9RkrVSVVHo
`protect END_PROTECTED
