`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sAeuj0rPJtR4DyYcXzZU5gI2XCyKE0QCWr5wDWBHyP8vrdlwp54Wj9bsvsjYl8We
xp2FrW7ju5d+B8eV3hM0CxeONRO6Ry/DdKj6A3aBwWrfeH4O5x4rPndJvzwdC56R
NdcheKS7wjsthKZM+5zOH7LGs3PjecU4yzci+h21BBnDztzQsvfHM5BTu7htSGh5
wXdDgoHQxlvuVSiD602MqKLKD2YeI2a3Tn6H3YF7lnW/4HiNRcuktBDZppv6zW7R
lBrTenL/9eVopyX9UmY+MCHogxLjMXNrJdqSkkFDL0RHIxZhS0HkgTcDTnbN0ZSR
lNVM67cFrDl7ePuOKLAfS2B9qcXQesp5nsl8QxF1su2AycRN8r+YkzUZYEeAN/98
HX29v+hoYOUeRItVmFFq/ahnDnewSpM50iINjy8Z0yrXg8olj9Tl2vlug9z9ED7B
dq5nZuPIvYFI5X9o7GUP2WEYw6wiQWdciOFR9MU1oEdm/ddN8iX1qBUiAqVUCTjH
OioN0gtW6wOcueMgpMgfFiPLQGsm4/SE77DFahnPM3xiJBioq9XvCIvZ3eDSWHyA
rJZQsCVd0qMtS/8NW2e+0w==
`protect END_PROTECTED
