`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5eNZ4AOB4A13lFqhEKzHEttTZQzjQG18HaUQHmnmFORIfCG20AE6nYnRAtUUyiDI
x6Pp9L3fpzW66DmjSR+CZTIfBFOEdzaOj6/J6m8YCsVkTuJpXcB0BDH+oVKPLYrt
uXmrIyhQc3KiXJz5xKD/3+RXZc/WMISfuAFwR5DawoMR+ShP1oC/fimB8WUvFdww
4ZO0m5EyifnfiVXUFOLFjX2Y4z74i0LIDH2I5MkJqyHHPtNNWJjMoHgatxs5yh6i
kzE4daR580WZgXoK7Ol6dmhVX0qWSPw/BsUnQkFTa21IbUu5gAB89fLnMKx11sTy
X5Xy/EAhuVhak5jydYYhEzAlyJmClkoa0gAri4fSXWQNsTv9b9S/tRonkgUFgwbI
I9Z1fG7nePZQdsaqo3f9xbvzYnNwGTNzAhGkYXsmjRBaghYodoPNqRA+jVNl6d7T
ysWsNvm5Hv8gCwyt7PFqLNdrAjJ9sKslyGZfePC1pM6t2HowatrfUsuFrY00Inke
E5hiWcKuZZuiWQ8E6XYh6ubgxFUVjwNgix025Z3JsqeJyCdNn1Gws7LE3B9k+7HY
5If2XLYnHMtLizPEZ7H1I/u38IrIktKL7F5vml/X6hGOH21Z3Zra53V5e8IwQ8f4
uJaNsCLc5wepikSlvD9CdZqhOuL+hNz9IDaAsiE5Fvd2xF5wglCFZUDCqXX1sbOM
idNcDbUvQ7zuww5+j2xUVw==
`protect END_PROTECTED
