`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qk9JxXEjQdYSVocz6KAkBjsrrBcN+BQtbR418yWr6Ra7BF3R5Q0X0Gw4RIraDiHp
8vEHEaDzXXdde76I6genDQsm7YPXf0rR658PPAODOOwoM0ApAwxTKEM6eCCaotea
4d0QwyvZG2JP468kAj/g/Z/mEMJwPUCY0JtG5SusBaMpUxFFXD21SEr4SnZt9la/
KiwWOEzhh3gvlXYKZENak1gHNI62u8qKZNCk0D2G62DDtS7uq0aGPicjTtJ9SjmY
JIfUQpEwfKMOxo9L+FiCiw==
`protect END_PROTECTED
