`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zLltEGWD7CmqV/p+uGdKv/JJauUE0xc1aTI0oSO43zIl881XjHtpUWgg2rdMEsYu
Y++52HS1nLoqkwaHmGT/5kjZY4ktRKDIvwVYv9McMDcP6o7eXLOrnl28URs1qtPn
cLjAP4tkeZZDSqW3/iLZ7AsMTJJSf5pzryQwpOxHNztd2tD6wuQq0wM/xcLZ0Bgk
jWdzzqrBn0Dv85PdikGxFVVXCU5n9n9A5Gee17Z5OQuU0soc9ayQzJIiviv3ss5b
YFZ8spb84bUtTrgZ3U3iBPyUisji9st98WJ5oLiLw0vJ/Lev7CaDY5y6aFAUmqei
K/AC6MWGdd0BiSNfkUeY8pYlhHZ03nQwrSx2mOiC7oK7jIkHMf72P6lZnmnFDL7/
t/I+hYc14iWmeJirgMXW5g/fncRgv9XDQLht2dZ25+QPFQ6GZVFwNbMl2ruRZsXj
7R+FcRwRW8Zjl3lOPmvS/Q==
`protect END_PROTECTED
