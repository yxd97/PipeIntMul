`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOlcTsTuk4u8TL+YTflHd1kYmHU4qzT/cHwAVzL9Pu51+ZYD4g18O2Wwk7avj5aD
QZ5zP2+7BAEf5ccKv0gSRXTWP7Z5l3+mPtS9GXI/jYxaLJrJEQJGUMRODuJTQeaC
gkaBFc50r7ZLOI7/lRFd/Qf2DlK+n0ELBLA3PeDsrqNK7x06FucAaGYhYYLT3psO
2ON3iMnldBgH6Eh2Vm5PdXXSjwgcXn+9xDa8/hql0lJFigkZ/3oEZZSni8rl7VGP
Dod487sD10bpF9yecjZ3jggXVCjSfc2huDgd+KxokuDOpzYbOWidyAVDYehkRSL/
dWjNWociVHp5IUSopzghtluj3AUuP1BNtpJPHZ2sYbrOWiYrYWFC4n8wC0/IdJsM
qeqK30bOzXYDszv7wtFfH7KJ4qgNnUlyOGaemDlXleSjPbV2aHn5aOKz4MBKm7cA
K03MrpI3VC2dwdkWmIdzZCo1zR0Mw9BFz3SD1tgdVAYSllWJBFv7IR3ZqbYjfFQA
BNbPul08XZxHdDQeeyYnQ/EnqR09cMGQZr0MCeSXSbl6S0lhC/5ilhGT5E/pctA1
Z8OzqmG0bms4y2aC7QV/qkWoeAj5WRNZxghd2m3wmCKKhQ/AqiSqBtk6ZqDxRCGo
ZyjziffhoMW7DqkslWhtIUipkTNMLMwkWpXzsi/64VMomsLec6akqvQkRlsV0n8M
aoxMUxgrUvMnuQLDjtpbTDSLfVFwfsG0XltWqzUV5KsPN05WUrx7dYUXlVOFuZF1
LaFBttjGMEZ12fIHGmXucp1JrDzanjE0Va3OMRWgPlLkfsnd+C44woZgj90HnmbH
thxIx7Pi9YcbMKkI4YU6jG/DgOrw0a1U7P2G4eZqDld1oNXCwCt0ObjO6YEO0nOF
7ycGdTfnTmGsDaXwqqlLxA==
`protect END_PROTECTED
