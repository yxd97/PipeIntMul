`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4nzAcrH/DE4OHWR4vYHI1VZ2m2piiPm7tQqdSNyphSBdwuVx7dFmCpPb62Hh8tP4
HGLsnUIyhXHpwE7RFVba73C75YAWMoibsGXxY8QE+l1JdCH+pgYr31Qmw3Tlg7Mu
8msBiW/eIL3MfAhbRHg4AMpUJ69FyD4NjlVOo1ue6DMdWeblCCYkB6hdOObSCMS5
I9kjicpbiavH+/+H7kkA7oM2/DPH7SwNs7tMVQ4hhdqfEWbbB+cd6UsoYnJFPYIt
+zzTU44MobOGOigJh95DzCDrTPt1YCSGNRZNJ8y3Kj9Tx6CgPrhM/Jt0RQU2pFST
7qnF7MBLe6utex/8fScTK/+v+b5GkH0nMMm6OQPg3Q37/IeDr+haZb9O1ogV4mCZ
OiSxp+w6niWksCAbftGNxKHG0Db/nsTb++QV7t+n0BNkfqqPDlfrWRPA7m+GLKT5
ZeEfCJsk93czt89rf1RbeVX6ZEEkKOIeYtkEkzDZmpWcQqYPRVMSYvTa2UdptgQ1
0E3Mszqs6VbOkteiFWcFdPkQgveMj0Ktjsm+HUE67HZyIztCA0AtzNS4ChUhvUKw
4XijBcmy25CXj9jn914mu2pGk9M8c6Zs4xgF5x0PRvPhQbTp2pUonOGwLPrLa9MG
L/6IvptkCVPfSEQr4GT322/rF2WLPWwS9Nr5V1RKhz2p3Tx9XkcnV3Rsx+kfT2rR
aw/p0i02G560G8jxOFS+pXIqBQyKa8gAulEiKrks5gQ=
`protect END_PROTECTED
