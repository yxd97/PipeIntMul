`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N/LtFppALoHdglFZh6P6c5s1i5eCY2qrZTydARRwSOn2Xm+/z/JM8Fq8wlP5C1iq
qQ35Ewk5D5kw3JwbApH/0/jUHZS7ocvINapiulPXg8aA6aPqcMSw921hnvtJkF2P
L2DydzPeE/s5wVGMRRebFnvdkQpo2dfKj+ykH1usvb55tyoSa6zzBYJZ6I57xY0F
FRjfKrKTX4SuPjj8XhzDBhXsK1bLAXp3t/gr+lhSKmdQXLpg4+0sC/GfCS9S88ew
lAXUmmnqSDELoUpIzHpi5ouM5pAphJmYLleVpZ1GmgMej37uPDmBP4jG4a3lTD+g
kfioBr/kLYfoyFQcAhuIVo16Ss5QIeRv99QeYvxXCinT3LcFW5C/xZkl/5zrD0be
jcn9m/+98O7PaTrxeAYVQCuf0j4BpjivdKwCwsDi2XsAGTSlCmgPWCWIEdpD9Jnv
wIxoZGelJHOcYlp4eeu+HmAOnYFWA/nF7Qqtd6l8bj4=
`protect END_PROTECTED
