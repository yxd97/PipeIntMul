`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4l4V/mEnJH8Mxe9kBRPzR6WN6qRKg2Ti0Fv3A9jkGmp1gkHeGadXB3YEW3l+scLl
7UB+raVYS3vp1Cjkl0Rkm+Pd8IedRcqju4Roxpe6QplRucSYB6lMmCaSCxtILdm0
i3Pk+j6zMEx4V6y2V4GHDLRUBSNvVBdO2nzZjpN2myhLKkcGhKFgV3wqDAJyoBkM
C4C86vznxUjrDZOA4ApWKUlOtap5Z0xeVX55QdG/G76sHLnHm7vcsIx0+CEd+3v5
l6fj8Sj+2z5Ss4Q0p2uXdt6GIL7kTjB/RLrwK4GAlnM=
`protect END_PROTECTED
