`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QoETEcU4prJIvPzpt0OX6lXPvb4EaB49kwLaewrBP0YORn5dw6dUhpavnV3NkQb5
wMwGYCjjgrBgekAjI3iz0Bo5XY4h/SSrngt3CqQBIQGqsWlSgMz5/VC8XYoXigVb
7gjfNXhFpSHHvcTxuW8Fw2DzJwuzVHR5APOz9xkEOAitDDs1LuieFakSf7FMoLuG
KvC9Qr9CeLDUE439QJ5GjSoE1mXpt41pHcoepvpY0/gW9Zw8pkr9D7kvIL7Punzw
rISZjqKgo0cRtn9sBNj9GyMxcPMDNZhOPWXHbgbQkHwdwBhwc8kcX2Zx5/hX6F/m
2CPwESK0H7sJn68P4+TWo4L4wpq1jzrm3wtGST3bNQSqsL+hXivKbuv8KxigdTqo
5v4/JqwiFUzIgJzqQ4YFEw2/N2Etc1ScDosECSSxMgENmRbhcVD6rF7hpIYuIqQX
G8Z94TlpXOmFAyve3xqGwcJR0CymvpPsRCr/nbF/KXqXpB4uBzcCqITFnUwIFJ2s
mqT84JqB2yQpVmD7UqbTzUuysUNUpS7G28hs85wvBCVnUGZJAK19cWY9Eku3dJ/9
lrxBc3m5kyLiLbkYF1wGAzbB0kEC4kGdfMT6yRiLdOyxXVfXk3FLnSrejZlB2MY9
xmvu4iQ8/vsflRC/tDKyiaY+p9KrxZ/GJqdrjL3UEgYzulomumZK3KuMtlUpyncd
rlYLtDkTTfBwmXYKbSGfibvurncgPKaeOTeF4z6UjfxFblPCtI8REj26prdbdTWf
Av/nn8irNrLqxmj6B3cUyvNwlzyjW2DS7694YdpRf82eHkk/a2hzFPuyCIljs2dH
84nfuYpRXinaSFf/O9Gw+aD9HvFOdcbvTN6Xmm4SsQO74uILLDnL01vZYaIwYzuH
MPLAnMDd4bxsbzugT4m3fF/LW2qxor+EgTaxTcY3euh3pIibhvhJad1o9tuS5nNp
Ry6X2Z74aMX1k8AXehL+tYSnvaVFdbTeLOYCsXUSl8XhRac2TmE++CktO5Os/Oi+
/qGO268NQh2a3a+j7o+1rQ==
`protect END_PROTECTED
