`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KtlYTNTO53v2posBdTVA2bh4fyDorDS8BDSEy52A9oiwoZ1fawvCcKP9aI3nafLv
7AIkdpPYoj2+innynaTv5ziCt2Rjjq3RC9pChQvtodLeII+1ao44FMYBMyovIYw6
CdX6bFT0NPzYJsaXZcX4PCwuX6ZZmMMPTNR/4hZJfL25pMthRNa73aGF60/DluDQ
w0eaYyQcWhO2ixpz/hJyz6iVTtE7kXSs4Gdw01sIxLvaXFeSemIQDPldAWiLQqJ8
XbficG1U2nQwlJg/LnKm6mYbJFj6kxfajt1U5WL3at4WrgvCf+p1y9nrN3l403PI
SIaJ+2/hllpBS3ywlXFhJhU6GHF+Kp1zOOHs6nRc4NYf5vPNwhoRbm3QNdssw/ba
BUBpr1lp+z/48pdd73eLTjjNhNhMi44i1apJ/vL++YTUaTP9iwWqUgBOniYKZUGC
K6Vpkxi3OthF7o7qfbgSIFSq71DMcX5kYNB7Hj6jajT19Z1wlyCRPvBBdXzvJb1v
o1LhrDOng2sBl+yF0ix8FPUuuvJG3hjR/JTH0VapFY981jVuu/1bG5feYWt8UybJ
9ru6A9l8cv5oWbqzbqvJyA==
`protect END_PROTECTED
