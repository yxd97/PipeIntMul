`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAnAamEoLiWyGe0UyYYpJ/IxhtSe3vyHwwoVvsDvb+92iZw0fUa+TXHf9b0u98nO
OOI+qGe1JA8xSOWjnq5aIm5AgB8bFYRmyTUv1MNhM9xl3lA1o3+v9m3ovgp3/YL/
a4Gy4loYokDbw567JP6dPvusRTVhJSMwq4Z5oRFr5UNlDW8+57/FvFKooz77oHnP
fOGENoRUS3lvZKYwAGRcODqMfgiVZu8gKjj3/YrCSqyV3QZNihM4c97Y+B2ln8JM
QXSbDjZVP+8fjqdR+nTahzYnF+TK31lj2/ozZ3PRZTmcHn11le1BdTnzG8CXzHbg
nM4rjgpe6U1tZVGBA4LFlwASPhnhgyi36LaT9y4KLCMPtBc+QhkExL/1C2O4dmpv
E9PE3LB308/KvfQwn7oTEQliwcN6d7J/BNNTVot2h+Li9iC2+YMre1CU0YvW7Qq1
mx9eQiTlEkIMuif4m6d1UrZRzOPYqvXdMcRWUpjVfnmmW2N7X9SCvNsP4dChbksM
0RGCZJtn7Sc3l0xF4e2P2wHCrmP4h9mbZyjTVoSlvXFu1niAySd+Dxl4ubLl/NeX
ShuntXEsxnM1xAJh268+7LUaCE5c+f9to/jS/VKtNRqexEeQPvsALb931/G4V0UA
mH48rHZrK3EIVWgN+8yTVek3n1/XVEItEfUOjzM3wIp/S4Irv46O5eaU3bjCspF0
q/6aWyNOX43VzUga9u6w7/zlABLpW2s3DLFFhTZZ/jO71u5Bjn0beTPu4woUesxz
2MNO/Cyu9x1w3Z+DGWLF/S+lXdtmjpUP48lPHJ2pJbEDO5QMdaw/TdWOPb4JRHYY
ecP0G/RQuxHOQMPvC0EOrS52qwAkt7w3N42TWmAewjt3mOKDy858l0rfy3tGEC5C
V+wiZWZfvBBj8WJNQdx2/65kz2jzHRTwv9iIfTXd4pvuGx691rIRLcbNWbFwZjv3
bZKyHnOlzM5nyd/l12/FDnW3QwxiO7WJ1hjsMHa51WZiRnsWZrlSCTBJVG9NbMxX
uCZq28GkMWBVHBLN8KLBvAs0NfjaYLMlE27l/RwjOCtXhLQwZbiViKVyWvJRoyQG
pzxpbV881nttXj50BpS6X7SHv9jSqv3myKC1u991ZCfxE4UoEf6urMDtGdQGwlOt
DaYJCUCgjjDSiv1hfS8AdEFMa79u64cEhd7JxAEWDAheFrlc/JXgMi2W4JcDWTzs
F0rRWa4LquqaGr+l3wQ2HhBHjFr0kyZkY71qL7lfHYBCztnYf1Sm/1Tf7mKS8VxV
0o1HMt7qYRvcPEZq+CpI3yLgWKfSsrMlZCmJ7hzpZWj9N3/WWcK6NG3r604SoAoj
IuwSO10NkhzcDrtZufU4dvjP8ImfQFRsgdU2YuqAfRrxkqIvlagA9rpRtBEVAGHs
g458UfwgYcwNfSnmM7xTFi7E7rxpBSMMtt5mXvfkCjF9tHtlJuQUsBoameweBjjB
byNe/RnWKHkJ0reyHaQbiFdxFqQFV5UXENUZno7JgAkI+KNngvrV0Yi8lroSD3S+
aFKtnhlzus266VCIF9QiBAKLKG7UMw8bBRN7IoXPKHk4uDp/kG7gSye1CgwnrMM+
0TIR5vGPNSJQE2xy5uymbofDeRaLIKIvKkaFVvBkW4edmKC4wF7tYnVCCiUhjAkK
ZpPToeCVJFpPo2V/7wwW1DkzS26LaWdy2IG7NuoIf4nBdvJlADmUy9IMdOkU+dUN
6ZCrKRc+Du+80fB6/oo32XB8GrUD0ZdTqVrMItnzmMlMzyMuDDRAG3P1zsO9pSrI
clv4zSV+471B4Jb39lipnV6FFyY7/RZOw66VmpboTpv4CBNotlSMJzc14JsALEvE
IsVRqk+hj2ZJZRAiTeQqxKf1271iaVroNjdoXL4v8bMvmglO33aRcK/CHpMFu+1z
gQrU8hxJ6/drBc9dpFYr8C5SchzYqF29viKqyOUy8Zv7xp24XbcsQp5wFdDMf2pK
bqkwgAr+vGQUa/poSPxzQG95Vq3gOWofmudzvlFZFfy0JRcVvD0NKcA3qr4cM6Uv
rUmcAWP2/H1fe9hsa4pQE46WBBO81MzjDeIR0n7bNzMrf9HGSkm3QY2BP7BoArci
zvnPiiYxJCIphjSBCPApMosL1s3zDeZYuEWgmS8XpaFisrjhcxECwvVYWJRvvwLl
a7TDAno+oGq4gCnl7TUHgc6952UatpB3AzWxAoxJPuJbIgZ6HEZ93C+ue4zQf5Ud
wSqXwXTMCco1JIhg7PgUyMZRidWfQ1DQOttmdWl9hlIPWTnEy88gPLIFR9/JZOhp
bXIGMtd21ERrhg0HJIKKPS1598ddFhxxgm3Ia4WC4CH2MSg8gXoMXe27C/maBc1B
g5fTZxmkVRFc2DGBOBWTJB2w6GSCtVJ1ww9EHOHk6+z3D3772sJvmq/l9B7k3BBJ
uzLiZPABDeFxbliLpn/LcpvOqC50IhykBM6vzOlqnhPOItTWOaGIy/nMfCEE32Qm
GNsy1ARvh0VdQ4mBsdH40PQyYXW0k+B2vxFYpwIlrdCmA/kXzXVdAaXWhEbaAHR8
QA+44JOQx8r6spb04HuDXtdJcXtqsdiJRl2yS8qCer+qVN8E6e1sKM+C/AB/CJl9
UDZjvFCiVOLEWtvMSluyWzzUy6Ppi3+D7bKMTIpTP7Jw2AueJsiF2d3KRgyw8JaK
1g6ydvZwAJ2WM/DvT+oe4N5igikqfDsqiHnlaPOFMI6PAb8zGyFki4lChmnutJGL
UM4rGwkKAzsT4QvCPpHs3l6Lw8rz6GIllYfUKQCh5A9uoijcd6vLbS6d/lji9ecx
P1KUPN07KguzIEHMbeGA6AAYzFQ3qYdRZ3wua02/TXRH7rKFUHi9eH2jdjq/5+VN
4TQsWkKinZB87a4HoGTyUgd32AhdXdCXaZSEZObt9Qp8ErGKsrd3GguyDzHkvTaB
Y7E/ZYgg1zYdAJ+8ZwQ2Usm+Q505NQOVLdpGkokszNBYgDzKGwqXOLLG1z0VMPWv
nMh/BIUjlTIjhfZHA5pHwM4/B0AI1ybNOG2kAbPAFcdB+qjIxv4OjzVSmXwj4n5W
0UgeMFzeFmjuPGy5kOZTXTIL6G0nMk2kKU9MUzrXqBAhtNTZHvWBbJyQpuwfWHLl
DDycm+6OKY6gFNF+Jk2pk6z4hfXz5zrDgSfg/rKQDmWs2PBV5UFJYLtpkBpb3+wj
vaRhPw5/BN6evbX8HHfIi1pDvZR3aicgeJFaTu58F6QPVUoFSr8fwFEFPooT8u2X
yX/1NndfrS0BzCRjpizjTgShzc3kpK/Qg+UVPpMipxq+QXnrAqVN8m+e6bdtdNn8
AFSCn/+EmGgfFmIZagl9KqeXNixu5Iz7Pr/mrKUm99RdKnsWxdJX/h7RcEng2/Ad
qtk9bM52UK+NSnLIRAWeaAc3RipueLs0ICosVZX78Jtp43lpC4dX+I3Fo/VGjLQd
NJjAnB/57ClrbrySxdDxuYzmWnr+5QHBAFodvO8HkUBtUsh5kTRsu5nf1b8myIU1
5BdSepxvLZoDDkODCCVV73R6aLsVJ7ZiiYfYUCkeFXgW3VISibiaiDWCADB1TG5v
De/I0/YWqM0X/jyP3GziXo6IVKln1Mrv6BSXVRQeYnPCHe7S+pNzkLtzA3O6pMZU
3+btQh/3sFKdgSwK3PC873RKYvl/6jD7YTeOMEN++qWxXZkQh3aOD1wPte5yt3/t
SgN7op8gND7JYTMcjVdWILIAox2I1Kf4YWiF3QYP6Y2f4IlYSpBlU243b/tqd8gp
5arJp8mwUSM7rt5fFHmXgItxrx6i+cWdNrPQAF/zl0j/XhlXOiKbLIniCZ/fqZhU
+TSCrUYSb06BwmUw4FpgjvvJARcSo+yfSzueNJ2PzaEAQCMVBoDvk3w76ywoCDoG
aIFlHWDxLKL2cdBfrJs6ofAYu+YjUcxgfaK1gRaR7ycEQ7z8tuDwHXK843YKwlOs
PeoXoUW+w7dfADex1RNTse6LyLHBSpU8MsXTKXajvCI3aR9sb38CvYFF28vwSzHh
V05ClOb2J9DX+Wkl5wginihtuVyTmUIOZl9NcX6sT+BjaqfBu7vkDoeV/BNYTqRO
Ll0hv1iTsgnRNXVhG23iBClpfyU5Njbn2rF8p98T70haPGsFhDA5OmNwI+4KVcho
`protect END_PROTECTED
