`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9dXhcelsus7LGLCGvqXeN6DIBZrSWCsrTEoNEL/m5LOx72daysNQ35fzFh6e0fuQ
akAT/7WILUEZGwNGdU+1bssVn8sOs/r6xhhjFOZIjl9oC+LWHdZfOWfWhQXp8/wc
J1ps4Dhdjdgv3l3Y66yhzsGsukFPnQczhfFSborQA9GrpKwzVJ4ZFtirc5ZrkJfA
MBOArLmmU9L5V38RcmHaMxSYEG7peOp9dIPH77E0/IPliHPYwdbRKL14FWXlzsrW
Dcko6aES/pCP4nhLgHpRrh73ZHNmJnt/rHza3TL4slDpJItSe6CsoyO2SUIx53jJ
IBBdJ0ny+GQ0GzBXm5y3QKeh7atzl619f6YrE4VVCPWzS9yvbV2Z6RiXZfV4tp2z
mIOhksUeWAY5uJlvKUoOgB9UHUc0RybQw272pFXQhAs=
`protect END_PROTECTED
