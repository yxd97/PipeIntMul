`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v65ISvLfXn5WiKFwyl5MfEt/OAj3rAV8fBONo9Egp+8OGfm6n79MveDWxPV5EEqC
7mLAKfm6JeFmj3K5KkuYK7E/UZ6xERYJMGMToGPTf3LRZIE/liPbtVSKJJzwC6bO
2ZlasYxY7XEjgK0uVeVeOgq9Wqqdjnyg0u9MYXZmL+X2jzvajya4lzqdeNW1NM5h
l4j16BNXRsz8ghUY6avFu7LBHHMWKsLBW4PKv5DkzeLPKilJAtEM4eFEhFK4Tlqw
iEe7A5U4Uir62FA2EgicuNJZ1FPBFvb00SICzMK59aMvWGXEBWAhX9DH0PCjzljP
8hXPRDZE/3Yn+n9MmVUYouk/oeqPUzMYyWZuvELbBv7HMeSCUJXjPNymWtJW7ZFI
8tpy2KwYxPxFMqPhl49UIQx8MENYBwhSpUbzOyZGGAYd9J6zbJ6nY9WZT42GCwgs
5XPLihlFSDI2PLo50lPv6bw+UldpPPrbehX0oekvcCvSGE+gSK/PndzyZqy5cY8L
JjFlDPR/B4eQwnG5zzSGbULQGoH7+7B13bjVnJ/goxKqmdAwQ9jJxCIbIlpom3jV
BBSaZckrwlaSQLw9D1aeOFvMu899MWt7J9xLe+TllhE=
`protect END_PROTECTED
