`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DOW/UL5vpjM2HCKoGNZLYMmOyzcl7cNqKpFaNel36sAl+W/l9kACB5shhIqfBcRV
GUO1IkE5gEByNBPjywU7f8AqRQ8FmtrQ1gmdAjW0yraVo/UFaiu9bgnX8QP1Qfrb
oXOt5/Dr9KyUZjCRQIasdGcAbiUWP38yDdAMKJKIOfNum9ETwa9/Zw99o+0T7Ytn
gEeGUSvRC3v5bFfM2vHcxfPv1ji+TWq2UXNdogRidSpSuJ/vjqysiFvhaX8h7g0H
JMDi3UVobS81mgS1BjEB/KmRnDxMvp4Mr8kECKM4YXDmbKd3G1TBm03TrPkq/Q06
qPXCV1XWljq5rgrZDjmbYA5GYmTzc5XJIzCPNW7B2HqLmwABQax9Tu8pqWjNRhf/
4bqx1tI+Yaa0yK9HyAnNQvt9ugTDMKmEx9SQzgWM3gHrDxkvWBxP9jspoUaCTEJL
FfZ3HvQzreJ0DKhzNXaxzfAPtYCc7sNctBJMqLkhvdgINUA+g29jaqzwubYzswjz
RuotgK0TWRQpyGMERZxXAlvtpUnCGCafr4P1FatMobPRcCzLBMbn7ST+x4igh8L0
`protect END_PROTECTED
