`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpIhYHQFy7+p5XW/42KfZ1XBRYPewv+llHsDxJsy6cTupVW50+a7jECsutzJXRr8
2A6DD46OfHp98+fdv44s8lLb0rI9myGh9TuDSBYzXts8iEdhaibGB0K0P9XBfjlo
aL7yTxIKfLJOg78htqZo+au4F9dSdsOHC5lxfaeXpTBiLV4naqg+SiC6IoPXMxAs
Od/YTkKU4nJTHif9QuITunxaiqAWWJLHKmpwET0VVUyqxLN42lKFpT5VIZW+zL3i
o8K4MepXqPuDWY1j0HcuqUHD49iN8acjef6QV8y7zVcssOLsDF3oktt7dBXuEGyB
i3wabm5tSWIIVOV2rpl/87/IVqkQxsbDvFsZcIclkf+mExkKvFElFWKEzho8Oi3G
+Pf92/q7XWJ6C2zBI4O7gwHKSvCml8fzP5HR3GeKixUzKAGMD4ttWgmQK0U+nBw/
ZEE1xaDrqeKk8EkMtZb82QuUUBnoO0MVWziT2vTqTO+v59DZ156DWHOy6EI3pqKn
TKoSww/rVSi0k2hd2YMqJ2bxp7WfpKbfZsohojDwazvDlvGkCtTA7l348q9eURLe
xY9J3CcUKjQ0HxdC0rExBBLeAiHogBYR8d4dhg/aOsYr7wBsbGnITCYT4Ouj0v6r
34BBmPLrweLnqLeKaYHP3haH1hIDXnLIlMIxeunamuiDJOijMpAKewDnj21yeJvU
y1p+TdJlvohfQnUPbL9i7+N1CJ4WTnC+kUhUt6czhdbEzf+GLaWPwixd9knyuHQP
dwgXfcYSYhgZI0ecxaAeN0/KF4lgHZIVIygXIARZR2UN+oc23TeyA20PKvYmf8OC
pFcr916i8XpQu9kFRX2+iFSEdF2rR5IuST8waO6F14YbBzxq0HyMMC72BH22Ophh
ezCedHDMgSDCYwFmMm6KSVa7MYjzhmzh0QeVkOYlU4zPu14xZP2+cl2no5KHlakQ
91ZwR+YW9n/kORguJ10lgr5wih8ilsqfpQya93gvRWYFCpxnEYVcEY4PMohysz7z
7ricBID2pymZ8iC6IWfcQinL22oSW2EGjFbun/nP/O7NddFzoom6j23GrvVfaAU8
zDfFc57WQkqU7Dr0ERTSMZHviLZFSTsnQJ822fYWccDf1Hg9CV1oxpp/zymTB5gk
/acDI0bQANJAtNeEYQM46cdkNDl3/e/2JMaHVgCT5u6ch99SBewtXoy95FODI30Y
EZZsEJTyNjnUUKB+wIu6Pg8J1A13eFOErP6K4Tv9GyiC1ZzqzpwUiIsjdkyaJ163
gL6KJ9YMFUzrq3sCMdfadp8v0gv7XlpQxmI7DcS0TW1qa6jahmiiEkdsOGMA6Hc+
RxmoxISoZNGxp45he7x+YW8ioo7KQyADXiXgbmDPvvBSiNcEQUYyjxVmD1BpvTEl
8w3FjYVKN2mPZXLM2PtQ0hqTPd5cHmxX7njKa+QeVNtB7fLIPWrjX77z3ki62o/8
tdhZbs6W5+3JuJ6W3/iLwDNfJmYSjeKOC7EGt99tDaWQ2QmGOcgMjEGHDjOqw6wM
4SGWUWo4gkRoblB953wrZSSscF+hJmNFqFw4GC4jR3185+WvIuBycUeRfBJ2Kehx
a6WMjuXBKx2Fobx8OSRkWT7Yauf/BrJsUwNLk74PzULXTqbHMp+pnOznTa7eAM/s
BA9/2wimgOUytgaNWnpbo5DATEMxHgSKDvuaGUAYQc20FbB10GC24x77Ne797hm+
wsgy+L6e6xH2tIZui8nS/KqsVX0E0AXjR4mAqk9F5GMGwrRaz5JZkdCk3rkvYMpu
K68W1COhCpYMchPAJmSjr0zTV7u14+16XMp/Ok3vKWWZeWWK96xlzzD6YBDtn9aY
xRG8Ax7nfzNQZoWSzrylfLbAuxh6jyhICIioQFNJpmzI9GoK3MAmjHYkOpsFLNx5
TUGJyBSaTU//ZH5v5T/fvhgAtg3qPwgfdZ6/K8at1a0Oum+qn/wpEM396yI1OIZF
YhyxUiSvBbrXMcVkaKgW1TszXNErfCpxR7Nizv33lAa/DwcJjKN+I7p2emV+UkLY
bDxJeqxzhI0h9shnEzXXV3qVz0Qc0huH51gUHSeL6G7VGG8q0tfJNS8ero/RKtLg
av49qL9v1EjQ44OKnJhC/EsRhlNz+FS6u9VqLUwz3bl3LX3uaxtcIATCWkM96sUr
n3oVgB20P8wlKFOFec2zlCA/3oEFkCygC0HNG/wrQDYWc4uG2F7HS6uUq5boxW6O
kNh3COoPJ88JoactCvRMAcJcy3UEFARYEf+RP5mfVzKtPBEfamgcoUXlgjs9vYIn
ncRx0IY45YCc66+chQn0E0v1uPzqI+kdNWigNjpY0hXq14xvCnKOzupTTjCGHC7C
bivPT6rqkvIEsJrWYl3d0tG5vZgUoqBBSBgD3VdDzqTWbM+Esc7JUdXABARM/8HA
xEg7OiRTBksxdoquALmOsA0MaluB87vQdYiQSL3SJIiBL4donFAB0/9jTxcXP1X2
BFdO5QFSUSjAsIYjOFN6Z6hC2rlcshkozBQqQUOHq5JBGFLxnB+kDuucqhpVh1UB
Wb4WySrSWiEQpB59T7EYAM+x5aYNRuutozALIQpLlV8N+iLTuT/5cD40QZQWLH0c
afVWf6paVRTfgWyAdlzUSg==
`protect END_PROTECTED
