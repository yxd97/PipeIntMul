`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SXmmxTC4p2iRn5KUoWC1mk1GMpvxgkYKeJ3K0l0VCqOEfq+ta8noUHA18jmYP7qB
GDYNl4F6QTXr+3cUq/ZaqvY0LwlU5VvPcO3a/3ZAlbTOKPshnwMH4MBAd10Xkzv6
WmXEWF1Cf243psZ8rr8kOB2HrSVQX+vkvKBiSVe+pVUO8cSStkhiIbfF9+2rWC5U
HIx7rMeOGQhCUqf0b8thy5nMP7hdoeiKfQ95Irj5lDOC2orvwVPs6Bevdp68sAO6
41jNtYsAirmssIRWR/fRdMmVd4S0opL0T8KYPOEzEnQi66y3GA0rU9AOTrGXumbU
3fGbTBd5rvxgQFY7VX5kHTPe37KSHKOB9ieTrmCBdIvGNypKYTKMf4uSKPUo7FeN
mhFUEbu5zrE0/c+4SLs2lC08GlcUs6eZ0kTmML4rw72ljDvKbimqLFcwiL4KJka9
3jwTlR1AeQGfkxOcseIy/Owhl+SnbzzNQcJ+1ubaCn8FzWxmgYKnlOuQZHqopI9P
pj1JOGQYqcPqduGxdxGCKbODg52+AGGei5tk1DJd77dop1ilmD7CMbSyJK+oTNvX
tV3RaOo8cBDb228Z97GkbQEuU9EV7eTFNFMah688GYZ1L2srN53F0VruPoQw/Z7V
Q28mdLI8n5/IlxVyvx1XXA==
`protect END_PROTECTED
