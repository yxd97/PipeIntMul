`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YHEIKY4B8hq9CFnq7xkauwVvQevSP9pptiAy+D0VvmTz6fIqCQzY4chvYGfHMqMC
/zNL12o0HzE8umOxgqRDd4/tlAKofOXv0M4wrDPXCTWHn2WXrJmtbQ+WB55/yPF8
TeIRflJY/agd6sUje1JiiNn8jjmz+f9/KGsnMDRu00W2XiYNdvlBURbir+oELeh3
RlcgHctJS13ALzA1QpCZdUsE6Exjwrg3fkEEZo7X7zd7jcOP00woSuwmF+yk/i4O
wfZvy+jt3xSTkjbm+ZlpVBH6e8EXrsvt++LxjKJTNVzC/Qt9pCYIQEHAag5nWg+F
aJBidzjmavRXNhNxrAT+OkrMse94DoSxcHzgpOprJYQlAyQRY+EVcrpKE+g6zZdd
0a2NMun59ly+dex8S20LJ6AuWhzwgFOnlHlmvtt1pRHgX4UDOb4gWD3b9TX86GJK
ngNVmZ4OxkAKedqpmPxvQ+9CMwOP6vQ8gOt8DuMauO4zVGMoJ9MSZEFJ+ihC/iq8
A+4rhBOcXywtTKUdTFVt5JG+Eg2BolWPW1N8tYdxQJd8IbHnQj9tZgChN5v9Auqr
tk0Xb9oT6LZhzDcjT65FUCSugvcqzQmnBjv6aWJxqSrA09UpDrY/C7W4UBuOSxij
gtgDlBD2ZkKz5/wX/xoPmZlTwEPnhd8u2/ZHWDpkNMbIdRaAC6roivxxeCSKXWZq
QrY5NsA3x1Cqvjol0ERR+gfYxntAZ+Vkwtp0bDoHuYDw9RUlQ40koOlh9e3kiVf9
rXRtFMa+0inpWnE+1+x8/uNZTymU8aZNo1/qnEuRHuX/c4BZ7gRnn50cnSm6TBsn
tseLbphXHOEdaa7j4k2MBzwu7o2i/eEXmrpLm383z1+qwasQB26b1LL+RcVRbrRG
FWjWzGbqn2Ul+S0cUn+KwWlNfLgOjeLo5oK0U8wGO/dd9q4227YiAEV8PReurrLh
3xiG959Nc7ekXBgEC3HDI8+kGRi2VHYFTpdFSJe8FfUWqWHpkmsInvFy97HBjGV8
ai61s58gFC6faBpRN8dWorUnb+SuRAELItAi5n8qU+IztIuYl8/J8/n23Y3j4VUR
M4Y2sapVmapt2tfM8lDRJTqCuRkRXcke5EoEZmkCBkSELD09e8j1B6MTLSOP/mdh
iK4qHdbn4fIhEraZrIub/mx96ndZLYCICGOuhZaekXC7BGDF4b9M+O14UgNrzKjB
nW8XJ+hg4oj0XC4yd9uDZ0X+pIru+stcSR30SA+hVxnHMvZ4e6SNFXE1IaIDMPJG
I9MW8TycbBGETTF2Bi7wcawqkIe8bFO7wwxiK+SpyREIqmRpO4l0hKxG8+NxzzjI
vPXy+DoOuDfIAiP8inYp4UXm+jSy0TClcQjmonMPEKzOJ1+vNM0zaoV2q0kFTgae
d7eiXlSIDLm2EMnE9wnGnMVX8Q9in6ASLKgOx+DPQ6OEIDcvxZjtHhtc+x2c9lW5
4SQCmrwIYkdwq3HeN8LLFZGXd3zyXB3c160fLCKF1wlYKTWkGTsNr1Ml4ATs6M23
z2fyBAA0jPP30rk4SW9PFqw46ypq/O0tYZS/ILuhV4eI8wUkclgiN6pwJlLTrYj2
bspm/aczHYfJuMjo0so0bfHw+dv6Qv+RcY0RFLU/3TK73M2Jd033+kZJ+JhdDeZx
YV10aV/rbtSPJrCZYLq7sTOQgeNpxrthf5PvMHUEs4uCbwZ0rqapEJGbcKRXb+AC
PZsp/Ov1xqWk27v73tlTpGhnfaAvRGA2g7PaCtV/RIoGLHMPy8bd43n7PBblxggf
OGnGb5ZgZgUCbkxR/2bSZ0A8A67wJBBMXxcCR6ck7ZEEDxROhyDfpePfxzjPRY7j
KIB2KHTg9w12gDyVypasbaEPZZtg0A5cR26cgO6P+6JLwNogMczXqV+iXdQXxTvx
uifV6R13Bo0dSx+O/yyuZEmyTCf6p6iz0HM6qF/QbEUNwYlLgJwabFLk5PNRudFx
zuTRZ0BZIR4dAiHr+oscH7PqOgirrF9vjt6ZKguj5UIfqhYWJo71MNaGzy859Je4
b2Aj+oeZFb2DnDeYKT9P8fU2PoloSjmL4Sej07zvLqziicvOOJX7fD2t1w84CKyL
c8MpgtnaaYHCybWLvtm+rl+dC+hgcVlFG29H35jmrs1FoGHcvEHnzfmBYJ9N+Ipo
xuylumav6L0UnQiTRGMLlwROMtL/dojSvDJ/CM2Ykc4IspQXvno/I5KwI49+pr/x
Pb+rGQSIh9y4H6h+c6kHEKPUU8SQ1d9pD/d+vaxeIiwYVs6gmKLy0ozYxLc+PBS8
3MjIBebPQQBYBr7QyIvTUSJ8aDunWdTn8c+ydBv6LVYBxfkDpQmRGK+0foPPTv/2
6BK25YEAxJxjKJh4Qp7w9hxSCgtPSoYQmHeWszmSO8YwzlO6NC5eJn6fWwtw7aMu
rUYBJs7VcGwnVh9f3dCZzTfa6pcq3jyZPCDqgU+I1EBFd9VjyAqYuua9OsIk/BFE
yxnY/OebhqIfQUMZhA+c+nZ5Y4a5n00rjlaPJeH8gnl8fiJ321fpGfYmvQJoAcGO
z+OLDoV/Xcr94Qy13EJIycLWtRBJfUpl5USjUMrPTk4FuvNkmgtL0t2xOEDp3d2c
VYtM/40rP52MGRxvQLaPMZOyifx2GRaZO/4kt11Ei3ln6Kb0Je5SMWKqzl/Tyskj
glbIg4blie3wfH7O78H24DzXQFG1tAf376OA6jb94Rm8J16mu+k4jhJZoCJmTtJT
YrIs/K3EsQBgx0FOD+O31siGSf92sfTiZNMS1SJolF8JQtiDNuJPtOOx9+J5fjig
jgHDsN9hxXqJh9MCWJYG8mh0xE7px6SfbHuvNJGrbt7NAB26UfsKQkMsPAReDMPF
M54T6GtEEco7Ttw6QjA0RUpBQvLeEf1TZtu5w4h9/9NIMjP12BNVQY5YLV5py3kD
mviPIDsRBlYzQGm/6FHWwggZ4Rl52AhFo3eToMI7d0OOSHrDpsLX8wwWwQWCptH0
Zfub4/OHMG5B1G6MV7CxB49xnKk7pBKCsRprCGTSg79JZZn3DrXmU2FSlnJPVP+y
BMppfDSstL4142thMC+dDb6PMD83HSQsrlxC9wac0/VJ+BRABN2EvLEoXyWPdedl
h3rfIFfaHMiCsKHPESrBHJYyafsfo/plDen65S0pm9GBNpCw/1O/9koY/YzQH6ZR
f/IWjxQ4/IWYFiiHaun460bf12ROUTEix3mUoGH26NhgZSx4O7gqLLOG37nJVqha
G1MERcwmywb+PrA8NtjAU8b1ca+zcH8eflZJlVpsm6llFMaYJgvsMEzpFUmuCWXN
Hiu/aTjK3K1Ac8HWPj419oGFngjhvbmVEnchi+6Kiaxouedl1/NDXRc7T/iYGvrU
/a4fduKKL7tUUd4sUDx7mx6izJUlGp7WVr4vCOxHk/70iS/uAmMmNQG8/sNZ2Wz4
aUhrX4C22P14yFVC+lLGjfu3boVMAlu95iOu7dyCN9IcAfV0SQbYd3PrBWOrVIHR
uFYjdTCUlCO+bK5l4jC2WU9vSOpigeLOKP636cmZ41jqeCPbw5yUyBbizJOQnIcY
vqMG/041GP/JsmNHE6LytXU+iFhsNkWw2itJ/OnGVXCnhF9VYsS2v57H7dFoD94L
P9Cl5JoFnudtWUNsX86tym32xKrpVuzRVE2dMns8i0TqNnLYzZuusb8c7QSzDlfz
7MVRxeLz6PsGE/am1fUbBpnuSnZnZtTYpRFrfhiE2Vumyr7nP1+bAyx1R5+sJQfa
/YcaAbNuWPjTegj04vuSSyK2ST8+uAo/lB8GPsPFleCoS2B7/oPNDVevoJB91TqQ
CP5i8iiNdSk10XKlf6Nzgij3D/OkG8no/wpzEgD5jlB7eFMMF5JIJqIGeYBLRkjA
3Tr96qynEcruOZ3LKgeL8MIBZKjUpWXWpHSxn9HRXXgzr5XvZnNHfzYiM3Ua0YbK
7+NMqrWJeRH1XSRRbRi9TRKqwGRGEjJSIAvi4UtJeDFJGkfIPhhhkOrvHuKHEDzF
07sHFHX5kEXuSvDbzSJe1eJIljKLs08lfaevDihhgLWTqhp/Tj8c3u010SL6vh9D
aQBu9y6h+prjf9VD3vHRHy/gSRZRlJeTFw0d7qsk0PrZFeQ0sKOGtB0w0nzNjZWh
CDQj8pmYbscATdDR4rDubB4ye13VVhfLSJxgr14Sx9bRb65L9CEB+uQYTkW3SaQL
Rm6hvgUIvRdnCcKaAlh/xjOvlOQQbEKlorqoVUV1jRUeHdyjeDp/JTz+QPUgGLyF
gDNHYm3ssw7gJJaMhhDg8daEBwsYlTYTMjr65HS1VPGPsTDuWBWHwy+XnvxALXCG
LeLOfWM1SeyKIAsnL4pjpckJp5TV4kZiziyLu95A3u9YibNyflo8O41URRQ21vju
ma8VWO8GqnbDXHvL3flkg3YF6wGpcd2/VFPTwRh+JVGRK172b9pcaEvF++R504v0
cSbVLxpMfej/l19imXMPeJP3xeZ+3XHZaf1/ZGYT1lQqwmK2d+Hdymoo8H6GB51k
5cquG9bP5lpj28Fdu3CsGgUV0n5959vm6GPRKsKLVKxTga5biKhBgdDtYams+kCi
phfcUwGaFb3XwqtI0FhQrA4bVvTMO9JAIg5sWa/GiIQxXVoZ2s+JlLw1SKX617RU
Z4dXS0bvqOdrHs7SfM1MxCPWP7w4i7msEuB7NMLrWnxeMSZLNnyjWo6PTQAkmu1c
K5WUx/ESSNhCssmXIEgboJSLDiuOzIkXIRtPWZ0zK78JhzLLjlNC0HEhxhn7D0oo
CWXJqBZTZKo42HDMs+krGoD0WPCFgWspT24TeOalT74x5h4coOYPKrc8XgKq6GOq
bRUtBTwQRVpl6ZSwnA/GZGIAcXYLxCt+hBysBU3wSCsNXsIslbdmrLf0ivmla0vG
lSTOoxRl3w9BZsX/Gq90qfTAJVjSsTE6Kd6+3oyn5wIfB/TyWljeUMQMfq+FmEBR
TBRDiZx8J552QK2CAvj7W888Jc3vIZREz4UV0MduZGEz3dmrpKgImM5PAP0OhUws
1afOP83hY8XTJ+aIUw7NjhoAEbOnPq+Kz8oblCIg2s1B1nKU8Ba8jORCh5WS23nL
pade8edghzblNmDYEDhCuJYPaleeiaWobR2Luu5jCSHXue7Bv/gU0lzZAolrhcTj
vNi51bjBgcN0UfGGUG/yt/pi8cuWSeP1SVqMIuz8X402clEzmHMv6hTdpAaLbPg1
sLAJA4948fj6DOHEG3NwrXNfl1go1HrWbvdEnlPOUYLSPSPUZlzzQHTl/5nRlz5h
NCwY4cqZNyfu1MzinLJMy82R/Y0beFxrBG5YX6AMKQy1mVKfCxsrf53Gw/7MnEgq
9fmwbttKbn517vkCxXkkG4/z/HGZ/6LCCZ5D/Vmy9NAbnBK3bkaWZhenlai0e1aJ
KNg+bubPVczJwQfGDMiaQwpKhUaidOUylE7d9Y+POu3ysY8CbYItehkIt5m3zZAL
+2bMeb5n+SzvgyVdGLR3L99ECancQYIp+sTUdaSTqxVhlQsDoVVb/NRF2KD/Q3L1
di0MjxYf/l4FRkt/0nDf2Cbx8hHLvd+05Cth/t76azhhI7n3WYwgHbZLZ6nBmJzU
wu3R/YwZlbrucr4DlAaTX6HEjN3x+6sm6kUQBMkblTXbv3N0uaXUXJjjjXspzDsM
kS0AzuaWfwV+/qvWNd/gtIdtNazbiBTUr+hsxRs8K6jfGxqHyQtjgPh8ihyw3xDU
3gLIVtuK+T79F6I9IV4EKj/ZDL5EDLsNRiHGCjD8B2Lz0TeoUPt6ia1bGiqpcpZl
T3dkDwQCHChaSgVM908Gs6oEFUz59X3MH4TcyLRa9N3rnfcoC6LeHgzkIV5thr5n
zgiKcdSRBva+UXZSaWoYYfo7+kn+yxv/A2UFJJWtcQjxZJ5hQh2bBS6x9V9CZcSN
CNZBM9VoQAy00YLJN71UlVgtmkE8iJMemIt4Rx66JRhp2poBcxKosGwf1iN7BYAE
OKRHnw/go50wJUcuswlz+ucXT/RIEp4/WpUnfnV3Qy5qrLHCrQ+ojNEzmWVMAqRN
cn+NAC8zKt73lUgBQlG9DFG+P4HLm759ayyUDRUibYJ/i9ChRhNYpBSH91AqH0BX
ZbnGDFNnrI4IWlZ6AsX8SjKp17/YBO6j5DMcPb0kvkk5LN2DbxqXyTYC+x3RT7/0
4XwDK+dvRg+xbPEoiOeFZOh0kZuCB8Oy7qoAY7EtxYV2kO258HmkJuc5Qr9XFlxa
Whz8OZfp9Lg70Gc3MCm83dkxSs3v5i9deZw1Jwji2c/MUQTkCp7NDpcEOczr143B
uXw1x8cKcwzjALz5n+PJBQk2y7dEbOltLvKdr5c51IZEMFbysT2lKyxtSDnmSGpU
RypINEMnDeEUyKM2bTuBE8KLofi2Z791WEUrgpzKd1TxKVjJczMWrzFVTXbliuGn
g9iLxZGhXIPTGR2BUkDGfKXbd8LWtdN6Ay0UBEBcDYR0Uh4JQE7YBxiKSHifFJ2f
IsECptUelYj2YvsvqovQKk4sHIbXGavn/71gKfnqb1h4i3+tmQhDslzNwtwZ3XQW
y6J5Q0tWARsU0tutj+cAFjgVONF4sfrxVgqSUhgMjBOFuekFXeeGWbwvb7e83BXI
oqga7kEJuANa6Yh8W7WWMBKmswKuFmjrHkwrj90z3fOyP7FxJjN5MTzXQaq/PeAK
ejaAJDaQdkmn3vK/zLGCCbAwRtfD3W6fxE14mVmCanCg2DLkZCX7R3pGrc5KmkeM
G8A/H2fmISNAnfmP3GvePg3+a74NswTw2Jo6FFrDrxFE+/QDV14vL5yTTuWY49gl
WB14UmjKGm2k7VUdn2Rq6eSjhjGx+dF/4juN/IaIkAD558IQsWpMQGqpe1L4T/FL
AiCNSL4W5XKxQUt/A+M6BB8GpyHKemwYUXKV4VzqFfyZFvEM6pv4eHgoe7mVoNWH
Opw39n4viiu96KV+QbKPUup28DS0p61AzsztRipVwvcwS2y5audzkMbOLu72DovJ
vGziqEMJO69UmZpTYqyKkM37U7Ztqg541cXrVsfMRqEjhfLcSNe8bq8RsiCHXLH/
OFdYgWLs5PwuT2Uq4jjpIlDsTDW/dh8U4S6Ac698nQwfYJbiX0fGx+ZmGxKQYDhd
O7sIaG8LyApMFCC+S7+0L3rHFB5WtFAW+dZYh2/Kw6FmNHBe2N7BTjCLTc/Q9+xY
YzXTtbjeI3zbPfReExsQMwiYXrQTpgmiKMLM0wUNbog9YOAzUug+AEFsWglxvQVP
+ECJ0L7KqAfPf68ayXxaxbQGwwWKgOkPf8//5RPi+JttSK5gDC4MAWT1vyyWmKnA
j3sYxAGlwHxN81mCqAWmStDiKZs+gP3dSa5et/sWaCdp17k/7PcPMar4MjrNGCyA
Pons9/DgXvakSvRCQFBDGrgnuOep+SfdQ3sZMeAj91Kib5RDnX/sm8kHf6bmup4s
4DuQlZ4C202U0WSLe5RrChnkRJyw10hK8g+wqukrsPECarSGKjoxqFpMlOpnfkjZ
nhiSq+s7V0MeHM5BaRoqkRGrpMwCwRPUGW5i8wH9Xr1mQzfAhAWP5ClbKA0ux7QR
sqVEGiVacvp6k+cTqyVc02g0zjHLhijkn1uB9FXXf7UMxo9ekrYztWU0dhFeprdp
CS78VeHH6d9GA6iRPaEV1D3mh0haYf1f87cdd2bN4fcRIdewG8cT5losbt6zyH9A
kEaqcTKC1/eIF4YU+WgYdHhDrmHAvYQiA65/dPi9cDnhFmUpu2+Rz657qs5oUSY6
RXbOhb1NpfGBIiZKDGcR0K/oEYrkhWBbS+c8QGh9sqSOAnfdsjqKm4s6//azWswx
pewJvzu9y2WNMpUMaKX/IJr/waXRDN2z792blibBEZU5pQfXQD03SWS9JlsXffOf
V6tA7km1GAmKlVzWS1NZg7cwMrPMruoKzX2pMxY44KnZxLJOxsFSHvraPIZ5a3RX
uM8jnt+Ug9dMlFutirzf6Vt2ws2bvVCwisqQvvO7s8JqarU+Nkk/6mgl5nmre3YL
PTkU84gs4rBdp6flsGMwpOurdal6s5/LUwLB5O4FaBjRe2WEVix++Mf005suzxlC
bS1nspMHxiMKtgnhBu5H7oQ/ildemGXe5DHGiqQgVZLh+QIO0qzy30UQoEK4wsJJ
sj6dJYzjGCOWZJ9NNcZI26+2C/xUQqEcR8XVgesGm8bbliCImf4V1dY62Y021Xpq
PgQDTcQ+9XK1CzDkrm75TJpyoeOO9q3myy6jcAIF+bEzbkQ3+kCFZASv7uyxSPD+
31MXLZ4gchUXECyg0ToSeF8EHaGUhY76F/8XjdZM3Th/5aQpRQ0mv0hRrzz20LcQ
zVMVQnc4neHRD3RXdvc1Ap8hv1OnGKIcL/+hWvpITN3Q2uHL/HpO2j1zEtIoFr4b
d1inYhmvuVjXX+hIDQI9+JsiGQluoBZIpB8KmGWjYfhyFEPfdk4wZLZ6vkyYgWdK
MvcpO+ATi6BWBSlTFcl6A+pPgV0x6KLBzXCn1VryVWYujdDCTN1ZP8kbZQnVq4F0
2Hf7N5TZW3Vl6X2EDqJ0qhCad5UBmwSEcySmZ45ZW+r0ppsl1+aH6WKW47GMs6yJ
K092xyWf7si2rQwYcSaFz3KcABry07oLiDVH3pmuvBC/JYFsRdqsQwTmdzXATYnB
+Ke9L2WuXbTTEa4gkVKkQNqN2Dz6nW65xCaRMx9SVGsjZiKuh4Mz6F1dLef3mgkN
F6vO1c9w7D6HHj3vJ8uI09vf+H40LHrJ3BdYAV9nuXJJ3ldU+SaXp45QJ3CfUVu+
Ep6nSwI4uHETK0L0bGWhj0KoJ8OP7XYtF20TirLyWIkbvlVfqCKYEBU6LJr9ks1L
8kUO3JkGtX4tNPTVmL1lNC3Y6cMWzN/wfkCNQzUFEM8oxmLl7jA0ptuQtOXkvYgr
uvmZs3ugmX7sQmbloOVPyIQwDK3VNedOEVaDUHlFSkBRTzVQufhhAxtu/2SNUr72
B+xtDr7oHzmY+vanwlVNtffcCy8s8pbEKSDvtfKN7Wf7V9qsxHp2rxwXU9N5IMLz
yjJIUdx+oKWFQLthd3im/DEY4eN0qcY6h4wV0BUKUkS9oZpf20luAihaKGdioUyu
AlybSiU8jgpLgYQF7qRFklo3BWqIbGA6udxFnBehm0ZhuGXXuCEsFe8PT66TSRLN
qnbszCwIIwoR3cZfPZRUYSiGo35zgqebFgPFhe8hTFI52aGMrOi32lMaMKdqSMKh
EzOE46OlTNG1OymzjPHAk/aJsKzcGmUK4yZHsn8Fp7aEPBhAya0q+LAVNgZdd9nd
Ffb0sMdhSvMo9hZkf25bMNHIJax7z53yMAmspGiodR35hnKQm20ac8c/DITqyihI
kmb0aaLwzaN/nNrgRvFzuNZUW+Llmg06Drd+wvbmEPVga9f169ygd86tfRPVATzS
5BXXUNaFEAip4gfd24D4u+M4rfo//6t7/cWaLIVpfdTOCT1lSh9BErQ6nrwZ7jrS
IRMY2cD2k6s/V/wP+aMa67u5GCQEeYkPEzxHGP1IVWMXwRG4GS4f7MeFoAoUz6Xn
zSz6beZnSJGdIHaTxgSnVhc2usCP0/kgU2DHRKmF6cLV5EGxZmJSY8VvN/udnlyo
pgu3YVwv1iCXypnyH7T1yJVAQ24OxMc1EzSVSK1ChPqlDOkRSt1EYB0PqIaZgSp+
eoT0NEAmDnOpBOUaCdTDr2sEhBFMvajkEMfV/60y/IP70PvgZiRssrZOoxCUi/Sj
9itFdbWPC9UkP+e/q4LNXs0KhIKYQautIfh3r43J5lhG/uPpJaYlmnLaG8p0gZH6
HS/fgedTgHC4qDk9vqCeq05ob0xxeyHBUKXOEbei8BWepUWq2q/SlgCyuNmAG9ZX
7YrVf69dejUDqO5XnEHw6LcBILalrkUpUvvzprnTHNEbGbfHDoKlOiWAPMEns/sT
ZwiI2bYNNpJ6B6NCBJFuDt2W+XXwUml1lMJQgv3TlQVDi/fOoEcvkyHkYvWZxay7
mH6zpb/PUNF6k4rGOvPNDlaFkPSGG6pYOxANJK04ey8r0FOOCjfnYhU6Py9N3uKH
FrQJVFpui84iPoCgxAsWCZeiPwsMvyqRzmaU09nA+00eedL9wyWuT0nUizNf6nmI
V+CTdvI8H04Xk1dVyo5sI6l4a7mkDKSpDKu4oFoaebV5RqErwe/W4XjFXkuoaad+
8qwY7fmLULIsQaLAr7V9Q3rNHRvgnIrn6bLLRgWvX4ohOKLM0FF7dRBCuk3G8ai/
lufbujLaHdAv3DEH8uRmnGywK6mC6HOw7UDT8wzDWfMD34vYgM8KtyE4KIpL1i/9
lESv1B0sLFYoRkDLvd5KF1lQM4xVEBpvxDvtT+1gRpE886EPmYVn90G6hH4/Q7fD
xhCyQmELMZd+fpL+yc/7VOrbVd+IDQAsjud8COguYRnt+UzUAItocolKjE5XEkQv
7vju5mjSnRKTA00mR7XjNrt9oJ66/8jL4ElOkNuS981nsavpnt/5sKY9HG1Yl/zZ
1kh6elvxmddJsSgJc51AcjmGE1VMnDB1Ul0or7Tjx3coDmO6gQhCCAOEyTwkqzMx
l5xN+Q1BzPsSpddtAmahH3P9kxfEsrFuHWOCSslhWpXNtQtmLOBP0C21qT+7m3uS
czps9pDd9TwvqNBvMwMzySX1NoTV52D7syrAfu31HsL0lEmAz07apf/4sTCUqE6x
JxcSUrJz7/uVm4hjM3A5luFMasru74o/EkDfo8vkaY75MkAQ7/V79KNJd6JdrhNk
EQlc1zDn7Ny9GGorNZ0BgywV5FPaxR0KL2gA8AR6BNXm3l1L/0+GuwPw/CHUgRxS
Jy5n+RXzVThqfA6ep9MN2iBzyad0nQuVjo04g1d8x1ZOQtwUpnLvHS8pU4WpzSVj
qECC80Tt7oXAtOpcqYclvPg/IKtUlbsc1VF4r+ANNGF/sGWoyS0YIy5gTKGkBlal
LruwIwPe4YNXUI2lUPq1OrpPKeAuhsRwsLEJrbc2YIfbXtlS+IlR0vNZtySzvDJp
yeGLqBVSSQxdhfgDVcRV7jFiOshSo7a0Gu52xxyhANAPsrmdv/Ao1V7XjoLAZton
0hHQfopJFezQeMMWSIrb22y69VUEXDNaajNfBL2PWh8WBlXDJr6DrxoPD0yK7Na5
TmiBEtLTCVf1ildRKqqufgAD5NtuMzemh5ciofd6LedCgq42QpFNC7U8OGU+3wlq
x8dgV71IHgrhJqrNnF5t7QL38XOpsUqdL7+RevAHUZ4xbiAOdJ17eQzgDp/l3fJa
FwXml+14oov/02kFPV80mcDxC0RWs6GMRMEnJuGv8sXlDE00ROsE1bAC8nCb+En7
Ek52d28NeY+3cVwLNbrGqwqsYi0dnM40UNPs4GiGUT9+KBNbUoMQXB+NGvwYB5Aa
5Dm2RUJZqETCIlujoxG9GmesXcWJOpIHYy70WKi5NZdO3UYn4q1igGvmPdiuA6p8
5CbvQuW3jRJ4OBMZMwY7qYYx6gTrsd8S2odikLbgqVUqTUgpT1riiqQZVoinxhic
OCWnM8k1kI5hwpx01pt2cC2MPQI7xIn6dQp3vFmmNlE2GYBQDOWBLPX9X6FMmR8c
vU4s9L0Uln/T482CJXGv1/SCcNpNG9hwM19FQynRPgaN7WH3fmtViCxS4cyXS9tC
8TgMkBSzT0rUmW4mhrNsn3TAEqfWE79fNPmiAXNSl9Wyr4ooQ491sB/lJw+8uUn4
Z0sbTia4OzEzDzfzhdbaHdlK/pFNBYFIvmbW8pLxkrNDc0jqQY4Deey5B4U3eaCU
PRM9LGxy84Ihlv/GRNblU9eX4d+WapnWCmoolwUX8YezV6D5L9PIibXGp2AtFqzi
jUzsGn7sM1rtlCFPlyX4gtney9ZwNfhjABpbMX781zqxwqETfOQKpIGQMaPk5kRE
Oydh49EENLOElOoiXFziED1rWtGgW1l1rkRAmz7dmg66THom97MmR0UvPIU/EfUx
n4LG6LHbsNA6e4fuq8Y9wHUcSzH6WyErZukRjNAsiT8QQRlHydNS1RHENZkiP6HF
RxhiBz69s+4JjUYZ/ZUsAlQcLAOnI/IwrprIQUo/Aht1f2ikPAZVk1zFzBh+RWTw
sCbE9L4Whq2ZE3UcwwZi6LLgJEU9G78EMgfiP7V6rtjZWcCl8tjhAjf55KcCtLm0
3E/fo5ljWzNcpGMU/7508eaKgGXsgesfloHq1kdC/hla2CuYPHgUVIGjxP9t5qUt
bc+rVxpqdV9Pm0wSbCpORqilw35TYZSGk9yVxs6wd2TXkIkRMCXWau4GZlMV4YZm
g10fCNTGuXGKmiU4FgtIq8G8dmTTTmDHOtG1CBUKVnx3VOrBZKaSYH5tXR+gvUh7
0MpR9wvLFxC5wVkucPDPSndtYTpQj8G6sWxPJBgvXVwQNG2WXRwgfNZxOv40Vugf
iR+Waqmnnjtk0PeG50GRZnKMbonCfG2W7iKklA2Ub/jt0atuioZIJKIgNPDwgzYM
nKUA+tyoOKavXJZfT9I5Axq7sKVcN+tbBr1d58m3Uspl8r+B6PNPIXiLW3Y69XUL
D0LGiW/X+k8zAPu3UrLDS0QaoZfKIFkfSd2B6zH7Sp0SzE+9q6gU9iczCiCFkweG
oaJVRDhtdiR9YS0mZQqiUfwz0kXlSbtg00Xp0CoizMctNN7mgV9XVoeg6ZTpJBzv
MMGRA0jvgQBJjQSE76uVtTeZTwLdq8Ovwsca4a8fbk3RaCah5tBgUOYWQKQapCkf
5EyJpBE6SJQKRoIVzjA6UQUE+kjAWpVV329XomUnFnJacuQvkiM2E2YCqNUx9/Ip
rUd9YzX/yI6ZOTr0+SOD1ucjstl1vtO+L2uqHe/dLg2s7LHRKvQ/nK4z/SZUsebG
9v6JGWqXpCphr5vPyLWIQSYY9/d4ifGQg/gkOfp5pFmNY5Kxqo+m7wuuXGyDrS20
ed7gxNXusLNkBaoAHkekvG+PENDtfdYCuo0EiKk5P240yidCsnEitsCb195Em4vV
8+LatHN0pyTlnRmyN7SZWoDRx5sB3Z8OsUQ3CagRO4chPYsILCeajmnQPULZ240Q
UsP5Jv0FbxnWcMDYapApLVCN+KOwZrxgZCUz4dOxYI4YPo5Pl+G0f33cjdj6KXc6
S8uMCYxdCRsnLKIggvh5LRHYwh9IZ9qp74nutkC9z9+Vk/xPRNcUjFFnSJGMaX5e
avR6WwGBhN+zaBD7F1vHagfA9hLgrt89pn0hZMZTRN433Bcq7Y/Ai7D80j3sFg0S
uvgKh5r88kpkk3toYx8HHFo/DnZwWbU0Z8uUtDhN3P/B2jRH2LHhnB73G+JVOee+
N5no0MOJcCINCy0uNG1KZ9kN+EAexdCd63UI0QEZHvOG5R9gzuxlpI3qfXNM6DIo
KKGDpF3RZu3oYVU21JTzxsp60GTVA8o3Bt50KsXfPXSOOQZcEBXcOSUvxMX4aPsK
aiXe1pWnV8XgSd7pEr3AMbNwinjdnu8loS+yqXLy16F9NR8r2zo77vQmutjbKFk/
76jAThuv5D7ZSqZIa0LJEgzwtHnuUSMYQOt1JDyFzHDy1J3pcKFX3ionE3jGggbJ
69ghOyJCftbuOegPDpCS+fV1s1tShjpmfqURdd6/nXwr7Gwp3LY3Su6V9XdDDOmj
q7owKaIbl75Js8KIN+qCXI/42ZbCetH2QMqyuX4hnkumBMeQOk8e7mQt3Bn/sC/6
vneZ89ZIDaRvZ6av95V/k9ZcQzAXas9O2VB+sszhmg1jD3m1+dD28MEI3aTiDn+l
u4Sc2Z3Huzk2gXCNrGT6eZUxm8T9ahaKsVv3rYbW+g6ddaZWbFfmg7v5sSR1JHy7
ferq02k8E8wt9qrmgNZTgwPoy36Y8YVJ/6U66WD9fAvLQ404MEYErtppf75zqwZd
lkHmaHVOEH9AMFnHlYp1WeOMTa/o/oP7zTkWP6RkGBu7M641or/ur+w3eGI8slIx
IR3wwCewm+2SBQZyt9SMATvJMsEub8JHsjc1XFULJmb6x8MOJLHe0RsPG1uB3oEz
GpeDFVhXZjoEiywq6vMMMD+wCjgLhc+rBUw5Z6n7GB9c1Vxa6Wt8ReF1WMpvl8qa
0yB2ah7IO1PolVubWNGRNvpdL6weFefLD9L3AbErg7tVH2IAH3sqklm+qQBb3GzC
cXr9c75b6m/sfJPJ4KR/FNEniixh7r1Wk441vZR6iN7Kk+/KI7bvj6scgboNXRqc
vlhW29L2POb4on02QwN186d8DkrSo8VbYJc+dwRDx5Ua1dWTq2rXgJgoD6Y/uVPl
f/JM7vTs+CRQmYWfAevtG7ayTkXfC/NbUgu5KXIWvJDJyhK1x1bFIYVwzbgwSZ7F
kMcuAAAp8TKGYFHSt2XteuxS19i3sWgunsVNFqGlSL6M1y5oTdPyTu6lVqrPRo9Z
GBBtYfdgY8kzFaMjKB4bhN/GLvKxXphh9itTIJBIzgW0EhtxmVuETbByz1vk4Hzg
kM4959KQoHaKTfJwEXGVtSPWYeW7xCDJa/9sAn95i3rzLrDfWFG/UHlZRXEWTndF
4CzMO88E9/GWk+CBwZIGy+L54BaxGYVpgOYvmm+wfmrSWg8pAlqJbmPUR7gSygT2
YSDqqSYaHybGMYgPI7Lb8nJXYOQvp40VC1BJ1gVJkJS+8nzJSPLt5jhXxpMzEgcQ
DDz2B+Z+RXMUTjeUPXS38jamlsMmcTa/2t6zG8A1eK8SQWuyM4FbcRRpIOlroMZF
+kBwXPEusX+COWJ26fuXN7iOW4piP92uMQJHUi+cj+5Z/qs+pkFCdutFS8+SQYtB
+lCdfnkA2HHPsFU5eRVyB4IAVZZef1ln/U10K5HG9GsgfFC+rYFVCmLXjK4fsYaQ
Aes7b+RsHoTkwzJrfIPc7xMfqaGVT6/uuxH9jQ77jwA3mLiprxQ1YARQMTNwxiHD
xsKVsgGH52kDuHbNr6j+iD5eos3NLnzAQS9+k4TKilVj133TaLPx0cGlpw9pHeT6
kmni48JVjZ9MlZJLQzCn6qR0Jei6Dl2L8Uwnv2Bq6fXGTNRy/eC4EPtqJdPSPASr
Z0d9+3o5eJvkAn1xXUF/3D2UYwWaqP4uxFMWG7Nn6QoEqWp57w740FYnWz/R+5BW
VrrWulILbc88YlsLSXrA8jl4UpuGZha7H97gOX81EK6l1SENrpI7VAzImAed3Ipe
83Lxvdk+3eCXD5skj3RxAo3ac022OxKy4fBmkv+iDckT2NHnuRqvJ+n4/MEeUG66
bPzqa6TutPudIUm1Orgx+93H+fLoaBvm6kLmbgW+C2m8rw6iWs7feBm84UKPbVS+
g7OhrtauLHvi9oFg3XgUAydUlIqoX3bN5F73YBlHSTJ2E7uR/+kAbfOvnMbWTWtc
iqVaum66ZpKgTtpV5RaNkwsg8WCryjQsWBKUnfIiIuUx+Sr2QJxKJdID/X5n8iF+
cugEGQnCXGFXAX87ojVJwaIze+z1b+hENBcopwV3p74R4XfArZpGRg8RICzrnYzT
uLBLET3jCOyTyDB0RM75t29vwAswkGIKdd1ZAxsTIjcc9NJuR/Z08k58aARI/rJR
jtP+ZsNfKIIk+FO7IcwkATgNZnlx0weBxnkALqDVfp08jje7yyThkL4ETcBa1DQv
4nIZQx3oEenZST19kdp6bxzK3bVnw3gkqJStTgBan88Hf2nbfCi2T4quIXxOMe2l
s5636gT+Bl/4NLyblME8SZQhRRhBOQDQL+8q1Byn8Gt1Bluq5zoRh7BAPLSEhvNk
nNyHCyEPWU+D7v4c3pIJJFOc2Hn7OntMj4+9YbLYNUosQRhUFt3u4fWTDGKWva41
i6St6TwBE4j+BIaXS+Ur+iiyb7IMbYR4Z1OmwAjYkRxm2KpHtiLm+kPJj+17QVHv
5gP5+D39EY4+mGXO+fHUYhi/l4DzYADPktj0125379QSwayf9qAdNyNpIylJMuzw
3ri+jWPO1RFD7BjJok2onXkABFUGSXi0qAovpQuXHgbq0W7Cyi7TyOxbVX5T1/6n
/IWZ6FKcFh3jxsjRBdxFW7DeiG00zn1I5Clo9rEMJqltoheLUlY+6hmGXqZZATnc
h3H83cU6EpO9nLF91PRKfRA1UE9BQPR7g9kETTDdCppIBbwJkMTdJUejgNzsEsqw
XSd3eTdGzXesWvLpdsCLc51i7NjjgpMGPX6JAYyax31jWcKWpN7wHvJM0mwjgxIy
G+2/af5jwCp80SifPmQu7N+o3w54JOZDporse7Yzn/MIpSYSGZ849PhHhBbOfkcp
F6IsTZWjyZn63gri9KJJiA4kKI4DMcdPhiE+hL41407aUXvHBxpG4BLAeGdsAvAk
YrmljK3/zXY0BCc5XurXwah2+a/ydmKzcMDakg0s+RRJM1hy/rJtIK9VsRciT6ZE
81QNdUHadR6Hx/LIJUHMhMU1kReIYD8srScVXTnF4/tnuVrZE3HhFH/i9SpSFH0d
Ynv2EalaPc4EtXxvkMpaJLhkf2bMbJUFQGCW5UY+y9Jpq3z8+4IsGBDZg4a89BHv
B2ihm4LzyDqXpAoj2doAYI2dpdDjskAHGAJA4/RXj/puQuVe+vxvB+se/GE84q1k
RJKzosl0HPyGLcO5qfz51UzcuQ2gfzlSmqhz0IiqYiERHNUcoCj5ernA2xBkRDXk
gcQG0D1wCWFDEqs8QjLB92zRseovSdKUdKWVPv+aPUbUWCeBfxQcWUFFkv2bqXIT
FjIzTR/Bh8hp7FXGn4x6dfT12pyrcT615Rh9uctCohIoTlVlKVDLBd63WfKhiDLQ
jBZ0QT8WhaFoy9i9p0aP8Wwj6L4Emxv9kbpGTRx2HTD/6gt6jwVVXLN4yJIXe6/q
tXk+yBWP03MEi9SBHd0gt5DPN0Fd9p20/PFBvP52aMq1yn2e4ZznYNTg2TKDaIr5
diqMgUnIMPYLFDFd0+gAFw9Y3ugUyrd1D/n1E3h/7k/y9uKDOXcV8WUqMUrvYMfo
k79kj0jBdX8Y0lPwfXWkBz0ByW19aJOqaYHlP2ztXV0h8DdL9kGAT1XFfGTFeTTN
n/6FXyFTEgbZfJKmj38s7xOCLNhaACTvWvkhRnFyCnVclEbkBp3aSZIVMbI/JgZs
UUXeXtOIu5J/npmzrqpCZQCjTQ/LOHBGCl7xNf1m1gNDESzKXAk2rNfqb/cxR7Yz
pwbnPDL9QAPYQf6fJs17LzWL5q3M7V6UYPNdJxoJL+vPoMHPPLn3IBIzdtJpnTtg
zA6aIK5Xigz+WjJCQK4SBLWrmCQUX5RZRNyKPUsdKRpfb9mIyVSeEXZljD4oa34C
d9hshK2V115qUkDuuytAsi9EGUgNbNwBkcZeCzq1cT67yjK/EwK3H3IftLpJx7Bp
4tXoH1ifL4NN0n9mGzuy5vomg3VN0Q31M8Pier+N+PirLzIfBLmKQve7UW+sZk4o
qLYz83Kgv7k3H4lh8Tr3YaAyuTFAUbGbRXHLNMujKb1CUFEHcTszy1v0miku/tpB
rFByfL+qOwbKKA9j1i8mDx/sN7mXHSc/vXXkSmsl0YhHjzCPTsyZtcuJjYWvjEvU
lk5MHn0sUkdy28e8Qd2AC1J64iOAGHOn3mUFnV60EA42EL4tEObCTCl6qQoltMC1
P/fFluB0b3aIj8BpPeBrbe2oTzoin1ZBY167IrUWGOnU1NT2zkCeFmkZL0ED5L2S
myZREkpQ/HottfdtSpODMmFzNy8dJJhsYSJlmm6cO8s2lA5LCndvVoIbxr5G/OlJ
LXhFjmX3Qb73Uw6xwEtzbY2485namDrgTUnedjfwnTh+Whth3hXGSdvdkV4yWVto
VqUW5lP4bF/Hoyf8YoriKU2oEYGeiEYwPKYqgBnkY8FX4H55TaF9j8bj43Ofa6Xx
SMyxxkP8mGVjrciYhqHKZbQ7Womqam2jGUL+qkIZ0Ygere2FIJy1cgD3NGSkErt9
Z3dopcEt6YWTUCNm10uIO7Lb4edONc5MosqQDk+hnYJJ3I4zTr85QONkxwwIZHIs
2bpbho6yBLba/gwFliKBdpt5Jepy4UDJ/NOFJy12nByWamcJ1YWQdb/MfV1+olga
UEt0BrGDN0I+lIUhDKCfPAqwHwvXf7HJJEVFXXf5oQUuJxc6bFLrQUx65Qaixvr4
y078lfTkP4btaWJbe94Tw4kHn192YTY93XPfwKKtYI0L7cE8mmG1MaaOzyplZH98
/1JwnGU9fle11EA6j+5PoCZe4M/jaICQXtxjDvj39fR7ws6afsooyuiPTyIgfn7+
kjN7NL8WbxSxv7igZFdI51DBFtLYdhaEYMH6PTHUpBFBDEJl58SGVJg3p4kkgW2c
dnv/C2PARrOoiFGpygtkf3IDtopat8e5BfzwsjzzEXCN7TvwH0/PRCcOsBmOUXTk
Ojigv/cKqlrd2vLXH5EY/CYfd72EjpNO8kZRz1hUMJkbDi6zYq24BF6xIu4hKWRZ
Vb8Ez7g5sYb/TwbTDBBuVru1g7c4uLp6oNquNPLPcF1WD0qKCpj0EWHve1kGQr7c
Wh/FtdcZmgruxPbAaK04i9QSodoA8j6VY7RNygCpqvuW8W50mPu/urI3B5j0auo8
CQbW8fCVKgomaHE1P7cL7hQbX2CJwOrXkRNO/0+L9CtVG3jjZdXASqOUDOAuo+4K
WrCkiMM+Ru3DiYTrMFwWZura0No8Wo1Gdf2KTr7G2IWS8DVo0GZ97dTJYPvWRDbs
zlnp/CHAhRCRzLD1e9+BJwcinOkydHntb0nz0fhAci7Zj0c02O/xpnJK/mEsnivZ
o8mbIbuiadrNOVyXIB/2rPkpT6sGXmZ3k9zCT4Ftx0oQ/vwUeFHKNplDU1ndTlml
/a1puHCLZ8XTtJ4QrAQdgQqYOkkEF7/fAJINXWB+AB8sP4GahVqh3JgYtzfiUqnq
GmQNX+rOG0CEqMSIUzq2wrnBtwtsox1CYIZQ9a0FQRPV+2O1naEOSnrz9hAw4pgI
ZAcTrUAuDRIKD0/dDcjmXXyaznPkCIM2culU1pQCsXpZ5+2+YwadlCp4zI4xgFBf
HOduZ+Le5NNUNNNxKI9+yqsKrWvVaUd0Re6s5UD+87YQPDYiS0LpkzkFti909bE2
UHVC1+O7nhiz75GwhSi5iGdOWkHIlfho0skc8PYv/COCOqAls/qfowsEEBqSfHmQ
kVj98R7+uOYYFiQvFwrKGf5TAFJRkayQrVoiUvQYHjB+CpV6JQs1uMGK3VJsVOmT
Vcl+DvEFVmG8pJC8gGyfpNqupIJicwVdOYHzvXZx/bOI4UQaDyl64US1bzOOhBwk
RqOiFl0FPzKzUHW2llGaVO31zGSDRcK7Xbstx+yLpjcR5HZ6c7jWaMedVKJkHiJA
WNSRuNTgeTGgWEEg3ptGcqJtdgtCcOyh6Q6mfNZ5r1mie7RLPmAgEaLxiV3XtGIo
dUPfI3+LmYM9pZsBg0nXTwGijBIN7wzd/3GAFN4x+OU/UFNvuMIz6VivbL5Rc4IP
zMadZYtQ/u1ts72wxvAJgTqMNg1TOt6/BUXSrQf4Zf+bd7TptBYHtWups2aH02me
MNPXtfv/4M9krzHIbtACwqBsIqvrcWLqTna7Imz0DZIYfDA+3Lgj0bwOFx/g3vl+
1gce1CdyYG3qEhqCv+2GpWCRcHDXdWbg4iWtParE6TF19KDNZHksB5maXKg7iiV1
hg6Ojk21Us+2LoftniIUAGGa+jp23z0BkQue9mzA4Y885pdGFjPJcYOAUE8fHpV/
+jm+5QzPmP9Xw9cDS52XdxK4avj0wRYK7w208cyuQQRcBfF67LnExgQf+DZjrFN3
/DWJWTI8gW7vklrDEg38Cj2TAWDAi4lYXtnTAlqY722tvHccSNN36mDJd9rHP+9n
fvrLxISogO006Xl0dKl9/e1eMJQxKm0/VVuVz1gPcEiWSDJNyrXFA856ql3w0qHY
LT8xXR7O4aG/aAvb8ndx7XbT8gldFol5/UNOO8C5tyrRWrm9uGIcN7U68YganCiX
7ohnKK/QNYqXD1V+Zb9aiU3gwxuvD9xtIvzRscJ8RsqhfkuXjb16gkWECVzb0/bT
gAx9C2lzy0l9NyUhtu0XQ2Sm1a4QxjiCW8Q4AWeYZjRzSz6QFMLoy20OlOdqWhGj
xOXynljPp8yc0NrDu0VPQYuf/67UlandrXbdj2uZnQu/eNZAU2nnZmbhdUC7LLYT
itiKMCzMbPj2XTNBrQalVFANSuB9OGRY01WgpM/3dg+CsEmiT4kydj9ksn0Sc+yT
ZULQQx/WRdzAhVeTRZ6uOdOb1xtcFo46qfWuA/TdtbAqBt5CvGaAMZJi6zltEJvZ
O9PcYgpX1Dxa9ITJ/Lp0IL0V9NlJGX2MG5vqMLnsvyfs+UiXRcheG7M+cSzYCH0n
rZ82aDsUQ3wbS1FNtJXmJkKnplGv25I74ZlZQFZ8949wvwoIqqJK63IlIdCXHZx4
Qrm8jDCVT+bmVwg0UyWuha6d9riHWwlLtPfdyc/OdammrmLgJ16RQyR7I4sk4D62
YtP/oOj56wDFeT720VBWP3AN7AqdS4te/7jL/quTlZzQMh++0bPWEruP6XEnwjbE
0GQQsfSzC+JhldiSAtbi6GXfpoT7xypI1KH4uqHKUvzzERkPRbLQgAg/ByrAjms4
Wr4culHt1TtXgk9vaLubU3eLbG/D0xSijKDUFHLvxHmWpPfvTedX/vNfznrwkEq+
aVc89eaG2jQEUmXEiPHZ0F6ktfGGB1SUXZplZh5+Zgw5D7mGt74G/748kufPgsxw
3cwQHdWMq+zm7lvrkeG/RJs/PxjYzTZT+XdqqZ+I92RDVXXEXRTOFtwCitYLkJIO
p4ula6kXYxUIyaUwo/O4Mp4Htef3EbkBL49B61n8lActlqpwu8JfeCE+pNA6poSm
P27sGg3gVg9VREBpZJBiDk9SyC0C/f3aqT6D+rDfbPc61ghWNFBDQ1/mT8nKjaBU
d7Uvrj0p48ubEPPeSQsOKYyKSvgXE6Pn1o93M6K4nLGQfAwfVjA3ebkE8AdiHs1Y
0iVkXWQhZNToTlHFG6ZsXUKT2QeEwdVn9kp1h+iZc0frUF16hJXPWDYIMlPY/Y4s
PNZLQRImmcCb0evavTuX9nTH/fJCM3EpgA5D9Bqbqk7jeDOa9xCN0uM/WfDGI79G
tsdj+HaGrME2vJgfy4ZL5trO/TmJTB/az0KlZnCbcchxQdJVwMVQKpciZihaDekb
AITm/KD5rbn8dG6dJpvhgEMrNVdKAJJOF1OdV/TS4yW7uZbjKgk+k/DCrcrcwGzt
TVG4PQSAHxiPf8F50WwwPw0EdwbxoxNy/B9yItrlYnlvZR7UbJFLHF/SYmIdXguN
CGmLx6mhejKM0xuPM1tF82Ro7Fx9Ywwo7btqruqAP6faBmwQarc9/367T8eyHFZw
VG32zahexZEVsh7nMb5gR9v3lbDRgwdefWeNDfKm/Amg9x9kH3F1NjXBtlsNH5td
kYzA8efJ6YVqEfzrhzfvKRfx07DZPQ2JZhqZYXAUA5xKMj6kAKpXxbNBuwa/Qelw
iqwv6sSLmNVGQzs0q9pic/cxybiOASfFr1GU03OjVI1t5+bzhEyxGiFeQRwbKXEL
o3MRUqAmqS78p4QBtCyS6Bt1YbqX0ChXtNA+AmbSxMcue0B3MzlbeaWSC8pdRHP5
LQWEw/rwK7Ixgd+XXw6R+xGUNl7bVb7x4qaVK/j41Ms7Jd5EYSfme96i8gKchFOW
rGfekMnJ2GIX6+16fHLrsnUpRrLu14vQ6NjDQIG0TffDpnlwKGRCeNSd2KaxYLTm
dHfLFoHwDvej3AKiz3IHojW8SGGrr27WX1114YIUngCXwJbPMv8HJC4ik0O5/roa
opE8rh0poQPMfR9QNVxHKy8pGXU4UqiyPNUo2xAb7mZ2HeaL4ZvMR3oKPJXcnbTZ
y+gCXs7yUQst6kALqVYm7Sp2kli5I9uuUr/LVLXnm44rldiEP9vgD4tyFJhpQKm6
JUH0nR6XFT55ufN9RULoE+P8fbuPwFOYAXP6d5t+M/CKrINMgrPwVye1Ljyij71L
VEYPyzbZCh3VzMBCedfUWIBc3Ylx+r5m5b5l+hcwecsgvE1lwNsguFGBXocMofQz
YZydVj9duVg4dAxojjWgw29o01o6xpVX1YauXT27RpwtHY4St9r9TTMx9IN8mcT2
nI48rDyexEWb+jg+qoSbRhzXmab5AuO4d+0DFhnEsoDzsj8MC5Yg6wDQHNv8OWOs
JfaavmSdNw84FIXMKN21bswNZzppjli4N4NrlIVlHaDUJ4zt5ZeeE4nufqcbWAS0
BCvQLKzrpAg6HuX4UyiLAmWNU57o/rCHp4UtiL/3tgXsLN7TYEmLyCfJ/4FZSVwm
pPmEvuwWMPzqhS0PE9zV2+K1SP8rF30QmA6CHj4MIY2C55qKm2gYil6i9u2TPOwi
E2rw8zMaObvbGMc12Tw6F3Li6k392ZD+Z0hKp214UkAqlLQB/VdiUs+JqAi8OgsP
xFb3D1qy9YPUUhAbf4ZhC8R/yTsQOvZ9cVOV0BshZzViI9vNvUq99CetRfTWCGPw
jjUQz8GxFOctRvvSzDA+rSz94eerpWZW3acwuZjG0jUGTSmSldNi0qEI4pBg7gPK
QemuKj4jqiQXX5YbwQIk3jnoos/rlJ1lTt0pyRWr0VSbWGocK4sMzimwdFu//Cjx
VlbS3SwOvknZo6NMw5GO8bggmszfDQM/gxXdV2DNP6qEQ8UwJh0x99bEm7CY9NdI
TwpR/joYx9PBEODTSFpymiJWa/eGn2n7TZq9jqzSgDe+DpMBUeYrhQ+/mzh92ZZj
D092YbD9suZBLUdtXQqNUencuh8KHZHdy84DTaiF+0oL08KMgJE1CN3jEPdx5aek
N9IuFHlZNT6L9t1HCLN7BsEevaLSIDWjBrYXWCNmf1ZB6T6YyWUnODGHXMHH+sX3
DagDGjz+h5wQCKuq5OMJL5pJPXer1jyy+uihtZTLsgsA4tZNiWK5PZtbbmXRJBr/
krprMxnILTyWa7OadzRzsS+BS+D4z1FU86RJdOLbqhB9pgyBcqd1CBxPhVZ/LWxF
OT6fIGyW0rtNg2oroJ8n81h8T+nnwbCp4gaDRqpDTlBQQIvRn8mJPKSIvzRaEn76
74otywMS6mpmCeJx7oWKM5LQQTcREPcwN3elNpsxRjFL/FezJI1WhVOf0SA7PSjE
1CJKc/58cJa1Onpa1Ss2NpIkrJnbs6uAl0c+jyAis8z6LMCarIHjp0JErwLjru53
s7sxznfnX34wdStLd8LWBCt684bl5DHx/f6ccJDD34nKGshUFKipRa7aXrZb0goN
9BRxTzupi43mlpHJQfI4LG9PKX/gZbQPsaJT82JcVIPhQWqeTJK+niVF3MX1pIoA
fVAX7UF7bTwITNjVTvk9bbWpoqd+DcAYmwfryhbN2Rg7/JqBCsOFU5MO6cj4mKXQ
E3NkfeDAc1Mv8O5Isz54SKrVY+2O6d1YokpoL6H6kd+brdIOXx5AixDymNimTJGU
zYmsiAYOburXH1i+6ycOOQkmQ/02Xx10GlMvid5F2qyjOuJmXCDqM/7v1Gzx/LV4
0FkBLPiOzE89YXqiy3h7wcy9CRK4Nyxh83KKurk13FaAZ8jsvT8kbRq1Zvlmnm+N
v/6Z5ruyTgWGZzCRlUSmzmy4MpFUon6ddja974+/WuFWVJDXuIKeQJyW0/fW6Egu
V3DaYtlWjDhhEzAfmj6RNCHc12uWkkxYwPy4XFuT6hd9vKQZDASJ5UtUga8x8iua
smHe49HKCSCydBqZ0VJVewQkN+CgxNxK5gWg/2ZePIvfDUnlt53i/rtp1hya3CRk
Fcj4VfaElaNK7zxHXyJz8Y+GvCVZO7cdVNCk89Uo8vJRbXj43/J7DWdLJXzu1B63
H39k2ScEAOY0UyZb4MeR8MVEd6Xa77w6o87a5CkAc2aLEi6Hyievajy25fkOwMFz
+Q2RZFK2WlzQ6MpFUUOKx0fGXU3gWvJxo8rVUvaLSKbLgTVlHNhuEbxsLAPncl5i
MpkO6bNJ/smggEHYmfq18e2U9sViFOFFwSRgQ9d0PTP+lBR/G0zuCiALbAdJYX5d
9gkV1bg+GBvhgM9fS7rWilLme0bfu9HZwmz42Oc3ptlL4+pFvr/olIXaqJNFFXA1
qfetjhXC3dqzn37kbsII8HSHTpStQrHN1joHz3LtJcUzn4ZNOdox14CIa7Lpvov8
kyRKJ/MEMtYg3dTiA68JEZ4UAt7KQAPwBgleMTOGoKn8jPRr7K3+bkjGpwF6732r
7Do5faeFwcb9wvyBO1F8WlwP7a8dCyZBfisllX/8Qp1JMnxaF1sSK5Kkuct+VhqE
CzZZoKRC0qH8kn0gcF6TnrtRp3R7KyM0bBZbFyWcEl6BBq7cUIWNlhq7pvfPCn1k
tCRLnFd9v9kldFEfM0qACOW9ut6kn1lGwslfQ6flwNyFLQti806gsfDv+FeJs+iQ
SRq21p5vE6xvTB3V54ujPrwun2ZvPtpo+whQXtSJCHIPS5egDctLYj2kAeZ+P+3/
/OmqK8AFAyL9VWWvofg27m6999nIc98FkGgkyBxgWbSj0vmi1g62pVKfMTQmi+h+
viR3iHi+aiGxxPB+06Fu1NzA0nF7NSR3eWR4YYZ7BiAQi2Xk11V4aEQd8RcCW5DZ
3d3BedpU8j+JocX2gsogrwpnHp2W1EWI4L2ZcJyy1aubi8On/j0cGcY4U73hjNQe
vv51a9wzFXG7qZzr3uZ1ymXWOTEq8FFfyil7a4Zpj/i7zSR8n5yGT9pGErJLfKK0
xZsZqXDCQr8kbi4sciZ6mZYIka1m6YWMy8IEE7+DdzkTQUYi2qFDDwqNBAF61+Dc
7sjpOjULrHf+7nzJnJB4A2zzyiwfPWGUXJ7luYMc4xrvnQL6V/OYUeerN00lKkXD
EWwH42aYaWlLStG4GrX6oeq6eXGoKCISZPynmoSZsnHLfNqLDKZNHZLR+vmQQFv9
tAi4fzw8RdszOgOQH3mGnq3vK4lPxS+TT0TCtyDnOJdNa4vmi0BV6qQB45v4UcE0
/O85kuh8CQTCbTn0Eh37q4ro6xhtcnu96cPCMYn/Z46kw47m3QhUKeLkWQne4RNo
Wd5wJlYmqoJGfiRUwe3fKOElC1gs7S+ei6T3SoVozmMfB2NfANUJEo8kMliyV2R7
3Bm8NsZTJ8eBpInjGLH6ZkFsUHQIhukpFi/ySbgOlphki5O9GgWB8LYUh9PYqfch
ET48eGKBXPNClCHfNMBpppUQ0UydKbi3utTsBmg9IIV7LTOT1dnQgqKY3XQEp5Vj
tgE1ZmhmNf8MzJ5r07arWDE7VsQSW7lO/xmObKQlRTgECzL6O/JnIMx2pcTSJsyv
KX+K5BgTp8/oIy6aCulaMXzv2DjliYTsQn+vRcfLDytJ4fw626qclVDPNYWpEena
FUornXUMEt8l6ewPrMXG+rnADEjgtQvytSuW6S6GfIFvh28R1cis+p9K/qObXvuw
lOob0NwKMxPBjd9WcP8JWE1pJOOWu5KxSIYkKOklG5QlYsuCENby0yhH4uViHIHl
G1Z2Rc9uBIw2w1YumVIW/Mz8yW1Xtkul46dPNCV38Nb5CpYGo8jQt2WplFLkwa3a
9HSuoxTHVYlDCqhNB89nZj575wdPtMg3rvjb9WbJR48fFsHL2nh8x0AXLUx2Nb8a
qag+ftoSjdBJOzIrBPOhUDEMzi3k+VdOt72fH+rPRXB2ws8pEg/yMLK60NWSHmVw
rj6uTlGdnpt5YZKrpKk9kUSf1DXfXmthqhUvdLKBgEU2JfNnZ06Zq7qRUycX7iGV
4xGJyoyRVsf6en6q6P1WwvejqlhGtubXfo7Ji45IwaIdO7dlGc4lYXnBS/AAJNKP
IJEKeYBePETdN+jB46lOgkjWL1Jssfe/LczorjivUFqYV6xP+h/KmVAzHzCTl1wB
yjGkusCPXVbnwTd5CsDqgG5uTqu4EAy6KfilFbZEVIlwJZ2A3Onb/T3odKDK/WBi
kgKSbzBsMJhY7vXE8pITZCUVdOt6YiETzWKk/DjOBm6K5wMU8Uc4gExh58EA4AED
/TW2lbBy/XM3eRti6BydGOtDnanjIucnyIvsNZBxMmLa4FP4QEliUfT/WUo01beP
yYkM7E+2sgXLkAdXUePkqZw2F8ojoUPoh6HYSjfMX0gHFekbYhPVsDxRMgUdMPCD
6rWLxTTEV8HTbWfhBkTV/HNHT18h/vhg1XKGsKTOAzI2w0KA/tMqv8CuqKrKhQ9n
XXd/jiiz8D+0faby55rhCYNvMMsPhSNPTUtZ1Yn0H4lav3keAf471M76oDJKIVSm
3f6UR1beT3ZCJobVAKguThI0WFTl+R5V+D7ObzOzWLkfBQcxkSkujGMHaXChwtZW
VC9NAlAnMxc/xw/aaQhKFQ6adbi3vPwBX8zkcK8wU0Dd5vKYNwq8+MrOkmJk7nQE
QYRk28Uemr+j6JnCbUJV6tokSE0kyNB1YxGm1Lq4/qVEbqlEKzNie2I+D/4aLBjI
55eFDBqhx337ZBdf4gED/iuZV8H6nM4WhYAEe6sdfIbdwq/gBSxXm9q29aDHZhg/
uUCSAdGO617rA9g+Q2MKZ6mZqMS77HG07J9dpO7gkmpuhfDBY73KKxPR57ZQSXq0
s5L5654EBQ6S6pW4LSUaU6HpEOlEWfRVxEpWtyjefbDbYmV9clRudGSLrCetQR+9
iYUCOMfCx6XeV+EqDrIO6LcUKXOCpeqy1NN6fzHjQX4u1/m0z4qy7ctRrkuWFh6G
/ZVpFh19iV3dLSP+P0w6rgrHG6cpW6RpUCUykH1yrg7bLot7WEhvrnRAWa0oeUHh
dvBgJRJkMevKy8NMCjF/vw0qyt+VtMgroZ6xWC59ACxCg7+iY45kBXCDNe08U2G4
Thp8yZ5bPNXg4+7ZqwIUnWz/yfJ2sCJPZd2RxlppdLrpVLYd4aR2vJljl5ktTL4G
jlx8vHty3O54d8TivRMNNUZziY1nndtZ9KfdGdGDlsSjeZPq7nuOb7RC/fa+l09x
5CRtJISIREQXW2ITJju4o9f95buI5Z7BNG+Kn4SE86BiANMoeTE402KiExVzOzXZ
r0LE2FLlf+KEqmyK10qoxDxh+41ebxsQpdO/aeeYbB+3BY/PuzKe/xT3mK/C4zWz
OL4jVGsEuUIUVPTqOoODf6GIgIOPI179tXc2ZyOCm46OXdBP6lroAhGcb2Nko5G3
L+cWczIXm91Xw4LcO5WA/jx0WdOSebHKKhuwCOxuNqasZO0QzNwLqvBUzvxCviSo
UhGPPceGckI4x9Y4qOXM3m2L9rdpVllXLg1XyY3PnrnviYWzhOv2YjjvXt1zsWvH
yJZQqsFVpMQC4ZdMsuatalZogR1MtbqQLgAW26wAXDE4cbI/fo+IjPg8f5kdaZHw
T9jYAjw+0aFKjZMIOcMzEeyyFxjrFvHZU4RQDmj8VcmxMIr1eLn5JX3ZZPbMVeBX
xk9u5jFLg6twJckMpVLHw6Oiog61U7neDdORXpffhM7hYQxxtoDTb/MebHvJxNrD
SqN0Wb1Ul5jQtbIHJnayvG3p8cY38X5lCUsIltLyz6nwLwLf0wvMl8txcLIwZ4Hb
1QDz6wgicz3gkHu8Z6LKOI/1LuUSjJfWwfCZ+QLytTcU4idzsOryFWlodVH42Zx2
iC7wWTGxyNN5ffkvALfmn68IHBR1549xINgstPR1afSj9DiBxAMLQYCSLG7wghfp
k2UlAI+KIl7lyRcEy7B+rpU8KNApvsg+fhUJe8dGficaPUHeSv/cX5xQY0WM3/0R
zu1JtmfT2XxjzUFoCTDOEzxK4dQ3DYDS2wkH5EJ5LlYouUYLUeuKKDwG6HCXCXH4
QoXkzOoKnARszT3zaB2U3BM+CfT6Svvugq8MTZoBD9LbOSsj6/CC40sMK8/4ca85
mzkrIUsvWUMWU6HUgYErNVTC3JXmT/ZXQLrtYXwVjtCwDuoV5LaL3BuYvRL3enCt
xYvKqr+Cu8bWdzKmW7H0kq9uhLXb+XEmo+1DAu1A722biPasMor3fZjbw8H4BBXC
WqluuheTPxfk78ikJ9wkPEHKWoGY21HEAYOWOLIuW7HdBBFRvlQXIbkJj25i7vru
swRKlZCEYKERZpEL5RJA9qrBzr9cpc8kBFCsZzuNjor22Mr23kJkbT59+tQZrB9E
gLbTgUujuF+blnT5Pm599n8KIkpjNH/wAhbkPobj/39qlPMEhkIAAoAvjFvWKSvB
lAtreaZjF4jDMhQngbltUXPhkQLYk4th9O4lLeN0plII2Tg++CMMvjdD8EcZdtaF
aQ/TW2HslAP1X7Hn3e0OzABDMlr0/XVzNckBNIMJzmT/dmOWQEP4oy06ON2XVN3F
c2fYjGE8yHsQ1FJq6V0kqk4cFFm61nCFNlWMjQedxrQu1t9ve1Q37y54UpPj7Aan
XO2Nx8YHrfOj9dQDnAVl07Id2JO40UuuRSGN633AcMy4alss3cFXBkp3+dJV2aw4
u8/xGvZULlwT6nZ1UiuzUK5HvQeqWpiOYjVjLzkGsY+AEH61i4CfjnN/561f04Ue
O7sT0QPQ/l8di+H1OJXOSeOuyNsjq5ljdVE0XJ2qE+0b5IvRrtO+NeY7pseb67Pm
0JE7Laa0WdZWcmKlEMICp0ju3ASz+a7RjdPJe1TNfn6G+zbB/v25eqYtBFcZSErr
Rx9vlcXXCvXtBgG61MtxXPCQB2ZRTd7r2xovfFiBPiPdYkTBiH/YOPnZVhdnqgqi
iuITZPWB5tlmbierPEWMuz5Xt9HaYPiT/el7qtPwQz7uXoYcA6059c/33HMVjyVy
GQQlyD2rsg2bCVNBHGLUdqmNdSIADo/IXvOC0bh8jPeGjJpTiDyaijdneV5YZQxU
0M+uwlPCExyMFr8IwwFl3LhCdQ67FSiPFEfQkZNl2BfBQuvqXo722AiiXaEpQTt2
N4w6xZToDJDqYVlgYif9H0OLU3IiCbw4vzyjEz1pBuFJeKgyPqKYIdzV9qVtT+mE
nIuWJu98tq65t5Qrob5psfosyPTuTfwfktsIzjgpcaUUNjprRnPCO622oQtPWcix
iPE16W4NEefjypufkk3Zyjk7/b+kXDZSvPk/3iUyC5fwOBXLy9+rK6XEcW1xtKtt
5p4YXM4+TCtZttBrGXQ0Y2Drgw9UcjnZ3bHt0vj3HgjljNcmII/XXIL1KqUhFp44
q9XiF5RByfRVWYXsy+HL0Vg619fvUY97zQ2LYw53ng+3J2KakzHUyn3ZkVvsCJXO
mQHralKxToaRbLwDiPNYlXw57RJkjBl2FDeKK7E0bxqqbecQQlFKayeIwPeTiW8c
yEo2bNBp++mugAXBTzrJtuBY3ApV5siuGXKgrueEd48SU0Hm20QS6+lNJVgsdLcF
5cX0j4Cl/PTzsrV6qaCxr+CxEM6V7A8ZT5UnYV640a/DeJnADM8JEG5mvV1/bqzA
BxXZHiOY2APr2Nfj/CgjWmp6Lz63q8J7TZcpomwPwOy0ILoSz2hue4A+lDw9iA/x
Tm4y7DIixTibOuJ6tX7AoXD4venUtbJXUQ8ntEAN0rgyYbQbsDyQ4517IJpLBlff
lh2Jcj3NMD3j0FhI+giVepV47OBNgIxUtSeH75fJ4uTrq10STW+hWEFX7+SFTP1I
/r1aiGW2dNgPzzELd5f6TBJyTphlWqS6iEBsF/VISQ1OfMlHZvIn20jKQJrwj9Jc
OzJBbpd70931TpRryGbZNLfcrW8sm5rYS5BG6YAwOaBipjrb3uXMJ1ztZLxpvB9y
lzKYGXWCgr73H4fWTlbz0HnJFqEJ51YSTr1dSSVwrIZhGkHj4OufYXPfq6cdx80N
G8XnKbmmfdbVNIARTiENcrtsZbElRQ/ympNLY6HYW4tJnGsI2gcxUKFNvmSBJHYC
hDCssg3hgcCOCDt73btKZkdL1aa43YqxL/33CYk5pFYK8TNc4eDzIpOg5/CXJVTP
ZI2IvLWzqHntYiFIYAFNNfRAClerktT/D6YHfcSCSZdGD1EvXJ4oqjiFsz0DJkAR
SvHn4+4A5FMouU6rcS6B/krhMvnj8XhbwwpsYPPvvHg1TGEswtaYc63HwfS5MqqE
QNIWJx6G2iLd3LuUqMEX40Y3FKin9VNuDfDY+9sI0IptEdPMZQ8P+ktans690Oec
NcISI9yDHWLLxbxGwkHP0NNaEpJQG0KU3+MneduUVLc1f49M6oem5G0i0zETgkHe
RRuz6NQE8xgRYMKsggcPHUUaishwH7lwixK+r9KUF3jOv6F5kjE9zg8LudBOd0Fs
cw9fz8G0yZei39/qk5DY7r05aRfu3UQU3KvaU4ZsCrxi1loLrjHTABqPRwbivgP6
CDiJ9N1RBeSOiqraxa6F4xhDWzM25osCUEWHrZTsUbsWa9Za43ng4war7PmA0jrj
eW5ZC8KLx/p3zcTzy70DRX2XrLVQyNIze9ZqEEs0v3JUW4T3tT2Yt25Lc42C/4PS
XRWjEfyfXkoaV0uaGnwuzDHFhUB7jfTXwhkGSc6QrvvK3LNSPN3JEb1RntVWmteM
ACQL+YzLv9L6usWsQ3nZuzSiHJztCHCcyDHyQIqS40uLY4X2qhYVkHO1IkVrJmb5
yM/9b9eOJDIg2xhJFuVssqu/LgUfX+Fza/I+Sg1kK3ByRMI/RI6nekk/1udqdimR
KOJ5+DlP0/8sTWGZ93R9tjCydbvWqd4+uZPa7ZblrCjN7hJohNajKVnFdHHWo8jQ
W29A+v/njlovDDTfb7/w6vPlVZpWkNu7vKfRYemfLuy7EDkbD3hnx2OknDt5V3wX
F8myOlDpduZI9YCecvX55zMFCegrygB14Ak/63nskMI62T9SKN3dnO2XxNHrW+VR
7VH2jgQYwcu4AYiQJYmYZTleUci60efBjotW87qC70xEc/ngIf4qAgQBXYoRdjZQ
ZnThw5Drzr2er8dZuBU/8f6nhu9RZsnc60qcYeu3XgP2K69Q02qckxKzxTFbuFDS
4qiMP86gENClTBSqCEr9ituwgkaPNwUh/5ebjDyGiM6xEr2Azu25QbWwcZvywV4b
kBVjntcYaE2VlaGq1yRuHsmouqg9ThtpQT/ZGbWmVw0uEvlNMcl4yvcd6sYWSa2C
1biZrEVBCjwFfqIZgotp/GC66f2FPZ4FBoED+ZYrSi0XC058HzjlbOGOfXHECDOi
pHpi6A1PyHYQEMh2vkGrTjH8WzmJgu8qkgeTx4VZMwYC5Hm5G3EydSh5I81sOTgF
TAsispgoDnOI0CtL8agjIa1rXdMMGl05I1Lyr4nltbr2nVgKEKZEaH7aOjnZhgrn
3OHqGTRsmZ2CXgU0re/a46btnB2SU4xjQHwdzYspNqsOCyASMNsFXUzgYhqVH8oG
jpbN1xwAJ+EtXgv7484jGwkp/4WJ4U7ewHh0/TztTiRmQkmsOEy//QxzElbKyodY
Jf06kH1HZ+8+62mOnGGqUd1IQ+J1qDP4s7AI9LRzUwSSIhshjKIaEN8KoSzXm4SU
6P1zCkN4LJkUScxxPgCYXTBv6jfH0/DnPymA2mMs6m5W13kVGKun2eS0sKI0bgol
Nl+8AluqODmWzP0U8fm7K2Kn5auOCrH8UvDFKVmmfCZyji8OfgyJP+g4y/mDQMm1
ob/IEfSLr6PoZEVGJHyPjnIvluUc4DT7vvhd1ZJuc4uceAJIwWLo2PaNn2RZ2ptZ
XGxl8cAsAbB/kJtKYE5mtcJgXLFIYaImAvb7qceaqz0zyTxuRHle2qIjJA2fAPE1
mAmEpxX+iAfw9LnTtWzToo+r4E9XyQkeqlZZAi8p4pNtsdacudB6AliSg30mJPf8
qscAxfvq6zVdA8nMc7bgsjwE1f/93BSm6sQjCjetCrOcTgU04GbHNrLku8iEM1kf
SKSK9LBD3fRAGcFjtQAAESjuEl61Po4BKYqrjKShSRmvChAx34g/nk1PuiLBthab
Fx3lZ8HRAExcDt+31tagSUgYZbmGFlNxnXDMKvYHav3we+I9HUlpNUvs7sbEH4oc
CArQ7fe5WByoKWuhOJVtDWUlM5Q2pAcE5hSETZb45m76odaCLIMLl9pw2c/Uw149
FbJG6mIIPhTU4XwPYI8jIQi6uq43zM9uBFwPf8zHZjqZjLiY5kJJ7HlIruKEzAgt
PVz3Ka3oAM2pJSjwlb4PWjBc2IdtoAiTnOK09NW8ltvqx67tok01jwHogJKeyxGh
Lbr7OQE3EVTRwpq0pb5A2xGSMDPgRyHdmRW2JAow3FPoB/Fzdo03msRDqKv7+3pU
hqFHhG9NyFHU1CUmYzRsy7m4wm8BCduvrGcac/x6U67JmCoPWFkfuulQDuY1V0nO
dMZPLtKxtOtTE3Frn+aAe3wvCswacivHXjRWvKLyDYij0Bba5TT06Ef30ic3OtrL
HMBsqnGT882I/wrl0yRuoWPSvDInmpQDMz4d/u94IHu865Q4sSPWBvVoIi9NGcsX
FPIB8oTVku8NkAQeoFFJeBKrhulDO7VxJ8nywsIXAasJm15o93NzdT/sMs6sU7fM
XWHf3eBNowM7JlEwSAgVA+7FH4qtQvD0Vg2Y0yuf37EXM2ShaDTrjzi/gapZynDl
lvGE9NdIAu/OKKQrcZJv8Ftzbz5WNOJ0VbHBD7ZklPbPfRJYysyYmwSisyMmLb1T
B6Jj1A2OrP4HQ6KWbaogRzHc+oc73VxcKJRn/KTrmwGfMSk1cxNEmaSXEiDLezvl
n9VHY1hV5aAAMZ5tncDroTr4WElphyi4w/HMYmWIrXLMFIL8x7OMv8aPzT6Ph2sE
NLlpxWnW8btKX+aKZTrssR4fVq2Q3mCFyI4/UDq+nNIeiTeMdcZUuUMW0Dr0ngHu
LX79nQ0G4q3xjHFAg9oikPVETKLar7SRjT+VFNbYquDVxJNvBU1WygxU+gpeV1+C
yhivAOFPPGxE0YQuplEg+fhqJGTCvSmSFXzIpvdpV6nWuF08olih01we2e2ln4FV
v0A2IwGvbTd2QxCUvP78ARjbcDfKI1KQnqg9njMI7FFNaNL+8bhkyc960ma+dvW2
oL+ADbcN+CGF65fHELVKbnQetU7gm4rmJF+pSZ5RaVbEKfRmZjs0H1Q95WfCqeBw
tIcYcXf+Vx297jnwPPLA5uXZPwXVt0YxlU4gaGXRRMe0382db5ayQ3F2GnEUNRca
YG9wsegaUoOAO0tTMnyJeptiEukpdwOcZfuHQW6VLeCQjay1uryIU450uveE+WLE
FvF2XnSl5lfQ8QeewCcXO9q0aB26hvu+bo/WkUmJGXzgSMmGo+Rn+B9hr7lT50l5
qDewdPLQDn+IcY3VTgCTmFMZx3VFcgSGVzCqFCt6bXKzfA6D70Osb2hry086NOS4
5JHT79+qFrHmXk6vmnmjFzUCno3bQwNztLbBSS1YMsR7p6jQQgpm7wDAyCcuqHxe
KoqSFUYLHZ2uqAM1VEl7cplpZrOejBaGcZMiKvTP8igqlznks+oKY09cW4nvGlu7
3graKmOdwZiE9uBNaI+i7MUut65rfgd+LoTxLRF/4F7oWtGgl3ZWYjx42TnM+m6X
OGn3f5QF0Cq5s1WZgS/PNSryNG35wR0BGBdTNuk3q2UTIx7ylr98AcTzvi5Vqcwx
QRRDZGIO3rw2d/Dx+bepEziPxSdoYX6UK9GVMrmsId5onRi3wxGbehgnWSsEQucu
Fkiaj+30R6VlGFbUUtmFXROnEqbMz8nKvqPuWmc6pxaVEYze5oS7pEVjBuG4euA3
ncRxPJAL/xOPur3igwBtwzuNhLdnMAFQqD/GY6bmXGExzwYCtBH0zztuqpMMs6BL
YcYf9uVrcOB3q5W43BCLeSjpZ1eEq/wEZOfe86BWhJUvqZ4bMQbBg6eLHwN3zUnK
Uw46YN4eVoKC1ml6gGd9rG5o/I1qzHcgixCwEVrtXhLvkeTv3GZ7m2EW4UNSfyDA
pyaOORJkzkbbD2kF63Q2Pt9W6iceaJ93vmdB8Biit3qEKH3itfGdz4GzvqjSxAUG
/4Irf4r0EyvxIln4Jsbv5kwXSxpJ2yFq0g666ZHFetEHPmzzAugvmGns5r7TxwPT
bDpank+uf7Jb3evsMWwQLSOhXGd0QUXVyLxYaeJsFdFwOzUblV+tJVeq31NfMcbm
rkmfKrUthDiGjD8LgGsD0ax/2MrHV8SWni2uc0NkehuE1BMEr8MSYsEGzEZDei0d
LURGioxPlb/LMVSbAjsml8OmHTSSCk6xGXpxDk9csaauhZip5BrtLCEXxpalcMTR
WB4nuxeW+VYNvw6rewBmsvzC10bsQ7a4r5Tw4rNFvY+5e4zTg0IzRUa36b2yoM9i
MJmqTy0jTIjgLvtvMol80oA4cxDTu1Gzy4eQBPf4kMUgj7yHD4WxLE1nTKm41CCr
CT/GhLmnbaVNmfrpN9lfGkMMDvMGdWKlCgZt4L6si6NkvgJleEXnyUS2WztXVvsa
63CSEp8uKhRz+XlxiALUVOo2TMdgU3T4ewz76BvhtlXXP2oB3SMN4CLfDzZznsQ2
vNeSZoTjpW0mIz41bGNk+IN+tIrvdb9K3zGwvL/oMACQug5VTkg/hoavhr1hkHnG
I+vjQM1qXynPuCJXcLHxP5W0j6RljIvQwnzZEgFE4gM7ISmQ5UOjvZQWXfdsYapT
Ua2pQXF8yRvJnw9hdmk5OiiPEyLh4XlH0GbokRQFenp7QQT84ky2La0hU7YXyNid
aRW0Hq35NtfQAw76PkEkDlsLCQxMVHo7Iq46QdbjzCoH76jIts7VFV5cSvRnIjgL
2Bsn++QywBtO9RJBvMbgpKotuNuQ3wCfxGRrQ9RVA2MoovV4fVLH7n4eEb8F0Piu
/CmHSUqxpuCTwgcp5sUs2BmxWFFhJyiS2LjbdEyunxAgRoC6ngBLaO7JLWeJrW6D
ybXP4fKrghi8oQlaMYObjDBAwhNxe1nX58dp+RPXg4SBslvK3do6TK0ob2h1r116
2xkzj+pK00f7ZctvpJSlZdN+ujoY5O56a5pdf0KnLX0wfAggGRFCfSe+hzHwSE4q
OS+lRUAYKWTKbWKd62SfMCPD53VCQADvD7bUs01R8dr/D5nK9wiG12TfgApm4gj7
PJ2BD5ekQFIywn2dK5mDZkdS5zEUImMlsBzWt+lDzFsRuF6na6FYy9RuWONC7vyA
jp5QKVDQJ+Kea4v2tM0iwGxnA3frG3bWZowRTVndkBq7eKEIU2ZOPj3hskjUym6k
HSUsVHzGLz45TRP1RXpi0Ya3oBChBBfhVHpeeErXR4oFk4zLf0X69n65FsYFAi5/
lL3+TiymJrNp/BpYYjvtWkZpDkXLx+tYp6Qp/cvi0e1P/ncZRpvgkBDKSrEKl/hu
bNnT3F9uiu3Hc6WXnlVOygONtnqCJ9ASMJmDmx8Wt/4pvgiI2xA/LU7hQylfEwa6
+wx91oxYYQWjWN5yJL6v3FCvJGi2ikoxJKL5GNv/8vU8KBnDrjAro8Ys6yQNaOPQ
QWHS2NQzHhXkW2wfLefjQR6CFwp9hbIwjzU43eX8g3IHUI+COQ1fEX+ZV863xTPb
twmPbisiF2KtlDJzbNtcM+DgZjlb2Xwqml0VJcywJOU+a2xyNQWiCjECKMFoIRE2
kLFRpAxlDYFuNsBieTXPyump5A6XrQqaxSCCg4mDqOjGpLVwLOhJvohYCFdhjWKg
HsvpAEiOOmj8jFha5LF90SYACsdAFo8h0A4UY1CSNtvDX/87fCBkkZ9ls8E9dOJk
YhuRl8v5Y8dSmQmMll1z9I2FFbyZW3FeMUtUg+jpQtSfdxrh5MKMYP42hYguiPD4
YBmmcU3tV3k2xdBCvBkCK5CdtZP8tNCEV6eFxJQfpX7rBp0vYNMggOQ40LN14Jhq
uPVNZZrozbYN4ZXnCPXGd5xF+NswXWBd8l3gXyKe6SBvREBY1wCgObg9URX7Lcgi
AyvbpIYqNdn6K04H4X4rJQJDuFAUek+IvFm7UsiZ+EYWrtdz6oiK2R7AwQmIvZB/
as8gxQOJlcyl67bvV5NDnisGB10jNIE86Mfhx+gp8/ilL877Lep2h2TlN/vQ1EVO
qo86jOF07jnvk0h8CTWKheSeTMbW4FeEymcdiyc8uc+C8EurTEm2cHTgGTkayObk
M8wE1Ktl6iJz//6A0g7ovFTsyQhrB8+pKGZjS1WFm/rCH16VoM1fMzfnYAVEGTj0
jusOJ4+Wy6fedFWfM4UrPX5k45K8aSzwxh8YcBlSUOXWE6GUmx5FtW3P9bYzsoCT
oYyLQkYsLrWTukQOTxIT6NxEhtHbJBQ9FIH/8vQqX/n9diHXooo7hswg4PKDDODe
UZpVx1cibbRaY37jvK0j1Twc9S6d9zQGFXdsmJW36zFexnHGtM7t5hINrn+f450V
DwmqbXo+qDKC8BXrUl1ldolGECnvRXA60zKEc88BmlnQxCTe3MaoLfy/hKemz4Cv
xPP+PqA8FVpRpluqQSYgwDtueYcvy30DbvGCfgBagEg2h5SfKyNhiW6SGcmprC7b
b8gQIJZdSc9OZ39pImod98OlQZeB8Ac/DGJl7yTX8QPr/NJM2zvjiuN689vnZjOA
ENM9vUFMfiKEbr3HSnMu3JOInSGVFBr83BDtoOrG3d8JON7tegWhwePbzxWTesJN
SQlq4CSfVa66ql7cYS2Kl/R5s8fLYGtEg9/EZVsKj/3Lzf+xsUQZmYbHzFca1PoA
lUrCv0V4e+mayoZmEDrNLNgkYYeuyeIc6Et5nI5xpQlycoXUr2c79Lofgf5o2Wr5
13rOyflDd6L1CWuoNq92UJsMzFkXDVQZ8Qr0of98jec3+SZzpcT1zrsV/sJwDGtu
pwbeK6NO2W7YnJdhHC4Ohr8eMyFpf6GmoUfdbok98ew2T6jJzjVVn7yVAyQ6RKVz
8NkA6y9PGb2YhPFSW7KPcrFqdX5rjxygiwSoQ4PyPpfpUaJCj+rP6ivwU+nGjxp7
fWoSqxRgcKSuxN2QVM5hESeFz3iK/yQ7JSXPbQyR2ArnJCThmgtYYDLg1SMQ629d
RD4V6JjtnRTlIhvTc3chAUmW/f+4D5pDyYn7dDFMA3ExWMJXWyhmUHgFahZ6S0jD
+4V6NGeLcfO+045u1GlMrdep4CQV30J6nZt6LbKW6hHya00nnocdEin6CQYWMCs9
U3n+FuOZStkQs8SFbI0YZMF8U5wHgwmFT7ltouFkATieZXRfYQY04WSV+JsXfwQ1
gwTW8W+hSq4QjG39/sfbRl0F+1A+tuQ32AjCc81g0jPLFH6H0/IgPFLrWiCvr+RX
9ravCINwEQnUMBDyJSX4+Sa3Ye7p7KwgkVtxEgGOQ2xVm2EfkjRCbm34KicPyQNO
fccr0+fQJAYF4eU5t8294gJHOKjhY6oz4ypRuWkanR0/tY+8L6xtPoM2hbDFuw42
U+Bk1RsmXVKqEMMGocsAbh+SDz+zAg97iIZBXn43WVePhQZ9Q287HJu2y+UK0j7c
4wOtnFJbXr1U1K6OBWnStBpWgTCya2uc4rHvsik4kf7/85AopXTpFcQ+IzFRZtwF
7Wsli0/kqMY/4wnWzU7kTheOuToQaTgXB5gls+0FrnwFxsnxExdolBFsHScuiezJ
+xNXun5spOQr7TQIt8UiJU8NFlXX8uMCHWvRONU6REH2/dh+DvfgUnNuhAVuJgGx
uxNzefqEr1cN8EYTN+xR8bh+xc7I5OpzAZDCi0lz6RiVY1LLXdscuzqR7Pqg1vc8
Ib8ih8HV1kz6Fcza/pjBF/Ym4lkIlVDGL9nZbHV0W3beZUWb5nQedI/AEbncvr6o
HqeJthsR5WY8ZVDc2xlajWOU2tGBV8vQFgDdPqaavZ24VVXVSeWP1uPhwopxHWUk
qhp+oUMeDEwIZe1xI3M7cXQ9keJu2a8Eg3w7VuR5MuD75e/OGTiIs75jSTYkWKRR
UzIyU4eqzQw716fmgJAjjA/+KEedcRvv2LbaedrA/a9e5qKry4vlTCQ+EfjKCkcA
dYgfQhCAYFuP2sMKucRPYUfUJMLAx+E6U3N8qcyobtwr/TZSMKP+nZ2FDn16uEB3
kUdCeZ31YNp6XKzWcxskokobjwuwEyziYALYIWQhiKsC3+U4Jgavrb4EPHT46pYi
sN6PWudlyV/Lh5k3/Sfv1oB6HqMtcTlZ56pf/BABzpU5IeYkwanm57fFfesuDiGE
p9WjV12zMd+V+/3zVL08jwmnwTf2pYU/xcco7YGSGA+o01lV97DIW1SysyxhUKIq
04kAn+gjj/xx1gRUOasG7vdvRYCe3tH0GoxvI35qW5lfhfN9NMCZk/ZAIUQRF+ke
6/lP+8b52wo93tx0eDavjdxd5H9E2p7z4RUrgHBFjHYVEZSaKZdNUrck0gmfwRyb
1zQl7PsjuHh0A52HA7dq7fFyA554tFkH2Yj6T15sVqGn7eSHKFJ1Px+I1wsKJv/9
5YNifj1odyW1oZ8Ne6Iz+uWO3MlSvV4WkxqIXEjTqjl5sFHggfJyziI5D9fWjuUP
aIRFBZP/UXWk2Oyce0IW+PeMUQuJPdOzMDlVOBvofa4IR4WWQvuG+Hat8U2X6fzX
pTgOH+qjIdTGhzcn9jIR7/H37k4Pq/urfnSImioxv6XuYVFblTMVQYc/4fVk1Lf8
/AfBAuT0R+uJ3uG/sEqwldJNJNY0DbhnywBuR/9x43p3FvLukP+5ehwzunnKiRbi
gvezIE6hJaiwCvNdn9FQstPJIkdGAPqcDcryxKeams1yl3FvVuFdD9AH2HIh9fWX
jQYkW8MxeV4TuXsQpgHkiYJ4FneHgLK1GSP4Pk25wsCeByUDKQ+hC+oaBI790qIA
XugB0NeEhOTuSH2KLj/ov6l1c+tGupCj6oWr/F8cjUtP2rfDjAKJk05sPuJuSj01
NWUX5EXR14C135QF9FyXSMeEfcNgM3Dw/6CLEk1Q+lhhsNcUZ3nxWKDJSrjbPSn8
+z/Xn/bXls3X/S6oY7ii6XfkZbS4+8N+asDjbtys7cWitnfv172iUjRR4bQlcae6
PIlpg7BFEDpiXut1kQt5Zd+h6Wto4var9pQlrG10uihq59TU3LZQQBKfgLWJxYP6
UkI1VzD7hKnrfwnaFtJeJ0U3kU9aBTQaWalzyAcgU9xBJdJM1lMC21XZV+7xqlL4
fFootbTrhpWgc0Ys9uds38BqBNMQ+CYtmux3+23Q4IUNPIm88MRIollqE1h3MOWJ
rmirUCLNNrasWs7NrlKnIJblFR8SQ6H+PHn++/gf1kvQaYEyFldjwCtuI2NCpv8K
EE3EN8iGL2weweYE7Fri12a0/3ZUd/N5CaH2numjb5U7L9ppIqbTHrFtiPUoGMd4
5ZvYRhKSRtc3YmO1IM51sQaAtNLU714mXLpkXRmTPbbq5uCm98soY5Ds45CCQBed
fIW1oY5z/yo9lXM2YghWgYrqUAPF/Deg/k2lj46ogh7uodDYwrzHAbDKpbRTUdem
jN+0yXcjfBfAXPv/W0u4Z6hi6+PmiWhnqgZ8hC2yjhm7g73jnaUhqgDlSJFW+Lf6
VL/msR0KJySY63TUCyp8ukXELTJ9sW2yz1jANg8/T22Z+vm67UEErEo1GCg0+NmB
dtyK20h0QzQCI2oGM3IHK9UgoaQmCFpNq1Zps9MDALAWMIO0J4nX5ECO6R0MQABm
vZxUHCkakq8wDziSA8RWisLha4kh7m2f1UUBGhTTiQaAW75OKN2YWSwT3E679qLy
qjluC3ZmDK+lT2DuJuZkGutcTN/acygRGM78Q4SIQg6eofp7ZNo1ew2UYeRPXc/B
C5W+p3K8fPLWpX1yrVhvPDN0Wg0nHuxciXOIRmSTobjlGP4Qun5W8yr3TTtG6+g1
3yrfdCXr1+Vj16RSgeojBEZGuv7k5Y2UHJy1B1qZ35soOpUKFJkjkw21oIGiSPTx
sDITs5HFGUOuSWAqgpCsloabClCLG/F0eLu8mqFngrIxvBQ3ZhTwaqj1VTONJng9
9Uz1KYFIubbLeSvUekASkva7oQGBomjyYWNziIjkKqrUgucAUt9Z8TfB3Wd5D1Bf
wXldEdkXgUhJVb+RzuAUP2Vq8lbzvIrlJnPVUJp1ZHC6iztQgWHZ3WtZksaL4W4b
ZC93q8jBZWHWlXL4g+d8QBHNxmf496Bf30GNgGDMezCAcsF2m+hROJm2sIjE0rmD
djV9xupJKMf9NOBf5uyy9hORxzfxa3mf1yOzXCnNBpD4KNUOXdJAOpLz82kJ6rO7
BYWocKFHXEJAMHyCjyZaX8hTE0vFvPWePoOaXAV7/i30gNMzBilbOuoC1JJeA+8Y
jOeIrYBcLsqWxTDEb9RcXUXTlclR3WYQ8qLxg1oR1ZK/nmyntIEiSc/RYVbMGFEQ
dgsSfGxKg5Fuwml+Lz0OqLHTstuB++BBD6yI4C4JW9YqQVY+qu5mbTWWBZYYrGla
QqIGV4lNouPydCwdLQt5fjrw3d4xqiK+ovJK4eCpobr6qg2j3kMntXlOBsi/S5xO
idlqEcePhtky5esCVJSGiFjoZoiC/oaFLJfm8lpJqjgdc3syq7eixYJpB830Hp2/
l0qylSeab6INW4efRHMMUfq0UqufngyHhp0o3/UveuUUCXHrqS7bGIXyfGs5SuGz
uSGkf3uQ91uBfxT2dSxlhzdGZBv/xoa1AWVJgXhfCQ8mf5FI10/FqdSzAnyDrjvk
kRMIs1Y0llU+Kp8njiKqmImvvUARaYLr3asI1q6uTrMEKw7wVjqNX9C3XlAfJfpP
FWxtj8j75WnGivQxwT5NzpkUPa5r5wSaTDvjQ8eGtIH7OS4yJvehSd5/SV6Z92x0
iLKefU9j7O7iSttiTYRidgNSpezXoGK6o/seLV11pM5oYLHDp4aULppzSdR1OcmZ
3bUfrT5E6EKYVV55LGseB5rAP6aZ8NuzQz3gVGoEyv7j0tUCHE6yHvihefim4fYc
ruSz4u9v46xRpULcO+hRTHyojF1hD9+FAopWVnQNc/kssbrAnEmXDmQK7pp5h12J
vDiO8g+cyag3PGstJhVgvV7L8RcR+vnLpagl6O9LrOuqUsJ4Tc8QjuOHZdLtgeVx
Zha5Cl+cJHOBrAn18P8IQd2FlRrIrUxrbhhichDHkXn4Hr0IIRCcZjtFXCmsE4Tl
Mvn+qOqUDBx00nG9BNSXY6G++L3KsZV3N8PDVCEAfTBVh7zEI6MPanan3L8sFoYJ
+mexGGJpDVzLbzIWKrREh/IHsYNuPmYuy5QlIzyBu/oLfbJRmorLbQLafv8YVqz8
wOBZtAGKkddD/GNP+TOpg0oGRh2KrlemmHixZDNAdqCKLUAvDwzSqBACHQ8nZ4sm
Om+LPsYKiJANHMLKCjwnZQFv+ZUgA70W9N/gXq0RHR62SzobvsHMSxmz3oCBKlta
GKGEfyNNI6/qwcZ0GS239eGKHNl8EqrIjl7DxzUOirDmyf9Hcrs3QTPJ3L9h5hRs
/GAeFG5RUUPWwGkjxZbr3tlrg0ZgxcNhQoUWU1bc1gBpBLXx8PedK2+Kvyfbv6EJ
JLhKW9QKtOXCT3SrYqdOUh+itQfiYhODGqHtFJN8DI1IwdOljEJdkbwAPyE3IL6w
eN+u26wIG8MHAa8cdJKsMMhM6w1cgfW6Ky+w9BYZJrvL31uXN6P49eMhwwYkCbQT
a6rUW31jwtspF4BA7Z4BinFSFDdFWcK4WhhC/OTlDWelz5lomsWIYhxTOKkWuvgk
JbP6BugYl/N4QZqt7YjC9uDieAfIHXLNfmPA9Q6s8EC22spFScOs2oJ487PDwRSl
9h5xvpPeSCnvbhhljs7GM3cKqYQ6Vo2M0K9H9Sl4gzeOP4hbCnZyGgs0RagmG5dZ
BVdcnqsTI3h4dHkCmttQzWq8FIf1105QHsA2SjK3xh1AM2ZRwTrVuzyP9UJG/44u
JiJ1ZgfYUHQQDS56qAff6n9qo1cZKASn+fHXidH8SjYy5jd6uIoFbaXo9xqpQHV2
SPUgYdDxFdDtkWAr8OPXybotDajjh6ukOWE6fsicAa/7nDpwr24q52FdO00pgoF+
mTpVrt/hrtiqsqMoIz9347kzxFxYWq+rJJAGORcWWOOF5YU4AuyPboXsk2jXrTIu
uwGi64U3jpNvGyhNZ1E9Kv7oz/etnOyqrk+N0aVpHWG7uKNWO25B0wJ0YrSxflQD
mePZQ6ewuY4oU6n8DnNUwvS9J6bsLUtsatHTxZTkC0pRQTG9vlTM3iDfj7CSCqWf
sN1X2cPcHLBF9X5uhvBUCVteecRtZe3PXJ/Axm0gNeoC4lAcvB2k425bU/j+FD07
cVKxp1NXuOCh9+5w2nsA0y36oy3yx8tzORz5Is3Jb4hZmTKI2EC4wCnbgk9Al/qQ
WJGG4cnsNyYuzto232lIq/22D0onHMwTXSXqdN6gq4z/dxORTl+b0R6JwAQm/2PF
DLh51dZSQ8aGg8AFAN85lASVn9ipZyyjxth0E2Q1WSQ1bvY6rylN4XcBm+n/mME3
yOHLqrlTWndNC7Liqja46lEA3oVCSCDg6rkKXENzNLbfPyNuOJAbA8q2v5eNtuOb
Du8n5dcXqE2fM+nKaBIWJFqGD5WSXcyVkJgeHR9zy/8TyBP83Znf+NVrpbg6QSfX
YXi+osX0tkuvdgiBUhPwBTT6zo2NBgq9nO9X0GLGUM+Mth0QkcicWdCgCf4APfkS
YxgcUtXo5wEJHUAb1VuxGuQswTNj9HhMeTGOufwFu8WF8KO+9F1qeXxUwovIYpF1
l4ct9cj22h1Ow0Co1fE8QjExKnIJlHuzTM9Lx8PpCgz/d2SyzlVX+/Q4RqwC+oqD
U1qFHDdzY8vN2IoUKvJW3I6fCqjU+AKDXrBHRQoPvUjgNAm1/rwXhH5QsWswcxJb
MSqu6sGinll/GqrCWhqDB/RuChMwt5i18/XMz5TU2QvthSmoXU8E4CtC3xUihhnT
5f6PoXuIReRlM3Qz+4V/z42dnDpGs0pxu5GHDS0TheoNTrx04Vuoyj8pXrCNs8LN
PCp0uZ07daPWN/Uq7EtC10BWNf9P7qsuButyvPdd+OXQPha6sIxcQnm/RCvFMTBz
QK5W2Yb9MOnshMntWPxYWy4ewS+zX2SgEUJx5rZTA40M1o6B3WERJwtqWyaqJ3IO
ju0cn2EotSc2NPOePcFtbDZjMrkKpF0Fy3lTWiQtS3+pSAFR9880sG0UPOGfBGN+
6lSvW0y35UBmN8Lj3vVk48gcZA/ZIh44Olk+9Y4fzIZ9HSCkM+DjiLGrEc7OVxpA
SUIJa+9tFoKISWxD5fbBMxBrQM0tnbhKKd63N+cVlz9KXgMGE8q4hRjqgsWUw7XL
eIpQb216b2yxv8oOaTPGqjRfWwrcHytpQViQ6XqqUHJdZN9IKEq+pb8OPwZb05xX
kL834hBoMyOBPMQjIl3b+uzXWawXa+/00/oH+cSudKCYl7RvdKGXqYY158Hyk6PW
LNJBVSscqY6630H2DnWuSRYGkhucYNqT9TywT9Oe8HNzUE3az7ttrjfTilYWagac
FZGqzu17R8SCmyGTkZi83J6Evbs48FHTL5Lk+cAlgzxSgE8S4mKPc7wgaNVeoRfn
Uv1duQt5J3z4Ylcuu5Za05FUWwcPjG4IByI9xQ3DZYRTekSXlLNXVnBmE8w0uYuL
Ze85d7AfmuVB527KEDLKTUjbQovXN6NBlyV8/XtoqwbGR354pmjUBJed40TMMSuS
PqpfpV91WpVLOsAnXH9y6pRXytlQueuucKQByBTIdHsXoqQvcU1YLlYS2NABuVv/
s3kkjVzaNBww7G3EaLLaokw3Yu+RXxEI3yVKJH3l9gHAbRb2MKuWS03AcKii4WeD
Zu9KFnfiQcShAkapeskH7RLaAl6lDv2LxaMv4vDLV7HgjnTiuh0Dxvxdq1k7456t
Gq6TRW+oVbVbazKd0cAi9jkPYgjmxCFWsNaK0EAiwuEjLFKE0HliRo4Cbr2nqOku
QawCuJi+hFIYKygLAxEDyymcG/X375W8oRAQiOTHkqwEwkIRhO90X1fWerT7Euwc
xkvmLeIHF5yx60ls3XFqIh5PDOEnI1S18u/15QeFQKeWdpXYLNAP8wC37DIjQHlM
NHtYu9bxnqxOIr/SUcAVEKpImhDUwSjcQyQ03R73O09RRJFDEKYIIy5Vfiq/NgqK
it7V+z9kXw2bkrn2yUIQ/fUs+7tuPK9m6SEv4SSH40VhxUvo7fAfIipyQ9fvwZho
7LIG7Jvy0bVLyHqlg4WOJiQ2uBXoGNWJl/j8jJR4sUGp/DPgRn/dRvjB770oZBa8
UhXgCv7QMggcNzR56OcyAaPglwlaW605NJI+VRTQeyNZt5Cf9EOF4o6rLyfrj+sE
a03S7bJJbjvJDlnemgKuswkjfaE597AXUzaFLcwbZ3HAqo7fgJlV0CcfFtx2k43+
Jfk37G3xISmCwWTGmqfPFfki0bmDAkIgznURgzfD6AMxCDA4ymLuli9JbmaNR77+
MR3aEJDY0miZOshzlwySwlM9k2ODPtBAwpn9aCr2s0MRLFEuPkFl/MQI23HRUjIl
ZmVasQm0gN9xqZvgOB82zyh8Gn219OBdXDfJgEoTWinzdJEqRy7ITq7LK/RWYaen
o/qB9WU3n9sR8c8k79eU3ZZEK6doQ5aguBF0Lttp3vh/Q9O235VC62Zg6mVXMMXM
zWAX6B94HeLdf2isqjbi2uxXsWv0GLUVcyYXttz9lWr4aZFYCc9O5DKRfZ7Jj/Am
K8SSC8snJ8c8CHIzs4Frii3LooJHA7riZYUOnslvt4zVBymdiHIOr990nULigGrZ
jiPOChoienLDBHnQxTBsNTm+Nn55JILNwOn6sfSExuopIYR+93i9inLNX7Dqvs47
hk5nwlMDgRGTWQNYp2Y14irJVWRvUIBOcKUoFV6j8O+RH6dDHjbKAjv41OFgb6RO
EXYSqR1c0pmtGUrCbe19ttJ1qbWHs+Fa1H3WlVfNNPEzAunuykQPS2lW/GoGTrud
uk4VieqU8U4yA2axLehjZNTZXxp+s98XRGKj52mkJDEqCygVPc5SlAJN+0xoQFkt
Pnz7dAn3TUDDZhsv/UvPxaTRwQs+MDRLIf2KaHGEkWatrAEjeQKw+qYzH8lm7JhU
HRYDj5rq45WukKqNzdUBX6oPHVQEu5AvXf1eijCXaPEiAha7TjsQh+nA7kq9exaS
KyWPLBWw97vFpek36wTcdzbLu7GEAuATNS+lY8CBz+iQJekcGDB8X0mCx02suDbn
nlJX/I7S86EJwsLo14V7CXKpoJTz8KG+f+Q3ZtrdIuBROF4HYOMZYJUCOkytV02Z
M4LV8qnvCHFPv7CFIYHpC2WaWp2QV1GCXhigF0r1Nr4IXBU3bk0xOU0zCShdiU3v
fX09nQ/LcC+ZgDSXi9DZoQcVbtg1Pk9frIvZF+P5X9+PQd7nqq/gAk+vtVzy/uS0
Bao2r+97hPgHWyURsaP4H2Gfgkk/HrREUUFcn/P6n985cRn7q5O8Do+ve4n/4duY
BXb1iuze/Fpxo1KFzoFnmQf28QYn9oxT5H5KcS2JdoS1JKXXq+JdgDwJES5AEunM
dFdudMzNTdS23Ql+GAYFwkeToVT28US0pjqdjRPK0EkiWKPWJZkj/6C27yRg/AK/
B0f9oOSmgkoiH0d78ObsY+P4g9BKcjmUgURAx8OAHLBXGsr8SBkYBCHs5q2QxD7g
MzcWGF+4w0nZsCxV7LdYqAdKtLuG58yCNrcXxlqDlDJSUSs8Qo3kLrUFxBH/jJKZ
+8cnrgrCVj8wsf9m4C2mhjFJhKA6I21QkTKl3okrnQZ+SEN6r9Uq3SdQuLRPridW
Y9KM6irgoLdiLoTwKftZy66WMSfKkVstgheki0OoGB3pnIAmJFswoXXMzPqRAq5U
WEOJsbm/h+9MyginSGoaWSLTg2+t7Tx1CHbHdFeAv9EUwS2X8IR106pHavhRgv7J
o4oJ/JxC1ZWVpK8uRZecKgSnKtygYU3Bf7vQrA15Vaoxh2E+NSEbvFyggezROXyW
qcTZw+6hTAZipauUOqbHRj0fbiuKLY6ayCqwP+Ddzd1+iqFl5j2Q3wxnzMWBW713
q0w6UT+1K2QMvwtAQPkNbPQSMzUPDy5ZDDdYf+YFPn1UiL1oYUYMFLg+z7yWx1ZK
L0kSRRvJnaVQ8RchTOd2AdcJfVPSJ9Z19BXs0ArjKh+VVq75H2hEuV6xKJ1pt1qM
1GkqqoA3EXvKJw1Hw40UxroLfyWTi7EYbR+lWNqrlEp0JYwe9MctXVbLV0M/NQ7H
IxDitvhrQ2i5mo1jLlIBnzsTViuuhhSLFXDO4IVbcl5QXZfeeiSA/Z0km+oJbrgo
2kXHrhbMlSxjEGrfSRrJZnl5iUNahuk+C9CW+R75F1kdzhAA467bji633vKngW8g
+ssKZZXR6XdrP8UNakRSDaPLhbQEDmAEerB0T0hiMCSmbxCmUrfs6ayhr1CKzhKZ
NV/G13kpim3mCYYzLLpsnPNZNyE5ibQBtpPwLn+T9lG165SY6fIKA4CLepqkDvfB
OgR3F8Md+76O6QBcc6CxqPGUf0Qsi9q5CvsSX87RzsR+Dsb1fBxOzLBzEUKHSoc7
AK9z6YYbzlF/F/+ZklGgvSO7uDD5ZbDQS3OcE0PXX8XXaL1gFKBRO6TCR+cNXQcb
2yRigM0yuYJhww450LUugPMZJvrhwbA/XxBwPr3mEKZEXwrJnHCLbQ9jdY3ytTP/
qKuQmdoAoGpFjaeDBHCDrMVSOnwhkR+yrMTz8N1xyh1ahjxWSPCgRzHCgFVieqO7
uI1JbRFoHmGPKjcAd4qteS/DQ9+56IpHFJ9YALf/iJjeq9q8epRvmIFZkf1p28+G
FJ/05E3bj5648iqtL0xlmLxLI2Tg7uD5VBYuANx1239gEFCCHM2Nw7T5OAkpKfWk
Xw7iJy4rrRvEYuMWxL0yzcfCymR/MH1d6xk3T7uhujEoHpL6WepXHR/mbLgvNLmh
NvDgYWvwem+RBfgdyGDA/opQXyNQ93Y6LNXLIAIJgTA/1sNll3p02jBKlqHa6vDN
TMbiAs7CWTCrN5kBEnw3ZtNqNcHJ/KycHTDg041KwKK4Tab3BikAMpXrEwjl7l1E
Qfoe8pPLJts4Pw6ABVHi4ssR7GldAcEHPnB3rtNKuPMsE2yc5PSjAi9Wzp/oRYyL
fa1fq/1oRnVHR0T5w2r2QTLblt4o3b50BdYaUVhb8AEV2FNC48aW6l8J1gu8+djG
JMaM3l5pKLA36GFfFYWztKH9vjjhpQ6ENLZBg7QlSltOyG78VDTiqAISCdfNeKsh
STFDuWqVD+eGc4MNqWGFWAHpl1Tm1k6txWEcHnti2khwNih5rhwo0YBIFUlsXkM0
29t4O215dafmvlmGIbZJy6PppjsJqfbhn1DPJ/RqEBCpw+dLjkrJwnn5ugYj+a+M
7LSvSy2C4mr8UOeOydpsZLGQTtuiW2O9/RyENxoebRuV8tuNOnu7qi2IiSadUuH6
fz5LJUIR31ad2XV2RWLt0dLRX0b1qNutvybvhZk6fhwsRDwQZ0CSOHEBnvOoZzmU
upzRQPSKW676XwmNlKDSDXzgehkyDjxBRQAMY0qXMXzcTCl1sl8dxxwWBxOHYpIh
OoGkUiUP5kg36MvVXri7LO4mLyFXSSMD/qV6ZvoQVl6hvvaSfOH0VtBdRiWCa3Jy
QAmNh3nGkO2ONKXa8+2mcd1T+TlDwsj6tHoH6SuP7A55o4hFDiuOS8AkA8ODB42M
MJAWv31Jeb7lFEGA/MJ0QfrtCXC/kofL2r0lLNdudOcLGRL0q4eP1wQjnAatVkOM
9endjbtNSk9t1zuuZT8TmhJzkiWCvjqb+sIoxWMNj15GBp/SbS4vFg4sqxH017rG
FQHSU5aCwLSFEW8KZGSwaDU//9KNZFGqqycpKv7CSrvTeq5BcS6UCcJncu5MPvYl
BmY8EJHF9tIA5u36oxmfuORKp4+waOTK2dx9QeYhcfkVJ4mrCHrHYLVey9hdzOBc
3aIBwFxwqhl/VGc5qRib0esJYNN/IvfebON0CE0GTp9tHRF4CVWvKw7s1XZ+y5cx
bFuEUL9pgSWeGYIhRScjizLFvxva2QD1Y8M+bg79NnXEWUwmiOOncYXTuIeUPh3P
EO+xdg2wqmBQ+KGhXWcT8uHudoX2c19KupW3ZX4rRl6lvSTu2wSJbGUfNtcjZpTB
6CtMZG0dlSIjzSwZ1BdKjYSy8agseFuauwNqNIsHrgTEOsO/7UNa056Qi+jmmXfA
6kNbUI8AidNkUKrNtv6C8O/dn03WYjS2mE0UYkaTzjENxZqFR2PTeQS3lO6OSFaY
tP8v1ciBN36q8TYX9HCr3Q==
`protect END_PROTECTED
