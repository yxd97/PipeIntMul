`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRQIYJdCFMQwCzPMOC+e0C5prlPCXfWlqBR+ygkShToeOpHu7FO46IkALw5qF1/1
pjrLl06h11fHv01JXRDdlACls7WX/+cOmCFuR6IzE4QLOPL9dp72RWdEKjsVbmjN
VkgLwrFgHRo3kO8GL+pqHdgV7AEYkKKdqsJpPno+Ps82zbtWKDEs2KPp80U3pNgt
R8uqkdVEEtGbBBRfcwY50/HQViei696lfDsBEWdjh6K/rEmKsond7WVbzWSuvD9L
uUYAiBc6jROJnXK+cPdSAk1gWrXAtQpI0681TzrMdcoZBjvLq/Im4oCHUdkg89b4
hCmqB+EMtNaSt3JWe3rqGQ+70T+z8A3ltJw9oskmegxIDgjK8bG2YeWLH+/Wp1xn
UazmFsKVqruSXlElOi/JB1mPb06Q5WV6/tUjNwRvaSfH5s1Odaz8D3k9d8QI7040
ovuyCoriBIFLrsaGnHVktVH/Wzb1CV8XqsuK8byJRuxDrF4zmRxv1KWCmTem0+6t
6GV2roc8CpH8qfcImzAew7PMQB6ZxH2jVZV2Lgx00O4/0HWjuCSfgp7pbA6tGjW4
7jHidmS43S2YoIK511uuKdH3/IsiGnhvcxi24yjLQbQCDJhL1fSDianje5vkaYFV
3VlT2mVVZRGnRITbrtF+U+R8+rX1KMoBdXywcw6+uq+IKKbcNXao7geyG4GGMQCo
/0heJwIYErm9mNWD+f6eVTa4ZN2pxsZjWyNYyjHsnB5qnjQv1dLvHB/XZiRLo+zJ
1iMZK0CY6OfvgrC/CRMYkhfexUDQ5/A3Bqp3rfj3UfI+tJa4/GTVKdNxBRpjDLfK
7Fcj844iKtGKzVKGfKgtzRAmkYx1XqsxrTiSjYnXRORyRV4XKr6dBqeIHf/OlUAb
Zw+/BsMFj/Yo5D8KoWfNfXaVhXY3I3L30Vc3trgSjziih+u95kzi0l82hpY2CMSR
rRWNmmuGSJgZlBF1I9jHrBpXZ+Dccw/fQActQudPlYr/h7ILhGPsyrMg5c1oSdgv
wOhAvcZqvn2e7YVUe7sbYW+6PVVZBPw7o/bOZsLkG9kxaoVMbNUdfE4MsoJf5wc3
Tkp1SoLS0/3dIV8aDVLDgd/9czFvy+JEFkU+K+f+HtlsQHWc6RQqw+ZL0XHz22YR
5wGsKnl8TqpqRAiy9W6FT+pVsnlz3UFUdz/9lX+TQyX7W/7b+9W9KOY4D+0HkgvZ
vXOT4KBsG+b2mubYMVmTlt0fvCYim7wAOPyd+o+LTJFKV2JCd7DGho2yqIX6VGqu
mp9RNWpLyXrhFErGPrXSD2BBq8+vdoO8tbR7e05VZBet0EJXzEgZPXjbsk54a6mp
uwsqM/oMCIC+m0N72uuwHppsnEnJc5kKE3BEQ7W4GdKqz+hrqk+VN0poCi0iYocG
L27NBWuG6yJhX3cbNRjRcY/dcJNpU17ivdyDB1ImiW3byWWbIBxyibyND3xvum2p
98/9OtNcvWhfgQNCLxCDmQ==
`protect END_PROTECTED
