`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b9Ep9oX4OgYClP/b8Aa7yeBKv1f3zMQ1//iLd0q5vbwquBhYk4Jw7OQ1CvF7BEu8
F8Ws4LhdQ7USY2eIb8NOHSyJEA5hGzKVPt2vTHMLAexQBnK6xHmFCgnhWXjLp98b
bCyg45jJLuudMBqXUhDpMRSLedZH+FQoM5MC5uOINkaSOEz8y5Jic8qWDUjuzdH7
J6MSFQs9czotk18YaV4gABpsPXmatTAUJzM28V2PKtWwibQafigHAGY3G4rKyGvs
gENi7gkOgAf+s7Xi8x7OtpeiW8naiGl4PvW1hhAx7uUuTqyv9XQIpAbkoqr/rwUZ
MZFjB8uiGhct3I423OMbocnqHfirIsPFpyeEDe649YaUaP5xeOAZeJ85NmLdaQr+
FiLCOMd6Ib1CPybhFtV48SqzGAVcEo3/Ha9R8CsMfnNNwXAF/SbUcJ67qpTTc7Qg
BVavGdQBIh5ZeD8Zr5ba9OAi6mhut4YcGhiIZmUNH/TUo4Ko3wf3S8a91BruRrJR
z2MRmmLp/CdlSGWrv9EXuhHFJm7DOP/0dP5J6VyM6zbiii/Pi4rAFZ+XS5OMUMuf
nUztjNajK60tQI8c80iEDRfhijufuf9CZkQwXaU1mLA3SldXfA/HM43v7PcWj6J6
+szRSJdPyzLty0lyJk3BoMUfwSN6fikBaATtlqdpG+e7v/gqUC9S9yBpTSV6uBiw
`protect END_PROTECTED
