`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m0YBV4c7uUSQN1ZV4RLlv6CXAHSuBO1X5vlzXLKS5+wFJ1GM1QaelwlCQp20uT6W
6zwOCONmT8U9Pm+qKB/s2hBZ9Ksgb2PpKH88qgETtW2TxXKIc7RrQht79k46W6gA
ucJKc9MZP8IqNOaZToPUlAoiY442Xy92hbFlSdrpizEfXaUDTgXInDr/BNQsVhUn
TsPj7G7nEkWLrP8Y5dnbrbnuv/MqFe/RNtAmVVcI/iooPhWn1llLNDoZB9NqWtxX
aZ0ETHop29ndiBVSh+LcxzDceJH2BMOYx0jRDVp7XCZ38iU+BYWSYaNRtw7PNR4h
8RIotI8kDfhu04f2f8WnD/BkdJgKO6+4HKUNHJS7KkJfh4CGi30ReM/eNRWjdhbh
eUPkM/6pP9tgJnoA73EAwiy1eWbEZ3dipapYNSAk7hIJ9rp7LjRLsuIQz31tgutt
bkdPbei10iDwk1AYbe52yrx3yxoe/vj5g2RfxgInclfC3N5NxRbu1nD148J+853q
`protect END_PROTECTED
