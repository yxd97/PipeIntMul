`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JYAbZ/HvmDitFWYYYe1rkKWyt5UbPz9EgFHHZb+BAbexbcSsTwGQAB3FdI2kxryy
rlnY67v45QcSv2cGIS5vaXj1l3VeP7B0UsU3HCK1u5Hj5Bpe/QLepJu+0ZZiLW++
Kbeo3xPMl65UBt4bSIz9fqGK2+vg/Pk/sOO8JdlI3v/A84WtG7ji2SbcmEtSHO9z
gJsuVgGZz6HUmnMQyOEiWnHY6TMidGYCkPaLYNcOcnTJV8EH8OimZ88dsqS0ZGzP
nbbvdeT0orlG7T1v9+vzNzzqk3a3WmeZ+06oOVP+NCONCvWAL8myK0WvyyHzH/vM
8Zc1tjvjkhlqqqMk6XRiUA==
`protect END_PROTECTED
