`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkHaF2toezASveOMP4KG4eXsZ+oMoDyXOgLdDy/fzmHqFFrIdn41lsOHJRu6KvHs
8trWrpEaWtdZ85mvRUN1KZuOlKJcKad3CBFXJ1f6/DWoInN/ms91FjyeEg0bbHh/
2OeJbUwkngMAEw5Ac1R5lLXFimdeXQLVhs3BTFywGlOv3015fBRLQhC35h0oJzkO
p2qeGdewcdzz+TwDhV/glZKb9pcfKZiuNGL7J6FUDF0XJtEsYSeJ5gszZhpKtaty
/vV3w4VcvQJfPzB41VoKl11UKYC0pf8KpAPIwiQtwqMsznIG23aGyCloXkto33o5
aBKRskUKBtQAXnCioMW+7gOFz3JAEbyIsII3uznJifErk5GYrkViXR0brYjVTGlv
wMuFy1fwpnofKF9b0+sGwLHt9aR/+ijNekOAlkGXHOTHy1DmN0/ULbTDybt3Vt/H
ppzH0L/tfc4dLe+0krYmCzlXYsm+Sb0rE9+d0e0H9RuKLOpHuHAk+R3os4FP1VPg
kXSy0AGKT6L5m8rZ0gMwITj5Xa8MkKkI4UGxqrnDD/sNx+L/FCy1EiUGoPrpOGjv
k1TeKVzaNhzNIH1EGxUPZ6aKfQFJT6OXo1keqUjSHynD+MK9vA+PcGTFpZhomW2R
fKykkrWlzSsryfK0gfNZKxbUb1QwW/EF2rJ0WHoJPm4HcBJDFSV2ryawEG9oiBq6
otNYXZZDdKkbdMDIxgAmb8uvBWI09XDRj0Js/fa/5HA=
`protect END_PROTECTED
