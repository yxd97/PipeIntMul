`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZDhQWr/R/C/py88mnF7k7ycG8AKukidHrJXhj7mffHZZz2rupj63HQw+8ROqQ1OD
EslCHboch1JBzqPAOfHtU6jhz8awT7N+f7AXE99m3nOPYqH5tm0PeM29QSG5doN2
znpdFoaWi6Ck6zpra4AF1wltAbAGpNJNeDvUJ+H0kPFLEyhTeOvQo3GAheIGJYIV
vjZfdlF4KFm6f/lSYhrREQNBTfPF7uaeq7HFOCllIUItMLwdbk4n6U2OitWm/Nkc
p7BATphZ5mB4jyqcsgpQ3bJLmBZQ0oPR45SbYYSK3+UdR885uNimBkzctCVzXUlA
nGwjdnA2g+3/j0dLTShSKnXeFlNSsD8CRj2Bsjj6frNOpXLCsTtcc4lD572uaP1U
lLk7bLk3LTJ1U26xtlK0MUKtzi5vNUi9WqKRCuucBnveeJzB43a5AU/MwfDp0OcL
SnjFZKzTgSauizTjBYEYGQ==
`protect END_PROTECTED
