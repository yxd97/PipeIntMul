`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gn/wn5OElrPNM1zW0SCTLQSpmLlfe5UubfaGlgfWbh+8gy2z2J/6h13q6SsVe9xU
UA9oOzkZ6ue2fX1HQJRlInA6EOfg5QCSIuhZKUsIm3f1sm1cJAmnkNscsMsY7I+h
BlwFmemoHpcla0eC0SkXKXV/LYvhk6bZgzBLoWQnMqnt4BwJIg/cC/uMkorqeCJx
j0v8cFK/pqDwYEdzSysgpROZMBpcUMzwvuqEtT6cUzUkvPjwScYlR6SLcFXkQJ84
aCMWCZHpSFH1qAchKgZ1hSdR9E2d4h8xaed4s3nI0CG8h0KCzBrhgdRwlXC3PIq8
4/2KL1nx23pDAKZBuKxt6DuP7ljF7S9gGI/pVF9xY3clmCEEYts4/FfdHmPYV08w
UFw7Bv6CgeSGWSsNcSZAHJuwCastTVOFKsPKswOMx166ovFFPcKgmlxziuJPQTEW
sOreo02ZdUHrpBJfE95dezSbXTAw0XXzL7uPW5tlyOL1kDd9Z8vb7KKDQDhD3hDS
qjk0ISZilytAyHQn2+A7aIt7gfklXPQxMofdLCyPNz3ro+bBi/8l7mZkSBpEda4o
rDC7xD6POx8QorkCiGjJqiwaI8P5rQRVizJy1LRO02wB/qXpLt4RcLa07JIW4itZ
sqTPAUY0efIC4kDHjQE3XKEEAMETq8irAXutiur0rIE=
`protect END_PROTECTED
