`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2S//slQsYoKE1oliovD6WuVAehoxtzDGgz9hZqbAqVpIqOHIr6vyovJxRzL1crQ
I+KcRgL5ERNXHW3J33khciTy9SEMQtF8i1OtakchIXo5E9ixdDD9fv5upUPW4B6B
bnY07d+3+kCL14Rahw44CCQnLR57/TNtMIkiCJu1H9TqlYux7+K1b1IVMOVNJFfh
muO164t9CXC/gg+NTG/n16FFANilM/z3utxBQ7QfdfXuQU+eOlbiJcSD7HyrnajF
o8iXqDKeLhMlsLsPJpZX3ZOnwfs1ZXy8rCuC8AoCcI9oQV2U6WzG4jGtxIfpD3XB
g05APZo5CHjIDm0aJQz0VGBkci/Cc0QzJaAgrcyUVXOTcGpv4JkPMucJmvPhp00Z
mHSEn1MR9A2wgI5nykAwmmXqZLcb3m184Qqbja+ALod6COsl46sNwmI/T/MC0K6f
zSY862/aSTw4xn/WFJbvuKpIutLGWkeFZJ0f3dq1a813GEqTrlWXWrGlsrOLztw1
CpNPVilqXuOQKe9REOjPdaK8pEeKp9AqsYcQeL529qNSZVKxNb9hWzIYOuSz3bxb
IYEwD/QAv69ggVJu6OecFwkEi2a8sEcxnppprGBkH+6kMLY1IZYXOtomh47jXotn
eBp22am9GjFXB6EncKBOiBz+RgBuHgyf+lgOxHbPJQvU05Zcr7cHgOs0hB7hBhfk
fJOTdXPCCK7awUQMQfdGbWRIPsf2YwcrUbo2ZbCJNc7gNKB09H/6KUzVVJixNVPI
`protect END_PROTECTED
