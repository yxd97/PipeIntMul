`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SaIK3DBrv11rfrQGHBQ7q6/gfSwaHlYhtg7OyqD8m+vnRLNvXW7x/Ck6+ry68LCN
b2H5oxtOuikbG1Yjvsdqv9JjyfQVm7gQ1rZa0p4ZJM15Suyp2WtL+hSkt3/OqaIz
Z5I8yu07adfFj4LTctiLr0jeDoRcjHaMc/RPLwVjMCRjM8dkl7ZvYeXLGrVMmJ/a
TQlxjK/pJ6OoU35QRteyBeUKy8B8ff8pCVf5sJS8AiryNxOsbMV0PHIsHurDjBLE
tcNc+w4qKjtSVtw1+d4TBfA6mUBk+TNmXcqtEETMiH81mMSV2UR/DiJEui+T8m0j
the2nFhISS5j4tWprPBYyMc5E6QTxPEnDf+qSNYAjdSI5pc2KaIts8P65rPwyzQr
hWlLViuLtJYnazVz6/oZN17a2rBUH352PBsx1/ADYv4h3eTVCgGynb+4GfyOHHyi
gc+DKGhvp9i8/h0EjomxejlJraEEbgPbfxyOib3YZbNlpM06X7WvUX1qWcJraBA4
Fdc+W/pfWI3f4zN18u1LlhFDCIRBAg/5slxtgI8mlTlSP5lS9IhttUdluLTK2ipc
sezspsoAcnP8FCGULnwZgamMwkBEkXwdhltF2lOWwJKd7aF4WbfUuZiGPMHHxEnC
NsToiJuGLeGkgZsDFXSjHGcCir09SvXTUeXCFUmRCrUsFq2nkBtDX/JdhqLo9rQ0
/oz0unTHtfXxRH+c0a4GbjnUzCZl8Vvsdd4EZlNeWVVawb2u5axYwMElbdcfyOft
4WQMkL2pFZiONlPfE5h7fs7MsM9WtZzniRr/Q4SWtrDIB4AywyrDaQAkDMMylTb+
bzLZ5co+V1N2w5So2yFvX0seM76B5lVtLiBiKCTULYDh+JFGh1C/LSh3S93TaNte
NcHADuFYBXyHoLAIYXbRqAYknoX9j/X+hYBnJNSt2q8IWmAaZiSWof+qzlQDDYPr
iFWnVTKScfz1EE5tedGKIDp34IouwbROwdVNkzfCs5klRURfXLBFyIs20IFBLSIx
7ZI3kufvnI34hSFijU9gbncACUAdw/FXPv2RrPcIjXrrYxQdGczdwEybRi02v8AT
Ht4v1A0hJtHP1+feMh2ePY6Lu10MVmDfr0NPSQCYwv7Iu4GEQilPclajoR8qG3Fc
f230BtG200GINbMGFu+LMPMq2VQ/gktVEIW2Wc9oabFAk8nGT1QBxHTHbDeSCpSs
vbweoDUIjjVdrxe/oLfM04/m9VOjvJlrh16imCtFuh+J+i+mRTbMkHqZkY6HvU7e
2l/05lCXOoffrrJIYdRuCz2IA3KZk8EYC2RBHJ0RlPpL+ioNmTJVzj5DbLLUoDKP
Kddb1xZgVIZhzRIf8QAyGEnTU7DdAV6665ka5t6OW1rSeCTfWDnOhylFm7/GVyZp
v7BGqdl6fanXryjb9orGFzvxExGgK8x/ojKNdJFhLUSNGj+wKLrkorbWtSauE2MV
7lZ6eBhmR5bmLCSQT128p9uO1MPuTKf/VjpNCnaEy3Ps6dDCHBJFDCcaZ7ICwkNG
z6NyPe1eoyNOTtghlP6eJ1tvZ0CMZsCJ9FVcpNRcXpU=
`protect END_PROTECTED
