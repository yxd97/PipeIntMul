`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNwFbU1M6RO81SzFQrJ7eDxCZFPa5Y3nfELTJEVvTd5/P386q55pBKbQ7xjUyubv
nHgNl5K1VoNYQf1Mu0mUzyyeAFVRPVJxMEHCuBReX9k0NBlsbf4fpZp7/0hgBoWf
Tqdkpqgb5R5TDRWaPfxbUP68Kbkk3AnicajGqCpEROIatoaCcj4OJEw+tTDKMVqk
zCkGvX3m2zbtt2fs1J7ZwBbEPeB82hn3AeFsbt7d7HszNkikur2k21G3F7tuKVSG
T+T67GBZhS5MeNsQXgW/pGoylDNaXgefa1jZe7rTPxW/8TTwRTSAzPIPWN8RuAN0
gLIYVPJ9Y6XNuCBhELPxjafX1onp585T5mt9jnXIs76hW3feOsNdWe+Gmve8/K6E
4cR9VKlwzJ/6llNfPzacVg8lh3BEgwEQWzoMp3MU20SvNoIo0vAmom+ZsPjtOUi3
ilq7krSRBYNnRccwvd8s3t7LL1XCUBnIh+4ZgyS7VL2/AzA5YqRw9BdISHGot4Ur
DtkpSwvkZa8D0XM6uDC5+Sa/SmucLT6RLzlZ2SfpiuVmBLyxSQYBmcE3LCHJShKb
SrAh2zQNvpz1zYvgVo3aVThKa9EAWnPCUFFwV+l8nJmKaJ9yr2Yu4L4QWSK7Ki2f
1rEXNbOkIgb6JjybMLL7jEXl0X9UwjKlye+qXePS/L+IhsdCX4A01LMWkVeMHyO0
HkVoSKbSBqUu1Omwz2J92xSxfaeHgLgUz79Pf5I8nXHO/Kz6ep2vGC4b3nL2hlWD
P5aDbK7o/G0EjLmFc1b/3sGECJH7GCBH0Uipanw0Fd9fRfh7c6dApo2WVsaRruB2
XGjzoDV+HWLQJsKGRJxJ/DCZLp03JWFRnDS/bAn37vtg6dXu8XrH0cAEOPfEZtka
lxwynkcYbDDPKr1m87FoRT8AqJ5eb50tdFfsNmhxAoC0t8T5Y/vgIdfBI6D7g/bF
j2GkrBWCfmjYfh65ONILpbNX8Z+HyfbV0xeYpdAC+v11hcOmVY8aAzlPuZo1zJd3
ntXM9ZrtUacIar6saRFO5BS8ckAPQMAvHC9Cb6SuaO6vHIbST3lLABgXia4k7xMB
WLhHFs6y1MXiWj0S+VX4UcKS/Mq0fNzhANLog5g0QHC3zwCi5noiUJEa7vyPynsU
`protect END_PROTECTED
