`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
57nvJjav3OH24cenJIRP/iQqMi4BythwC3G4MvrXFLtNndPlv/yBxOrR57PQ1Jz9
F3tlAQkNeFMmTIve7pxBMI8grEBdUIjelRtDb170PdFlvhDxuxHd4hB2edWLRcl/
wQop10pNsKdghu6NzsDp/ARSzP6k0BGM7wjukB39I8oCDglW+IKx9iEQMjphBlEL
Zl5gPdgBL91El1iizm9z7dBohZ5qvFsgNT3ZMBCf7QU4cIK8GhuHXBGw/D1uECzz
3UrDUFSLlFaVGjDyYsgRCm1uClFE2Na/E8mbAW1hSuPnTE8gJa5r7kjVyE4qHAuE
3iwpzjwoVqSniJ6SY1S5i8ezIQ+cH3mul8RQ5toXhVEomic985f/+txqOe/wtO+E
WUYF4zlcmsj6gAzwi6gSbRXy1WE1jPJ9Twt07L1IS4RDj2HPY0+eP741O28S7zij
ZjNBRIw3ZkIfme8PPycTPsLwyjFkmBornGZeHp0S6K3xTHY0WqHbNo4rtfDV22gx
Mb15b6jmNdV6zXSNB4cJqWUc70wWkBHuFquMvxicDLBNnT4GNbO9kORoEVzs7mkI
fk2GhpYDEeQeMHBdRiCkGYVCXif9uajk9kCcF5lmBA8AHToi0n5jviDWCkCHIj/j
MgydGPBTnnL0VZcveu5kyQ==
`protect END_PROTECTED
