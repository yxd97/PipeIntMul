`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8uRiklW5cIZ9NYrzbed8iL0jPjSFsOmTpjwXNru8mW9fdXZgWIyQhg23WHNIytqw
LNnL1kXKWFYoTfVaFFhopSEwS+Olql3kIQeYjZEnD5im6zy4FScDNPWRtq2Sp8qi
B9WhktWJBwNYB7NQ2x/5Ry2VJVPDSo7RdWEx6sfXeVYJLO65ZeycvJLKu/R/IOVr
SOCTt4z3+FAwdPVtzVzBw28Qx9cgh8CIqVd368FUIzcCdVdu23L+iM+Tt7I59nyQ
gLIL1lkwOlRV5WY2tjUa1Ft5EgRjsD9WdDUUqb00ocvdL8Y7Qsrg8XjV0irTcl6M
RmC90uZc4kvY23shYJoNjovI1f35Hq8S8oNE5mys5qTn8asrE1n8TLlv97P2FJ6e
0uL+7pYulLVJiveX3HsU5BURLknrUlBtKhBP154PzhccL+0EB9maYjpV/IZWi4cd
WqsrSt1dTObvxYyMsoOHRA==
`protect END_PROTECTED
