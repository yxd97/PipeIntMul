`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htuRmvpExeg0U/CT3ij16UmKfQUBcEuRj3NHcnlntsQ+YhCoEGxg+/6t+BJuqaeP
yQr96hZSeZyEkqhL4+aYHJwY9wt8grXQ7ITL9Gn06RWlKdFYmRvlJMGyAVcKhd2+
hMAr6NCvXhZ9TPxWjWpFBgQ07Q7ufPRTWXV8SvzB5biqoNryyEU0PjgPGeWPv7fA
25/mhgC5nQ/OmyUAx+a3T6GvkXy/njmdxBQYFurUblwSl/XQZN+8mAYhcEOD2S6T
GfvqnCcpj5Z+j83jVtmG9WguVUS7t+YGRn8Ek5SgQ58i1tRAfp1S5wz3/J8x2a+J
TYNdcmfFfG9u2NFq3HbpC+su3f+bG2/1al+rNvHq7kjchwGWTLJSFKSJyaeATfPC
SPgoMK3icIt7zaXL1GQm4KSFle+qw7lHw+PP8KGG0ZDfIQAbR0ni8+ZR8Ud0EZGg
FiijBxqGS2/uGnjx9Gr8c8hfryYz4d65zKZ0qkvCNsv1UM9/Gjs1DmyqgaR1oihY
ywjZNZrf1ZJMJkPWiQxyxZAFbPw2ZYetK6aPnjLMzq+mKgb6/41iwopUdYA7Slt6
oFejffrZPpfOyhp4bZUVI74opjivXP7lF8B7ofh0cBw=
`protect END_PROTECTED
