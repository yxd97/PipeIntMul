`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4AsdTaG7aKcRX3hEHhklfcQI9tj3AzQnHHXhJ10Mmdd0r8sYocmwe3KD7AkrSyW
fwnRnIrmknIYsAbYdRuWnPV54exgD8Qlv9UhXAUp3tFQMjy7zm1j8g0SU5is9x1Y
kMi9FJhH4KkSg7y2bl0YtQ3f1bAjBLWFe92oog5+f2vMWUiqrMA2COcpbBnv6fO2
PL5bjRxYtYbPGZ2Ww0rO0KTfgXppbAjsa7QXH6welHcvSpi3hon78WVO+kfE6Q4g
mSGioGTy56/wzQCgpgMrCwyYylXrD+g8s0/BzL7mMM8Ny+UF7eDbMCgm1LdxYfP1
iUKaylNa/iq944xfBotOrS0lNHPrBpKmRGezXZMUU4nAiqSE6nM0WzWcxM8MK+e0
8Jab1YKsLgBrDpdHpBdJybrxVYqA+ZLvA5hvBpNLMX0B7xJMMNIn3gG8yhKv7pYj
tKflS3QqtPhjGyAfNR2e9+g8bUAtzULBSlc3y9WmvwQbUonX59WSH85MYtm+1Qlk
L/40GBP8S1GROLPWNTyy7VJVcIGs0Bd/Fzp5N7KueVPhKJKCE+7600BgG+Bk5t4W
zyhO9CeUVUI+KciXMZVVYQwy5eY/8GgJKOP6Fo33GokQ2JD85ITALQZGJvHL7xy4
FZOr9itZRgoLZriEtOrIivDxUf7Mkhhc8u9eJXAUJsCxNtq1lHglE59vtRACTjjb
8KwH02uhp+J7x9DszQJ63h/2MbukbkV9NBKzdzPJTg+ArAZRgS9Ckmy9oJqmj3RL
TWKjuy/alqsQpJtvqavIRBYNBrRSGfCXkGk6NIMhrn+3ooFhC2RR2akjAarTW5QJ
2TC7ql8UztCGzYMTrZbs+LLqIC/NIXsb4hbvCw2E7A+MAKflQ/Ic63nZN8b7GJoL
R/ZEmWAWHk0R+sWVpIHI6rD2gNnSeFmvFvLh93T2tv6z9ab7DT6KdmNWKn4RFUhE
v5kZAiazV/0GTYnT4nMibHG2zbP6NUhwFRmRmCi6nr0qlhCMoxBvJEZsVUFKN53B
NhNc90K9e4Im6huPuh9B5xEKMeUlUz6LQNoMiI+CgtBc9TbBPP8pT9UQ7aOabO8y
sfK0X5rzVOx7Ghkj+SZjYabDwNni5tWimjJj/1ervhvwcZmNibH4aWxGd039HgU1
zBGx61cBfwExJq4VJ+/jQ53p9pCedoM7R7fIxIqzOCIpFy2JphJ742QsTvMhz1TW
hvnWJ9IK6EaTjzYb5J66lUzc7cmdZ2B98IH6ddpgPQL/gHr95e8LOrB3sp36fdI3
Y0IvY7r96kfoygT2He1/KDkHTp/3mWrxPdm2M77koM0vJFBJR2JR8VqlXPnI5cj+
`protect END_PROTECTED
