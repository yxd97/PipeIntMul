`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKvKc4sWknASnkG5vsX6hSyOjHNVJbICu/tTM4F9jd2gvHBvHxgpkKKQBPH0mUwT
bLMggviR8VtDPm39NRhM3WvIxT5lVJ1pWAnX9Cqtq/JMcNJDXqHk4i7sdfo6eYwQ
w2ae2VYI5r+EoDkHPn6+vw8+R2euJ7Z6bJS3ZRg5fFz2feOJZnxyGKL8XvMXSM2o
LRL8Sjs3utKrhfblPKhEOvsmWO+JwUSpQYXCElhQmZ7rKIEtDpC4W4ltsi8iruwH
v5/7vqsp4Gd1B1V0xJbLBv8T6zU2I9+zMY8kulND9jv3JTsPNkLkDmZdGHv1aEHw
7XZgZj89Cp1kEqWsfeypX+l7pR6m5meMpnT/Y6wZor90xhNr704i7344KzX7O0MB
OT/iMk5B95agHAqsgm2LOPRt26+yZjnoFb7ZlhX4g+PZBa2n8iHFoZOfDIsiQ47W
zYq+hGeAVx0/H5m+XOMH0FpFpR1EeaKKvQEWxME+zWknvwnMO8xOZ16+5PzFfdgA
PKA1J0NSyZ2Dfhe3yTjNO/2M26lD+rIZOrPKFMOAk0NmEu5wpBxrJqw53v6GZTzr
3gA25zfxERrvQeeEHOI2onFOvOHuClCUh3g2FjokDqK7+2dwBrWM+v0h37C+nT7V
99tqSFC2cJiDHw1MYehiy8/gWbstKfrfwxk/PwhftsE=
`protect END_PROTECTED
