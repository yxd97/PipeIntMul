`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yb5tFIkxZAjD050RB44CHUiqRu0aa+otc/BFfoLJBGRQoH9mtCTBWXMtwLk+BekN
Z3ETqTeQ3tD/I6SJUUmFdBPJiGlyn5z4hUm891Rfq5xQZUGho8EizgJoth0scVAv
JiMqSWcXyVHNmv+/dsA1iGdoMZlrReEfnviMPkUqdjR+HSZM70B/7HWOty299n8r
1XvSYwYpV4nMIJxHI0+3KNSapEFb6pEZrmQ5sUcQ0Xo4l9yt8dAiBvJUaLsmLJ49
jezoBB6opRBP/XBT9cnRGg==
`protect END_PROTECTED
