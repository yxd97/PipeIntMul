`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qu58OteJTr/lRS0IJJ+LqNDXpxm/uX8ajmKQy6art+x20/AoIF5GSoQiCEvXvUse
oJZUUdl6qwt4Jdt1Tb37JzTQEyS7JVAfZ3H8JZRdDDpyHnLsRUb5QukJo1VKhzso
GhOSDNUYbSai/NxrNwWqcJ8y2WL++9e94zheDrRVwlPJy+gR0FXZSp5SHBZMWtZL
7FbASspcR/zfSjpGLdQaTGFEfRDqYZVpDCgltycA4j1Hyrq6VLhILYD8rocMr3ON
+P4cWD3OqXf95TGCQRRGkJiX+YDRfd730K/Gw2vGqTEUJxqxjZf4OGsoKFsv+HWr
miq4yQJU1MGe3wA5/WjW4EcGSL659mim3Ts3SwR6fH5Y8iLG4Zr/YcxLbxsYDiKA
L0ZfJLkxxIJlnM1yVkq10w==
`protect END_PROTECTED
