`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzxptdDnc830PFUGAt73nYwLhb1GfyA0Az4zZ4YF6TlxoFnLWqR/UK/FwJTs+Y1+
WKh07fj2WuZ1yxViYBecEOfrGN2i5Y6Dkt1n7HZG2C8DflxT62Sb3QmeFGS6vPJT
92oBo1Z9pJuL0wFvXXB1P+TsOxUjTVy2F/senzGvAZK86bMT8eZMdi62n9AQB9MR
PTK9S7fsAIqbPI/eQlX5dLUCxMAIUNkcbRil+zHRk39QDIOkk2olaCGg4LhQynTl
7sMNRCZ4DsCEbmUdVH+hDE2sOir5+KFy3391c5ZNrT9sluE1WoHrsv44xU4gCUEk
d9Yhm7EZOjqSntq/kdpD5wtNRt8rzhJtsRCAmFoTPpWeC1mVRxe8oqcBDVJVOsbO
9WIkvcz9+2pGEewJuZQmCNepNPuIIWrlygnRCUQ1Gf3PpQWaXCQMX2IzmcBAQVHS
1fbLuCdhhHtzrd78EIki8iYN5X8dZ97QAvUMqb7URNEmS6ce5EebjYejzhaa+hv0
hxxINQ5C43rjxNER2BbIW+tBsgfG4I8abdraos62C8VBx1uT8+zE2e0CSg7mSDFB
vMSGHU+YJ/2BoTaWCgBGN9YYyRXTIprlJ6/Y/VJr1Ec3kRjZo8rJBpVpfyG9bUhw
Vc+n0Z26c0Cmj/gY2oBC3IHwUolCdDJNY/S7KxcrBtRVQBJJE1MlrEc2gRYN4qKL
SJ5sWXJZVU5xSl3SW5yyhQdYuZLFI/XAhsAc79PjuL02WKkAt/+0j44cWw/aZ3ro
SIwbSQamgUC/jHOut6PFll9T7FcaP09GYwYOe2TIyUDwS+K4SOvXrrMoJ0VunfGt
ylP+afsBkKPldGz1CrNgR0U2UuUeREQauAlhZAA69erGzfwIHaITc4aQGD/Q31kz
mtqMr8yR2kMs6L6MOa0Ebsa/e+17H98jQtoDzfuBLz9yZcmnK4fv/3tSZvqPub0K
MFol3+wslwcDlbzd+k3byV/jP8/RT8RtxMdhobAdsEiIfQpYrvLMg3MPDRPI6SI3
B06YLnQ2SXV43HjKYfbjfWPOMRK+raegxt30Tce3W8NkCHxf3C9c+0+J3BnvGtna
1WYov2b0/IbUdFj+WjnKVxkuXMJ1fe3QocYiMUPCMwg8LuDXfndo2ekhOynIoGiy
3XSJtftsHZ7T0eqjajqXd7ZPeuBzh94j5cMDvTqP8nNDPHwcRjChMIc3A9gNfQAn
N0PzD3OfmaE4J29Jk1cpD7OaFhp+Sq2VpbTghPBrou5Ib0Dyc6AvoDI0BRkE2aZC
4cy/zBSz6uya99Tvq4Vu5z0j8jjIJMgUk+cnqbsaiP5ZBUQpiJMpKfXByTpk1RlC
06JSG2JsrWJGLC5jQDqG3LksBukLQOH2Pk2qfoZShDkDftmkHAYoTp2DJeK5Qutn
GbgiKaaDtOWb/iJYI9TXHjGIhx5tL4vzWqBgUZUNw4LQl739B6pgxvrNUON4iAHA
a07xFrVJEWVw34FADP4rrEBbn7x0/o33Nhh+Sj7Iswpf0i5kKG39jSWco5k11NiR
Yval5VvEOiJJ+rs6KWqm2zKZYryCsUySCtmRC02Dn12gx6A/VVuNF0Pet3DCC8we
CF6fgDBh7mDWRLWHICkPZ2FlKo2v9oQfPFpcJCsOMdFb+HGkh/n4yb7JSc/nnIHJ
wj/538ymQe5g8dQl18GSEeBxhI9LsWoxROSPo+icPPrS1Ik98VT3iFchbHQyIP08
FgtxiCZculld0HLNM2fWS1k77CbLyZUrgGQSw4vN7MLuA/eS/KI5ScVltVU4lDB/
jj/NQHJDcT0tRKpfEKOGheY2xkBYbM3oCgFAAZ5VbT2FjS95K1K0RPGN5E9K6t/L
y8wVB0mPNz2ioVt9KTMSwCP1VeRNwh5aAV2KlBw9oiHgfac7GVZgUkgfFTgg5bD3
vE1lc9to0RDUOgGm66bpmeycTfUp7oiqLVDSl94P2hniIjuu1xULkxcWZvCSwZ56
R8dXZbJ9R1U2hsssDBRthZfTuuB43y+y08bx9rPmzingHlKAGeHW/0p2kcJSpV6g
o3M79h/4DDDZus2JUfJXWVmC3DJqibLf662pp6tvWnOzgpX0zBW8tLmazFbpgq66
WOUoMe7JRnYR5NjAjiA6p5RIIzc+oM+QEz7SzySv+dP2zJEMVspfjCfp0JrkKTzj
Ca61dM7CcqspPYSI1AzhxJhvT94T9DPWUvhB5rEYD3R/qYoumgHtPuFKmhfE6Iwc
EvaGUB4lyvXLl3urjDHulLfLQEk/H0is1IaGmSZmztTE9KjOr6rVxTucWhhRJd50
udr7v/JbwNPj/HPvwrmtHePY83XAKA6oTxLzKzNS626FiN/GI7HN+s8ESIAr69Kc
id1Fgx89YZ+TD2oOonJQfD7+yYJBcyKcFmP+cXVX5qvFIz/lEUl8H7L8AI/QySvU
4T7w50WKOX50QehD9niNl8b/btcqt2ouKIDlhJcn9seH6muhDvdqw3A2rHZxFYdr
UdWRtu5NngMW5R1PfFm93ZUYYTGlkbhCb+0HXXAwPp2+U9mU4z+Sms1HdMAx25tY
0pKy79ku06mlwl0fHVbG1FVVZd4S4bLGNCCqL+RGlMwRQQElIqiE5AoVG9ehZPFG
6EaqwlyyPgrUSGT4XecRBlMiJLC92fZPIRpulGq0DLYoGmqmNdSYf6lkEAFpU7+z
azHGgX0TIAgys3yjeyapsDohaJ3j+QzMJriFPmv/BE4N3bVHl+PGyMHfDYCxYlw4
fwAcHzPar26PzY/2wLiZeW4AO0xmAGigeF6hCE1l/DY+GWNugoLx9SMhxPgvondM
F8d/OlKwnuaAIwsGPPIC6eqnlCBBUnk17bok/imAwIO0Zyt9hjDyYl3nqIbFeeUU
5qTrdQ3mzE16PlW6NKIJ1JdqUkyhkwQRFRg9qXpVJI+EAW5by8a/1x9XHNPsLTFc
lfRt6mQWd9gxlipbE753JejkckfP5GoX76UAY/8//RmgOQCPgJ0zmQ0aTnDcyAy4
tpK/CnI/mUwCrWDrAMlBWpSL6oi1vs040jxIYwLLGlv3jjc3JF6PBZiDUNdvhhV8
YZVHqBx/CaTVepFBbv9pwEUFgOVsbSijbbk3k4Num5v4dyh5CgqTQmhgxse/vk4I
9T+J/5gtp0sQAfEAUnl91H3SETXVkNBuU8mmxZ13hLAaDgEDTBvG/kLNE0lZ4/Mv
GwRTOCplpaviM6q892rhc+tFTyrL4aVxG1iEe8oD/02TpjOr+OdbrAbJ6OapGcHM
xvkHT0J/yi+IgvaCJUV42UAWCkF6VagxizICAHWsRsZc9B+3KtSmEDGCAtsZjU+A
KrHsgb3YqLhn7uRMvPIqRXw1XHhioi3Kq9wA525Gaz/P/Wcg0U26JLA3tgZnGmDY
P9t2uyWT3y4lAGfINMVxu/y4bfR6OGgHkGaZjHH1VNpeq38JT4LPzJazrrTfNcNM
wKMbViKP+Ax++iZpvR9PUX44epCqQFYUK2g5lAOnO33L0hQYziazSQWXDrL2mYEa
hwoYlA5WVDDHb3DmNsjEQuMTdbt3z0GHx+njHoqMm97RBLmXQwNkJGgJzaj86+bF
tHpBM2sEvKeG1WMzUKYye7co+prMAyMSklmZVQi9PTAdmgXyKgpi/WDgVSFXunSK
ndvUbX1ySZ04vtFRQGSHxcCYPDnOKfTtADnLr7lbzp66goBzju6ywjOFKo2bnchf
5dmftcx2BS6pwmiKTv7l06d2Qj6XHtEpQSMEUEOJlBLfuCkmblPJ3659G/no5RJB
9MX93vuQeor1tGva4hP14yDNEjXaUqne9XO7qLOVVPbVct/lvT+ePN2HA4aVhrtZ
Vux7sZ0Cvmf5GqaiMoX7gzti4jlmeaH4tq/Tid6qybyNzyjZjKkP46Cz9NOHHoOb
3sQh8CF24GEgR4GVFmwcnuA75eFLIlFonXcEG7NwvGUfkqVWSZWLtgPV5zFDPY80
0I38EmxJYTW33Ky1UmEzrNff68GtjkeFjsn57Xrs+zSyccmImexMwSWAk/wJVhBQ
yeakMKcEeOnErvKVRS57VqQ2yiMqswmrHuM9DbhJ03IaIOi+5FOMuwJUJQ/OxeiA
lOZi3ooQ5I3OCHMkpEbwdMMoghqyOOV9FL8W0S0lySbfJOdE8Mms3gcaua3ZQygd
HH2OBHiXnAUnLiqQvbg7llbQzsEeUPrYV9KN65E0tLYeXjZBVO0S5Met96zNpLw/
s/qdM1WpOf+Uj3V9Ddcnw/w9x023jfzCkfjFYsd2aHCaOZq3icwvR0t2YZDBiSFl
Qlvy/PCNq0rXqPcwC7Ll7MKSx2up9OEt9Hd25S1la+a2upgAga4fHuLqMZdY5RLo
zqNX65NSnjgZk083Y94lfZwxvF6v/BMXmE979ur4ib3dixuoNZnax8p5LEPBR8x1
Yydhckbii/czjkgJ15HxycTwR1eBoKU6V+klB6UEG2D1u+To8u7Z3j8CdTUBMzKB
pa3i0CbU/oUOYjxIiZup7zAesKf6YQ+79yMGmwh/j5Z0PXx7RSnsqoK03/X9qq7w
n+YRqZpBC0FDN5qtCNJMHpHLo9jBb03N5nbkfPR0RmCRgMf1b3OfvZh6F/5VK7eT
5Uc7nrvdjMEYhVFuG06xb/e7TI8E+ZU8qkDsO6lwAMKYh67VKObhdpoaewl209ih
`protect END_PROTECTED
