`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQvEYU/gO4joqvBxlugRI0ObvLXBHiQOTt3GBbqNg6BXOx5muGlmtbz2SUTwjK7z
6LvQb3rj6pvTqg8XCauEXBsdOplTA59E3sxA+gsaqk48oxjsMMwz+gNpeVBiNem7
k8ep4AAt0azViWP8kHbLOJKFm7V0IQBdS/iQXwG/fn3cEmgTDvjDKC8e9lMy8OzM
T6M7fSMDoXWRJztRayKgUSw6Cw+v/un98uqOFBxVUhHiUICr8l2RL00IO6tt0g4H
WaOZd2oDhcoGy3Uyx8atlElHEUl9hJoa7QdR6zTdWYeTadie6kg85ATome3RP1yz
e3+PXmU5px/MBEI9ICB0ljioR7MGMV5nBd6UFJapjeDxpFUc+pHeggzaxJelYhiY
SEZ1jm0aaNVcb0uP4pdtBh1yc211b137NDhEx1AFxJfF+zjlqnTL5Qv/KAJdOtSz
HHmpOBVABkrARsbr7VY3Q+P9JFQzP4mAYh2291wOLVw=
`protect END_PROTECTED
