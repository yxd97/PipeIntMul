`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T7kzCXYhnS7MBY8lk5uKNNEGs01ktugptdLufvLQpGKf2P0HHKGl+POikXUr+tB9
teiZ+R3Un7sNrdfOzmOWFs3euHyPeidIZ3yZ8SdOOoEax7Oo+jDrlT1DwB+Ws2es
/QcxFatgPaan96Op7Q4sC5Ta/bmLrQoQppC+2vWYgxvssO9Ynkk7kSr+mBeBndZJ
M9rWyxrq1o7ehCFg+lFQMEm3iAPtzJdZ5FE9EbB7Jku/avFVrMX1CXvSuS39BKTe
U7ZDFOk2ltjsfHHWapk5DcyF669nsgVYd3pB7ySzgueBZY/3vZXnT+ZZoRpb0GBe
st37aUcWHiaYqthmrTU1Vg==
`protect END_PROTECTED
