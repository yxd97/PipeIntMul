`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1aCklAZzH4qc2kjUk3jD9Ahr676eXH0oQfV3p0aK9bhMQ3iZ1/XaihRKmw9iRmp
QYe5w7XsjaG/cJljoB0Ne7DyKGjuPAO+xoY5u1hd4A426AYJFhQu4tsmhOecHYWl
cyqxwSWQXKwMKCRtr8BBoPtLBYK9A9qC3YYIQAqKHYPW7d1Uibi3GsmLK7A1JRfL
hOp4OIX10BGo1Cd0LmPYmO3tv3BbRzK8ihCkbudNKsAXUMkPHd/EPgsO15hDFR5r
Qb4xsqyMq/YZHOPjGAq6DA==
`protect END_PROTECTED
