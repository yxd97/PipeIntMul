`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jDJp5uIbdllWiRFzs0Q0L6UElOlGQq2Id7Jxtenf+wS7GgyLRfewn6cxGVVcujSn
vCRaOYQgxD+IsdYswEAIE+c9movP2tkpaBlchxaWiejTh+Tnvtf/MMWsxlRLfiEJ
Nsgn9D3GhDNgJtGd7WBNEEOhBPoPzIS84zzrRlC6iI6jjNUZf0NigDb+yo1o3Ggw
qKxzGmv0qkvfL/jIoYPv3c4udCYdY598yQYotsLN8qG1nxOyNMvpl3Q/2yKz/i4z
3GEvVqc+Yvyn3oi8WpAeS45iSKrnKuAgrkV487HFp+vBXn1BkXI9bEQ61g7tKsdj
5GFz9Za4VsWGeGjL6lqrnmagF582E5uiOyDirEWCcg3+e0m2BC3NIcRNF+ovJbCc
7w8GwiNMvuWzouQKTx/UmUwkVwGIex55bsCROvbKfAVQEZuybvBIg2POlErOLDmh
QUk+wiIwccFmwhrofexbThtPYvrb/xnDpVBzGM9yhp7X9wrvib68UUDp55xxC0ob
DpSPwvKbhwm5mXxkf06VgQ==
`protect END_PROTECTED
