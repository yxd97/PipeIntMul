`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIxkZoE8DIrcnZfxiicHaINidCGwm/2Nzf5+KCy3eaFzPgTaNE8dyMbs3mxlANoR
c8U0x2tjwmz+HpCJYWayaw0UVEMP3jjhqXRFjADQ/GytokUVYGjII6OfY7IU1waa
FHuFwTRi2FuSapzG5idp48JMhoWJOMUJdors9XSJi5wG4+iuu7w7I2xaECQ8wMcC
RRib//cM7jucSWgkL9eUZxTKo8AHNPPEglIrCGTeKBPZTjRxCafrGzabBLL+2dn3
zUsuH6J8NXB2Z5eb+nP9KS2a1vmV+bVqON1cw5rFXJNf+3b2sKh8DnhonhwloPZH
hjqiMLpWs5at9hxDVkGQLjeyTQleI0qIFg32DmiQj/Qwyoi8ir9Ve6ExiJ91/39c
nHujheeP0Mjm5Bc8lMFysZFQscdMZbJjOvFI00Hx/5nMilEijDFwgvDB1drAaHEn
YLsFdUceOdWUYA/TIfuyETvwBE9ohLpZ9C1nMMPU/qgzywhKwtAUZ9CDZlYL2sH9
xWnnRQ+K9ur2K8oMwjRxcV45D+ssQtFvxzYPGb+C4WZNKNqyf1EqWWmV0tptrkzQ
SOawPvKkqplRwKTGIBGLtulb2tYV5tJf20G2i+cJPmW/H7Fk822k2PGiSHfEwCVQ
CfwzMNhYx/RuUpWlMpzTiGKkTFmfwYRrJQhof69LitgyYBoF1HySCSqMmhUwn9kn
`protect END_PROTECTED
