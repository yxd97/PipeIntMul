`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mX5BAb06uUFA0i7zuofSmkpnr4bGRP32hiSOZXmdRnEMc7j3t74uYsn+cC5BNpw5
55o4LKlHRQV1pMWs++LP6bvzil1sId6hczss5z7U3Swdx/GPDSeKPyuAvJJ5r52i
36IE1sL530xUT5iLnUivWhP8RBFHGR7wmORmIVyCNi+4JxMRY1b7qYT7Pp+TNLAc
PIm+7XwAjKTFvWmLOu498Qy1ilD/Gq1mx82pT7frJ7sOklk2Ye4xJpzxzJD9P3k0
mp9nBY6S+cv0x+8H8oITzUnsodm/ltXBcq6cDqio/jT/qmXDFsA33VUI8CGMGr3S
z3t7/CZc93FJtyhI8502R0OvYt/vyPTWRdX0mTVSdLwzuT2AVp0MFaT+8HQTWbv4
1+Rcd6pcB+jLeBN0uYFMwMRqqb3J9BhNguAs3fmxKv6dhMKWrJJtLuUQY7oxSZGg
`protect END_PROTECTED
