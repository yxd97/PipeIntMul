`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ytx3Ol+A+5aTw9ARN6EBNIhbEYBiMcyepRwFf7DX7g9GmeG9JhCjHxhXauPfGyvF
QlCJsddWx3J/b2KiiRyg9Nf8nN8ubbQSlKcDi0VWZz5smymEQoVOKQW9BogKSwwk
J8D61QyzYNlSb6NAN2jQf+4ZEmnUjPqycvQ+WLrIFQoTnybtAd0tAo0DzDZUpjve
YYZVGxPlUzH31EBpHQdqHGyGa+W4stt7HnJ5JOVVtey1a04Yhdyfl4r2MwdoQQR4
jEWAJgr9SCM4Mdut7d1x3HOQhCrT8qjq1Kuy3RJB6ivC0Xrun1gsH4k/Klm2sKV3
2PYph+z7Qkzedjb8X1OAQAbzeqHu12hTKhM3/mSmkQdfsUayoMmfNXM6bIreN5yO
Y/xpJYvu6A61C7EeGTWcz7yn5a3uM3Mxmnkxzw0vKdy27Ype0KPF+8AtP3DK7mNO
8kskd8tHuqwJ47/DNJFLyf118KmHlFK2q7xdCGYvIzjJiM168WATws2v+WA0lirj
yhIbgp9O7MGkSv50lMiuIRInxubgQnQ0+LASMBDq6gE=
`protect END_PROTECTED
