`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VcNvmkzXf+UwyK/sNtTuExCG1Dj7LFAIOv3oXYoLQZGJJEQb997sU7Q3TNQffDwX
3Xq7b/JgdqKPEx5gZDMjDMcaf/sFgrAOVPyCvKqkNhJKi3e/HFXADtbMco8q9eV/
4/CHu9ntpVqy2OWxXakMzAht9R1U+ZYk1BS4jtd0wHAIm+6STvHYcHrzvZeGCzuA
D5SQEbMUr1QsSsR7HLBFYuBhfXSXfL8dMhxKILlFFTr9Ym3xl4fS7hQlPPrCv4LG
Qqgshbil4kaCJuW9fIazGXhH1/hJC2QjohI0P8sqQQH6vR0E5wqMDOsk7F13uojm
f8xIs7ZUMstzn4xmZtqs63ajOyrB8h2Z7qJzirMJQN8qiSXjjsA561i9xj0GzyEF
hbIlQso5QHr8Pjrzt/zm/h/dBB+P+uNxS4bWk1qbj8+0pZtgGgZPHdfji96abH83
6tPraDqEDvU/HogGZnjnGobPF2f/Qj5qDnnj/x3rvRZ0pFfqihqLKw+lhvw2FBoM
sDHDdZ26kCzKlJ04bktWRKh5IW8Q8hCCS2x+y4XzFtCf9+er0XMj3g3hfMI9kN9Z
58qP7FSv3VZ3uv0gIaMH3ktJsRi9AAuUw2XyGr+F1homfFcwYAPuJORH8bMU0LYy
vwYjjba7lCP6moCkA87ShTJnbB/gAjVEAEq4zr4Ty2i8cmAVXMXMVpJdcXZ/MDm9
XPm7GtcHHqZtiW164wJ4qGOerbwWVHqXrVWxvq88TYJQf1iekGHeoTDznTXKV5om
pUqIki6effHYHMCjKML2HoX01zgPPKKSIh5n2AcY6qe599WV8nnD6PGwLmffoFAG
1cLTqrAAuDlRW0SVSqW/s5yaPA8oflfv/bhTXSUtVaeWX1P2qVGwnSw1HrYUQxCk
2jePPVkhMsAh2YX2NP7vuhIgxR8OnG2bTTDsP6Bzuv0o5o8NgMfnfDBp8WIBO33S
V2oExHrT5NhD1gs2Sbx8A0Wlt3n6+SeU6DOKOEsv7qlaWFeUO95iLedrkKHTVJNM
2ce0e90PL09NUzCXcaqNebOAjg+Q3XB0QYPjivc+mOTc37oXDPjKGjY7OztU28Vk
+p1nWoV8B7CiD9Zak+Rle6k1pA1bG/69lPna9HKz200XAPRtqloErY9SG6dS8RcK
Zol/G9LwtTxsjw228xFFsufys+glsEFqk0b1gRPebXi03p8NFbw1OE/nAmdjkwwe
pLltduQCGSjh/MG1xK6RU9vU3sAZY4G6I1aWpWXPDHjn1CcXNc6G+WMzzympMn7j
sguQOALA21U+QTlbpeBagVHdx3NFaNbQA+ZlD0zRGFNoBYUQEh42WPv3rdCjFe6j
ffjU/AoLwr1RhT1Yvkn2bpNwaAGioy5LSusdkZ1CcFunN7QDVTtIOVyWlH5Biwcc
A5QC/V3RoH2xyjs78bfe1oi30FHG6ekhFI7SxOP8y9VKcUZypt5C4IF3YPXAwIho
0z6DvFugxwXxrzjRd3I6L/w/ymSy+tHBaTIixtm/pKlRFoh+nXFigdmcwDggRWYZ
mhF0DS9ojT/WiNGSshl3c/HrXDSG3camKnzmTcOK5H70GAGwe2rPl/MXDYA8491N
hwn36XWdWafthsu97Bu7+3GubbIgmzA2OvbbDh0Ob3CPr/lGzY3b35jn82J5mXkU
8nlcwy5WnKFXiF7hON1qCRfDtipcQSU64vNXWbEwCesTNHV59sL0XonTt7zOSxhJ
P1j+lUTqfZjJAadhYynNnt/POxP7cjPFPhtT9Yxwgb9SHCquHlNFp190Kl4kN6zB
ByUf5ZLzFnpGdAjCli+NEJbHUzwsIrteHkE2DsnV7887aWfKh2k5RtbK2/eNn16e
qBG2yo92NE+t6aDvr1auVF+mWOY/CnJ/89pzzxoZzFKJMni9LrV8E/oJPma2dg2L
MbDY2zRp6BqU6L9bUaFlS0/3jDjbkonCmxro/Oht0BaxLRquuww0DaNN2hxmI1f4
`protect END_PROTECTED
