`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5mScTGbtkOd2U16PMKWsqVb3e71DTEomBXMee14pTnHz8MFTsl4CEfgUv2HH+CU
Zwp4yDINPdQ5CDQromVpWWyQR4O6OO5K6foX62nL2ozokF+Az/bPIHgnVPbImt1x
emI+MOraGw0L7W4s3oCvYAMrvYVMgZ9TDlpYPLZIeBZ/+8sV1BdBoIVFoZKPBhsm
GOn7NWeV+9uzVU35WyvC2gk3Yp0m5XuFTafCopgKTG6M35BjPNP/MiZXmD4fddnp
l8NlczvblLcbpfoLaurBglHkDriIbO5611mBhdcRTAplGyQMon7CIsJoZ/LKUqO6
LWS75QF5LLujsSRbbk+AGwdG4dmOPNuqvOm2LJNsEN6JUKR/vdCaeNLxq0ChaTeo
r5du9TkUsPdxFqYuzkEPy6EOecU8//KSFuYcV1vFR3RQb6WSA74g5zpZd9k/xYLC
msunSad/pEbgpjLlZaCZQ8+rUC2dfO1jLSsQMnD6hy/mLSXk0EJim+rtWvO1f9Ej
121NBZT6R/kIqadQLvILjjF8zARKxSlAajsy6oBAlsWyb9wbNW1TAlJAL5aMxOau
0Vv+1Lj+3xlrtCmlOD5bAWtKkwJ1x6OQeRBTPFSWK2TStapCW21enRyVQ3xIkluw
B486Bj0IzYArvxlUGrn7SUVuaJb1pTtl2LN9qM39drKdPCIsXhcMKTfoPx0ncVXd
M6ZHIh6BuF0mpfHwJtwN2cwjZIph0iFgp8GHl+UV1IC0PFtyWk4UZ6vb81WINroD
EZa2j7hb7wSvXUfKdIdbUGrabrci7iAMgi11uYxbHoTzmzQ/vt98aLScsmWu7qO4
1ckv9F9sy7TbTpYw1iVx4qh33LL85sMlicPg32uW9q6AOv3wTzHC6pZHLhSz1OyO
R+aVnxQX4u5l6Z3XGcWBhzGBnelMlaKEOjwZPsaZmPC+LgeaihR5OMKsu/6OYQSG
3CALQRwhUt9P5nZmuw/kkDexGmQgH1pf145bCOiHZO0=
`protect END_PROTECTED
