`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ECLfL/9iGzGzsxQwR3fo6nLi9aogsFaIsrkHejyIg6q3ilEZAhJ483tjBQLkHqxV
GJc/l72DAMLtk4kAJ4l05JSvlVVWWmVR6gUX2rldkLShfuAIPi3tGJ4XyWx9Ekbk
dQ7EoFDLaZMo+m6HGlsWWBP9HjjvgrggDPetKWPfndIHNr4k5oZ2oR89ldhrHf35
zO5pGPEnRDwq8PgHepGwN94frUEyQh3+PSym7htEb5RtjRWFKVL2lqCKA/+iEIpI
EbfFz37eGFA72K3kR3Hpu0hmpPPSHdOJjfj6zT7DdjtRYn6oxGyM+OBaKDOkhb3b
eh50rJotCCw3oYeMB3+YNVLccaZy2LynOx7hYJXr8E5C+elWfk/wt01Y9WX/ci2E
ZjvvEDcvWxUdS/0sxX14+P/pBSMjGU2MLul3I2UfZjH4kx0hdZ6OspfZROLmn6IY
P//v9OfEdM/EFmNrjStkT0f4kvER8Spep2ukcn+QFKUNc6yYTzG8i47okd9p7PI9
i5ksetCCWkCGXFYhQYUtQ0iJgv/Ly+cvqbcDW4Dg2ThHoTl8fygeylCSREVvFw1a
uJo8GUZ0K+aIMW0XzbMfw0STjAeTiFjSzhMTb/lvDY8Km/6EYemmUmudiGAo8L8v
Aw83cWfDPsiKsaV1fkKxuBCynIEBVHarlTFdVRWOwTb5LEVstLXnXr9Bba/JdEvI
VQqVOcw3XKTbu6qjdH95QtcbguMXnTPhTPF1hvLbVIFkT9Seq5ECjvUyRCSDxjGC
TierFvJl6doV4TQeLxWb4H3LVnyUWUBZ7kJqgk5v9Px6yaxkUP9hoPblVAj7cnY9
GaK0CFntfk3aA7KIoO7huwgJPYJ6Enb78cQG2pXXdjjDPm2DGOu69c09Xvt0L0NP
g1hUk01+XP+Z7hcIMYY0d8eqJ8TcVHSrOSk3vDEIR03bL49nbCHdrC999r72H0NU
dQQJFZl+TRZoAtpHvRZCvkw1oOA96vbY/4pT1yrwgLPMzsf6okDhamp0B0PMVjfR
LVY65XkdxLMFMoXLp5fTFWpE75oherlodWkEV6ctRj4rov33YuQpFpOa3sB/1Dt8
Y3l4d065YNBLpEW/sKpGnJtfd2Jzp6+uNSMOyXb5r3v9tW86q+dNw4ISNly0Lrjh
GfhZVerUePBAy+xGZoWkLeStdrMYrWjMY1WKFphEZtMQagcC9J7UT+svT2t3XOWG
Fi4Guz3U1VgWdx/tEcrQ2gOmjNXNbSNJlb3fzwECkeVGvGFTlPX3BnqJjctMnEnB
CsMHcDk3+oBH0K8bsNJq2BJQkeyPbdUBEC5TNG7rQdtSBj8oBSkBz8UHMWfMlXtH
/4rrTq6DMapceZDNS6slBn5TpgP90JlWrrmGUgnFOtHlTSjj2imEnKcZ2CAJMYOH
qug/2toZjbgP2468sMmn4nf/jE1u81+H574YsJt+xA97Zlnnjqh38AmE6Ytho6ZZ
`protect END_PROTECTED
