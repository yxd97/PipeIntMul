`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBsN3HURzvv34K2nQNqeRft//NTAEosmbi52IvMwK5mYT8tbcOOvrbMqW2RmOgx0
Z0S6PLO0AIt6pg/KyH9nRy2DjI+QQmHWq0suxXslivRaZeGQVuK3qtUxpEe6WYYd
Z7ZqQngZ08EXmRP5TNU2y42wm28mv4FZNEEmeyMfCMCgoVMoyIc0YmBwPYVhai4U
nrmsjqWa13wTiOyRfK0SV0QRg3AgrPndL9dgOmUENBJ6fVYDRhCl2bom6B/1QInE
hhJP6JaVrOp78nIjSGB9GGarwxXQHl6T6nAduTJb3ZRmnktWSTBcY31W+BGJ9uYs
xa5pA4NEN+FoYREaZN8XNQhvi5fmuZQVICIZQKtIGriwOEAYpzA51f+4IopmQ2oi
9JReEFh9PhYamjhQnfI2CRpDCd098KwvtpSj1ttIHCiFIqJZqFdbkBUKGg5kyyqs
gkm7OkJHs26QpleaiHTS5FwDVFB4sRThE09EICkBYmrPGYxBpDGUkRDxOAluT6Ee
hZLHflRYFnwmYz7OKi4Gu0vBhM5P1qAQyDznqYXRvVrfZFWi/rxzQ5F+yRFjXaJ5
u9bUdAeqHQlHWP3J8yon1FVN0ZUC1arNKutY6cBSx23ze7Owb2JXM4G1mHZvlsIz
Oe0XaiEpDjJVUCIJCmEET/I0L8P8X/PAnivgFKU4+ct1a7USg/QCQJtVfnwBwJCB
ChiV23YBpcyE0VNAwj2pf728MkcriPCGEOXwUwb9QIX0+sfv2BT2CIzE0pxEImwH
3CRR2sQsUsh/4KTOQFFiAeazi4kLbf/hwD5Eg1Q6K2Eg74EKVrd3KkZ1CV7QRqD5
mXYSAv/qj90io+lCEiCVKwDRvav84o6dnHMEgEn+p0vYaeuoRg8yUfQSTM0Ux8hQ
DN12INo9ACfBml8gK96BkvxaLv7xeQG0/Vse5kszEiKYu2uqtoxJKdDK10jfw9pE
/F5X82pGVAN74hSV2JlUl76d8sqcty/nHevvuisuxZzFePL1B8wZgm3qw4TQjDOt
2vR31mN7ODPy12nV/Zs4UnHomtB5drLiBx/e/M6pckZA7f1lXiAsUmTzUxvTFbfe
8ZVVMS7SqkDyP184ExkvClk5CwFw/r2GQv7W3VhQ3JIHnLsAE4gycREUqTbhS4Qi
5+Gs7LqOZwzuHMF46H6EecXJMinj5qqv14mMn8IrL6SaPDWwH2I7iB42I2tW305Z
Ea39uokzTgGvEZQl0FsmPeWmPlP2Xia7ncDu93XnCkfcgsbqSHtdqEZ1MvenMYKq
IBAYbYQbmkgnXOqWuY+3EQtOjExjt3VSoErm9QL81otstzpKWQ4x4+tf9zpbE5uB
MalMaWQ4U0uwHf6WmR5Senof0bZ+7KZMqVUGLjXiV22oq3sRw2VujrATPKo9RotV
YkWH50iCzk3whohtCp/AZogOlCoqFWFkdEkVB1kuLXqJg8yHADKIifPUSgFJql7C
gwM7hBmYpsV75km05WWg9vqREHZPMNbN/Cij3aQ63f9iQ+RngUGFfqbs1Wgcsl0R
ECHilfhul15WckT56euk/lpa2+QkfIhqW/LwYY+f8cqfXfJ+D8depuQAukmolaxF
a+/imOx591iSckrQtyj0zpDBL97GB1DBPp+G6yABSy8iVAlIc9a6EsHnjGSAnws2
UUuLQU/dZD9ucktBdg5G2K46QyBHqUW99QIaaExNts5LDUs8PlUrnylu7NBB2J9Y
i/e9yctWHASDVEYcMGO7N/AAZLR8tAQ6N4zW8wdV9tlCjmM4iAbOFtwoLJ9nSv6r
TNavgmz3jv4nbiPFkinDs7d6UCDBEOUARTZcGyjyrovLTSyxjw/xi7KkB9AXPbcI
QZ0v5fc3xlpRFhuwKhh2VQfW7H37a3w0nnDw8FBLDptfPnJq99oCH4gcnGo+Kz6z
22EqxYVtj1DSG9Hm71YtTjcA6YQAZvX/piq45Xg1DTR55g3BdzbfZRxDQ6XKQbp8
pYgFXDq2lZfwj36Wx5PXE6GdOojzbB1wOLZgoHviWJa5z6GvbBVDXR4GCLazG/vi
2oVPuSTr9gUexc1jICHm3oS4a9ZLWU5OTEMrp/plN+XFkX5iNrP8y60+5tOue4Bp
cQ+hqTO8epOP8racz3xZJ5eXWCLhPKN6pY6CR3XmaLUXIv4CFQSvUowqoDjUjfG6
rihjOtLNqq/LwaeJQkHaZO9SNMPsQc0Yre0XZvNE/TCRjwMdNRilZVav4OT7ArVZ
NOsZMinz9kkrpi74h8gR32rJFVYNUlW60pyhAOPaJ8XscRGT8immbp6rY/dZTPb8
phuLYZrTsj1Cmzm6qZIb1pGR+Z7XnU4UOOZfM9cKPTmmjy9x7hHZwLNuyqT34Aqo
Ric73Yrhu9ObVOit5oyy+ekqyuaag8IQTonIkJ+kHC1Fu6SDAk7vIvJ1N57YC3aU
1bbred47vmexHL94KHLeXthGrSG/onBo2XXMAz9zYfz+rpXEwEPI6Mse1KxuCPwm
HIAvcpje+qPhvJ5CDfeUXrUO+97FTgr5kQbGzUaiVpXdCXW4ZyaYjq0ULh6Tyuor
z0aJhmZk8p8cXJEYsvsoinq4M+Up6JIdBRLH7nwDG7t5eoj7dEjKiJ0PGxL6Pk1e
rHdQVVz8Vrzk2unf4oaIEFU8rAz6GUg88RuX5hFHXB8Gm7y1aTAFI93R1GeFlzBo
W2M+dby/iInTv2mc83QKtga+47mjIx5Bm9v93HzxmCqPYl6Qkf5Z2TQuepGPqmUj
RGzp0Ot+ZdynNhM7YUeCF8NuVSTYotX68s+WN3gflmv9P0wAFfXDZyGLq/Vuv7NU
R35fqzi6xebMHuO13h/+YqffrwRsCbKiIn4LxfGgY7rQoU9vSfLm3SHv/wlwZF3Z
wTh8LNETsBnN8D21Ykcrin3/aCLqO2SOEBVdnUUsCXTxeBajGzSPycxZgYZFRtNs
9GLnMjbKVwE3ADfpW7oWAMIWiGIEdYqnkaJMKL7TLZTMuhMmFFFHI5oPVV/TlPbf
NnkBJMqOZTkg9UxOgdCqSMyMVuMF2pDO6xpQJCJ6Yy+pft0EE0omnYScQoNPZl1P
VRJ6INOO+/uXM+00ki7RwZodTc1pijg9cWtW6HxY7UOMDz0CC427/XNKzfCdW7LM
wUaje06BbnNizlTimYZopgjmPWHWM8ZdjKx8NyfGnY7tCZDnKFBpoNS0KR9YcM7t
7RiDfWnK5eTkQ4G4iru28LkVFQJZ3zfwU0ryYRJE5VGHtQbSXPFF2P6r7PY6rm39
sQ6c8XAguqyhdAprd5mjrhoO5ofnaUERhaq6vCb9DtX2TdqKoY2J7b8K8t2J9JMx
uupWfyT0kTPgUHFJj45igStyhJI5A01XbFeGtF+XP8iHTOkzU4d4ePlMnfyoxgM7
/sbtxvL0ZC0L9je/3IW5re9SeLthJKr+K12i9kjVSEkRBTwe0EcXaRJvBqVPRBGq
7xUy24dpf5DQWf1DG+QITpu2NFSTAB+AIeSgOvj+xkRNYuvTw6WcgTRHgPaNyDbs
W8skuoUukeiHeb+NpABeYyle4uZgAwhwizlk0HLnWOslpKqxJ7fXl5C1BwKxkLDx
8DsMI95G/MIx5JXWjg97sBmSdKn4S5jqFsdNTQX8G5nIGqPGVIXxwhpdr6aqceHo
S+bXnNl6wnHp0E3KOSNdvuVZkdaxD6SwIHlJ2yxBbAtMEW/Ms9MxQ6xLlN4d1ife
OqtX5/8dhfWEI2jE6K0bTBg0AsiixDHzyHYw8QLi1iS2tnPDUmlAYROEv/EAVIPu
J6N9VheqdgRuC+Utz5oRi43LDzcnfxWbyUc9JNrzmVnmfs/gypulJ7S4ais0n5C6
NCgyN2tO1HjxHoKK3kG69DvTiicHs81to7CbqJ/Ysqya9hGjB8fbeuRnfdxd5YIl
mh74aiqW+D0mD7tb6mUW6nt/HmztrtVY9SChxsZ8evFG5/JQ0/uWMadXQJpY+l5k
rRe9k03uc1HHhtZXds5TAxILnVE/b3AzPRoNtIGoqdTnyHfdD0smAwNM31BNh/K1
//JDUuuZI81m4+EBZq5ahXABWSDbDw+3/Gci3QZC/iMB+PKMKSeelheO6k4qn1Dw
+bX0uKGXU+B1f87vBuH/7j9jp6+ue8B0DJGiw4p33pEtWO1GhXeKxhaAfEQJAp79
wKw3tJjv65I4WC2Grey5hzQ/JuH1DBT3/UkuHyfWuhzWoQYg5soSgpiAX0cqGNbN
4N7Xv+61w7IuXWqA4eftl+caCL/dyK6igYF0VD5x5W2yOqvP1fckJ4AI7YIdkcPo
a2TSBRwQ31E9gYQ5v1SogWUHanozgng170E5hM3rHOSZI7XQxv+mnZWTDb4kmUCp
ZbdpAsSpJtCF0yKGnrE87uc10oXfm10AsrIwnNdi8qMZjHbhsq1rPdeNAd7WRIqN
IHRrQ7YHW+U5BHNQGkdnMU1XI3ddPA8NRmjx8Ns72kvgR2li5RL5JEMdAz342hmr
ZavsNO+rECWYtY/G4nFH8/fT0EiGTmVM/zIb5TvtUfWh3G7wNRprt+dYcKsXAevr
Whs1knYq0kaXVfvJLiMvx1pteyIpUMUeiZ5dVa1zzWXFDPiIFwAPAAUNGrDpUEkp
0Hewd7aoT23wHsxUWcaCp0fk272PGt3y7HBbds8JZOs/P7VJ3XIMjyyGGdtt7V1K
UWVF3ROkBK3R53hM5bCGuVYZNa2msuXvp27nDMQoyi8Ahf16l5Lb0C+nWS3u+0tq
8fLYQD/3TzjwOAdqqE3RRO1ftyqsl3debtdpB2C48coE6UjQu2wZYFy3E2M7lThU
v66g8u4Yvj5JsXdL3Q5cYLUql/HlwMvT3C8fHUzp0xra89ODTiLKqcCdvut9k0JV
nntqR7+DcXL0GcQrL3yxaQGpUj6wDCBPKMLkLfapnk20VwFNW0MUZL5wbw7ed1/l
cElZ9DDO+LKOSyk8Y7filnM/t40RQkQ25+xZrKlfWEBLCxhR/hVzOshsfb3lAb+h
wnl4CPcIwLsepwOiG++nDkL4QDIkmFrxhkTW9GxUUPjXFn77ScyrtsF71yYCxFuy
5u4x6OIsltsqWde/FE26JrBSORILrBXrtQ7+/Jpy4KtohQ9YNFxs5amxYKQKIvum
4f3IEESqscvsTdMIemGslOF/IGE6KfwKoYLsgQ0n6Dmmw+6kdWx5uyh4uqN8k4X5
5ep0Wu6ZHfgIwRc2pmG6evlPIX3STxNgluf3UuiwpE2a9upM0eTbJMNWVwTjQpKO
UeHwLf1vIdosovJG4d7GQy/kIDdhVcJCz5a18attZMEd/xbj4bDF2aOj0p8tHFna
f1E55Enzh7fN8UKCeFSOtO+Bx1XCQib7XwaMqtfJz1fvN9GgLyZsnYkSWcd+MQb6
crD6ugtslPTXIWXJ2gQuls9dR5bP8m9YK4EOuyQ6G5w5dLueVcaavsldsKtU8PMT
jPNk4+8wueoTwW3xT+475S+Gt9Vi6CJqKFMUg4WKfBrp4WGvE37JD3e5sjk1BhQN
KxQvD1fCmZRQNRcQUpGOgZnW/Kw3HB244mJPlyBnJz5Q3qBmthMUhbsgWASz1fQZ
fSfdnNKYeLD8DJJ3hNzdbyduBsCdLsmu3KSMxx1NtNgTvyfABs5nWvjvZuziyL5f
x9wDLoxY1JhletFU4VkdcF0xDk8Z3CnOwc4k1g7DoXGmxk1fDnlSOmG1ysWNksCU
0p3jGZ7dL9d7jbfDhDckkjNTQD8gvXygY3/u6J6TqmkCO0ZnP1FgrvDgmv8Kypqn
XF/a6YykFhfhDHDR3agY4l1aleORdN90YT/hypG6ADAF9Z4Cev2DeShKhJuUqXwr
Kg/jn0E8LSa5KMKx/kDsyTsCNyLn0xKPN3OyZXxELlKWGsAEt+w65Kcye5Hhk+rj
WWQut8T6NvfMToSG8gs2v6ne9nWG5+eJhzAern5cxbGRQ/JsxCoIjfywhQ71ia94
qZqu2NQFRhXrOds48cDGIsASeInQrpsw6P9Hsn1HVAvpzaNreKC6NeHewO4ox7zZ
w61J/6MKu/d+qCl8jK4nUOg1vBCcQZyKHfcbIQE3p8qpOmt7iyd1tl8KFdyNLh54
ohb37FNYc5Cx3hoRXvVjqZHM06sd2nf3mHOvehLbltgTrwTRMmQ1KuKJrf3qiQv5
2ZiP8sVo6dRIEinBiu2J1IefkjFb31WUk0fWYKtjncvpA6oRctCSquRhkLe6S5bg
8uBGDF8omKT1+boDZNO0Hd3C1AKAR2T9VKDmfhHGpzM5PVkNOH8xqXoinizWCW91
ZSdf4adgPqkivmBlL3ovRRoYcj863XZlwuLf2REkbyzgVqLvTXRbeT7Y54xDIgEz
z/hDfFO5/UTxNoLYLE3S4T39usBXaN1AqLVYPjZO1gdmd5/l1BJEilqa93EBH1Pl
9YrAxMQpby7yN1kJKR/EIQaeZZ6I3Kt1QPhv+TVtWTtMDyzc7zIt5lrBGUzrOnkK
KAYMCIPLG942os50bd4ZlOfSsin0mUOy5WfFPYItyRw9RkLsacmvyUpHyDH8/V1k
nxR6015FwB2OAJh2gqODbB72IEo9nl8RT/gctLP295EcAnaqFBa2bBTJ6++NAQwR
8pJUDCg4RmhTkumFFXq4cL05KOKpgSriRK3wBdnlJZc6rdxskdUwdFbOH5zB2n6W
j7N+ALGiv3ykNwFh4ks7q7Lk/DAidmJ0CtCYc/ohl7blAfc+IpNXXXRdC65jw13L
wIJoGWYrs3wf1PYSbvjV+umG7W2igwTsBsoCr4JgjMXm3gnpWnN4oHw1CnKjjjZp
+nxLhIAeCOBc9sXEkM61nIXdIOFRsHmGZKFjBURshoIxrnvr6ygF8zoICHU7XBKP
d+uXQ0O0HYFO31+obEOlV6Vyovt0wGBNO/equ8q7XR5QfFciIKEtIdL4xOpSkPTh
PBmYGXoD0K9f6R2JUefVl4gymvOb//OWhEUZHFQT6+ZjF09UaTwZYiuKg8n466wA
HOHZw0ttvNB30552J/yZcrO81xZgI0xadaV45uf6Xrt6KVyjsmR+fCCQVAnlzgBR
JT1zW2vD9tqJGGlnqcPORz+6QTGSMrAgUOixzEZno1TqCyMecDWk2WflIktKFRjc
uEfksfkmDT/bEMMVvxG6AdrAbwssKbEIEwPR3R5glnyMsvLjWWWkigV+ZiWbyh5b
+3S46ku0fM4m4VMeQy3rKQGpIwbuJG2nvNUsFi7T3PfQJPE4CwRsyA61c/9eqaum
h1gsMAM5qJ3JT6KeRiClZmHyNTfcyARHf6VXifXK3tg4HDQOs1pCITL/K3sIGV4m
KEMe2EAmEhJTQVwz/7G5eAv1ptaT7Kkv49bBguZMFNH0rAhLM0ylMzBT/Wr2RTUv
1IH+zTpqMmvqxea9A7Csf4IXhp3c/CJfPgFEwGwFvfBQFNlDCdqXYvvx3r/8y4fr
H8osFSP9KojcXE1JR3aCXTL9hVy3gtBMFmNsRlWoOW4/DtMRgrKcyPVU22jhN0gT
LWntUEjmeIKQncJvzEPDxu5mVtikETJ8NGT2jNyGzhO5fzX2727Q2i+KZ99w9Gcj
WSqU7KMInq+Qsm5HBPGzRJwW9BBya7xC0oQbb/0GQAUJE1jFAgxopgDp8+Y8WVVI
5Ywr8BAazNfpk62opgq7J5m1Eotkfg4JR2PfnxO1qzUWeFL2U08qgT9ftINz8dLF
zP3ZScUU/4adlbgoFGfPsGS2zFknJ+tQQ9f9RAaaX2eOaF8JOzmBoUGzFom3m9AC
Bev2R/fGnHwJlRD0RrXARbCVjyBM3YAjhOysJjB/LrfqsmCWJm4bkSkVBZMT4bvE
J1FK2azJDzPOqZUR1AJkpimW9zTaHuTjTB9UR1suvysrYO+03AUefCcggnPzA6on
8tUPn/WQYgdNppcaC5O0WVsSZGe8hj6XZ+aIjByJMalpcRs8KaCh96tDYNluWXe+
cALu3aRKXE9SfEKBQeKH3teQ4pA/2iM6Qa6O8ZyneB4ovO5vaCuU/Ff3MD4DbxMy
dqZV0+rFkJKo0Po/XePYp6LjimCAZlDeeP+FMtB85iD+/MaZT/jwc2//cQs7RHKY
DwjpyYxV+K8k8xOFb2l9570AvIhMQoDT20JqKnpMR7gMJ/x2kKWHcD5fCSocM57+
zW5I0MduzZGa5WkVdo1bj5ymUo5BgLMFZDZOj7mC1rXx07jheZLr+nX01owhUnaE
0WCaNcT45TliRDGh8TdoJGJdCkmtEzJoH+WT9NHU2HXzUNXw5mYq58VAakJUfddF
e0i699I1wlpdkxKp7o0xP7CirJ+txA9XtuHxojV1sLM2LtJ1loEJAKHCArNkj/X+
btMLSehrm02QGbh+a7ZDKzehdMlZV3RPKBq+VoIO5AUs1TN/hMITayPf8uLhEU+H
XKCUmYwSbupISW8n7VucDB2ZpzKR1Wu0gN0HoB/bWNs7KlAyNsdqLWj9vft7D9s1
wCcSiYDi42w+/bsoBB3GZ5CcMqyg7j5z+SvKNl+P/lvKM0hVO+NB7aIiQwgorVM2
LFivWAaRov5yKJt7dPSiWyzmtMa5oW/a2wmJ2B/m2BTmXZAwXiWkMB1y71IB1TVE
oJDgVEfAyXzKge03cetgBJXKSDw1WBLnpimMpuYq6J/7z2x30FJ9uxFko2r5HPB4
04LGGMeWef52ZIgH6P4KV6EB45W54MFo1t8mTUU9OpPbMg6ekoSdD7GKcTFiPzdq
2lpwIRYI96ZTIPZkSWyXl1hg5mFMLivSnTUGzi/VeJCxYOyKrWy48/XM5z2ooLOx
RGmMg8HQCer0oPdDAj5xtxy4k9jUEHHDOqofaTdlt+oUmwStii4Dx5pqfC1XbSHC
Auvhjjn4rF9GdAO8WaNY5NKo0AozHzSDSr1x3+809NkQyGA/VlnxmwJB9Wkucq5Z
DOnVGAfFOc3ZZuEt2NZtYBEgkDQZs8wJmgU95BIaTD7wEo8YJtSHKrbhAIUO3Jgv
XcXVWVYpI7RBlEjFhjGtuLgnpx7SRHx7Cb2ogKt/zgmrVke9LxLhlRuk5i83H1yC
jVHG0u2CLpwETEhJm2i/gjx9IeMwiUdWOFcOzl9P3a6aHf8MXvkglpmoUVMEmARz
m5xoOO02QiZj+iLIeh1JOY5EbSeEC4NlTwDMUBSMDME56Y86qYPh9siNwmkz6yPp
ZfntFPOBmI64uyduvbIoEdzOzEYgvzsuCqj9mEGbU/+KowdYPyF8tNjXcfULsSGo
iHsKAC5ye0bodMNrWkr8X4DXEF4sC9m/GljDeIG8Oj3AF0qoxrv7jj8M2IuEOtbz
2tTDDlXeHH7tFNukMpmB4DUAno1zLwLOZy6JYhvPFn5K2Exe5E+AQPtUelzNZxnU
zhzAdiB6N5lTVttAKv5RutcQ4GOtqdjHQ18OgtvEdB/EiCDM46kr+wYIe2B71waR
k9vgJ/YSZJVR9CJH4yyQGb6VB0b12dvGQFVLcitaKS9+aRqZR2XouwF+mzIJFlV6
VtBXndfDxZS9bVfEakYuD0ea4DDIs5znOFEO7IfzCHsBjPxIjNY00XY5cgXT/LPa
B37pb89MmJyRsxW4mcW7u1eJqC7sfBwQ9yvO+e1VJBJEH5+gunqYc4YORzFfep8I
gxq8lLHbtosBaIar4NHR2CzrVqZBNzLyR6r7xcYnLyiljpRmyRRmiZq2Lx7mP+0d
MMhtP6Flj+FY+yXiElWg0YIxtbyqsCodPfBbsdErT/pqGuWgW8HoXcl/kqU+6Z8V
sGa/hlwss6Jt+WNvfKuvEb9VltDXPn01q4/7dI5Qu1XCwSGOnRcGr6yoSNtw/XsW
Fc1my0gFgGqnAdhDEB5p1lZ4E5YOZ8Xjqh33+RVtVbHYDXBkDezHQ0flPyy5X6jy
c1yQUdPj+DXLmzaDKL/3/WCCGz29gGkqGhrWPXDJO2O6aoydfDN4kNhIzRkFz8R8
IQtibwjuhpxeNLwsH2AJOl9kC4uc+qR771g/yk74iUKknmeIMQ9kFlaj8xB+UJrQ
l/ovhlizxob/lBsrj0bqt1F9taanks3hHVKxqt8qW+yhz3id1jd3Wo7qiwT1feaG
9GNdWz4Q/4P46HZBb0COTUNu6JtZxusmVfcO7/M+U+Bqq9MvvRQ9ieI4rEGs2TBK
FrmWhz0EvxrhwD16be20as/7GK4OVGK5l27sPWcWwfTk4hn/8UX3zU7z3G/BwbKe
UHC+nOK1q8G7TBo2AV6pB8dUy2eeAPKVCSzDlh1RBJKE7996bdGq+P3pltFX07O0
Ef2yZ2AxudfWkY06rEhWlio65X5LyII9mKyp92xXAq1YcIDAPQRS2faHh07WOgMw
Ku91rnhxmNfiw2upi6pTlUDuSudGV3dWbboI08tgMizG+zaJs1aC6GoC9at0JWbl
wUTgfING75PIIJIWld8xO9h0Lcr+05l7MnGPGiCcUtKZg2Xl4KorvT+dIEXHM1JG
mDpCYmTuqtmzZ7YVS0pAM0ghdsKcgGXuEy8ouW4C/VzIpon4AT/10iu/qH3Q0Uf+
KVCFeWPJM/pkXPecuzAtUMJ44CLOgtqIGQ57tQRgeO1SoroHY6ksl1WVsDnbxyam
oSiasKL/nLUMRcNN+cS/991f0zvLoBI+Tid2XHVdfG7K9JYq1bNRvMolgW8JHTHp
EoSof8IBv8tUnFmRN2qVL4i5SCF9Fal8lHMz3pQ3dzWZxWhnTb2BZClLs4IJeXxF
n3p10ebfHOAZ9vCqdBwGu7neB6NlNC7Vq96wwaEMH3921GAjXg7TFpvqSGreDyCd
D6h0TfJ4y0Xe7ylIgX/0/7CXo+g27kQ8K4XGWQ/ZgcvfQk3CtvnzuceFaFT51GdW
1iqjABWtEG3N4t8dbL9S7vZe047cKeIrXYOAmhULKX1cr1r1sBYh2tQ8I5Hw7gY7
oOrCElpLwUSOgga2ANkGNOqtUJzgNzBqSe6qgv1oNRlmideFJ3CoMBehjgtFumhO
iNvUOHlhATQa95rV/ueHok1vwu4Sqnpl1BAztiUtaJKSpnaKC/qmryAyJMS7vGdN
FfucciUBbws36U5JgEAXE3yfHMZTluufOPIILPfXtcRD/6/Pt0HIp36RwIcNK9Xl
x8iO6s4I/f8KaBpQzv/FOOIprzKz2VMjwGz+U8unlHLwfmNhyGjlShKAqVq5NSub
WCFRSNLj8QAXcN1+wT7d9fEGC5GK79Cols8Gh7I4X7Wz/2zUaIpx39GXfBFLt9s+
DoGoP24xtZNRuFwnnCIp88Ez5vmrYJAIt2fAY0BJQaYxdiR6YsNwYYPqe3Hr+Djk
myRL5las1kyWke+TBnKh2PBw2nOSca8/iBDDPgMjPrMqI71NZzuYwqDCOjs1qfll
+4TkFuROxpJIAo2etP9SzZ3eMjKHcOJs2B9MdE8rMaQChk6Y+BFrQCRRqLSLeevc
2ODx4cPOgMBCqqK6Dtm2/hrhKWCAlQXrRWsduWkU9Upva0N9EDKg4EOkmIQzo3km
TZG+T/M9/zgBgRRO2bfpjEtkreT9yWAqPZ1MYr4i8BJYE9clofUtxAnuOwKMETT3
cGRcabrfLidsgpm2M5xm+LSIC6+bAiYCQ4Tcn4Qwk+g6xJRxC1STz4M/xFMwLpS2
kdPS++gjjnmeOlE4ZrN+Fxu98QePgXEH7ljRorMXZrGiBYx+qggFGpnMitRr+bq4
2AJOdFtRBvbXBWDH89N0Wu4Kc8VGCfGgP2oyRkdkSErWzznkspFQTfe3Qz3nm32y
gztZ6/adxHF4IpvW/OnL8mU6QbGdrOP1r88Fq4NZ21X+0xqUNCneA9XQE3RgyNcn
hG7q4EzNO8ks/JN5kdzv47cptheNor+8CauDFctCDehiYIJWPTSkcnk5GnBDRFWi
yyRHRG3UkV2Zhy6+4E9qIQFBYJDN/NDF/V9oCXRa0Zf+67dmAZ6/yheR2WsZIL4d
DEVp+ziJlmsg3vXDV7d/lUSJ/BFyERsdOKlgJdbLk09M6IJBqPcbX+WFxGhlqi47
zdcOR+33JYBKhEH5J5srApns2IXGa2sUFtASfFpezO4xsl0hAsunzoFNhzFP8saS
wqLLfi/0ajM4/3wVfhcs3f9lhhjzMB6McHKmIGzeKKMv33HEq7C7dAraa67WGNQA
lIohLXbs09cujRMmF2oyxoL032oOEjVQviTmhevYfJzPVW4AoJ1TctHO3jLYXWo4
QFcAbkbV7LVafhinW6mCSC2kPCt/i01lEyk1yXkAQ45lzVcaZtpaVw9wkY9J6WnT
6J2s5DCK4T3f7lPa2o6Q0SLGNEmeF6MOQoGPeMYaIfwZ+dcZLO7CxVTfozmVSwFl
9L4ve2XKFAImowuDh0p74Xkv9wINtxVJpvAO2wGQcaalzH/y9nsFV3k1XdAg2hrG
l98PP/vqHLgbUAWJWVkNxPFlSyI4dMOjyjoTWUTGj5zFjulImwLFwAaz9NhGOso0
z/HCFKbsS56wcI+r+OO5FkjouUkHwG3fDTcZLH9LDfOk9w74YHWPeBfUm+iucYdi
gpgIzQA42Io6gVK7+yVRBTn1lCO25QVZzkpsSYZDzipZNiFdRiQ5OGxd5HPCvFoQ
DBaRL0SI2jPtS3deFbf1zBwGgX4eVjUWa9Za+zJsHNt4Mn72RQ8KOs0BtuVNrTjF
e//dB0pI+CgmZPLvyZJ+MJ391gfuNNQibUDYdyUa85bNDRsaj6hcf1jyd5o1BGfq
qH/Hn5koypnjEPPCayRtGqzQlx7IIuCvmDwbbD9AamPVda3ITpzZSt3jp0krvNdK
0XglpCfUFMy1jgScrIZB9umdA4Huo6C4iPdSPRAok/CocWgW7+qP4TrLGcEsse4B
SnyyK0kQ3c0l6JbrC1vSRV3UsT4xQSbE9FNEKt0BE7fUhdiIjMzUGO32wvCSfPwN
s5hQoa4NpUDo3I6a5yEY4tKNp6PzqSMNV+RmbJqVHOWKnPqCNR0qqbVM3Mkble3v
fExbbVx1jBZUStFg8XFvbJl3F3eanoHyNIfQZ0MQMqX9lY8OpGXhi0jX6XE8vGMU
FY15Kxu+jLiP0uoS60IZyTKS9UOpOp83dyuiFS5AQGJSTcAr6pngQtePNJFJDVim
9NdV3z2En8H4zQ47K6blGdKRgnl/ebZJzcW+PT6390QBfzatM1xNP28tO52Vy8Yl
5RAuOB6x1kA9EzCwEPvxRvLVDQOf0ghpTRlm8jpl12JvpBR5CCC4MVATVnPBGPue
fbvzp3Iho5q6ksbxy2o+ugls2WHEp2ZfzWYHhC0XgrXXK3T73jXAzxmQlNaaSeqX
988NzDKD9zOAl1G9cj/cZf5Ou79znNP13ceg/HTfTXYJMGL0sqdpuIqlRU/d9m7n
E3BAyttGNmy0I1sOClxMkGZwXu2W1I8vXmPu9E3qqHcgDeN3sxUb38g3cAVQynKX
Uui0xbudaYzWeOo2LvnhmxXfq18yJiXopZHd6Tzc4Gt196y8ZJroVZmp5oo8Dvri
HbCVgx2cpM3fsFxvoecv4aGfPbm4a0LxITXPHLU6jWbvFZHw/PWgbLJvif4kOukz
`protect END_PROTECTED
