`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeK8jCbkJatHOI19rOXvqEDr7+dfowF88kbwMDtgHOq8szjnnC68yZcjndsBYWf4
I8p4hYxCc1WVkYqWNayGNlZxookMkfoEwu/2hXnRS93yld7xMsainw6UJz6Yf61S
NvczH1O1Tcq/sWZ48qyl7LIOaD4DdcwNvwRFDYYTbYJkyUj+GilCvZhw7JxQN9ne
4LUjWT/rTq7iRZswg/XwLxVaKAyCazhNgzRvec8De9JFtIbx4Wtbdu/QcqAzR0zK
MjohPeiyUUDrSEAeGhn7nYJdqdzRvxIA+4KWPcjqssDUPFwmrG8lGGChbd+1gVI+
mr+Ftp/PVhMWa4S9MLC6AaNhDAY2knLs84sxR57DH5ZD52JaARQRgVwR2TC6geE2
pzdbs+P8cdj46O8TRP08A42Oy8chvc7d55UQMg9yJWcek/2gvV7V3nF6HERawxt3
a5rQ4Uw0uTO0r6rMbp24NEJlI3GPkCHrtyeod0nNvP3TdoR8bwD88j3B5cjCafoU
6nMtrCk3/HNWhBL5GB9VtCMUa26SbNGAssbLReuEh3hxkmdiJuGlgMWNM8ngfrAI
eRbONAMSiCR8eWN/woJPevX7YoVrt6MwZC8Q5IxP2Txau+lMXUE0wYZ1rVfbJZ/f
oSeymZbv9FJSsk7WJew9dNLVuYymjqhXk8P3QYFz3Tyqt8WAsj6pDSrOmbJohVq3
2/OjGtLLB1tuHv0LfFrT+j3GR5w1XvinMXn5O6VIfbC4/cpXFPeTbxV8FRpvngRT
QwL0jP9ep1uyGReEGV4Zoq2ySxZQuUvaDZeugwhBKBKzBr2tEVPhcmsqnoxF3yJ8
jlJTLPdYNamfhXZkDuyn03OAqERJyx2tQehlTWa24bJsATpYK89efZL28xjQ0aId
uB2xUFPznU2CBkwAGmFSyAXnyRCagKWrDNQwq+3PSFqOZh1691DFLY50qjALJGem
jloWE9TlyO9fyqtq2ju8mx0bU7yFnTMiQ4P55p+iI26MfBjS29grs2mKjixCokEK
FgubVOcfhXOUbk+9OIh+1H3srZjGzJy2OcVCfZbaH8xugn1e5sf70GQ/T71IJ/Kc
HR3DqvL8CzOiLswD/kJWq8zy0ZOldbJKrUUH4hVp7joi4JrRsuOUtuPfYibnkLWf
71X3VkzdcaP0RONULtKLvwhKsNyHDdN6G5GXdSMtIfHWiMuf4Icw3J74Hvsdmehb
WWBtvRaATTP0w/NGmjAEinnq7ugFA47hSc3Izkl+cM3VGJytNPXD1xWZ7b/7A9yI
`protect END_PROTECTED
