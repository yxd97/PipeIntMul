`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
smKvMT6ojLUZKe1Wdec2tR4G47tyx7pJuRdcFP7pOkobkxBqeWPw3Q0gZWcU1Qyf
diaZJS2TzWKRb/1k/0Oj9oSwS2HY/7IWa7VBpaBDRffEG3EiQB5CuILqF9h6ROt0
0dVJeYdLw0NRKaniSSQLIZwgzjBNq3cY4jfrWXdkFz++7T/oTlRO1Eq+QQYwv6FM
sg65vkSXI2nhjzXaBXG6/ArIVqS15X0vekpcVw8svuW49ySJQSyfHFOTEu/Vm5OQ
zakWGAdNZT6jXEsNfepL+rHlEmDL1iaYbIcwkmfGu2aHu1vmjxVZTiRbXUF/Uojt
eHdT3BzUoXTxmCee7yeUVu3gZS0EFSlfsPnw7hFaAsCqddMajPc8zqY7pX2daVCX
/pm59X2aLvHB4+ah+qF9d6iYTkPkTL7eetE39I3/85FWIN8BD/wmSnzMeD8xjDXw
kDtxzUtDVQBnyoTL5+M1OveSjWZxhY6X/I05IhgXq2gwrUOXF0RpRdN3CtP4QPZa
i15bYCLKQyyONJoEu8eEwrw/wTO5ZrGmBjG62UR0VCc=
`protect END_PROTECTED
