`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TemG9e+mSi7I89yRHddobFMgx29ckO2iTDa/70cjIcmIdugGvwa/0Z7O7a9DyKFl
tWvTjREZwgFBQGTO0Xs+Tp+P/RPiG3A2zM29am3ZIrtl5feSjxaxhwxfoSts7/Tm
lSK0aeuFJh5GQGrwHb4lbUNbyueO/lsyUlgVT/MGmT6ox4qh9vaAOek9MkaqlN5w
1qtfZTdSbBbkkF51GkORlkDEcK28zzaZeN4RHSpuCUy36/KFTRbLHgac4RGQYu9X
m5sCOOQ5RgrbRqF/bGcwsuGgALFOQkJWYAIQsDar445vfOPMjXGw0/6XTPammAeu
yvhckWIGiNieEWmUro16/w==
`protect END_PROTECTED
