`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RObvx0ZWvAuu6JWByCcgG7/BVZhsCX+tHk3TgMe+J5/RzZLDiyFjrOKNaSsX4Ntt
dOElFXenCmqKLY94HERbjF8/RoqKGmeahNflior5f6uohPL5NrwYTDpOwWWgrgjE
vYw9iNjmB9sqPsFI6sHSlfclJxRxbI9VtSkk0OihpGhgP+R9bReLTjvjk3pEN0Dt
sBWARlg9esW/gwx8/JcnoUWyr8rXIlQWyTP7OfpEamq7QuoC4tscA7M7z9McuFdh
`protect END_PROTECTED
