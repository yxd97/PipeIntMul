`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OhzMDcOZ2lzA5zGp2c21EiKsIY1PL1/Gz6gK9CQjdslVkgAxFD6R/OCoqYs7Pexp
vxaT2vXeBgAEBvxg/N5mYEP008bET+zrSeEtsyw2FwueOkHIpM0FVmLqJF4EdzjF
kA6aUTd3xEN7mUmzqxRpSznjRCyrp0/1crYIeqiyPBaQL831CbM1qQr5TMljaS5D
Sc/Afw04qmD1BXYuqpGeQwFALlD9G7So5VZOQVC2/oermEaEjWjYe+dxzn54W9lW
wolWmQAfdrYPWPOe4RY2BRAR7ZZPiNdnNgDU+lFLLiIkPb8QLIbzXFFQw6MuXK8U
WO7qyQfEbRO+4BiIeK4q/DYbqLz4mIZa0dxiSASQQH4JH2XloMgEzhljSYbKjJCU
KgAoCLuWcmHpYHWj6CBekpypoILoXL80ymYVaqb7QUq7abayktgj1Ut4bsA+DcMM
3ttsK6Qyo+K34WVDEKrPTPPGtg1hXEFrW2urU8j5OGD1lCK4Pi/nH47/wc9FXOvX
FMtgUtQVtI9nB40aKRPYEtYTsWOYVSHvX/Dz98j2s5wamsGReOcqVX0fjU3MB/S8
CElXZHV3eleX0DfOKl+DdqE2O7TRB2rrQTV+zNV0cS/lTZ6Jy4zJf9J9qr9dX2fD
45bQD8GpFb4hchu/NO14XK6XS0UoUgqOlIeT/f9VOXKRKvG7+m+3rTxEy/2Gk95i
Ig+F+LPvYUTyxf89z2g+q3Qtw5kTxXQBugVXdBS351oW0FdvSlSYHezQ403zp5AM
vJaJeZ5Zb1uPnSOlISq9mZOZqrgGIfBpDaKNJoh4ihAfoVDJHaC+M/9nHQPYJnG/
SujNfpTvN0Z9nFXIpZNVQW1PJCrl/dqVdJW8D64DnZx7QN60TDamRkV7uxtv2usl
UWvb1z9NFYhWniqb2iZntgJAjzz4gi1C5CoUXog0Rv9LKN+vGt0PqcKOtPqTRoWB
XuDxMoYg5WIW93ZPF1G9OMh0e4KWZ/I55nT8swn2CSKoGVdL0QOVmXp4VgqsfsVm
wCzO7FYX5J4y4zdqDdS7k/ukvlQjvjubKhiyJ9InK76WUXxPlQbZhGR04uShnBUw
9s2my0NXXkG9HMsse3Fr+VouZbFYRhffUQk0UGSV9apO3CFKVolI36zIJqTdUsnn
e6jlUaKESCysZ9iFOnMZGvvTXjV/WjV5xdGaxIuywl+YZVJ/KwsM3Nt54CEoQ1Uq
LEHI05eq1VQiC8BF6fuBcAla0P+iFIABHCt6QyMqVMw+e6sBbbXui2i7J6vqqceJ
qgOdgxrL02kZ6IOZAddHCVmDZ7Wvyy/s0V2kyupAMV0uuLqQo2EnIlbYssGK97Ve
/NtxKTby+jGsif+4Im94FHYmcLktqmMlb+3l0mGRwFIAu9rzAA6ItxD3FjtPCgDU
Ns3sJ6ApGWueYfveUoD7N2ma999+BGtMFyKXd8n3/1xCLEdbaceRGlOEl7Wl7z1P
bW5y2dhVZ3hftUnZwzKP+tfFd9+MaDjJNDCnwkhVzspnSbk6N/D+6h4fvoTKasgY
g+UPLbDgOJ+o+IIWEKes2IP65D96hp4JQDSNOSoztwHnU0dHn3xZRVcauwntljIK
aVXXRwE9Jrf5Hdo+dulxVsly/S3KI9+5r8PCL4jHOPFTAw3kdV7h2z8BnP5jXB2h
OHbgWt7W6w8ZkyuXZrOQsH/+lro4tL2AxLJDiVsCNFaYOyQLr6vxrEILuQrbRKfn
AdaRcvCithNLHjg37g78WQKfGUHrXfWoKMZ3YN+eG+BhnZ+ZU19WwjO+OZUV1ASC
djjAmSxaHll7KpJ0T1ubVmFkcEVeJUDcsiyXG7b7wc4wOzTlCHr66JwkURUlNBjX
cs0XcFgW0gNjUGI2Mmb/+DmjBOfqfPsAFq/Tw2sdaR6boXI7M2h5Uxu3pyAlKsYp
KJ0aBsJRU7AYcZ8LUYn24HQUqxqf4HAZVFc8mKXeqkGCMlKXxVO1dbEsanQwr/yd
Tqb5sL3HRx20DBMBqFjpRu2Jfq3k5sW1rsbLlfVpmGjM85Khn5MIJuQDLKAYLqBi
qelZ9wMFJCKAj4wKfFOjgYLjGJi+xxWk3yOPOx7ZIxw=
`protect END_PROTECTED
