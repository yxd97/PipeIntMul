`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0+xoPdiT02uKglY3NaSHHoKS6BNyRd8FPD+H88Tvtx/zLK7fkAyRYWDS1DcDBGDc
KT0b6fU6fG7fYljQ7sI5ykdjoG7YfoWMDYVIrftbuHF1smUtX+6Qm2YehPtSgFSL
SF59ArldkGpx/BQxV6IG52cfiPtPoay4A1asUjlI1C3jnTbwpbemQSGDiEJzOP0A
WXThcJ55g9fLEwPoXVzmamW2jji7WM3ATEebDFW6bGWLgxGbrdQvsVPi3dTG2SSg
akTSMg9aYjqAeJTkniYA8kaNyR7A9BqTIanR0tFUQbCVwtxZmnFtT8JraFF1CWgA
6aZU7iOjKN46EebKJ3xVJKKypngW+QsOscjDgTWXRblX65fm5Bk4OfIi/3JFTu/P
iI/TA9IhycsEjncOnLRYUIkXXjD11CwdhMUuS6Z6pbHZZFBBWoPD6I5YKIn7nJHM
zTqcrkOfLu7Gx3IAHqOvmpLImkjqwjtcSkIYK2k5rZ8gLNop4KU8ugbibrl3YVAp
s/cQq3tPTwUXgMdmwlDzVL4NrGFBDtSTtJln+0gY9vgppNIpuM0Wc9/Mc6QVZjj+
+sgeSPgoXzT5JYgGRmwCPPkqzrY0t4KTAbURA4PvU//acbNpcX9h5uDjCGCFEAwe
VOAIhjlJwI7tT6ndbDcSgEbTEYKAPZiVbT1yl6HF0rQyujG8LW6DPTn7EdJu136n
kcFMYR0ipcJHeqVvuhdmZ7PnDfKrcQW6R+uVBHFuAWYt8EbvA0grINBAspNe5Oq5
auMVN78up/IHtcRSjQEB7XnII6EeMnxYpkqvzMRqaHX7UA5+2wWAY+6VkeXgauEC
VUt8fFYc807l3bgAQSSj2IWkoeolp56M1eRZ9P60qKt/mCE1IWLF30C4pjBxKuzg
5FOflz1B0gY5qvE1qL6ynqtioeC+ADkF6Rx45q05TycLpONYWbs03Q1kBNg6JtK4
zm1eOGLwnCKpUUgY4ifu8QNBZd+9/DHMbd0CH48d1fOG+iiHNDV1e9PFRHbG6v5z
ffnIJIvy2N0jS7YNu8dmrFw/LEVb6pm0GpKlIODmLi4YNhf/zl/16DvHyJasYCIz
StSRVLlXmGKT7UctPgGpYsgU0zRbrKosRcvcUrVoJfP0Oji0G/274UpAWE9nvBh8
Syz89CZ+EqW3OCznaNagz3zp6UFLhdi2YM4MtywgEUC0grsEK3HfpWZZLba1vjrq
o0KUc0TcFTa16HYrCztEl0VAjAcQ4fgBolOovE6eN7CG0vVueuFI3nrMaSabEgu5
OpLp2RNahdGZUtraFoOvZG1tivt3Rr4FsuF4IxGoHIi0vyD3RNKntH4J0oXksc+B
GLyLht5B/GnCoAsXG+wekuqc5dZHPd6UHcJpWc1eFLDDnEeN7JMevmwHLb9fMAUM
JaouvhWB+YqMS86iBmmRbgbdobvsPmcAXWEwK7NlAq3DePEoNn3x+rOrG77lLt98
`protect END_PROTECTED
