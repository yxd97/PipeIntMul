`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYYDo6CAvdNPb0RVPs2LxoUBcgDGazOdP+K3YdTuZBPB+k3xoHpPw6LymdMj/18e
LI3wxlJRFWRZye1byq//TTsW+D9pY8BqQzU87RkgoyJNdgf95KS7x+nOGYwi416f
sSr7LxgpnlBPohZ1bC+PGRLjmwkZ4CuCSDp/5CZESB00NiAfmYZ5NC3qyh3V55H5
URxpNh7Gk2C0p7cGUCkGqHAAULAY1K548zts3ezQKY0PC5FkkMhimYEGDdhR2UWM
TW/apLjQ/ABvrpxg67q7Bg==
`protect END_PROTECTED
