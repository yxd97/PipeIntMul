`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNcAw+Chn+PtJUGbeN1zivjdhV1/m0MtGl7plXZTAHDGu/ZvqPitC8LP5PXDbmBN
Cg5I8iFwX21y92ZhbIBieYGutf95Ix3ljr3aXkok4nQselQ2hD9Q+0C4SIBwzmwj
3ThtFEmADlXWg5SZWtv10+2GFWTYYnLtvCA+L1HvlBMcljJbT1zDebM8Ip10xUVF
1JC+LLyGJUjCYRVfkqX4QMoT8lKDREvksDkfGfSIh0OOtDGK2LrCMMMUXsjvFtZd
XoqTdPjaxw5FkJEAI+JNXwHHgrYBSGcM8RL/gW2uw6N0KY79/1tZ4RR6FFW3l+ib
fwjFtbXyAeocldtjblTpC18lE/vwGcwInTmEOwpVG56X3M7uU7u9as763hF0QCV4
g2dieZGdmT15WCuKre3ldufUuPmiNV34Q8ERvWnlTX5zJViapDw9w4EtsEMZBGCK
smSuSFitrDV+QLz6KyBsCnFDI8wZE+X+oFWaBkypgTxleRRcmFb4HKwNRNw6hdPy
`protect END_PROTECTED
