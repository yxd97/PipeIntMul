`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYhtXS2AWJ1+T5AejP3MfR7u7kXANSuslKPpCaGqtIUS/uzjRVGrNE0E4X5FQHJH
hHWPIfrP3eE6wxioFSKWHhA2XLtMoGTNj6aFuzbu58LxBJZzM3pmoF2XBUGW7p9M
WL4YRc59VPdVa/WFqXTDu3o3XhMvBkHIofX9EIfWnc+9/0xmzDIFKE2w0/KbYucV
9Bk9VxoLEOwIv7gSKp1JQefMRNWAmoq5sb31boJB1xmCuauRhloPLQF0i+dwV3SW
af+gXwi94j4B1fO3zsvt4k+4ZxQPt+m0nc0oHCaEYjteK3tWBDwqTW1JScGU2LKY
YrrEIgHXbqR2Vlwjouq/HGtWx5CADH17BNki8QcuX9KfVCt+N5FDRiUp8yfFkYtf
R2LC1SlHUbef8P2Dw2v15nWEnNinvvKpn/TdQVyjxp+KonZIlXM/Xk41A6fG8ihG
2YXtVIivmwZo+CDI7YMB0qD7EknLS28PDiBua2velpQtjusYJOiOSdZMQCyCDH6Q
TFRiNm0yN7w7QLTIGLuoKqVvtfFWqRL88l9DA3OBSOkTAWTOcIXBvMwifJ7BRrCi
3/vzZEflKrxrspl7nJRAXcoz9upidvaUi5F8f4O0WFGJpuSQH98Qet+vyWs8idIQ
1+OSK3oYKhhtqShzfE6bVkx6W+xoPMpTn3z4Qy+N6Mc56X2+M8kN5nDB4VQ++BVh
uOj0r8YjWbwi+WyVeyyI+nfC01GgODWPMVjUPdcI5f/YUqfboKgeQnd9ZxGf2XoF
JKwzkKc/fnNzbVXhGnJgFQGkMM41G7vWqDVXBPVWSPUrrfE+3TZsVkeGi4599Bvf
NaPH+xCM/dJLaGQ2qhOnBgQsZ+XOchQ2tfkxGHL+rTmevWECJ/4No/huWct/RfgN
MyOeksl3ISr9rAFkNCgCP93T3NSyiacXg4inMM5QjDIAG0V/eSL5cVuCtRjRkjJ4
SnOFZeOISJyMRi5vY9Q+lwG1dcqnsqlGulKXPsJKFe3IVuGqjl5RUq8KTbeaP7za
QckMJGbHHnhoA5DP/wXuQ0A/QeGLrtouDmuTrD3eVdI2GRBSThu7VCCxGmfbaJdc
woSRJrIpWzSEIWVob4um0JNIyqPl9KhJfxMr5UEKlXQZZbbZc8vg7Lul383KPFNx
mkCk/ohx8MkTPIp0c7MsjZGhsl+Omqsu9p3N/NM9KSz0nY2Ro9KZgokLQn/YsLa7
2AZRCEJVyng+un8f7sLP0pyHBq9nq7mlSJP9hzIe3QXwb+cT/ZtsvyVCxUuY0Qif
r/0fbmfgHmfsMD/aW/exZ80ZexPXV+bNT8tolHXzkgNi+0AxW6ziCrR4qWbOJQGi
vtF2muLbiuoUyfh0nD+XJB1qQwpyeaetRHVGFRyJdW61hgEGOHpH25X/AG7PyRHc
T7oWNtnprhuqnRRnxPOnENYOhgzS+xfZ1/9OsZN/yNokw4Qni2lMVPJQgoXeEr8E
nKQlfxNeucEeQqRTeQHHkxR8b5mv31Aw7lU1TR+g3Epf5B/66pZNMI4m+ySs4eSp
YHrugvuE6gPCjESs2oj2gIflpMxOQLBBaCCUVuvtVo8VyVYKw+xYHR/UWdIudxCZ
ac4WHEME63kC1M+zmL5+fXiheyI9BVRjP3UDe09SxdU0u/+gVL9N5MkKpkePs56P
cqRGupVYmER8l74o5JmUTxiblAsJ2ScPrFxjPS4bkWljvAVOz9FxfHEAF/+WQbpX
6gn+JSd6vBrgtQtagq3ggDabd3ocBf4aSwS+VhzHz0WfWl0onCnt6NqtS5iYApue
+D+CU2bbhw92Vnj59qDXwz2gOtZc1Ten2DWNJBwgvl8Z0Drqyzk5ELObpli959ry
PufSjxMKFeWcUMnxm6dnyyXkOgbIiyCIjjA4H32Oj0JrZ3Hzu/hSsXerlHLA9LnI
D1gXjVgZjDfY1Ak1I1+MknlRrTe7awE1iHMAUAtitIikTCtXOmJwBbRqWnf/lmI5
rP1DzDyzvRAwkfphb3Yij/e5p700trQI56fehZfEHfgrdJldwjPiXVrcRaLYHv7Y
1IEpnfSbp0O+521kBL4o8UCIvodT5ASZGtADWn/7euPSfpVL+5buDITAr6zG46ms
jtX3qvxOrvRmhkchwb2MrnnYBJhKjEblgS1EuHTTJ5oXu6EzsnKybwO2negqQtb0
kstNDif+CKw0ceYgH/3nJsyM39vwL1SOKyLFSvfi8YDBQplOr0t4sz+HHeeMiGk6
mSGWvyNp/wV3hfAxji+99FnLsXc5RS6LumnAvLWMXuboGpUI4NJQB6ob7+QEiIJG
/9xDuB8xWBIyVobIMFUyeyxbpYICn+Kv8oZVImaHteSJkAWuRNNVS9DYfWhdQjKv
lcMNMnAYcBOZEvBMNr9Een7iDSUTTtq+WWHJvs+5UQE+c12BMPdnEq0iMiObL7rQ
aKP80rM0/gvWEI+FXgO2wDkz40SwbJkRcvccN4AajL71uTpJ6ujD3/78lViKSVsL
dtwTeEXwz/nr5QtYUy625RZYStu5Mgy3Du83OaLeX8pc4FI8KfzXeITdFaCM9ldV
1iZO0ZkLr02mhGITjtOAHNda0E5PxovKfKb64h+zLkX5a3jwM7S+x3nEwimgEnAO
DYOFwVht/BGRKHRCUq5NdoT3gjZ8jPU94VpvoGNZ9OXpGBUxDn8x1d5PR7V9xVWT
67HC5rWAT6sSNDg/HM/yqiFeKvdR3PYVAk1qyJ1GQ+PSVtPfwajeL1I3NIVD1YDu
SIU596rr0K6zlZZa1UC9+8ZNgB4oyeF/NNpPwksy3ADdr84d54TLWPlHQMm1PDkt
1WwzI1LGizLxnsEWwT2noA79HKtJtOjPjXH8e3K51IGoEeyfrxCml5m0D8jSdU3B
MGHku7e3KFuDBmEzivFVnk9jwHfAox63ixqCk/6Mhio0KOArgdLTdcD4vTVUuod4
MA2raEZXEcoHI9/dF4hYECMaZ38JJwkiO6WuDglPggnB1E6cqwaepiJFpgSvy2Dw
pfc8sfsPeF/sEz/MMGN1VlaFZuKWulRnihBpQbVqLUnlZQzzFu6bnUki2GWsRyU6
MLjHrvdAPxxS2ASvS+L6VapwKZjtwpZk/yANd9guUupIVEss9usm48foQCU6B7AB
UhcavW+qZQFuXXWqyjZEnjHyBm3X8tAkrYPmBu3XGAcXT+S1UHq2kpdKZaqCpPMS
KTXXE3TMV+qhMKkTXUfwWN6IaJ8+NQ2Jy9J0GE77XameTRbOjA/dwLy0AqAA9KqS
hd+xbEfMqBGQmpihpg+3fG80YuH1KgEnvQWyxqoByYLMr8uVqFaTpMyXFCBu5Ide
Tpx8jgOQk6Fa5oC5P8Zf59FPKVJqsjC8u1tDjo0B7SKLjks+2auV1/0+MztzZLaO
JP4gkKpiPIZHSiBkiusLHvmFZxbTJ3gyfiLh09Iknrk107QXSlI6Q5VSHt9hjFW1
PkLPIXdZ3t0LNbctQ76vJB/LeK/dloyxPu2bAhat2ec3Mf7CoqseDbCEV2c9Sup6
A/H/7rclxJc1DGw7zTBNKK0LhT6EF78HVnT2auFuQVxpx8WID/a/q5nbohHE5k7l
g5s9EX0a7rx/HqfDIlPBLI/07CrEQVbhipBlU6SNqITtURraraU6JNRWUE317i1K
i0RbLgSLwm8f2H1g1EFQTWSSlGwQwy+0PeegfKOHrPo5dCuR/FacXxFrPXpasNGc
xaQ/h+gmYN7OASjz+qcVKNc6daF6j6vMe8Ay8GbGqITRftY1nYqxJbNhqJbCgOLe
JjCwHJCebHal+9R/4qa6GgMruJkPkV1r2Nhc4eCatUXhcPvU6Q3qxg1Tm7y9z/UY
uTPEh5F6EWTnjEoSGKh95M0CUUZw8CPXS3J4tNm6p0KVZadf3iccelkMpxnPdbqK
RnL6F0zl6N2fh9HPIS8kSu+qbJCABeHBq836Wm1kRIMAyXpveFU56YaMGobt8HXg
cQMfnwqinJq0p3BYRLVM1y0AehP9MOcxIY7rLDua8rIlEOv1/3dHXCeVnFnZ9fu4
UaXXUHE9yYQESEnKxssK/g9fZpCpEhITLpXFkIiDoaKJznAyvJ/UtKFhnfcgt534
c/wzfD+INGtdCJzYLKSo9Qre/bOTJ3U30/wPzLqd8v9FUhVZd4Y6BV0vFtHYgAS/
0WV/nX3znnYsOMB/j4n0jNx0U4LAVZ0EMlhgYZP1I3VA8KXGPp73iy7dvkNPx+uV
HjQ3MSL8CltOqhdwaWSlGmeD1OOynOW7yfl9XbK5MgOszqdEsydKSTiJM0ywjff1
FYwi/FEIWTg063vp1tk6uzno26l6ZN2GVK8Qdg5eIZkDW02dVBALSJMlRmeF6lZr
iMzewWNX1OY7J6VE0HAoIPvoTya6Tnv6za92PZb7F42qKZIc9R7BtQq1AVdYLvP4
HXt+IiPYdXmvUEJRr/dIYhVcmRGm+RMXnI3ECI99LhIV2kMQCJEM2RjUE7T8BSGD
p/0LK3PPpuxajylCyWMt/mj+2rlBYwuiB4FPFUX465l0r408ulGfWolQUxOcRprN
n9doJ7qTQtsFFiNNyC8Mzer36XhQpkZilhGm4OA1dntK+mqZKwRDfkFkOOnsARb/
se5GRHrFXUgTk92RYmkYz9JtjNUnFCyBSP0p7eh3dHtkbdn8u32fYiHVaOZZRul4
1xAYNKcb9n8jhVslsaHnQ+eKbnK39Ae353hBMUrjhfcMaa8FbT5eEWsqunx3TNk/
B3wg7jbUyU1KMJugMTzm6wjV9CZSlRqaawFpLzzBW9pkc9yHd8mGldE7/zgtQtWE
ZbTZ6pdSvlrfTaZXBmCirv3QyY6bsLMEs3C4Cc4UNLdcNB8fZdHZsiU9tWrkPI/8
CLuFljRR9D7zf/UFWRMnd7XlJnmhK71nNvW5NBVf40EUItaTvVrltg1eBa2wjFkj
egEf9a8/u3i48oej9LdkaYX/SZ08z0XRZ2PANVChathC3Xz3siucoBbjS0Z8cU7D
LMkFhy5SS8amz+mQYlM3beuNVzRVbPM72/qjygqkWkQ8BImSGOE5Hri7kZ7BjDKa
mmFz6fbHIpzLWq1bEe+L6QmgL5SvOh82JQE1wf7tt/lJ1/LgP/RkwgvWFWhwrSw4
dFZo5moPkeMhoqVVc3RyTBJzdCQH5PMMgS87aVGGSj+qMW/cS4+sDeCYrlKN21lB
yXJUOlW/WoINbn+b6cLz/dFUpvMmeg74JUIKuzQLfrZ6Vs3iLzMLSe48Op6elh+4
fB4Kzx6JzVYx7jlHHWzFX8QRph/RINDotOgRaTnpFg535lNPtBrm+/j34pwZxYnK
Y7IrSorvrArx5H5+pukkHuiAiD6eMSzsjJbouT1b2PQinu3Xumuelu2+QcZFY8Ct
bfz25iQNP03hntkkJU1Kbp141m1qJbLVajPS7167fl6zUveAOzz/AxlNZGywl2P0
/LEXPqrU0T8hWfkj5maDV1Bhwi8sI5mOtIlkEGvglCufaXEn2IgjQgACxIugGyyT
rqPOt4KFTagl1PXCm2+sy3qMolcUIoJisHjk6upjCx/esYjSiS3fmKi3Gv0lpg/y
jNDz53j5uHlHf+u4W35F5RsZCMUyeYqgrGCbArxj6tFRPIIRJRed0xboRGLRSp5x
vG/9XTE6D0mwo6wd5V34zCsll9rv2kh9oHtyFkOfkEJW0E3NY3lV0P9Se6/voupS
Za9b6K6pWgCyN9mTffrAnj6e9aj9TOgrbmuVrRIdN1jwE49Jhdgw9EMYWM390jQ6
hwM6gtHS+xldHjne182EX8Ij/pCycfbHv9qid1Z+abtVQP8UqZWHjFddTHLTbieh
UNijvAwpqYzZmXFjEATWEVRp2BkHjB2b77ZkaK5d+nBonbcONhN3+Rsj/KkniVcc
+SfB+GZvu43x1Lv2GFZeiNA7feWD36V4QRPYC4EvkmuXJ3f6+k/pU02w8jKsrFov
1VyX48qpgWavQlbJckYNpWDoFJU54GIxvw1N90Og0eA72v3sHhBkONP8DtdcAtP6
hfpaKEZtCctui1RD2J7WaKxtEf80tuBj1w06tAaCwh/N+Zl/qlbZ6fHCwgWZ+NWA
0F2tAH2aiIrE/UBtQPNRXV97p3nZV1xjmpL4JdOsoUYn4/+4fbNz8GqRQkogUSs8
PpNDQSWwQ4c3Fb8mF7yqJvOufdaEuOmpsmbYG7pPZ/u58nJq2CRdZQ2BifboqhUb
XzZl+FRAEH0xKl4OaI8V1fmk3kmSjD/VSN1siXKp1emoTMQ75OyQZOjlGCh88Dga
85wkZ0P9yGc2R2OPG5aZ9JYHVHOLcW6GRC8tQnHo6d5yaUY2vEdOfj93fACQ4pur
LhjEXfe4aUwkwGE932ZzhZDw2+NvrmjaiHmnQBjpN6Qyyg6MbC/YdAoCEaelJBMZ
PU4Q60WO7QpZUa84FvUNfn/j7EF/ZpiCbff1d48Kerf0mwJ74xM+5YE7TmjkNVLc
QwbnenLHg8+G6uiVXWwWyRxgpUBq3JW9hYbP1LJpHFp+NJK+hqQShq9qSaYF9eCR
x9+nVCcyY/okZUD/CeSrVPDtD7wHUDbkOIOf+bo6V6jaWlr/8kuTY3UjE2+mhwoM
7fecgDOd1ELiMimNrYIFf/fgYbS77kSq+hYwpAx1eGSL1VhdyNEUfEEHQlZe/RKe
Y9sMisjtqKUSJiSHPsxJhn4qe/cu07cAU1R9RQ2bVwaL+lJeTGzfmzEF39d+oi4r
4b46F7uaVxxRBXsTSR+gWcGHBkk3FRzlt9plviJ7scQTwSVq2dJtpdDg81QBQese
VunHu6zUOPUjDHgNUKvxxs2Coht43uKrT1JF18cic8tRHA4vpV/1Yk6RhS3ZyjAT
hGBazveAp6iFGlPW4WH8U998tDRJR2iouAOONfgpruo2Jx+FpXbDMTVg2IUNI+m7
ShDlLtIPbEKJaymeJujGQuDUcIhxF6Nn1KToIfkGMBv0DX6RvdRo1haXOX5M+s85
rgm8qe5hrKeV1+Me3vpI4sK81QzJA8q041/oVe2KLwCdgDPnv+7prhlwrbvfkB++
SrItLQ8LSObp4oTPbyP4qlQVQuTBtpXZ6YtkxdZHnOb20XQYz+A+uHI2X5bKHBsl
XaJtR6sPvQZUQBekjCx2v57L61iab8TxWpxDksLiqN3rmHSIhSiXVN5O34Il9dux
txG5m/1Ucwbi+lusMwA2/U2kumfecxn4G3QL4sGCnp+ym139rw4KtLcZn+iQmavD
qSKyM4OBoi6K3/kR/OpVeQ==
`protect END_PROTECTED
