`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LcBV8Y4qeBMpUrqLNVEWlJUyDge11XfpvDbAOXzOI0nXt6JRAJnUNIuZRZifOeGb
FLBuyVluOz0vNgoVn7LoiTEZc2X1vhfnIfHfiK9LktDgcCEezyTL+pNyhbh1aioW
coepYaVm5NiCpJ4EJ6jiglezoOS2SajlnSTQvS0/q14mJ3c0GgNN9KgcoIUoObl7
KjpP8zFJVnXF8v6GtXidrYBDbp0uubf4CvfGp9evzwglsk4jRAMjmpiLZoHdOLzW
Ae4x0loH+JOalpsYK3rltuAg0B30mt8NUtfq8tyJgrolPh0nbnHNnYypSfZcqTiU
RSaOVp2dW9Csmi1rjNQe+EgkG+4ypDD6Wd9Ot3BfHwQMq58gWHtac3MgXf2ho8OA
15ZFr6CIBCKUtPDNpsStHFDfOpJfDKOnTjBEhYVJsJKQj83weoAgmNs3efULA2QF
NBooDsfOPLGgs4Cd7a89RW3F9SbKr1T6ND8NdDvAniI4lWp+puQbl4cIRp7PcSGV
icE8Fe+/BEGvcT90vfr2oLEpVeUkIiXSkDUxEA8lCBwcC8zK/ELy5X8UwqHeEHH0
D6x0HlFV3uvEHu29qMlm1O1R8jWIj/LKj262kJ4t75k+3HSzJJ1e7hfFoYR+29VX
xbnMcgt3Ce7JqmQ7hyxOV9Eq+HxqzBS+8Q6Sx7JZk5eMtQuWRhGpJJ3qQdmDDtly
O+VBn1TyT3mlUF3fV8NYAoRG/a6yMpxfcrobWTa1uDV18n2LsmjcAgq+U/AEwfVD
X/HVE35fW9pM0noGzEcu4g==
`protect END_PROTECTED
