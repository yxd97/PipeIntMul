`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqdstohZG3AFzT9dOSJSJjNSyRCKtBuL2lnnpm4oQVgnZuPPlQjUYXOle50QOYSQ
hB5XT2ZeFWsnKm9RZMVoA3PTk+6gGNYLZjhExJ+hW3xGSPkC66LGCDJnxJGaH41m
ZItsFP2QuW6yexc00VTOBCqv6OeHYipSTcOwgrhLSu/dzZfKOx66PEnxRQllnZOA
NL0AjsidVwdvj83VLf/CDtBOZCFUk/GCqeipTclvdGgHpkwolS2ZDlWp4Zh4tskD
eydsbVlxvzqS4QS8n4Bd5GgK42v3BVq+pfmFtXB1/b9cw0xl9RQTV3PeE+mJ3H8b
DfnaiQeMFYqyqhYv/DbtmQ==
`protect END_PROTECTED
