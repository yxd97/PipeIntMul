`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JU8MMglPVCLxIeVx/V7wBIRQxxhSV83bNehcqzecvgPunqz5z3YSwcfIp8g66FN
e/gYz9INZ+1mVP70QJr5Z7WpSflmdxRge+qAE4kf68Md9IdHrkfk+Joyv6lf4pYP
H7vLsCfBmXxljjx4VvFyyeLC/OTAcUgG+DfuyzBONV6L78gYtxbWSNX4DWuXQd7J
NBmOQfLZJvOQVvGntord6pNFQRO5FClMUe41FOCQLt+11qBgiT0hIfF/I8Uu6W5T
GVCC+61RJCEULzUp/9UEpYQuifxIAHQ9JzBBB7MvoF16a1mgLG6ZsRs9HAmzIVnd
Kf6X2RBO9bcdZJpQk+uoshGOMnkvt/pp/F5pOljlQEl0l3JwJVjezbFKVzmKWu4R
eOMxsyOsNjyd1wBEjChiAUT/gRS9i6QSrTQ1UX+WxZDGuZQh6Sh+DolVy2Ixn4H2
`protect END_PROTECTED
