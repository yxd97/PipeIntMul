`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6ktyFBt5sCnLadapDxSS/GVCkur8b5DVuBr6+0nzx8d3Gt2KSy5gRx8M5hh4MLu
5kirSBPAhvEtS6imEz8eHVXd2ZOvSoXPLyq8rK0ot3MwR4tDNrkDL7Yx5rpCpTMu
1Wergmbn/btqrmmeyzM26XmKDXg8QpTHxUzTsYZFfTwkmzijtmluDUPyE4ssyGir
BeLd9sAnoly8wbMaFhLSbJjnCrEvgDlHvw1s9TLRSNgol5A7lE4gbaGSCJU7Sf6z
MOVW7EicCPZukCHokNBdfscemyuQX/gk4O72x+NwfCze5n8EUQmmEfJUG0/sv0xZ
xomugE7QURLsJsFypH19DA==
`protect END_PROTECTED
