`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hDpzJ9UEvX1YN5HjKIo2HxZDJJ5FtkprlVIkHi7DW4POMvtMYhAA5OO+d2LUimsi
du1N5tB6z6l6mOdllu25ibo/wc9WHg1q6qQbptJp2EpYhHhZscVvyde7beAUxjfd
Bnl6lW6P3VznNHeh0I3x9cIfQt0zUHHyBjppxfqLCRRh4mOFIMnXWoWHu/jGZQcI
753Ay0FNTxAWfTi2rmWbi5JqCsbAh3W39KtTSXR4Jlu2aniaBY3HCx+yHg6d3s+7
neOPcH0/08NIXGpC2y7XGhRkge6ZMxAgXtmyDLjH8ycsTAQypI8+SNNoY93Pw7Zm
76qkt+LTsinuxa7wlvGpJg==
`protect END_PROTECTED
