`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEdLceu3OL99qnsiDFbKIAfR7gJHWHDQrzeYSABsNarGYoGGp0yiTq7sx7XmahPL
4q9DQgNYKQrthOxC8pZWMsNGbTZmOUjU/BDWtwG9ika7Wejr71GNOhP87Y+HqymT
C+m5mkjTZBzH7lRNXkf1OcfHs/1nwNFL05m6IwSKObcTA+KTiQuvPfZ3oDDEcg92
XW3xQNJJKdkenved0+UDC7au5X+209ceK2WugIOuV2ceBgqfPjYL0pV2SnBtDa8J
WnaT3lm7xezpNH5LD/IHdCQeBDjAqKlO24TAKRuduO9WXXywr5RMn10SVjX3Uu/J
ctuau3MgKdaTMD4JvaZL8BwGoouJ+uUPzwzqjAzSiGjxrL4if3Le6giUBXEKQ92C
nxi0iDy/KHnUv5vPzivBRHDUVvwh4JzefqIRS8oYgYGOgDZX4XjrdpaOnZc870aw
9BsTs1WEz+ePhJV4E5bes1xA1Kjq4I0+AOtXpKTPqKcJ/t32AP3Amrv/gRdFyGnf
ic0c5tov6Jo466I6mzQo88qzCxLH5AYoMXt535eM+9WzHzz0P6JUR3oGJAxaGYIU
NiM0xnnI97TFUxLBq53z6yr/HGpDc3JzRmxClGP6hAyY7tOI6tl78KX+nLSwWMIL
oRw1srh1FrYFuFdtm+V2IpFMw8uIf4XCRVxcwBgV1mvYGxR5R1nMP0FGOQdUQrRx
jP2VVQToOieHPwcHbBKXouBGCQSwTlO9l+t8Z5ev2qUn84U0gWOu9xxHuw9pnryd
yuTwhh9wSl/kABDCECTYMvcDDKQ+td+E19dfe2AYXuXWkrLMHzHA2IEn0Dn4CKjy
Wi1ohpMDEJRvzvlGLm/etTGXQJjnK03KGJM6Um1HaFtSOgJ88rXx0oTEzJi/PkY6
RBIo6ovA03o6U0Wojez/tpLp4N6vpfvH1d7sxCt+kaPF2F64mxV9MEqNWDW+s1b/
LPz7SgOloOWEmeTve5ZjN/dYkcqmFXpLDEJywFu6emzdJHMdt4MAStlOPhNForAk
LKPcGZnEsvnMgwnkUbU6a5dcrJ/3YXBgVXtgwLuv4IPT3SWtx/7oxwpLgaR0n4fd
3GNBLi5AWCBe9V0tmOTFqfu6/908iqmkYNyRDJE+VjnXiDOFMrBXhgz10I5VhvUz
2XGJCrKp/pdUG7xvYq5RH0WhQS//5WkadlaKMJ0tbMgJJoVCbdoiiHEekv7klTc4
+iz6nxpaODQT/x+k+SOGU4F+LnTupYsE23sZ266elJCuXr3n/KdCZd/j+YrgE7ef
k1h5x1DuQXNscQkqLrBqYJZcQFzqC8fNJ39b7ZbhFX/T5VITKGTLmqmR5GuQJw7j
FFlL6iciCzEiAewRO0IEB+GeO5WuZy9XDSIe810bDFtpCsuSsk6E2bCEiDhpS2YI
qkC85ZqKTGJuvuAww26V2P/zElixZiYh/ELqQFw0zemnDS+P4RZYOXTe3SDxaorp
yfUn6LifO4Nb9HAmQA2RUn6QGpwmuue/JHlCp0Gg7zoNRl+qC21/Ukw/BYVIBtVn
H9wauCQtlOn3ieaJKOcdXQSFLIEugzBA4eBOEvobKiNePfvQRq5FlZv7vL+4EHLB
BDz96I6QqWqifVBe3Pty+kGmnltZ9FJcezX+la5BwnE5XuEhgsd3IAXsAQ5OWeDP
xqaUD/7LEoximJbjAbPS3kLiAQ6V+vnvzm+rxeBzeG+BGhl74qFP8oyCqWc27XZT
gwLXn9Q+TvYE0SGl0FGi88acSUSGX1PA6stDZZkS5aWAoJwaWNdBKpo8fgeijBAC
Mbf1MAxM/NyVHRcjH0B2s4fmxsuKetOxezIo8DT+01S8+0Mg0K/awjqsJ3wW5X3n
2TJGXtXYNfvZnUtusIX0/xjFdxG78mjTEpemA6qCvxGX4/MTBrjdND2rxD8zYZ1+
2aRJYbRYF2PHixD+PdF7qrTgdaDTivqwlHxx9XnUbjVmEeNdSMeA/KYewNClE0lZ
msu4gozrrwiwR7jwN68MtCGWwjPCB04N+qOkcNKKnpMW3tiO6xGAWXQPBQw6qH9E
i0pa59USlXnUX2DrsddXbhZXVyGOluK93KlwaclhO01KEJYdlPkufljGBwvwMXO+
KTWFyseXmRXBgCM7qDdfKyPwMY7aI46XyaVHAWzaZp+2gGeAQ7WOjr7HjFGG4adF
QtOdHmc3h1JZFiLigP2fJ/WyWbvQl3Ob4GAthiR2a34dw5dIXoOzRfvhfzd5jSro
Vj1FvF5fzTkKD6/AEY2249lEtipsnDa1xuSEnFUZh0bUEaX3nnnZAHyXZB3n8I1d
FxkR9e5WksptBIzMGLO4Z5KjGjamTRmZ2LlYzRCSXTgMOxktxtrXxkURoCMePjUd
wN3i6Zb2PmyajB6PM+8pzMhULVM9uZPeT53+OvO1fLidAgq4t640SKoe+Ugh3YwO
kLbROu/YKufTYQfd8tYQP36Qw5zv4QHDDxMEGTjv1HdcVB8r65Cf0vJ2ne5RELyp
JsHI+RLs8AQnT6tSjS77IsISDOks7WPxyk1Hqltm5X+7i2npedrLuF+VdoPQOREb
NUI2EIZuUxB7r3hOkG5zhcWUWt7g+F1J/i52+IqyvY1ecfdabkZ8r35YTollnyjK
BKR7LR1IXS7J0YlqChLIE7HdqLXIj4yE39J83OrUpRD9i2v+yVZq3dmRXut1LzSR
ddokgJ/fj9ax9CY24XKa82RnJo35ZdVQpe9/GYkmHER+ggVBpJ/i2U6dea42qfDj
oohUezIgM6rU3/X4BnymbhQURwhbiWBMQOZAS1xMYWs2vLRbTnlhoqP8ipzUyq+T
n5Q/HS8tICgWho9Q0sfDBTvv6S6s+Xrk/g6CpLIUObSGa1mYJjWBUfcTzfdQCmgK
gfg2rrvEeFP+plvsRlzHt0TbVDYTo8IqxjNvmH2O0hxb3XP8TI8tzuIH0ojtZRCl
ArJ4E+tG/xHAqneaoTpjEaNb3SGErKbTi2AY/Ko+H9nCLBqJbMhYmYxVnzZJtp1S
8VLrfYiPMswjKP7SGurXU6MIMJ5lbznF9JBDdjgbcfSPAr4TI66aBJJvGhEqpcE8
QfU/Q6JKwd78vLu9HBKGZTjpab4wi0YNjxCMN1uqqlwMnJhoSmu0byhJ7Sc7cp/i
Kc9zxvT24Ql5JZeOpVsx3vKQc9RwmsF5hQkHX2+zRyMwqybDvo47VzEFqCOwxZ9X
kZkv6rjUKWk0AK0Py6U6n50tIk2VdotROu2ftPvAkZTbT2wHp50hmIq4GkUzJ4YA
DvTb9Xz6EfdKQVGfcfbzOPIHfndk56+ntBHgOZ4gLDETX1gVa76xFDjmOWIKA/OP
lD/WfnyLrB9TTUj7hX8f4QtDjy3Scb0QBbLTEygndVuOQKQDOxESausCgsDYHM2C
ZQQSTtx8cIRxWKoh812wmeruF11wNWWo/H5QVYG0jjzzi/4VW7qhqeU2uPtFsMf4
AzRvLmLxjct8HsO9DhkFGqM4Gpt1MuAxKTn4dq7E7uiM/XTxoTRdGhC3BWEdgZv9
z9wxrLgcMrDIiQmRS3oSSSPzyHSpCfFCrHDC0nqZHyzxh8w4F0GN5lV1q/V42ewh
j8TXesMV8e5VK98V69GAGavubpiOC0MMuPf4ybdVxW2z6PSjyF1ZQvENbn/0SJT2
XtRvflBZi3u1AjfztMFBl9EqNHG03FsWRyGoa21tTws8VRx4MEXZD5F6OPs8KlGV
T4BxinFj4sjtmrpWCxL0/KngSTyxzmnV81iK0GZA0LwkJNce71IyQfrynr17E0TO
oHlhchyXJc9vNIXND7vcF1z/CQ4Ro8ThXOmw8L/kdH7PdHvkz9JJ8wE38cA8eZiS
HsMF5EWfmIjxx1i3FlPgC5iA/dCpMEejkh0shvW1iA9N4obRmmyrx58MeAysMh6l
xRditrdul9BJSNkcJVoaqaejfsCs2X2lFD7CW10TARuMIRhJB+/ozPEv4cQH4m6d
RX2JXqdmA16uZz2m28XPKMauo4CyxOpeyxvdmLHhMnvcevpe6tWvCm1hfzcjnKEv
wncddl13sB7dst7s3Ju25STGCX/zBbghQSPiYNoIanYxao9Cf5yd2yxVo3RDmFiM
Jwe20Ji+SuvRTJs2QVW6GlKnmgcA7Oa0WI5p2TL5WkXNjhntz3EQF4zsCxKLqAlj
lOvvJaTebe+Zs+Do+veo4T9Floc4nmg/A7H1jNlizJJeGj1gyJJOGzl2tUO4PqL7
GfUKr7FXSUvccNo0hpdAgF9i5DggUPXyTqfDt3LO+NPVxzdQACcivQE5AG19RBf1
EwEMO1qIvgrp7TokvGNvHmJog92NcITdqYRKHzJcN0TIMtfrCAPsflyHWRmtorLJ
15Gh8Wl6MBuAFalesftdLL4o4KwkaBI+RwJyvbRjm9WNb2/TxclcHXt5/puvkEF4
WGdtVxqJTHYgHyB/PIB/x0MkmLpH6MGZpJWWL1iiVIdpZ84AitAI8oJdCnVwQQoI
y0ISPoEoo91Rq9fv6PUwqN1/tg3snzMYnnEBvS5yO5PocqcnXHBa1kcR0Em6W508
yZ/EBT1UP6dNLQjJyffy1dKA0Yxn7U//BsMgUH1JPIJd9Y+DpvDimgSIXOAjpEun
8gNzB17Ui22mV8QnKt8SgV+Z4KMTAu0XdZMnLzHye3kNJRX/uQrSRt14A9qnC9Zl
3OpXkK/3FlOysv/90xVJDUQZwybSl4zGC5GZ6b+9o18zB+gh/NgxGJaq+MUr+o+k
tRyCVGkXHbqcswPd0uW+IsqavzEBAhxeV4ghUGLQZs0hR1YGb5svSPxRuFFXqASN
syxkQMc9lBM6CcoIVX6mh671ZkJccTCsMJUhNZOvGbK6P0xp/S/hXPht1WavrSST
wZSu6pUWe2SDMBYrFymjMUlyvITCRbMdXiv1IDik2dBQGowacYh02usz4GFe1lFD
f+QV8h5Q3B/7pohBeUXuyDZGKTKZ1PJQcO+USgz9az3HeP5jLXPnBvgn6sEKYaaA
Qz1gKMR/lSEyntbOrnHjdnfarMBpyUvANHEZv2sWDn6eyeNmc9shQRUOOx/eYCbT
sa1wfjjaJtQGLt56L0nllTtw6qvocrq2JJ2nqkx9yiqG8tNDcSXq/dK3hCql1lUH
Wk8mjRQ1occ5/5OyDbTu2xrOL4vf0D5Wxv2BOXKEsPv00WDcEcNwCP4zHoYNQKmr
iP1svQr4mo0CaCfNrvIzP1+V+rL9X7AHL/BZanH2khysfmIgK052PtXBbWSnWjKy
tBzXttBfYFs6yvX3MyvJJFgzuyUMNTXwKRcTMz7IguLhDX/0X7P0jmN6X6RbQaGM
sTYEbL0FVxBA5hNAtuESwdAcsv0cmF8oQRgXWS+XNgdwIl98wXuqHycWRhdaCMzM
qd9tOLlXZbQM70S4FavEBys8fWk4EsxK0UiVTIFHexeG3WYwojzDU6o4Q7K/XyoS
u1L3CXdwrAnxRp0hhLnZjRJQsrMYbBRT+ouXaX/jO5mdD8HsVF/5M1yD4Bwdg3Gi
pdLDTJqFtFCQn0HJEb9ufKabAnARE/a8DP+1Y+fLwPJlzWhJz9MQaEqgqMe6PAu4
cob/PFw3wSgSTTwHFPHJkDGPZRI4cyWyw4AnOlzEv0EhJNVHiVnRSD0p0AOYrcvI
jh1DZlTdu99kgVtwwe6qkre/adycnsaNbvuAC4wQQRCwL9/WOhfeJZdgXKT0d62f
K3IAwuhFqKxV7g+FAZYmNSI1JvuvgYWsNs0HQFuXGQ8yEX1xU5nWo4d4M6Rhl3rR
VY+wA014DO++3qS9DANgdbiCLjU0VoEH3ffCQ31w7kJ3On0Rujqf0qb118id3184
USRrv1wSOZQE9uCIwbIWTUf5J1AI/n1F0YhyjBWGKI5sGfO3zDUaKsI/GO7fwwEW
QShGV5Aj83fV3Xhi4Ek+zYWuXQ2DMfpvZmvmPbSou2IqInIzdtAQ/bcjjaARNvyT
7fhLoFwhf93nZhZSKP/VSVL/0ZtZOWEEZqazrbLjk+0tuLgXm0FGueHGp5OaUOqQ
kkUI1qDVmSJWw/qML/qnUDFJrz8bM356f5i7QRSW1j9bU7vLFVg8UWpLit1rbciC
9VElTvoiHL7KYpsbqpyzRlbaqw86fm20D9Z5PrieVRMqVOMwt8QDMI84cpRSrQcz
Jw1AJwHsuGFxgT9KCPxyJ7mtHcKEo6H/BU1z1iR0PfF+X4vQIVwVboREeXAnjMgS
03ODUGN3ckzDA3IyvOZIphSsG921Tv5+v5nxjIiJlJ5yyey31q26SD27PCUpn2PX
6zrVjJe1KSKwPF6seD489OJPhGv1pi5bcjPzUpMRgpzl1B0j64brLTaYSXdvhdn+
1pfpmKH5BbAChMUE0RZcuDF0V9JcMOTldc1VlCGHGyC3SPbZjHWFLCngf8bsjIm2
eOFApnVxQzj6iXUvtfBUrkHeIPiBsG8Gg0AcG/LAEUWxw7/ctnraBhbO4BD+ej7T
C7nKDwz8WdoGJUAlvAXCmw==
`protect END_PROTECTED
