`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0b08gRmuR7Uv2+5VX5OmlJYMQmPvhM/uHu0Q+itRsAYw2eZ/I17nYsmZGTqbkji8
EcJ5Y+tYQyTMOeMSMSqt6f+beXay9HcceuP+2shf0Rk3sg9hmmOSCbB9i04ehQDW
4qRiWrzh45AjEN5Al1k7pQ16TIw+tysT9H2ULqKPgSlZ1AMW3lZyzeRSNsIWRIRQ
6M3cUd06raj4jnOyV2CcPs6sUBi2wN7cDhd37DeVYCliBdnPLrJuAAvksdVDRJ1u
AlPE2ZUTNdDk9WPONMG2KrqpcsfkyS5M6pus87rb2MNlfHBtfGMkr2DEj0Mbix2I
WJ+2oQxkosLK9gTqMsE+tzr/Fui+fmAe0O4o1BNjIiR/K1ImaR2rzMXnn6DbhJ2p
8u0DDTsUGmnbowZVcX5Lug==
`protect END_PROTECTED
