`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3JBaOfpTvdLj/FbQAaqBpfhb3BFiu8IQgkR6tf1Bja+JojqgJKfsPRBvgfP2k5t
4aQYN8QwDO/QcnUkK1NH33rvlstqogwmEeleIxs/+DSYPhPB9S4vgGILO0a29d5+
j0KeeV1tBUFrJ0pIffO33PvODQwPFTZ7nVoxos4OPJZroHUhRw3un8/IRnowrw2z
JbvcrJ2yi3FXKizlAKC4ZBlJfhd/WjJck+6NSSdYc7+bXbo9/UCuTafIOenNg6/i
llaZNBVbWb6wA/gnhoaW+p4hz5Xb4XIwx8uuG6AoC7LxoidubBMDpvqLUhrOlZMs
zs56LyHirhUXq1+oEGNCiA82/YFOLgy25AEwcxcUoccL5+MHsPyRLEnA9LxeYRLk
rJnzLzTlSyzuJgwsZmZD6HwY/Y7DColPiZQUk826gXyRfad1ZWO1hu1es4q903eP
oZPNtfqZ+vppFSEegJRJ4OiGuTiWrbu6qhcoUfNHtULjZ0EJLD06PQeS2fQ2njnD
4sCF1+Egf6VNZl1HJsCKACJ9KwdV8e3BIgzOaBIq5m5nzZAqE8zJOPlHwPnBAOab
sJdX/ujKHZcWUSliRQxYWk5gM5DifUya6UwloKVetjtuhwr5XCQ+3PTTWBNiwvHT
yhdwpkI9cvZ37iVsJQij96aVY3ZXABcY53XwXpBkunmAlmiFQf/4NGbd+Q8TJIMk
x2QwtezwUw4jWvNQmdseJzqePKzcbHEdiMBIW5mosXw1VPXEe97J99sElNCYiuNQ
AlTqV3UJOXaLDPPbqjdufdmoaU7lsKHldtUJ6uIJFprPA5h3VipS6QFWlpRjfD0m
tFSMxAZ1sWgBLao45h2jinE44Yjl1lo0JY4+yX+Ogn7rtPUHM9rCyT4JmyiGlIAm
yLQDxFX3obe2BlQ/y5a3loC+P9IhU/nSl/6NHTM1elWUETZ0sfySUYR7YHnzrk1A
ZJ/JhlLSRDb8JyRUf/7n4/1PB1xlHhVjRO3crpfbC3Ka56wC3RqmzaeUz/bpQWaF
YGRvd3D2TTJFRqWSLrw4BA/pwQcJFSoctH4JBPi1/TEz3wMrOITNlv7qGbxwjiOo
PtlIEZ/x7PdWoBvEVvy5maevLLYMS4Fg+rCVNPU94i7i1c4c4KmPJBbMINXWgspR
eCOyxTbp0YgEoGqF0I2Y0ad8rk2Bmf7W4lxp0SLicXtoMWPuid9Pa2cojw7eWkY2
EL0zZzjUtDCpQ3uCJIOZl2pU1GHD+o6W67zMFdTsMmq1HBKhzo+3EK1y1/eIYK11
4Nxqj1JLeShbl9GxWNWPKXwlMX2xjMbWkrC61iijdM4Ko7+uFCqRLY1hVp3AByih
QwuLDJGCvl0zERHI394YF7WJioySXz/6wa4M4A4nejKMnNVmcESZNaup4t4SrG6Y
dvE32AlJjskRawPS3NAH8t5b72UrQi5kMnfRHvhZma4y+PQjNMd/1lEmtFuSr3KG
IFBnpGmSX8RXJp4wRHgiBfMFWtfKqojEvPGiVR5+kPVERqgchq+1JdfFzK4PkPMw
lQaPAFocRstchRUFJScJic35FxAypiE7tl4/vruouAISIFBNCwvS5v8nxYPwXH7q
ztFiRQOWYjsKi2qD7WgfzY0WC/OIFhKPgHf2XMklW9q7DCv/SD84gVtcaTjezqbH
tRk7mtA+HW9qqot/4gFgguTGANuQh64bTakE7nayIBotVJY6YhwOyn/WcGbOFlSt
BNvKFGMFS8jR/s3xmXlR6fMvjQr7YNoqc8hctEPFeeBA6ysIUYndYh+9QeYLyrdu
rybt5RQ9mv9HZSGIhnjHddtqpVdulNNvB/IOIjD1OdXEDynNaWDKNr8saieGT+eF
`protect END_PROTECTED
