`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mblkj+P4HUO1T8FRefpprFONU5Ks6jQgfDt5+FC5WLzutifqYVPqVVBva3bwDP6
wbI/ysSihVhJxQhLHoGDCTcpxenWOhTFeFF260chtIdDVIS5fK/6jnRHLnmV2JOJ
gHQy55+Dt9wqHd9aoSGRJxJgX5NcKuxkcGI6wpRjcGUaFFhUOf3/nutrGwokmLni
s7n6qj0EZAC/7/9GuDn71EovM6MFjCJI+lPUwmnf8+yVsBm7YLp0neQ5IzcTlkqC
vYyxjWCVST/KLj0VLVsol3XkADKeZhV14D+m0+R16AD7H7xhu1IoVumnaY8y76da
/Gy3EEd3x3w0okLmy6hsz2tTUqfopHBOrFJn7DvCsRCXR1R77VYkBUmIFFNYNxFI
t3XumsFhuONASpKNi3Pkx4mOnVt1e3JG/rHVNGumhjOwEdiV/XhXHWO/cAnyUl4P
GKwtgXnooMUNC/nXOjm7+xGqyp1adaEydyBxsEMEhKb5DuHV4JGvGDc2gCJ6CTjk
WcfPXi9qhqbObXm8XsAmVIfgEnKB7xfrO65jh822qN1PKFoYW+IXHH143RxZEe0l
Hv2jr8IR0DI8mlmzTps358RiDjz17OC3x5awFgfHFwmCyypZsBjMODm9FudjJywE
`protect END_PROTECTED
