`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StBoM23qUEV0rXQ2Zzd/XavTZELLAFeROy2pmcZF4fYFStlunBWp6pvP2LPosMuu
p4iMlle0C0p6KPLlvtkHse64jY9ZDiab6KwBU2r8taPnYNkNTrcSfUj9dBNigcjx
uy71hN7nNAlp/tmmWH344wbPSNP5WYskmKhSLs0f3512+STV0rG/x2qjEmPI0bgD
b0uh8+2GX2ThG0OOwkokEOfAYwEp+krO+KvAfFaSqmcVDH0THauXwgjPoB6UhLU5
3rcjzwtGelahl4jkHaYQm3bKeNgPEdbwucgMJH9VDClAi4lB5klJiifn3akTuHzQ
J2iEMyA6s5yJklQ3GLTDSxQT55VNsgUDEc8x75VfDGQAjCJlISnWFnhFkksoE2KT
E5Q1W/zBBSCooRlwvCmwOZgtPeqswkBKgBAdL+aRLxeHAjeLmt/g1DW7SA8iK9Qr
hA2dWelEP56hEYxQZJpnpGNWJa6MG3Rv+bQBnUfh0P63nB83uvNbjZtGdQfD8zF/
Bsl3npbCXPCRevmNzhOfAAnWWHsqe/GU5QXAfbY6UW6xzzgru/0pMH49ju2tP4sO
Xf2oBeqCogeFdigPPerXL1iOHONtEGSE7cohfRstO37e0XwsIDCbB/64WzbZr8yU
26PjyTl8dmhksFkI2DL20vEK428jEwHKvwlHgmPqBfU=
`protect END_PROTECTED
