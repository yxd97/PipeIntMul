`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DNqAlHhQLaKa2bEwn1NPQYxJZ/Rr4WNYiIaN2XWpZ7qyUi0hiT51rrlKfACWI+3A
zhBnUjND1zhnk9F449b3P2N9O7wTEpLTG8adaLBT1+kLdAqI7pNfxUr+SZugc2FW
F5CWqaD3S3qAS8jCBv9ZXiL3BDLGtaSdwuSoY3Yu8wdccgJU1Hc4bJIvsxBPeuVv
MRiGt2dcKwVbylUwzEHZRPQCYYAZmaVrb4xaDvAvXvuRN28UoZCuOPiAcUdXghkX
80CdA1z5pVcLb1Z3/v62UwV2pjTch63xxzawAeBvpniFT/2f5QemekKMAaJQluiU
vcQG+pTNUOuEEZLnAOntWjeGlZouUFszItTqVhCgsQ2wvDXLeldMEeV89XcniEGg
`protect END_PROTECTED
