`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16Fu70XopOpANL9kDJ2pk46cRzDEWiqSPYRme21OyApUzUHWS9v7xUUXOBZW1rbT
OC2bm+sUUT8etHrbM5QyEqNEcKfqm6WRl91+jiEZ2TMDe+41Adhq7eNyMGHNDDZN
pdhHAtg6ZkM0lP4vBwemQTBGBg3574pTclyQghP07iP83Tx8bj73LIoSiF6zOPjp
I5Bl3wl2bucdhNs1VoCgXc/xl2sm8qtXc4DBwuExYn8/hWkYLp7gcNGc1oBBrQOw
NvFhC5AdibIxGY6WDILZ6PIF4Fan4c4R7b+K2dl6OHmpsYmUHpRUUlXu21ouKt0g
kWiGgOO9IUiqI891lWKjpMJDbt7wiXAAnMUtjt8DOfBAT3GdO6YPinQO38Fvyvvi
WnJpXRq91uQV7f7o/8LE/ZFuI+7M8q2znRocV/ykrcOlWKgRZ3ahnTYywvjPKH57
WORfAXpFixNnz2WFIJNu0GKg/5OJuADhAc2jgkb66smuT6aa7d5Uo3qOruRqViOQ
jKGV9+IJT0TolgVkCcl+MTXKyVLWtPW0Dr5mlZC31SB4yWLXRPS8jj1rNBfSL7+8
n+9RfSzjp4oIuka3lU82hj02+jOkBhPRysIFnlGNn1VtXEiAV6+FZmgKLRC8ZOqb
12a658SZAfIEs5MUBqldvsXWz8bFA8NRHt9jTbsiLoEAYn6TTot0rq5+tGMOO/RH
hSvRMqZasPSYqICG99Lq6+QDnxH5eW6B2JETmvpP7xN4TrGmZdkhxbmgMGDoA38z
HZkkc05MckFfQTK+HmfA44XeRNG7LKRUo7XKf0txYni76KZbFdClU2j1pukNejE6
pz07sfgmDAPVINEETvEKhF6CW/mkEEvEu3pVPSXWNXDnjZWvoK7NxzRKpwACMIn9
rOVRWsA0whjGU8PS1psEb9ibvkrzPavub10dxDs3uGrDZ1kE/K26ch9/LyDd0xfO
fEjE3RzHyQIK0hxuV/XqEbc3DsHUOYtbhF8u4EvjCWCcGwVVkGu362gHrB09rFtb
w+pXZ+16hhuz/J/CcYQUe73QwC6kiJJkIPaZyuCrcSjut5tzZ0rczeBScWGY9veT
4NTgdV5yfMVwuIQ6Bitdw6pAtbVxN8mwVzsN07+Vdewo5b7Fy6A8w6VmU88uA5tn
VGTicI53iDnw3/TbGucP6LCY6HwZUuVNowU/PPV6F8/BaviRucKLFsv78yhMbidv
Ej123LhJFun0UjjLvc/jOa44tQh8D5XQTkX0XfhyErp22HeeSZlbwA7TAwYaKUzI
KpNh1SafsxozWvFYNzcLjPB9xwRAeR6OGCmvpv7a8DPUR+YXWv6/K9PRffrdDWN0
TUbAz2NiRdQaN2Q5LlzwxiceAdNTI4sPYLg+Wk8pd5lRbb0FhE60F00ncGAtkBfU
RzhghAU7vcVprjMw/yNu5bLAP5jPkgK6l/TZs7kH7YfQucxgLCGr0R29KEiRzQT8
9GgGvTor5o2jiL5hvT3Lo/OXb7Ve76UxVIaORQ5236mNVrCX62BPeSP1tIjaA2DI
2Un9joFyZ/KUgSLJCWl424arc6K470ia+k2vc8HeudZLWYj7BGNg/NPNTaxU9Vxz
YEMNi++xj9H2j2kjDRx6YchDC5eWlR/BLZGs47TgGKm+AwRtTXHdpK/A5ehu8MdQ
Y28X59iGJO1wO+TsLzAQq40JmDJU0vOSE4pYKriJhEkd7MqVLvT7voF1Rla2nsmA
UyY0BpGV346r1KgZ+D3AVjoOD5+1a5ABb9BD82qeGrON6+e79hf+hKztkR+jRVOu
dSSoYfIrGjiEOAaIR6pE9BUroITptXkeDhOUjaKNMiNI3NQRNH/MvxQYOG6ODAn7
X3YRRXuOFq1AK1k1pZvD0F+tiw2BIfY5BIMsSu6DYUYCmAHpwCbonRxD1m1KrGes
s3IR67k+qzAaCuk0zG4cnBa/140q+HHGgAsT0zo0VWOMAKADGa6JRS2PdYFGwc1g
94mWPBL2Pt55uA+UQiMOfKYk4Tx0XFHrXtFxhVMgyheeiq1yk+HX38nR7OQASKHU
FaPnrz2S5RzldOyfNFX9FGyVYTZROPsVY5QhsHSacpWfCm9dlJ+dbp1pgDMUZkQq
RBC+RQJtx7SOD7IyH/b6omb4gWODK0g/6wMXqVD9iwkdKePm56IwYgwctqJbI/DI
PWNEErtISvB44dWLm8nmcCyeI0dxBM1FYSVnjiFh/kK0ks0yNM2pP8KppVmeMF7L
IcK4y2+5SIXkgBGTab+m8jTK/tOLVGu8WO1fHFgm/VRr6JzKVOtblYk34lNDga0z
cKPcvIpE4kl4W1lT67dx8NJRloLV4ldA99MjICYCjwJNhQwliSFk7HDo/m9QXlMq
yZ6BZqgIDuQ7Jx9N7WuuSQh6y7j6aHuWeVH5T8KGtR6rckdD+woMOoIle/ZZ/QoP
XLXATW2XPJri6haixc1s3Ldwfj1r1G3PakO4UXrRNYydPkS4sa0UiG4975Mx0jMV
C6/93kq0r2xRUXWxvVQzyFivWu/Uhy4p9mizj02FTxH6ZXpuO5hgyELv9tPDfPYo
Fpg7iFi1wLcz8ly963oV2kUPuJolM8FG9zmreLH+BUDMBF29W6t5sOVuwGmDnkQQ
OPNufIyxeBw+4JBwBv1ca2n7Piih4EN3m8jaesSoK9ReaASZfLfPTGTdko3wPkb7
WbTKM7oOeENfkjUsT8pxQM7V2fdAcSzV9Bx3xQ4/YfvleUYh6gwr9CiZNXR4tpPg
UyHE2YJZofcTb/Ct10lsmyEB/1kCEm0I1gDEY9/JSh+BleiCA/V3MUx3pSj/fURw
myAwdUZWHk/WKFOa0xJPSQjlyJC7Bfzlg+6eP4zwMgOGovRVH7MF8z2b3h5KFITg
2xSwjBcP2LV6d9O1o/MOSozEB5E+C2pqIiZE2dVMpVhoqSdfRvWFoV0Ye2nyDqAy
OEVkDe0hSpBvwGatC5W8ZvhqFQAtYABNUj0tu2pyxL/mSb5NsC+tLdNCbyOb5+5G
K+Ymn3tY3+exPRn/gLmWnCftFFI7SNrtw3f0BFkd0O2J9lTcgfJFFtqeTKVlF/Ig
eycdcOi0PvPG+WnviuDHD4fxmPFo6vBAFga/5ZqGwKebUMpE6A9lPw0az+73lEAO
1Sdah9J/+o53pbnqbSwPXAe9o5bPddXdsjcTsYwj/6opC4ORdurL13qjNiEjVc3I
84Vrxlb6bTbqcXqrOiism3SdAPUcSkqqEfmt7sCMtbJyuEVkCgSQA2AYtephSKfF
`protect END_PROTECTED
