`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K42iiwtKHN8Dyrv9BmdYJr3uyKQbwjORDfQUZmyQUycimKpcIT4LrWBc7aUfGE+Z
FLORiKAVyi9KfaGT+xSiOd9LnY5OwageRmateH4pfPATD9r4Odu0nN4nBJeP8F7w
MHN57kxopljt1DJgb0MDtWNtTY9nhO7/9b3vKsDLMjouEGXab/OfdxP4zqvR/g8V
QFrT+NU1MigkKNLCtjjxI42GwmZDJZCvmDUKQZvdXQxaAnyDoBh3v6aArX0xm3Nu
DhcuES1ZIiqlSWJlk67mwkH4ywMgl0j6bAcXY323utbiH6u8rP6kL/Y2j8hdUwNv
FU3oDe5xnbl/+rjd5tHp1LFmjwY8+3e5cRtPyoXKA+/RjoPZIaJExTBqFrS8Tk8k
h2bTxv3mAPRoylJCV6Ix+taZnqSxoaQf9JPmIJUgtievzWRckqUFcjAZhUJYRP+/
OeEoABKLLNBV3vZGW/IWz3JnvCdIFoqSk8dgSldRyed0gJm/4aVq9kw0wyqJPE2D
J812PIVuplm8HfAbLjxCEX7Z6Xz1HOezbffPKMIYMRe/qBAe/+u7iw5knGQ+3s39
8VFfB4n4GtNSaXx3OLeSkka2hZOrtQXt9D0AvyzmgW7ZdqOwKXOK7h5L/oz46A1X
QDw+ICblGpK5ZEH1UAFOQwZ1bUTKi8ZDNXrAZfvaEvTmKtuw5P3/fZzduiLpW6vp
1MubKjUez2Qy6eM1kLK91tKpXXOKTiFhPbpYj5D0uniMhRhudlppp3XLAgyGvixu
cPBCq0bkb6Ni84hFOAoQu53EjI32feRt55nY6RcWPGrLM606eaJYlVizstpjQTHE
KWJJ4uOzKpUq/10ciadX3M3amssz2VYfm9GsXmkQQztG8eP8MmAVS2WOfY6EwVQh
MpZQZxCuByxT2LOiGPgKr6jHovfW5GC1zpAMJcYjWyk2uFeUIkLStAqeGpsOQLV3
UYwQCh1k/kbqxu2KR03oPORZSZ0dRM4qSQOzFIOO4HQVk8MpANoyXl9rUO9TLnNw
Jd8oX080efVSS8V1M9EIKUsU2anhF0MtAl7VBQxGSsLNM+glGjY3FBn5qmAb0ENW
Nn7XenSoAzRNgX8y5EfHWbpd4nEHK0LSEeoglDI2poBnOe3RYJwBuSVg79FEec66
UAdtcdI1dGxkCu54Y0UrS40ssL9GcNf3Zbh2cVjeb5U5UgqM4LDeYKcmtjqCbLe9
M4rfU0hox+62rT4G8mDkt2Gt9Qcu7G43rxJ6mkL881LviwujnNaZ/Zsskh0QZQmh
z5iJ4jPDHVG2HRFTV5D9PBBKIhsz8lrkZpw4bHw7NDMA9GoYrxVik+kfSSpFV1V5
w77X5r+UUYNBQ0rVpy61nfbrtuFqIaXbI3Q2peM7wL8=
`protect END_PROTECTED
