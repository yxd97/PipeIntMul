`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/RSRUO+b1DWgr26yeeOicog2ihjD5GUE1IZdl3gCDfGptKtzYDIC4+yR9Okaa6/N
lVPDXU7oiRkK/xb5f8UOTto/KkY+/ilf2yxP2qlRd95xF/9O47IEPniEnOO1TPJG
jYW2QFClH1k/Fo+MZ9m7ka4xSEmUTcATFeNZCBN7kaiWBjDj9sgR/8TyiA/Qgo2x
EngHD0QD9aIYdgqtutPJs7R0mBO//Q3D8UWhq1R78/ct/W1VRS0jCl0WMYXXiF2O
WI4mmB4KyhFPfFbwKTi+oVKWp5XlqH7NGNh893a4Ej0=
`protect END_PROTECTED
