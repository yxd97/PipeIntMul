`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vp5EPE8af9LIph9WwlEnKekzFbbk/yybFU1HTew3FWsLmi2NAplcTVCPqbsmhGmq
EjzvktO4k9oDLzwjdr/tW0MT+4oVfp0nE294yebaqd0IM0JGOw6pOOH8hTm7QC7i
AouUb++PIVBR45uRMcoVJec/dA0DzoDRkX3M3CdaF2TYPPN8B/OmfkNpSSsCQ8a0
+syOhEWQ2CxMNQcDYn4IZ4AY0bIYEBELHhoS5//+wjcaFrAGd9hZqvs0q3Y2U1t3
+WnNmrR5pM543hQnZudJFPI2kkbTCMBgS+Rfg9H0uKrFudK4GX363xE8ZyhxAB7W
bu5DlnP3lj55PYTATpJxCCwafOur8Ni+t078LxT3CqNW9W/RNZjdHN7IDjmF8e/H
z6KQyN4dOtYs8KEboffykcSv+ML07FjEGc0DfzZtOdpRP0Mahq9RelVIm6rPKcs9
IzTsRtYUeZrRgta8U0/LR3SpUyP9TlC8HLTGea46mDQ6ZOZEVTKO5jpTLpJgBKwG
kiGAT9akDi8Rr8tDS6TtNqNOmtTppPm2zSFdP6ToYX6vLm8kK/RrGjVQHcfiAXIF
Q26HfqdrzrP5tMQVYBJpaAcxKMTFK5yy9VdLkb5HSaEqo95ryKIWaYRDpkypZrEu
L2beooDmkc+HDMuWLGeH0CwafyrHKiHfxvqgDoCdOnDWby22erpO85jDY1qpe/ws
W659riHz80UsAn4wSbxFewKgWwytIFMIeKjBMUv22M6e8GQq54y5BGf0S2PtqUUC
3H3XC5YBeBvXbL8Unl0loOlNdOwlgSnE4LTGGBagrzXcov7D0qLcU6zRyl5cWntG
`protect END_PROTECTED
