`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hetQpKjIZ420s4Urqt8J6ptMlRh6xzN58mbMg9a85tbYG6c/3bT8ingapZ9FYbJE
WsZC/1efhEZGU9JZnnWUi+8LyO1pnzUUObILu0C/lbIGTZKzg/4ywR5+212EYBTE
l+7vt1zEyeAwq+4hfhzRw0G5DE0TuJIdJYx3r4rDw9JGepcnhSgYQ5k+63tDvNLR
ILSCoYj2AFKulL6tr+emVIT5ni+ZVpbVAg+M5TANCvggmQ8AU5DFCsVaNMhZ3KP5
3LI14IaiNYs19rIb5cFyOI2iX1XfzK4EqCDw8z4BDaox8rCTpyqoXqcqvQdGklbL
FZmDlepTWr9Je+V1O6Rj0VaR4epdWW6Hag/BLJOmafcJew6rWtKQEAoYYWkuhsg7
mprakFvbJT/NEUTyh7+3lN7mnK/ktr5t+sHnIsQ36h5vgbpSmWdyH2SrfVtn0mZn
89/X+V5HHtIIt9ydhPQw9v31uB1FQWT+p2TjvyXD5tWuTCj/VC+/yY1Kj4ZLqUkZ
bxZjODw4odgAFiEVZGmndDj5jMbWmbVoeVYtAYyHllcmm4z+700mEL1oRZLHtRwj
7qnRLEMLxRwDwNBSDAujdYBFiuEsnPN7PuYUaA9OsNzx33/6Vj4OlbJpF1w4MphT
`protect END_PROTECTED
