`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4c3gmK1oCevgupKhdPK4aeM9+xVwSfCApi1rAjGf9r8v5VRiarw3m6TJg2rSUaj
CiVYNqNRre8MPq8gh5njLn5kAiB6zhnIu68DX+1R/wba6p/FjdxmzzUdU7Knitp7
KExDnHEIghwvqDkMQC5BqQZ+9PYWJLLDOFa8C/7Gab2JhU4S8OrJljwNsFcVxjqF
wB7AfgKTkh+a+Nlnhe6UzE60MgaxDzzqjupFG1Q7HrAY0kQEHCTJ7odn8XAETjFq
ffOrX5H51VxIE8W8MifH5NWfHDnVpDo7Uwaa0UaNFDHPWb0CM0lZAP6DWiOL6PCg
cOwagBOPWN9HLUZESbZPrRoNqQ1s8kQzm7nAayHy2FHBne9JalLeGR+dToLwTsUE
H+2LGA3AABQiNZofyc6P/zp4qJKCVRSmdvmRGJKA6gc=
`protect END_PROTECTED
