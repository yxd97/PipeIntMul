`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3NXixek9ph+sFQTpETTXSBFnY91Hpy0+StkYI4VNUlf9UccuZsgvD+STsS+DN5X
pqjjWh62rbBAT6nNnoiJpS0B/B2oOHUoGFsPGWaAL4HIRwtmqxhG8nP/YM+Yuqju
427QV9ZyuaslIqfKJ1zLWbCxycovrlJe/CnXkeXzB9fa6KK93UGn64/K70O++Lyu
V0jwR8kkIH6BmIa2CvR/dRm8wX5SqlTjP3Ahq04s7Cdd+ErC0U/ZHNlIScxgw/He
FcdWOZDTB6O7ehTz3/aqop5LwPAUbAgD0xF1TBQ+rpvBvgNB8bNnEIG19gxJiGOA
PY6nA+VgTFbTGUgE5DUz6dUUNqdVkdEAxWpBIOgI0JQ=
`protect END_PROTECTED
