`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Oa43Orgo7sNI93z0Mk9/UmEkvpQgGg8XEv2Sx0+46u+5G2WRp7uonx3Z02hMsRY
SgdXVfn+1IcpXxNi/sCZ195EQE3+VYbFcOd/q8/6gjupHTJXEnMQsNAL2fHux+Zl
3JCdrvDEr20Qst3rGBD/G8aLfOOuCnfaxucfxX+KlQgoAUfv98NvtMcz1mw81sMR
UazZ/pIFhujVr9pBWqYQJEFc+bOYcDMITza2dyVeuKDsW9iG0sNllDakh0AbX62c
zhFJng87ga53h6p9VrJVNRbL3BXguw//oCetPZhSMSTuvBatart2ylFroHIGOHb6
r8jqCkTviBdg7XLLqjjwrA==
`protect END_PROTECTED
