`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCuauIJ9oB7upQErg+Ek5YVgTsg2MSD4aNzHRavb7t7P0JKCH7mjnaLcyY85Mezr
y1XeZqfMDErgACCS1v3vYj2lNpgTHNJJy0SRf/BpBAqIavTDN9AD+iijlE1Or292
wuauks5MsB7xs8XYjU0h+EnAFVtiuY+JMs7p3oHffrWEItx+hQfZswNbgpFnnHe8
T/1HqRNILWB7xLUk0rHSPa/cqHyKSQAVCzRddjNsYuMsp68/ZK5BbUtKBne8J/PG
sYLjvt4GVwDzqXt6LDOagmaothLSTaRlS4kRLCi87wpu7hjmBrV6S1Dr9GS4+Rr1
`protect END_PROTECTED
