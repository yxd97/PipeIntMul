`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOvjPhAh+OcaoGbaDqdrN3Day+Ocs6LTnpqLCDmeJF2Sl4zCMLoMLXTCmk1wXWwC
PRXb76xwhTi5NMDkcqxcesb0GKVm6ISnKgxZlE92IZUaI4YroKlxsUZzO64D4+Sq
M8TIvu4BXFJr6y06KBs1jdBpthJcyvC05bX86ZGc30t88AJqiInAaT4Uhgly+m1S
gsRkwvFEgbO/A23/9Vsu5uPuxZo57/vFbmuSPOJoRkvHn2fiIwEC8yM2aFqwLIFD
ih8rCxVv4Y99d4r4OMYNf23E96kZSE+aDFb4cUKfjcEtcN4dZQgwVpGoMEtp1VuX
x8xtfVrcU/DkQuRySNFYQyCYOvH9uJWbGq9QUHnoyawbRrISsHZ0hO6H2gUWexwF
HFctkiyQubtsmABf+g5jl8k7OAbkF9xeUjmlhlosxAy1APJfogHWvhPGgBEnRTCL
aKOUtjPpLKjcr7xW7uEILFK+J/9xFPA8fUpqIMbLtZXC//z057wwL6DGPUzS9XNy
iYo8C71OIFvoEnzEdFYjWJ0IqQHwe8fMcgXeu91PKu0S8NIYuD/fQidOq+1NOae3
3vKjLQb1T5y0NmHXz7VzDxyEM9jcn2uu+U0Z3I7mj9oEKv7hcK298dMctVEkd7Wb
/wrDtl2BKmzLmmr57yDMG7Rzjl3ub+kZvDYG5iK+JZa15U6tvXPsDLtN4BjKYaNw
ThsmtjxExHH1OpOH75oxPt20qzdEcVi1s/Zd/OAgRSXNiv1NAnIdB/vWiWEOVh2q
NrLpezwNIH2EIRAqelfz9mAGSkARamFprnz0FnELIdp49W5UKByQQQ5xC7NMV02z
o+0Om1GSu5YGiPfglZOgV6xOITxu3b47aCmh7x+UqlEuqjLvoeWFwUDFjoCe+t8g
LtdHzrAVBq5N3AzMYQDEANjr02y8GDNpXaQ7NlpkvvBT6eEKgHK0I4a6tvCdobCt
ywkmv5Qso3Q9/+Sy0sTJSdtfOVUCRc/ZAdyPu2xr9yz9SoVV7dEH7hSBykkSxie3
qTakjwQ/I6s8KuRD8pg3hzmOcOVeZG0qnjnOptGTKxbsUGbg8Q6OZa5kLDm0V8P5
6VhB2r2nouuafhLjCRwtuYoewyDqipRiyvbbAFr+4qrzG+DAoYgBCXzEsLuDAEHm
3PmFPPNibCC5joS+OD6zwQdxHbsEoU9E7+uIxF6ec6d3qdX6oOEgU29P/ECBkUrR
PzX6eQY7tGQLmplgBI+55i04H092b3+Buz+hH1cMQ9196ToI7R0LX0NFPbfgopPY
PgA5jYX4FPlUCA8Efop83JBv4Qv6N8JjGy9dk+uC0vl3r94yuZQBQ8wW8UCKtaPN
7dN2xrbquvg801qfR8H2KpD9y3JST0Em1sHmPacGz7W3vV6e02bncdS8aAZJVRyl
lrJ0WuV26R7xdzUbCUn19PHS/urNnsDXmU0um07TUsY7QApp+ATKeiQugO7xY3YP
/2is0AmElnrsUTolWcV9NUNbQUMqNBJ75IUsos57PhAjhTiyAXac+6lJ+O3Tpz/b
pgwwQ09pVZy66oPZBaPwn7V/G8W5+GO7WHYT33kaeCAETE8qpR4rrbJVuT0DFzD0
rrUbhjXD6gEz152szWHCcXrc9AfJuPmW+BHFQiwYvJg2BrT8s3mVRgN7BZguHHMq
5jL083xVoghZLJDeZHZ9/OrmUhMDLYwoOHQ6gDtwHPPKG1uTSZNrDdMCYu7JjDR1
eLFwZtEXv5MiY19XAF196cVadM5BZ+RbznwDc+lrl+KMwZnDEsEy8i/juTqcLoeH
hwFLNYSatHzQ7DS137J2VMNUwRQzmjuSDLZbcVjqvMYNotAbb77LLuzDJVE3B2wU
vPRE1CqeQeBwpM/cPJsf7U/Vghpk/EFoGRxC20rQIgJRBwvPpGoNJE+P6oPqMUdz
HuzJ8rERC/qQykCntKphvCXSzXNxT+mQRmXu58oMazynR4kjBrtOn6fpFqU+xtfR
0uadZXkzmAcEdA6cPXFEu1/WCtIo3aqw6PSP2P1mwr3CSSNTSKcK93cIjhlzcQRC
tFUgWE4sxXpCcO+yQx7o0A2nSUqY0IImRWFBRBunNK6NUDc+HMNEPlB02g+ML5Xv
ZxRvtzyPg6jUKRR2/uMahAzCQpLEheZTJJRsFClfa6vErA7TBAUhj9qk4wI71Nl4
VNWcX0x5KV3D7SjG3ow9I/fhdgStlPN9JSgWFSIiepmb3ydmR6f1EiveU4mw/nNX
krhYoHGxy/rH2OCHc0TwWn67USSYrib8VUp1CVzF66wveMXuls4fKXM0JpVs8gM3
VkUwP/LJs9NxqhW1ZWTPxR1BFoHaPGR90zWQ5oK+xUJqEIz+dCyT0a7n3j89MCTX
kIl3vagiMHYQNr1Ad6Ybprkws6rPXEwXNpBMUoR1fPyucJrXdnQeYfJ1oVk+3ZKE
z/hnKkQFt8B29G3vykH2dL9NcdYJLI+sKvDwb9wMCdSzqQFOmP1C4gLvcsUJNpBC
Xg3OBm5ClIFyXL1W582N8a0eq+mKZDwNcghk45Tb6jMAhqyod605i28dyliqmvEu
XJhr38EuTV1RlEq9zC9AY324a5vxNBMH8CoGYoYUr+Hjc6alFC54B4qf9ZQo0dxX
IzXXOlc7rtaKodCr1EnLBmztYSM4uAnnjeUZ4Hkf80OotCF+xx1R1KJ18zO4Amja
Bp9IVBBQaYJosdltrrv7xFN27QQnT7rS/n0M4updUqGHAYIOCArQxfckDyhLXCws
eyIGCF4JOAe3OhOMcBThQ5aI5uvA1HT5g76XyFjQLLX6mZdTZyeSRsa5OczmQ3Kl
OeEZjiJNeGTZ6OZxIheFMlg59z7FDIgEmAb4sfYpGW1FlBEw8/m6cBqNuVblXyYE
6BBfNPSmC8ttQVRWGDrgKsmEDi0BEdgt/cqRLCAMYBgIgBwZEtSaANHHTTGbjGWF
+QRmNOfNm8bapyG0SXv4BUNhv99RrTVn4oJKcPh7KNR2fdst17IdNqAFXug2n0G+
raXYzOBPdk6Nw56ZXDGQJ6Whgzv9AKDkU12g2BscNXizDHh6oDsUBPrCsvL9RFVm
4sOeyGMNl7ry8lb8WXADYnDlPCXk845RZNozPWjl/ldI4Xsm16sEHS16TM+Anb7C
pUGfCoMj/ALk5wsRn7EpVpgZEe/mC6MTmRbjXcYNWqB/KkwPo2Y8+4SBJyWFlLLN
lUIUTyLXR/dpRFSN8EB921K7EUUy0bS7xf2F3JnhxGNxnf0nXL1dcp4llZQ1AXte
EUtOYWAZ0gU47YaMmLlppunfvK4AyFEoUKtLJKrWCgC0LdxVbQY/Fopgg0dpNdiZ
Enl/MYZgvk83AoTTLwJ2TZdVjjt2KqsAlbWi592p2BUy8CCVx1d8qzrFkY6+EXl4
Qid1Wo/WIBiCvhREOV7KAy4/oAGXqtqeb/CNwzt+L+8Ee3mry87VXT/3mMTUQc9I
7QAqt8D38jPqjbtFiugqi+29jJIFltpjKfedl+qr0qojM4SEt+JOovBbNvPlaoG5
jQMBO4sXKGB6jlyxj8XD7/uGFpI7tOZjcxfyDO39ksjaAoTZg00+23A5KFSWrX27
xgJF1xRFh8E/gyfG4vbswCQpBqzAFTlyhpjx92s1Phrtg8tS0MX6WTbIsJjvRp7G
zPh7Q5CQYSdP+ZxCWybjZqM4jFOu0pFIAu0xZakSfl8tTX7WbIiTssfwGHRotks4
Dtt86SNc05OLz3S5jk3WESLwfv5iZ7sa/P7SJqUAMPpLwJ/Dy/AKCe3JB5yMKyCk
joGqTE/xRWJLCAysQg/l39pXurztAGQyL/Whf4RRb6Wje5E5qXvp33ajdw+SjbAo
1DeslQRsOC9jl3k257Fh9m2W6fegJr1eaLO6V2DytuXs1+r1s1autLHwe/wgIsnS
hh6sYNx3uCKtD4oOT4mRJO6ixq+GqIAZ8bKx9GCE5aKDNlu6CKPaeimMbsVyx6r0
dPEIqsdhQB/3qSRX0DOdD8w0D03OCljnezsdyQlwoEyVu1UcMVOPNjyuHQk8twC7
TG6s7IBsq4k3MpXoKTBNYRXMzbsolotif5ozFg8AQ4ccNOHLDF6gTal/eCwjhnIb
ij6zaaOpjb6gY07F98QFs0SbfXKRYypy65pPFPTqvsvtqwK7mK86T8sg+0ODfler
KphMfqGNyNZOCIpagpR7tA+VO3RMcy8i4rSsBNy7/2issIhKajiHKobU+wRx3AGj
07IheVQaU3rH5s6CXGpekUdrVMsEcmZBbfrmeaKVk3wD51lfLoNvBOVK1kdX6k/b
/Pe+91G0zjK2cAW7SkT3TqpY25BvgGLcZSrKe4yNgkhO4lbxKVipgWiXDSVycxzL
vFvkeGGpVd+6YzmQH/e9kCfZixAQpo84pF/Jn859eKYP7zZL1i7D+SRQoXkIIwj0
wKoJpZ7FX29kW0RPu9nF4LfKdx5hw5NXi8TfYXBxV6fzb7fRwHoqd1SKOFQphB+z
qhk/rOrMklS1DEhcoYpT9KLGVlIRDyyqFJ2yV5yH/zjkmwoe7ZKGsre6zzpYgEXK
YoHxjNLlqvAzmI1PJbfA145m6hYuw/6aop77ob4xiNTjL5tzsIE85YgrAbTxyaFy
1SFNPAD97dZftwVeQyvhNEWdpJ0uZrQTF8CN00rP50DOOAVRtHR2aqLn+nTexLUE
sHNbS40l02Fj+j7XQ+Bgfuzx0reYXlpiQfc4lMNdu075xUZNO8FVPAGsyhCqzjYC
+eIBqLGTXtn+MHqYaJeBQUsJFFcj1UB6zao71UB8JzOD8Bl5jIiqIakfhDBphnTs
/HouxVl1dMHyqRLYKrgzGnxrInAsXz0vcD2j1mdkDLJ/DhO/n6TShoRi2QHKPSQN
WzsVZZAXHH52gzQIfED8FdBuYhJUpnckyA7mVVPbnfHc/2F4pb7fD3Dan+pGYWvW
PrAVKLbSFrCctZByH0jK4qbrW2BoIljnSZwikDY538WcMlEBQ7l+PIH2F6/ssuxd
NXd0yP7CDI55CH9vmm3kFlTaTWmUrYGCXe1Y07DmquN+KKBNgYMoMmQ/ZKr6+AKC
L9kGP6AD3Zyr2rh8FY5Eov71QH6yXQDCuIKm4jNjOkH0163DywkoZ9/bItNYJTS3
OBp+n7VDMCTxT672M02R1khkeb+ppJ1zoVHJLspUF9B+wXogWwo7Na+oh7v6Ins3
rv3b5sAJqo5lgZTUi6JhAgJWEP4XnLXNnzTZLEV+RtnfjeSzl8wYRvMW6Xrfyneb
zzw3kfy7l7WkK4RmgvlilX56bL63o90G7inij8wOE39++1Q3H8NRy31zfUReQAc5
2Dsqct0i1fz9TD674TUrV4q0SZFFpdDaAtp/G5fyyb+AVBW/VPGUZAsYTmJ+Sc8G
B1q0+7cHO2RleNn+npgolrJOZniS5BHFi2DxFNTg0cD/2y9+WywwXZ+VYHENIs0+
GTMmpUUviOAl75cxLZXNJjkTloEw3DtPMOlN6RXQJ1G84CXGNOiLrp3xE6kDxoqz
1+b/UxUNlXNiuXCxQN6dmXYSZvxO+sgwy0SmdFaGDgyu9Ib4CXw9lzzZpw2y+9Eg
GW049/HP654EEa5YVqmOAZBDisfDZ1xD/HNsIozObPZ1JNFoANAbxyqjY5jcw1fl
bJCvpN1cVl2h/Nii+YUw/QQn6B4xgTaE8gaMoaRa3fZOmopYS2Tb8HcXRpO3/2Y6
o3PwIuGqCgVlsMct2yu7n7tG8s1L9Y2H5ZB2TA9+0NE3DkMk5FMNNJWzWblEcbIF
s9O7CRLSE+I0C9GO2W+O/32U7rmqDBzw6solde0ZdCi/cuabqTkuYwERBlfS/tnp
ZGjn58BETGYbu9pkIEuejoDLkVBLx76ZW2jrUjXwSwu8ozuLxNm4t7ecT6tz9I3T
oew5UWY3CQF/y5tMMkkSdV5c32fW2KrqB01mEhzdR0eOIqeHn2t4MJAJpBdCT+lJ
OB/MuU3OyggBHr5rH2p37IBxWmIhI+UyY8YohtIm+9CqlGrftJZ5M346bA4001cS
3j0lOH9qsZaXpVY05r1T3hJVdfciHxj446JEbPK7vp1rKoSgCCj7zOZ6JTeDlf6T
qzi2HcEB66yp/qETG4cJA/AtoPtFEvUcbWtJOM74GYx3NNuvkOXZFUoq84LFMiCv
EPD3LWhM7czH9psFchps3v5vHzoIQ0YwYFZFJHMJPw164szzEKRDs1W9k8nk3jce
I7fKgsMpQhKzTSl5B2d2GrC/84gtH3DZCE0CVctPTKkJbNuWWBZH+dFYRU6YwhJt
f//UiL9/odWscrQC52jt3SAppewj4RUKd1QpUupBDCDrigW1aOvXKo91EDex5MlR
7m6a4rcK9qB8Z/jHkfXX6seAi6H+CwKhU6rz4ZYk2Zn5TAMO9ue8yHlLL9eQr6bu
IF1HOPaf1hFF/isuPpVyTRyf+kMvGwo+AAK/nCnqyonmxwVyDu3O/FZkz0Ctux/F
siYOcrDRjaNMmkboEvCI4wtgruoFJO0m0OZhUwi8On1QIKAIM/xzXLHeVNkuR8yM
hp2kMS/ENZ9J4kIHbOEe6Bmo1ldRGdAvST7vJOIYExBkUdF4BP301R4XQqXudWpQ
hCaxcXChiErM2VfGlbHfkkVjLzpQLTdGt+4T4L+oesANfjxLSsS5FcFaPtkooKIl
qM4uENGI9wIHIjbi1wSqTDQ5obzVo+hK3UBBmWfvN3BUwP55TjF212caCimGpQ13
zNsNIXpG6+WnwyIOxK4nSjB0Sm5JtJf3nt/8+HePNIQFbFDJQEKMk9QpPpo1tGXf
gcleAZwB6GP645HEpXOJsT9W4urtqxAzlDZvvOZgLGubhTuF9ND1+k9q8j0Dj9iq
QFl4uOO7r3gqhG8FqI/YVFxTYUmMX4nL1to9uhUfL9Q1cg/JISI/GHLW/2gVe0BB
y41RNUdQ3OTnROczU5bIM7IZhlL+ZqWE70YYDkRPPMgKsLQ675An+olPiXUX9WM3
gfU8mwElO0SjoqBXPIVU36WB/w+EyKqK8CS5ZyBz8kdymJ8NENFEWYWKlHouvYiS
r2dkauy7CvUWuiX+ZRYqtCHnAnkoEhgIACDJCz7E0UYARRcVsd8C3cSjb1E5zYJI
gLXyXBGaMx6jdUNMSXJdfwJaHxbmtZR+icjLSqxcHo40YofDnmCwG18uKQ4xtw4E
oqdQVyv2WDVjQ2+8rbkMyVWUHR9+zrmYdf7pmvbVG9VBi/S+eJU7IdIImAEf+z1K
Z7whQqfQrxmlBPuV+xZHFAk9hqg3QBEqxJlwbhqe+O74A8tAJaFbPRgyA9hsN0YC
+QSuzqfk3iwpUu+qOqoYXmNgInSKuF6zvGGZBD2hQSsYobuaKk/4KPSEofGXs+p3
H5oi0u3LnIqIdIWj5vHTzYakSK7sh18FDlEJQDXtCuxI2u2LkRS2E61P1LE7rmIH
1kSA6Ga5XKbCrrO5JRMzv5tDWVOon5V9Txrk+GKv0Csv+Tgqla7fyP6+jjGrTAKl
kEjFL63b8yT6taQqTSOMQVwPSv1lgndXzEcxctOuwxKPUsefjUvKDGdXppIbDgZN
mWZmBsEJBp5s7RORA9Ww2GRdamva9WlF9SEygfmTy/0yT3Xx+sWiZG1lEYVmJWK3
Op1uXF5sT0HR6f6KDz425Y3DJD2ObgowIRz4tnFo4xHdp/0Hm9ncRAFOQK1QTaPp
iY6dv/HubvTUlf7NtaF7qywpTJAsvPVoTcJYFCrYAm8IvKvLt2pjK9pB40trC0Hn
HjSgze8GQ36m2xEUK0kdl1+oQafP008eCa/JN7ZYObJzMWfCaa7l/yA+8eEEAuhC
6NLlPbd/VZ5pMD4RfQkeDItjgBTGR1Ygtbm7C+afWEFSL/MWh9BtFeHrmIiPuy4A
FtF8nqMtTB/00n9WfC7auAY9YnIwBLu6XX6iKg+5kCW00kkgPsga1E0V1YOHKf6I
FZutVj0BkOr14V04HkDLiuDXELXM++rcVvm/ai5+vLqaaRI/DrxqYPc7UTJ+2fqg
GCXLG6EqF9fApC9XXVyL2Z27uJvmDOf3sGe9rheCZ4wNKBPIfbSG4/dLsh2I+daQ
MqYPMdxNGyScuPOcXtwJHZrfVlHYT5TAfqlNHE8rF9fytEGOyFDvf4xFPke9v+RH
I8I/BAt/SXji8mvW7XC2Ct5SX5H7p9hSDMRoxKRtAVD7opziMB2zIejdzDtoQrUP
eHLoSUPj0iyWV6xI+Klz8dNI5046AGO98zwT6TkJdSR+NLyRgHX9BL0308gD91kX
+08zZ9AiqWGvg/ce+PubdjF4PUOKDX0fuOeiyHpI0nma1NW3pe7pNPZhz8yGv0hH
KnM43nE6CSWMFlmYXCmUFkNY4gPoBHdmd4yMC6PQcjRwf6eAvdXN8SUc2PgUfTwf
XZ97gMdhedxvZidljnkiPPgHMKE7AMMq8rzosZUAPWS0Orxo/zI/gPQJOZRP8bZC
KEzdztnhRBKyqAhYe3imhTlunBeZwgexNL7oSbAFb4SaHJuTxVZv0Bna7gmi/Drq
Yq+vctysTFODpzbxMBWDHJxbE+/3CHra2wouymZNGXT/8eXhiere7mc9qyXrlTbt
6/2GhF434Lwyh+R71tksF2MiyoKF5R4/OYiO+zRAtzkjsd3bFZqitsW/zqGFPdz2
5X7/qKI0NBdPUHe2ZDf4aTBr9kSkaKj6/xjyds3sjtyZaLSTmHRfsNPOELFt2TmG
tEliHX378kxwAlc68D+1bu1GdHD4KMJlNPcYD/3kxHPAP//YCWngUFOn7bPdxfGB
NrGaWB+TmRqYlcsbccGp6eyNJ2gxFh0sgQB9l89Ps6ZJq8BHbD/IjGL1Ih9ahi+g
a2BCQQo87LIRoMFNHTHXuosuaiB9oUOprejHMxeS/Iev5i4rc93Xr5Ev8plN9Csq
nTIhd/Uj+x6ArBQdlyKvFA94P1MjJJ+Pvh4iFgRbX7u+SMOjdrp8cCnTCF+6VKh5
1ZddAviZ33qMr776FrTMyelFB+zEQkMf/MKy3cUiwHQdoUsdaCtnv3WfPtPYb/AJ
5/n82/6tAGvzOgOeFUUSsbbCyhXGnEue7CSogD1SpVxCZJCQNfnaA+8lpqkmOlE3
eIF207AEKYfoD7jMrRj5p+xONh129Q51ofxbp2S95ndJWt6H5mOcWYx2SLxHXsvE
e8lH6CpS2/5s3mLDM8sj8r5CUReusxFENNjf5aQKi98HBWZipodefIZ+xYzTCm34
WpQRHZxKJjZj8Puqaq7xFDZXZTwluBx5RgrF0NY7f4MVs/xupM6JYEt1c79oJvUG
lDx8Kim3m57LGHD7DxmKCzYYx0KrqAuxSyVKtzWteJXn0Y7ediTItBb/iIco/CRe
Mobncac3Qx1F1jdeJnf7mkQA0p7BIwAy3IKWVORnL3c54asKlKsfSi50v15x2l/K
oGNB+tyLpZXVzOlsByMdMxGH0+ilppkhMIaF0KkPEcodSXEnBtKKGImgdW18GXeE
NUFFHxkgV752GpQ6jWUEBRYRP8evRiRQjAihb/S5OfMt0mNOORmED8Sk34BE2yDn
Ji2URjagjv3EwZ+k4ueELqCHhXGwGVQKy9kZQ9fZLmHwZ2dObIte2I0Usg8BElkV
5bMSZLnT4cSI8WOr7JVEGhGoTv3i3ASHddf2gBBpcslk14UIqXe0bMZgGShAQyb+
4L6Osu9TjPJEExPk+LEM1Rcx0U8ZnSvoof/Z6MeTJPV1wOC0M/BVDp0uO7c3idpe
BbhV0pXKTQgH+f85J1ixC6ZFm80PeLlDNCblpDimjWIQ/TqjSPu7Wxq0fg2Nkl52
YRYz7+pEN9rNZ1SCBStZScDMBLHliFfyywrA7nV2neKvGG5+SnJCFe70qM7FVutP
xr9rKetgg95aOY/+RZZ40Lc+JUWir43oQ7HXRzoa+2zHvTOttEabaLM8NCw1U2x1
zKRc4N7uIHFYRlU5wRkKCccsnvXd3TCgSfGGO5OGT+I8PDhQNu956wiBxC9QvQX8
xnLBnS6ziA7PJOf+IMTGKOJxIVlX/R10uFYg6MIH68OIwn4z0XMjlemlRcpOB1py
Y4g47Z75boUjbPYMsLFCKP6gzh3HfDfGVR42i7lffhvWbV3ns88OF2G88WDGezur
RplCq1ZVRcrMim0Baeqhcnz+/b0zX5wfsfhDQw1xSs9Ue2nGZPF97qkZ3pTh796g
jhWh7Q3EgkCyrIPbnelpKONS6VW4tBojVB2/vRqlkYa5rsI2LbLrSKXP4a0btwV2
Hm2+lZJb2iMBOhyCgqRlZDeRKEwNvwkZbZOeUClxX/7M6IEDWeS/QqkIAIkTqzg9
ithdx2bdNNqFlPVby55WCkDkKQQpNH9o1UrTFyGVwm3GqkxxrJS9l4kfiIW2Ei8h
elD4QVJd7UDqxBPzVzBbUY2vfR2wimXPX+UJA5TE9VbFLjZMOwJc8JE33AWbHk+u
9YRgDCRLcKG37yW3A7zGeVMrTLytKK44gtERNXa4VTXiCz8AsFcidRIUGo7pA6Rd
L9W+KVKDnLGPHEAY5uCGbyqHaMgoIgjCVeNg2Ohe4mMbaOPzDaigkQ4cKX5eE+i5
iwL6QjJLBNCz5I2apC617wtABnOhuZwXN0I29wJO7X/hnW3dkwcus8hEvcjlyik+
xiELuWtBUBdJAV0sfmEVZYM3yZmxfbRLVJhQhQa18SVLpxE82ylJaN4V8eWVB+Of
45+Qg048RAJM/243pFTKxQqn9GsCUgIpFVbvHrAcAFuh29fadd/nVfYaeWi78MF0
rqgeI5FCPe2eokhdCe4cmY7jMfqTYqiMRGqsQpC/SNwkQa78Q/pJjIeQ2DVHbgKB
UW44hzScJS+fj88keKduISNEcnJ8mQcUQjSeOuDKvM5zHWremYz2PoN+p68u2P/z
SxlUnJ90J6XiyWGa9MzWWBZKhone+IXVTdPdvrV1WAu+ad4AqdDEU/QYW2AJbukl
QuLwKVCbzmIHfYCkYOQXxxnDHZCiToEt890RIV5IvV7fuRigrMPALogigcTyDMO1
W0S6NzR4EzHAnM46XFJGTUFjTIr+9Pd+kqgOkxqH25cpS2eOVychs2OzjfZjMavW
stdvtSlAypjSDdMJ2tW2fKJkzEXl901mWSk1wq6ukoEnUiT1CeaDGO05d2hMoT8D
/5LbVY4kGOHhEcFTBZ8kSM/ywYOf0RXAWRukBbEPFhoa2sPSnN42ukieWGRSaKfd
CwFK5NyfveGZn918VQ3wZIN0P5b057V3/sSCLZ0ElVPbwkDaY6N5lQwk4++l17/0
y2br7/1VEY7T2Efh8et0GZkySQb4RCD5BSBXjSMsCaDOv+2Tmef/q9F/iBFWrlch
xUZ9aklmmLckR1Be/A9B3w1RTibmGZJtqQx8ALt/CPns9gWdDGDE/AZkP4PCUUTN
L62yCL4zvWBNq1pc2UtK7wocR9yDdp1F0l0RrQGbFPrPsOsnt0ZKZOHGKCuWKSry
Qlw3RIFjUBEodlyShwz3MqaakjtwYzWsePBcz3+gmSmepd758uKVNM8gXQGQ8Cgq
FSsuG7pwU8vib6kVfDQyFjNHexQ/CIdkkgt2wEUdJN3Cf2wXvcK+59eBDuFHT9zt
6PN4ngCPFexv9P5n7m7RETnL1DHaqMK4mjlEfLADAWa6gfB5rQXCgCQeWXEcdqnf
WVMNuLoLJL3gVrVmjl5cRW4CUxuyLzK4yzss71Pj4NadUNhSWUaAMXlOe8yf1rWM
BIwCbU6z9Dus98WcQOq8WksEEwS2rpqhA02DMqvmLMorL6nCtALMfGttkKtbP0cl
+25r1Y2glrbXlIVHnm4ntUO5ybHQNHN9hSvsJSLzxz0vDyaJkBm3fib5/m2Y4KJ/
kUyWQ0KkwxqmV40OIJ8Nz1QjqwAedlQzW6vHxfYrCczb1rrqxK3TrsMDh3y8+bTm
SjkuK39c5S0yMBDHFglGyEpm0PZjKJ2QtmwQFAd/xBn4gRMgMcpNvXw8flAV9RHg
A5sPH+VqSuEQ73QYMw44d+rlFtshPZ5Z0mc0P70OBgDaq4eatxzcVtaxLXIAw8XS
WDBRGJnQvRgkOpJaMvIkU/vDCcxl5mk87+arMQDJ72lMIffXCb4BvIta9nl+1H6D
Kh5QAVookTSGLWmd10APH4qZ2hbkauTeQmoUmM3Arun4XpAdDx5Qn15AnpyiAzEK
0Z+Fl4tU1GeHDGWYpTcQzMRphzAMXtZQwy+LEU9F6H1Fw2BxTeNyp/rtvZokqgZq
GRecoi+5ZHCm4q0TSJYSxBR9n3lkYNlevGlcTsrInT9Q6gaV7zlSJfLchAnHeoYS
5SpzdzdIqRbzKTt9Y2smudsSp5lmmmHYRcFw2hcz4ygiHBxrKtreurqsZtFpxzpn
h/HT1K3UReUv0Y8qH7Bu8iQDx4KdlRMMdyJWdVIyOfUIwJMHsDz/+blSToL2XJW1
vLc2yQA7+vbzlsYavEwu4y3QhAEYJPPHk48R3aAAVtAMyaq7pqWo2FqLWVK5FRac
4uoPg226KwsDBMYLSKGg0e67qy3oSq1Qf9F3PAl+TkMqi/HUmgbyOD7JFa6zfmjj
MvSBeADzwgpB5ta13Ot27EeuvI0Kh97gg0Q/MiELnWqVGW/coj5czauIiMTSRVWD
J3pidtTot1aRdSuLCgqQg30lvzmT28M6ahtDhphwDQrz8hdbmLPTIiS95Sflv9eP
dnCIcMMclTTfo4o/AEASGTcSOeKsGB3DIZNeZmoJL3I1OSIFdwxp3A0WYtMXi+jf
BXzL1axl62EOvLINk1JEQvwlVPQ3dBBSZ5O9/blfFzkNkJOjn2M98/Vp61N8l0Eu
7rpU4heK3AjLnZdehko/YkEUIzKR/5qB2hTDldoX7OD4qi8bCygCj4t5NK7MC7JO
WSni0SfNR/P0eUNlYwceOUlT0i5Kl6JZIH43eGqmQoV+/Uzx7m38iBEzbJZN8234
gZ8/SAkQyE8qCVUnhMB1GfEdvVxUUyfKDb67GoY4i1Q42z7C5v/dnxzQKAIEFgqV
q/ogEsz13ZMXqEb/T1OAS3PEusRapzaulN6+yRPHLw05kth+a1p9ihacd49+GDe6
nULm/Bb0yfSXB0HNUonFlohxFy4TSNUCVQpm5pX9sLTAdsTgarT2OwfZqSbfUDd+
WohMiLPA3jFP+10MqBRp4siYwU9yx+HzldCT6i6OgtLXsBmmQZQIE9o9484mT/xT
Fk7D9EMad0pBY09nm85HU64KRMXavlPIwcU8OlIS3kPnr1j3FJcdfOlUzXmV58Uk
Y16oU15nD4LlgbIPzO0BtsXnYfIObQ5COKpA4Nb/eWY03FJWPGYarA3acr8od824
DCZXFIvhD2B2rgNsdpKUg0hA30TNEz98xxHDkwkilzuNfYS9tNgQK+BUxmxRJS4Y
lzuw6ldtR8JUP3UkjW9KjY/nEutdkkr22g+Y7t4q+0Dvi9pNO5DI1rPYtCOqyAEV
GMtkmCZvvAcr5LSNHzQYYyaOtbK0Fz98M+0nR93sc1r9lJmLgbiuzr/I4Rs0UWDh
WhQnAh3gGmAZ1mYQ+n3czPisuMeBPDygfGE45PRewwV6ysQNuzdFW7a44wgFb2OE
UQGMXOgaqUz/Hahk8MmoaynQ+4xc4p+/t/2GdA9GJfcSmL7n/FsbOikXamSZIsSv
iuI9zylrsBaDjhW6r7OxO7/EX1cl8iK9Qv7JDItbwnESfYWVzVwBNzVL+d2UU82A
KsD0b321fa9vypu/PJUQErk/mS+LLq/HnNw7hqexN8SfqdaOQYAQcw87iIrfXhxi
hAN2J8yeCOrzXw1K+00DRWyGeht9BRGS7G1vAe0LBoYrbaicYDJbBj3ApeyY4PMm
N4iCzZdWJnDpl0iC0j4ttzE2irhCPkT+oPXo9119h07+Tvdn7jAT5cQ8sOAthniu
5ZQn8rSNDvKCA2+IK2B87CVKJ04LPOLgzfzPYEAN3H2k068PQUjD+M++M/wwBPem
X8uMwMYHm8ZZYthff3cnk8y1/LbMywp8apYpS4kPgrwOhRHOPLFsSxtyySndP1W5
XQ0eTd7MA537x+GN4FHH40tlluIyu59/28NeqAIBqcxgnzrGoE60yG9cWsCtc0Bp
TRPs0CYw4ah/9HajaSgZIVVRXeXvLUTPcxFPN79kwsBQnUYPgjGfm1b2spFOt/em
HJYiAohije0BD9KZpxgWMF/WuZCHGo8foeLK2H8qsebIITGSdkeeqpp/AJKqQ8Tv
miIcAbylf48wtfx23SYnyNs1cLi+/nv7dIhe0ew4LYszLdFTLdZRaYOVLC0z2qG9
w6RyS8VAKAYwstOCgvuWhQVUJSNxNko5fWwcqYAlvFasJaJF4xuIq/MCe1IYG58y
J+UV8clUO1Ikud9xhERAPJa+nOrdhmQzJ74iS2jV7GutHe1giHAQV4O0Lze221vF
qdO6CRF7qUpqRsZ1DLBdpVn9ju8HSPjDO62GP59IGM9Zabj6vdknnt+Sya+Ldqbv
otk1MaM5IeVqBUOvFqyHCmJV3m7rvq8QaBjgiHyuRmP2lbrMoa5lRBeEytpBOkbV
PO7EIF2IotIfpU3hf+PrZEd2wJNpBD1YMeKag+WKFyUZGAW7Zheg5U9oPvo2vxxp
0grqhP1A1uAmNe4le3rQrgJMYGg3JsR/AorJk8Bdmrte246q+qMvpz6MhBn1ByBB
GzIz17zyTwuFLw7ZKsW45cNM0b6xfl7ZYrYG21NIFyu8y0tJwFnUKrqFxiHYsCHA
7NK3bzIvFxGZ3kqoNcD78SJijhN7kSCJO40bpi6D2+Vd9tR7JPl/JnKdB5Pqp/wN
qLs7PMlUzrhPesEaJrm5MVxssPiVjaUbO4O3WYokQERImI+8Mqj7kDBRYnk6pvRD
R8oB2dFSstgGRRKDXQCMFjX7U81lMqXqvk/D5WuxK1nPg6Qlky04T+bMZ/Bs+ut+
sgZxNSbbwOiGzwO2YTPGa5GPjwYTxi6PcM1HLpdPYDI4/ekpKluR3srFVJncdZgv
MBniD9H+qmcDjqNWKf3rCQEp0NTN4AyY5lPAhhY4KCqEj4nYJIT4lA4NuFZZMmoa
86oPiiUml8Hn0vAEK1hur1MGtODs1JFpIzYQ092/dOMlwEyvhxCqsJFtTLLvAFOk
Bhr3r4FyFSJo2n9h0Rxp8PWsJ/o8dlgp3wLIIdxMcfF+OnewsLQjW3G9GFX7HZDv
60sXeRvkm0feiFJ+xhQaJBCNipuiF5WYfadvh1ggr9X9ljXiLJhqIMDb1O8wF5+D
Mkt2lb8fmr9BJnJ0haKBNu39mke5jMPn5haRw5zL80Mrjg639ozmdrVaZfMuJ03d
iAX28feqo8knI+E2dB2biz99iHXDgAWopUfM9CTljt+2RZ0ywb99xFG6zzUIsUPY
GtZCGbZTey4KMdasqCiZp2pmzAZLW58uZb0uHoYU1EhcnBn0IV9ADgHEfdXDJz5b
7eDgNNgIqFiI3WSf9WgT8MzFBRu+K6nPBrYK/VM0cZFhm1+vkK8S7opWMC21b3/e
rTMeDYcvioUWShHc9AaYo65gT+dg9I+VAIwPM71z21zOUS0icbfbSroGiV/FA6w9
eyz3KuFiumQdOu6cnFCOKfwZWVC1rwFZlxpei2d7Xr4GU/7OVr4UtKscNxtrnQzW
u2GIDMqPhzI0xe0vbYGc2UL0xClpY1Zeubnw8l+MpzNnLIPiCmnm6k0P+AIudUgT
rdOzKiAFc6+Qeb+xDFfH0faOXN5EPI4C1xYfqvsHH41UPiRhF9P+44oNWWQc3fFn
uxDSfleP8e2IEF0zTFn8tDzaAAyePC6RBrHHm2ecn0qzKvTDNqF3lDGwgQmVxi3h
oSVbhkrQmpbtGtV+VBgXnoJWplyqWVOaGuj4B0WjaxMz3IL9RqDIgFjqedGC4Gu0
EYwB/bQQii6rVfMyp4IhSLxAcwiz+8M7DOkAoFWe3iiqW/wAUOmW8sBVhytrWNik
UX3mWk/F1/1h7FKUdXwWdyn+hRLIdqR3EK/6cisjaWnRzv1dvIfjkM5e9NIq0Hj7
iWFymeCUV+TxU7+YKER14Bxn1JK/849HHapXD5Z+VsQAnuvtxf2kOedTSkyPXAxU
h1J27ms76h5txNkUdUSvlRyBmsm67WbCh7+p+IWMujk8OPjXMY/jW3Afj0qPOWs8
5IwcxYC7f5pGBEx9AJ2ODqVk5cVKWquw7ExfgLHKUSk+2CkTSYLXHS/WED4CBwAZ
Y3T9oA0C0C0K1fHubEhc1eHhlvUagOoNs6LP1IT/ylCf+KC4deMZRNvjvjhAe3wp
7BMbgYrOIcxpcuzPtdOygYsstkxEFnkFgkg/V9jXWl5Bq2W2fAbiuhGHh36TaPJB
0t8L0y3DA8n2tW6ZTZOjhy8gGZJ4xQHZtpvkrOdEjTeZqLzutK4mUGPMW+YuFsi7
ynWwNHboMWp6QYQasY6nGfYFSaTBh1jppzJy0QiuIipHKC1ScbTYX8YEZAXqCaA6
IXuLPhIsgFknBfwMzCcdy/BtIPZGZnZ7D29neibANpyodnuTDZtXrfilz63b73GV
Wq6dOK3dua/3JAguueXf8lIeAUNR9x5kvd1Zh2YOv0e1zPNkefneiJWFa8jnSwhr
vXty7FGSZNu87rqz/dAXqjZXOa3XMKQgwNDqT5i6UG+KSgjgewGu2hWaoHkikp4Y
Abr6Uf2QbhJaozWn/mVCceCFAq2jeliWQerHq5QlQhnzTgvAqSMq4v4/8q62dOpN
ZaTp7DF+DV97GnVpNW2e6fuqud3IHoD7TfDZUkIMEMwUGgd0ziSpyB0s0qugjMtI
oN3V9uQcYU78VKd03bdGl3ekOWNd8j1pJbqclMpibNtZmiAF0FguKDHTmQ8VP0Di
V5gtZsOfHYtBth1VfL+BImmj1MEGk22wKqejq81vSlzjoJVuhX7QkvY2nOR5q7ha
VGCkwtOx7WMDWIIc/UDQRX+l6Z8SLsKhE4jP/y/+ANR47hzzsgeUXquRv6sDmhoG
KXjO2k1cX0V8zIxck5Sa3XYZ/ykDeY25oLuVcdNVuNoVGla8LI67dd6pZ6MVo+6L
o32RqmJ3x6lz/xm+AkW33+zeW60eYxvDxA6VqtWy/ECOs6xJhuG10F5VxwLuGikV
hFWi/f+Ybt8T2Z8e/HY6ALjlkJkOTPAmp2SPkVIi4ZxKphu9kWUAFxXvLYli5dhV
LC7PPAefF972Yoxkdlm4hXe6uwFXIq8cNV5zfSbbttI7l0Hq9pItYfalxDD6oRlu
rRU6tYxS6MDpMq0gvcwULeKKja7qONQSMmx1iFUmD/jVcriFkb5z4iB/Nvi99aI6
ZemC2AiC1fmf8jKe6NnejsXA010oqTLEF5OXOu5N0uc1u+NvNZImi4y9iFnvdxi7
qdP2XzPrzzpiYkOfuZaMh7hIeSwYdfRmCPjRSAMMLcvsnVpx+/OTRDj85zhJoVW6
v5lhlk5yh2rDLrlhAQLeWDSBzzZkF9SVG6OkxzcDH/ySV4cwrDwLJaL9t6T+ZNbz
T97TXiuIIXupBjUIoHe1WV0iV3l5Jvwbau4Xq3yEKl02P7hzVmV/vWY0mDuI3xgM
iVUgnL1maAmC0KSe/M0XgajOIiw3kVBsQ4U8CJxGMAU3VgbPdZAyJlrwGGlZsyL3
2WDC4rqz8yU/qgAx5fENj3ylEbWyfnSIba3gKsivDqUSD3K22IYWjLPh1G72LY21
9AdkzFPN0aZ6bRE4sV2jYSlMkct1SJXYzTCLVryvToPLBy5IgfbHcy2XIYwsTaeh
VEYdowjLfUkFYoZOycKUwP4P9yneaENm+WGvM3GqOmVDqKskj0bwpGjzEkAGZd8s
LnoLjFDn64u8fReHTG2OOrF356ToFMxwFKpLr4PLSvgtRwe2HvYY2eHGVGDru2gS
rdbUHk19cJ5lTYSv+BLZUReCMTvlD80diNt+AuoRWmdPWcmR3M/isvxJ+PjREMxj
CaWUU7hUOywLovyZgx2+BS0HYLFnddWAU45MlQSKbO34met5LUoSL4CbsF0YGpBI
TZ0Z+7LkG5rgnysKKuFeRfnAimKhIjlxFt6ox3NuF3NW79UUf9bhH0SSS7tQIMIJ
R4GYA6bf9lzAueLjXreZmFAGuJmWrCc6gxwHJiiLhywKNaAA+ihVIH2J/uje2akd
hHW3ansvJXPRiW4lGdTR+x7ojgAn/s5NPW8fJQfAXvBQhiARCnYyRIpJnBbQ42r6
3ztiH83qxGh6P17CDUKAu/0dOvly5+h75JT8JDjHZ0dW8xS7wzO6Zo9Inu4Tl9ev
+IUTtH4WjE4/kc63go3C3LVjXTjCAP/WnhONsUj4QxYfxlixHgW59KiDsTzvAxQG
NOtmhbz+szcnTIHRk+i0WzUCGa6sPiOJi8cn6HIagOXrZUG7AOTm3IoGDRzERc/K
IfoTIrjX+EHFPuEt03OfClfVsabD9wImhZQL5CQHMhejbEbGXQQbz6SVPR0BaVKe
66L0ARZkLlQFuTWJ78XMO16gjk/ZoPSnjCZPn4GqvXZRMROdCyfQ2GLmjElBcv0U
A2SAmTgCBRCseNmVf+guhMLxBe7twc+N/6B0LdtXW8yh2yrLTsOoMaN/bSafqNZ5
jqWbuLKa2l3posC8c44q8jFkd830onECb21JXaqGxIzaglm4GqE89Iigi+o8z8DZ
FpU4g5fLV7WpnSxq/IfTfTI3naWyeBmZnFOmndJU0ozHlHyv2XkAwXLPMv4WKMg1
JlzYQrTPtFD+jDxvnJOLZzygavxznrlzHR54vokhepukBhh2Kjlopu3q2ogdE+Zq
HkHY/GBiOekT9Gqm1JimfPVEPNXiHMzyq+XaTeygrQCESzim/RuIAOmejh8e13Mj
lxxlW6cNJYjoXsNp4oLCvRA0UEVw6/AjNYv9/CfTc1hqc5v/tF+Gz86IIBy91WjI
KQKTmFlXCzvbFCVPSxuK0TszWSADMxPVB3y53zMj5+yysKDm+32lFGJnZM0pBJkn
eRRbrgSJCooLS205+Etfvl4KeBMdl2uxnftlnf+gKuW2/U/sLTzLPaRaQpcH6jge
WxtakSXV/a4EbhzaCNH6Mbb5rtlAoaoSMBuAu43uRjGMX4xZbEWM9KADVY/Pv9ZW
ZHytbHtO0QaRpjVwnIpJJKwMLc6dGr2/GMRVBwNj4njo16pnAa3biGRD4iC8uG+K
gEHT6t3oeMXT1mG1L1KwvK0c7Ru2iwIUSnA5/2NpMZ6fvf032P7FGZcv1j8nzbNf
8MZZZuVTMSkYsUQg2dGZriZhy3ocDAf3kB5HipMzTjuxZZyXPEErs7XGBJkeevmt
/aoGV7HzG0fzXKzAIWp0Y7Ms3dX50KWxP197r4m++9y9I8+EQwssV4UhyYgGHMki
cYdlpx3ceit9//vpr407/6TmMprMJ0KPfGnscCo02iL+U51amGOG3XZykpYq2vhC
QDaiAFBcwTmPbxMJUqQGTb4/5dEEscSRhFkYnmFiu1g8qcuQcDrHTy9UCmYOCYMM
3hYSBarNZ7I6QoRKZPGou6WvSIE3zaUl4xl7lbzWhmtwMsaojYJHD6zJqc9PC4SQ
2a7h7dKtW+/6yENdbSQgE2iIIu2MSCA3+Ty2ReB9ykK1FXDK7wdWIpIMzlGbIORH
aRBjVZLPvHwqwp6r2joP+abXCgjNLOtDybFdz4Bg7BHqL5e/wZI3I6bh9I6jhQz/
krBXeG8TcXtQLLhcLQgaCc7lmDVeU1yf8cQAlVeRYo8uuHZwlqFf0P5Uuyk1kKqy
WgI/jvD3x6rzJKqw8t35Kql9RN5fqduPlgz5fLl8e3FM/6pltNS9NUD+GEaOWwSj
gf4+LRCnkoZWuuXfKktK1e55chUlpmzQWauuWWhKkupXp2/6vv1SiXjR+Fml+MBh
VGYzRf882t6vJD35lK6g81t7361MQ9yTWGhlttrzsrgGq3YL7IilsodRoLbPOFBE
CWvhpSZImKVvc6+xL0LenDWvdHcovr6CvtmUOLvtt7IUXp1UTEYnwFPzgt9YqFMK
VJL1Ic72Sk/mu98sPplc53WWVJkPOCI5uyah3cCADnX0uSSop+trXg/10OZIlyLv
0SSP7eD4KCSvvcmucF1yEz0HhgwGFysaidak/V0vuGkre1u3LUrN8vax6DClhKCY
Dgb4Sy+ClfPBHv5bZB4mSuyd8k8DtOMCYrRDGpj+SLxLafotTzVgmkdtmXNlBWQc
y++zQYBu809C5aqGcoXLZevuh57ccnGJRg9zvfF589LFA5/x6ev6lk85HTHnUweI
EKwcK2XPxZIMH7OVcZNFCKO+ym9r/6w+pFaZDig5Iv/Coe5Mk0atMS+oNIVFmQCu
r4NvTYqDOr7vxNJGDhbUvaNOQv2JsFGYUkGgTEiad+rMA75Cos2ieJZBy9Ad8neh
hgFasJkMli4EvpAWj+KMyeeB+A2eLUTuBv8fhyvZpaqnXhHrqRP+XdklQAQpilvK
pgdqqWC6LeSQ1T7hUA9QNMZlWarAjP1ioZb21FMrVJh2RarpqEBYE/OfgmKJHxrp
zftFd8CEXW0DZOWIl0cbhYpx/q6SMNSC2fwZsvsBihOCGxv11gi5QrNuRb8+ta8l
z9ciWulET5YaBrEwiUxhOTINHrQ6pxhlNKwxleMlziBmg35z+4OwJv5MTdNzxv2C
nIhvxRZBNF6duu1+7ko8AKE5KOABJNigmk6P5pOXRtty902JDd/6AMf5DT6X/cAS
PdJc3qt088X5t/np/qqcZ490CAz1AV0pStY7NuNkpxk0fCeM/RwBVrFstJMS3H/6
3+A7z8ReGQwnYnXiQnQbTKxpQ+44+KCeNzpTQ6ygQ+m30V71JV7BT8IWLW9L/WZQ
7lXOZAcPtagUKfs589v6lUhelBLMDZrIVIsR+HkL5tvHbMdAWwnd6GsyQAJ8Z7UV
dOjenOBRm7MmZYdJef0xCUZboAaYJZX9LEWtlXJaEk4SxrPxKx3owxq6JzMzHIYl
uFbs3N0Fvme60m+bK1vFzVJ2abci4tamZ4trNWv1tVz4pmvHaS6HnqquJkHcOuuf
m96rURv68rTeP514jwYSEdKALB3Qj51+gY1S6UDO/ueo71AQN2DwEqL+ZZyqy+up
GDvVd5NYXHwi3dq7AOXs7PzM3sAe0+ABk4as93XVBWtFHFXbFUx62cm2C7PWfm7o
rv/dm7fVGLc43Srd2WRQE1xDN/5YClyJ5Aq6s2FBBFy8fO/pBamn8npOZtRhpCnP
C5bRxMUGy2q0qgWXEXWLUwxv8ioKisn2bz4nTFq0qwF6TxU5x3giHoVCE/QoV4Jj
0CTcnu+nWpVeva0AOc6Vewsy3VI/OSr2tT68K2NdFH2wih5Gc0b3gPMtEE8+c8lk
wZLbObPdYOj9y+yjAw+qyc242iye6eEyH1FuT9/m8HIGVogwzELfXWe3G4PWRccW
H9BqRIjOaHi/87gBFUHtUj75DRKfKYGVu3z6vS+fhb4jwHpbN5mlOcdC/8G4aXa5
ApUfmc0qyX/I6iTPE7IeLMXr6TOskaMYk6hreRN7i/6eJEsA/Ym/zGgkjsix0ys5
A3ytUSmbI3GekEYRAqUOUe7o5Km/z5jit6qI5tbtH3SCjd5diweYpyN51Zgk3tu7
g4DQzROOewqrKIGjjDW0zc4FhGJ1JsjH1p4Ncg+F610rG0lh9VIh4uIYYiDZ6NU0
1QLkx00hfOUaoxmGMCpTrCiYD116qcn2AlJOILfLA8G6HL6e7C/tF7osjUj1JI/T
83mocjYetm5XVKZSRBvHbQDPwuMyCHIZ/jbyLuwXAnZNkGEDuiJOIKoZqyV30S3v
m2qWBrFVcVNno0fx+FyMJKEzKHJJavzCjEWfCjsDv88JEsW8uvDuIv/jq8yLYoEe
BXGyRhyEgc8v++CY2bx3Caurp/lYC+xCwgPKY+smjv2a0AgGwfH3SHje3oSuZMfb
T2IPMdLC8TLxftAKCOLuhH/vc4BVQpGQVXAdW/U00eSI2up6dq+1jUoRbgqVEZDy
kHK+/5RU2euu82MQL/lKkJe89bYBZ7t8JOK8vYN1QSefw4e2j8DZcwa5JvXSqEZ6
r+i3V011KwhRevlmLp1FN5cyatGLF1wyolKwTDaolemME8hIOQQwLmtjD+t82usQ
ygAPLQ12mN9wBrsGvRz9PvpBX4ME6dZ7eFtDtpPBbu9kSkUEFssmOZoIlJYbgZg6
xAA6bzhtjuEHHVtwAnoRWVNmawlEkiBtW0IWUnvGpaHm7ptpkrFs4O0piSezf1iX
0IqQ6d7UHbB1F3cNvuf8W68GePyd7dUEQB1JP9N753zpw15poSrTAq0qWyRxH2rm
ug3yI86GplZJaYJ6Cs1Qad/Rk4S8Mc/oP0wgiJPD3lW8nNVXS8lLACP7MZUjES9K
zU1UIPeli5WpKHnQmugqgH5mpmt7Er4KnRfEkgUBmkteA49cuFjpm2uKrwO/hK4j
Nes/ejFSRbClAnxBl2vEqmWJmmosYom/1s1GlkTh8vZJ7UJ6KJ8bcXgp0BD+mNqW
/YqDBXZPZF/GUU+IEAJKHeCHYhuIdd6slpTA+le36fEwKueWLb1Wyvkieavb0Bm5
5GzgnvMaHK0luP2+1Ly3PtNmLCx6QjFubaMfYimBcspUOADek6J/Xmy26KuFvUam
KhkuaGtvRqyYn7Khxsh/ynI7Kb5cARZU5sR3vzJAIjQblCBQy+DDV2yU5hQzSjyO
hIVi2EXs9UgpUScNkRWBUFiKl0bZj6WTmkTuQn1SgS5eczhLIP7Y62lcm7dZd4X7
kEF99aRIfDh2BUmbtbAyd4NxEtJ61El6ZcOsTT14tV9v6tl1Ne+gbutH8rKG7vQn
q4CUe5A0HPtkPgrsiQh9i8iG/MVtVQQBq2Rp/87dblW3+2gA03kSsxncsoBIEne0
Ac+ehlUMrzmpq7ffH1JZTdW9xqRQ7HOCcfYiwWPalZdX67pp8EjcYmx2Zn8Bql8D
SZosCLG1xIXup/N1qYnsVOudp5pgDvN/qmz4sxYkW4/H+5WOW0sfrs9eSV206B91
9VbI0VxLagO/ESwI/HRvJ/3plTDOvLaMhyamnVBeuXkDOHbry0QK/F7q6yFLa54G
+z+RIx1JOSMkjZLNJnDxXZ5SscRlaxGjZSjInv7ad64GCiNB8GaIEBy6dcFepIDB
4WVxGFk7nkKFdhHCYpVKstyXl6COhhgU19Q3ptHlWToVB1pkvj8r1k9dhH865ytG
cQ5rz4KFT9dEN+zUA+BYITEhX+GxUpVvTCx+MsmPmSrDZbxOIMz02pMsfd6SZ8V0
8CubblyebQzqU4Rs4KlRa7EskU4hmIIa5gfJvOqMlzKP94b+2z6bjgdBCeriyfwz
ZnZxSWUJW+3zHpv1Fu4oOZma4ogdueIQxczn7rxSyrRdle6fOjCYJA9nrba6CViz
vq8F0xy/31nqvvEASmOL3/Bcf2cawiEQ4khROgy/BPsIwh/Llznl/0PCOQ1Kfu3S
g0ifX+8qWYngDYeq7TTc5PoYeWKMOlLX4VggBBJrmtlLU3BnoycEMQ1bz7mC+L2Y
+6QqedX898eniSieRRZuBAF6dIPAQSpF1jpxfIXncVhrXE+KrIZHSnnUpcM5A0Cj
lvjyb/Qo/REu1zwZBmgpOkPRA27lht8LP556sd+37R027i2co3aLtRLeK09okw6Z
B2jDGVkI/I1wNk3q2R82CJbSP7E2Jst27ieyxYTi7yZqnQ8rM5brBvjKS7xA6bPR
N85cxg0SYTol4BE3B7etGmyQltz/4yskHqnc6UMcD67Mniq28/M97ySR87hmGtxt
n3kLfK6nL0um6fLZQ1c7dRmUosGZnWHYsg6etGgkeP8TFgjwseh/sYJbq+56HkPT
HYkWJyzgh9w0okvcL7CvlLpWSBx+SbV9KbHAwwbPU7QprlvJehaHvhW/QzJaXGs2
k8Pn8gdg6PI8LKhmdVnNs/C7vFRibNrySbRHHtE+VORkpBEruVOMz4+NqkQPCUic
wM1BEBAn7CQRkQuTVrM33U79lUsONl9zwXsNvqVp+uqX4Z4S1K95y4GmO1/lnypH
mSdR9zXowzsJxIXPtkWTOtSczxJvVqgP9KCz45I5pRbjlf8qhcrzta43l8WyT6b7
10e6gV1BId4FKicjxfmAgmR3gzUQpIJ+Y7WxHzL6jMOGQ0t+1cNbVBLCwaB1SZ8w
EwX/JQ4jOdaGC164VPx/YKBrHfnxlS5aodGunJPEdO4xYU/3TG2+Crpx6/fwuITo
6qD9r8XZUcjWu1ojtfziDSAk9A5hwptZkagSrFPV6XW9oXY+sMUXm9xGVVfqRRIW
9cMznXNyO/e5XPm7YeQAQoXcv/9QYHxnMBprXNcq7FrZ+agwHRW/aV0wKCC4qSgq
+Ot5OS/U2gVlZqjk0tI+uu1e2IG6zGi3BvHLsLDX7PWY0ArbxkPFP8T/1q+B2ctx
vLJAUhbpksro/P9yjYZs+XhHWdb7luHk0/QA943tgXqBYewKXoBYeWne/OEAA/O6
Ew0OEkkD8ex/NPL2z2SmQKFagcsHg8jhA68uFninKM3vlhvZk23ayE90QWG7xrK0
mMpsenFr6M8xkhC07IFLs8p/i83OgKao19L2WWtOhuM6xgWaUQCH9ZpBi0i82C62
AiMXag825geFJMa7wuNZ0BfjA+2gczTE0N+8PhDFbZtkbqU9Fi4eEpdMKE77lpm4
mt5q9RSyr0dafg5FjmHZhjjZ1dBF2Xed4Yp5hrPKnfJPTm7MO1MXRVeG408j4h0/
F1eU7BxzoV9Bvw0TtroFl0gGS90Rtkp5YnIShZRdLQiPaGfyxuD5n0sFiou6fhBs
Gi0ru2SvR8MVQkU9rlXy41tb3Llr+bzj6f1l24TKSIQsZtCeHf+giqCD9nIDCkSP
BsRstqALMT3Kgt+wky8LTIecaBrQN1lyIOvnNt96d1WSpsNYA3j/LsBjzIYVJQ1k
gjX8TmwQzLPyjBFfbWIEUEtklpX95OQjXCIp1IVCx64HxCWgeLFTWCxopAl1HOHC
wbxkmN4QW8so5/hdh1zlHL5SP3gtLR3ziZWLMmTVlSobTe5lpfj7HXvzfmFaihTf
Cb9BZf1hrrjazaGv+AXpJSI84S62AgVXDOupHVcJow86ZBeiRSDuv7IAKq3yNezG
nhXswc0iFsFyKwZovZfAQxWyUwS84u5WfTj8w/umgXr1k2Z0N0GJDoNsJeD/ta54
VCFUx/UFUpR6SRg+nOGSYdrs4BGOZNjfdIKpCQh2UfHT8Reu5cG5o2WPFoK62F01
3wCCfu+isY/eSQg8Rqhl1Td92rN4OuHoRXJEX+Ef4sNkFyvHXy+jfcqVJb5H8od0
D2eoq6Rvo4/1tcDl6OJA0lxyaSwF3tgrqsu1mKipGXXh8u/Wn+OLPdeq91LXDh3H
RANJWRhDecdR6naBZBcp1jS57a0HkQ8/oT/4mGOxbvE1tNYF9m5JwCcDxALJ55bF
5Oa1ghWWQJY6vhvYwl1Ij4+d3n53p4nwn84scJAQpp5hldFBmcNLZQxA3jvE1KPS
eyCzuhd5qUfZi7xH+EOXeRWJo+dgObnGP1bqfsJkOfEcFWF1Epr+l9fND7snrw52
ke5e6xNIwOqza9G9W9fcHlK7UOKHrCBm4rddSrlzSwVgoEI5CP9uH99y3x7lvKAJ
ezzJYQQJYR6j056K4Q7ZTvhBf+Z8tXU33vkp/3R3fq0mxFNQDF0dkMxmPRHUODVW
3zJu4hjA2qGO4qbfzpbXP+G6EofBO8hmMbAIvgcTlyASs1dLSPuotq0x1zmrGMSl
tOtKDYTYoPkXPcQqPPBo8xqDG6hk7JMRC55cyrVqann8B5fx1cvqIg2XjvMPJZ8m
M/2Il12VDrJGo1rUXQwjO9OESbfdxOC4/amaMLj6Y5Xie6fZdIpaNcMVLAWgas16
BawzezRexhCpmoOqr07QjVs08f2cFOjdeUY+XdFjzZ4dBQs8elEalQeFfHzehwYT
8lTcUlgbyKf3G60WxzPYZHTwkjYf9id9cbqKyYs5WCoXGgjtF931/Hf+Wg5P1h54
adt5zGkSxL+D1gTlHCs+zQ==
`protect END_PROTECTED
