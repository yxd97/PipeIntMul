`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4evNw6urikEiJth9FyiTZjpKD2TngNnMfjvHcP97WphCO4ecYMCd8HjJeTnJ119s
fvbGm6DoN+n5ggaojzqpnPTw2ccyWpf/ztbWpBhivJYUsSusWv2gODaScL9/BFFJ
RRXDFJn20Ag1pHZMZofg/GMErNZBNqDFccxfdytKxim750586a39oi18EYwaFGke
+NZFOGhF42igsxdaEfFB1fpeRu+YZSF62t88g326zswZinWeEidZ6gRMAOM0xbW7
8yL2JbsGZbK0BKzQEDMLJ8kDH2NrV2wRSR28iASwpe6SFcXNvvF4RagppQIHXR5g
QXcJQB2NiHHzVsQrZQhDzxy1N7QiaSQ6YdHJHuWsKbgzNGJ5rW32VVxEZbylRrVc
bkDXQW+Vck5cBq2Nf1+dky0TdNYzgohYJWETNBXfenQb/dFFNsbPE4zRoWcz/nuZ
UWGZ708YR+EHbRGsoC3hhe5+vbvxnux43RSqcougWYjcuQYIi6xzSQBIN6Un4waU
OwLoAW9VXHLTJOH5g+86/t023nfEhIQ8hFQ/AIcipnOatRaN927eQ9ZT6I2IEywJ
RHqmyMY58m/UcUV18Bpxag/i51FiL4E/8XLIHFxLFwEq8PhSwz1piGze+ROVMxt6
JbTmAMUToL7l25P2BscumTp5zpN+xCxTw6B5QeGnAB6nP8yLGn13s7YN41nllnFw
zz1dfTZ8iqa1IgOppHvCvZp8gxPEjz8K5iNkwEw1gxTYTx7Q/SmpRc9bLCodEL56
nbyiwdD5KC1NhLqJcBFkwJbFHO7V63QV6SNBSOOcr+M+EPZECEip9N9shUuweiyC
HF5pg2fjFWeTAU5cENmTaveSOGqbHPq/iQpOl02HK0f3L85UDIJUspLqvsp7aCuk
aPCapM9GjO+cgV9QTgLl8xqd9ojmDPT/VmVA6XLnRyRPURFx+Tant4kWfs9dcWvU
oaEt6IrUz2lQmTsxURO8ST5nAw/mGcw1KCAydiiVh5eskCDv+jc6gICPmh7j6d8N
`protect END_PROTECTED
