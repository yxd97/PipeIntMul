`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qp4eV9Fi2PGThJ7kteYL6fnDsxGS5mZlpSdvQ0RGeviDKkNywQ6sHKLT0+3UZACj
UcthkEOMFsBuFWV1ibzKqSKG+WT9ooSHxbFVpgdQifTUE1B7GWQikTvt+ew+WP+1
PymoAKCQ4yVvJg7fvkEttSU/CWBVqPOl5hFaDcatUFefiegG9XDmh+sMqBxeheXx
I+5RPxr3meXOOY+1IL9iVskOfbsWreXcX7bdjwMN0qtBtjLZxGK2FFQ3g3Ii1eEV
JGk1nDHtSXdvzASgAm4/5AHlnMVuLzrdZnRsRjLlsmzaQ54kMvEH1Kzn6BlR2pvY
3TWVLe13EPqv3BFJGuGdlSHijsqXJYzYg747lEsaYig=
`protect END_PROTECTED
