`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P83w0nFbXlkTUnVF5bKzR81f7qeP9ZETX+4acmsJUWWQ19YEAhnCsK+8PfjZBDVB
Dd1LXd0VUcY3P4uKgVl8QYp410Rj4j67niUbx1REE+LG7XMPWo6FVA3up7O0u2LA
Dr9Re2ywl/m18XIrEXjWEc4g2WcMvdO/FFvZvC3G9xT6VQLURyKMwN/OY79crJ0O
OQ48IeW2vfTZW0+Gijodic4lj52ZZbIO5U5+FMgaS2HosMHz/5H2Ldw7kTkylYZy
0UYpAabYPhi4V5cZpU0bcJuMRJzohCyGM+tZGCWJUV4BpYCvHW5jsN/f63HpM2Wi
pxMeyLYLxs1CrmdZJ5v7Aw==
`protect END_PROTECTED
