`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuEnRuq3gCOhZ3CTsjjiiq8ntZskyDPoB05T7OokK95qBg3c7ndyKs1rXiLM2mz/
jyxp593PKptYrrNC+WIgkUWA+rO1UwlIMMBfG8qtzoKZkp/BXOuY0ZXlQtlS2IlT
J1dIkDZdQzCXpEWmoUVQ8VrVRNwW16faaKgcEDs33KXnBXD86BtUbgYQgZmEoaNh
DKpD3YsFskErr1YFOLoyEtRREgqbi9/XIJyjZ4sgdYwqO4Uqx5dZ/w+Nedr6tkoa
3pufYxN9KslA+/X9noAYp4FIn1zmFWlBHaHvrJePNJnJ5C94RHM3J26TxMnRoCzO
sRmFAb8YcalxmqNlHQ4csX6T1l6tIg+QsiJsi1U3YasVzk2fy+HD+nQNFU9e7ewt
795CTnpK3X93atYkNaKnGLbMrWqNRPm9UCupTIOYbs1+yrL0zh/9fa7P8085fytC
LdiDPiZS0Rr2DwsMNPn7ywgYeVZ6cy+no6rJdlaxsPpE2/jPViJJ6KiR+9G/SH/N
L1ucQY7+EpJpbt2gfUocB2rimrjM9AU+0HeoGn75DuWsvZTmF4QRbPkzW+2vambZ
+qG9/VlysWt+XSluCtfEWYN0W4ahOqrqS75JVaZcNLW+m8trbb/4LI/5c0va3UAL
C9GbtIqj/hiNuGvp/xDmJevAnVU/jdfIT5+THk06JkPCChFBRAc+tcCjB0W7T5Yg
iGqDqNVrpulgj78XYjuJUKyVAu4BiztAXYcA60L7uDabcv6oS9PWux6Jy2B5VQGB
isfR2R0cLiq5WJRMjImjTv3lXKi5HQQ6ixZHdKYQSRUpYLFGNPW3CqDw0VZ42Yax
g6UXgSstyvndn7iAE1lHCT7xVuWNn3dTErJNjBNhk9Ru+Xi/a/O/KpwP4EYxwEQC
mHDUK2rDybBurTE/JIYPwgJHQGsv5FEgKfbDv8ptU55T7hJBsPegad9TCE24Ln9S
ATZT2tLG1E1SazmskEe+BBXCgPPLX8kB47lRBRfX0Ne+VqoZgjnRbA234ZSGO4JH
9p6il1LhN8hecc9DtGVEjuq/8eUnhuczdpJTnsQ6CTWNtbG5JWMcw2Oe39KiRrl4
bsZndtKzM1qj6BnHwjj3S0tLbeBJvgmC2tILNdX6yferhCr8mmi25BDaTiZwbWJW
oN9kpMibzOVA3TkTcPwIwemzPIBLXpvCqMiwLAoGTCS1HVtKXjSuW8jTGmHDcW9u
PL7jKjH9p4F7t+TWZGxAryH5v3ZBBCcGHXnoARz8ccFK7cK4FtzTGDmCxBANV8vr
JEGEzn6pwW04SpLKi4qIIm4zUzIg64UUgP6TFcn0lijN2TIcRKj/YTcB7i87PNUQ
luCcrzAXkDKKTTZiNzCBIAzUCZKbUtYPgYmpwUTgmSR1pl1a/79OwHpNJJelSoPk
pMjFMdmqHSt76oRPmFxual+A1ZbbrRUTU6atSMdhFZAtYHgnclpyZBNv5NAa8op+
zfFBaVwqJTIkZlBj5stVw2MmZPesox9Y4nStT79KwiOhSIHxjBT2ZJbvtTBe9sdG
/s/I6cozsc+F8vCT7T5ZRv3dSWAGJ5eKfb0lIPmRypmuFE8+JvRB29aNkWbAqwni
aecsRvs5bFTbhNu/Z0iv70AamTE55Dw0u4S6dQePVKrqar+lNH/UOWyY1v1j25EQ
4wqnvG7avZduxSmUT5MKTedVG+Ps3yKQ+kFbQDNZDYZPJEPk5C9Amq/L07vWhvQm
uXSvpiNElfVWAS56h/ohUSS2fF380qvmveyAE4KKt6MRF233Y+tb0xUNEPHh35Gb
0SAXV7xX5yLaNbHTTmUSyKdjr2w12uTxFZ5adPEmQZIXEtTDUaiCBhQJIMqSDjyW
qzx3sJIz2gkw9MCR/FH0uhEllEImnrUN979WYyZvZaV47iP2kldIlqulfkFkPHdT
uDmc/5J3gcJma1u5yZeelUo5xegzgA5u54jq58yIhHHLKWMzeUcWksCtdvd8YJ/z
CcM7pjGrj0/oMaC8TzYpGXfiNy/ScDTbuGqerainxe1TaXhUVe+DHWyMkmsc4LBh
+Mv+t37pbm7Mylh2ZKCLhOiOPBDa31dy1FT/99fyOa/FkFlmWmCrOzm1gC9NohVP
3MU7n6zwV8LjtMQHJ5awCpIPrlFSuTK0hjgI7pLEXcb43CQS/PG4NvBOstfsCQ3s
LkUCCNKgOZCafrlrlop6O21+U1pVMbLZwKQkl4rD3wQb+ySsaK8UoP2p7Tiu3we6
eLpLtXhUM+bFSHVwKfgJwqEIeRnTHi7cXXGIcBpp2sW5kXmsR7yZJkh3H3RFUGmZ
//MmeqFg5Wn1gcU3qPYnUdWFUuIZ7msO4wGcfaxqOmrT6M+RO4+7U2oqDlu1+9y+
iX4pU3YVEgMef5efVzqygU3T6E07tkGoW+PwRmYaxGQx/WbQphFvy8qpbb1gYVjk
IEXgntHdIIfaGxm3g/3efsj/jsH8EMQQB/ZJ3B7CZDskShSmWcZ7bEgz8b2KgtNl
c/i/lh9HRwAYVyIDB9HgkK2wI+b+QvQjXOM4NyqnGvjtEtW9q/mIT/vohqtho/Ls
MXxFlvAWilXILCiDhnRc/kjApsvDOHnjkPUJjSIiO+N0g7pNtrh577kxyZOg7qbb
Wb0DOoIWmByXmsYi3Vy0V7stYTb+XXOh6VASJKtNyPMP4Q/bfECdL6VHijkcpwvs
kHkq78YIod31/pP/TLXch1HwzI5GY4HnNuzgrTk3VerprqlSjD2TvfEim74veQ3y
1w9pI6DiNPLUzqdqM7pgIrLcNBqoJSE2rkYlurHuSgy3tvAo6NK9JrGHmNtkzNC4
3zmuixaQws0PBipKcjukA6KhjnJaaxwBMtjD8I91F+q8Dm0uyPxDTFePLdh+3SfX
a2VXhkszLD/3VtZwbjogwoSCeTdoUp/7S1ONlWgLnnzJ00876GJ5ZnzSs8bmVYj+
04SAXzEVWRaKvkDGKHxF+/q+U4ZlYgLtPBP8chZQ0QNeMUWnhRX3qD1PJImvBm+Z
U1Gicy/CdW5jhJpBTuyle+5bLxno4BLRq/xjGcz0VN1+jKgZbwggUgvTpifra+30
PveSF3eWdCZsPzn/ib9ge0/BFp3abHdzqdu6afUyDYw5eVKnkNAKhMiT9zufVUFe
6Q8RobQGbhL1Eu18j1WaojWHfW+7XGPuyOgY+7Qkxn3Ismi7oVQ/S9EX5fxm050P
`protect END_PROTECTED
