`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehDIE08EVVKqmNAKK80LXtJDDPJNuZk6iFBasF+b1oZANAjZqE8jDBoAy5PdQ20U
sXa8MfNELgrR21QZe6eQZFWplN+IY8yAaVTB0YGP85Xtthb/QscFxlQfN+iXbWM5
Kt74CvPgzJwbrFn1Ct11VlrjAdojukEoInZWcc2aSY65dYNyCKQuq4buwnkW1oGa
vhsoy+cG2q6LbY7eCJAzACtwmt5nZle+k/WVm0dcKDDuAsfV/1XYBMAqsDslbBSR
pT1blk6+Tlonl6iJanDf10as4Vppr78x4+dQsRzI8+sKxDw73p+pntHGPk27osL1
bwlF7D+n38+DAdFYYB+DvncSlKab5oiAvJ/PNYNO0N0yMrkSvAT4bfeoiansbMr8
Qlbogflq8kCAC3nk7r+dAhckeRG4XMOnVNCDffBe8LU=
`protect END_PROTECTED
