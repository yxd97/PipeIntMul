`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ox+y6yHZqJD132NO50pZg/vzgUQxCGacFgGn/gvMmkZEuO4lZSAtIfkLUmNiiR+f
Xlehsbkm1u92HcPjp26a/kRia4pY8phGt1oQPpW9vPHe/7+LT5d9cELpdO/Ajq55
aoTvWHPmpbCbBV8EWfIYJS96hsFoPlJz1FozoZotvZr0rMzcepSeo7oVg9JIOcC5
oH5xRyQrjUFCSBniKPHA5gWFtpHY7t+EY2IwjaGUQBKbj8uDhFPFURC88ntnflDc
U4S4S8V7nefJzivYNJnlio8sNBPdotCqYoOd/qeLkcrq90SJ3p7KcypbMc5k376n
x+29KuWorsYNEYIyJQmn5a7dLsgdFvi9gowcqTXzN9l8Z0I0r3gZn8oggKA2JoHS
gha+x9YqHMnWqnNMqxNlUG4gEN1ja3sx54m8veP0Ymcb4MOthCAJ9JHc13xL2FrS
T4HepzRKfPlkUIrmsG2nAwts19xLP1A7s3Oct0cocLIibOShu9KHAwiCCb13o37h
`protect END_PROTECTED
