`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1PYTmg9Gjabb27TJ5lGfxjaXe6UDUSUsxRLPgPyNsdfKI8qdzMYwK6DZh16kl8e5
wx8TkWTDXlddjhmr/jeDdk3ZHtG+BUb9zzyhmfZSVsyLOHVoTMlklNlwuUXY8bRc
pTsOzBhTtGVQyY+k1jwyAL0T25uDOQbtFKGkASpa1HJhW4Ugk4OAS0gZbVhMq6RU
zQOTY5dPQg1MX8fTFAcFCRzzcCDJUX9jE35JeGFcTzFJfwq36oOjjjJMyM8Sjy1b
6pHn5r99be98+92Wake/BLAhh6aPKFIaOYsHEMaQIgYaldu9RS8J99jwIUGMDlsm
pAuQ+fL2P6n2/Jav5E4jYtwYrN7ehwKVJ9z+em8pzO0TvnF4gFwv+nTG29Cc2LQJ
4F626cc5wg1UZQcNmDS+54shplx4wPAlWWr6z8kApjYZOTM1dsifYgjaYDIVcAU6
9f9nP+qdTWGDrWtJa4MFfovSfHXwDqh5ezRHS6CNFA7fsvlce4aLU+ik7+zKzCdM
`protect END_PROTECTED
