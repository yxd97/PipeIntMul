`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JvbI2V0vF7z0CWEjCg22Bb4TI0WBiS43D1l4EgSl0uklU9z3fv7NHc8u+Gbj8Dtc
dPVvCeqISEiFzAiZ/MnykBOs73wKc3bksq9BSNJysBMNC8XD9n2FW1g4sCaoITzV
H1n4wWnkERbL4aSdpg7zZalz1Uz9BGXh8o1RegCjsteePdmdrSlTbGr/WOJ5LW2C
FM2wpkHFYpgbRx7JYVHUo9wvvJA2HlX6slHB8vABPzda2Ic0V26pW0xVro9F4Rs0
lvwUp0wujZFTBinNBrlPTWfllSaffk/liHNiEA4Ypasd08XG4bHhq6mK0C8VL4y6
aP0GuKv98r/wQxHZn3VCGH4BylKckLcPlf/MqnK4wrctBbQ2VQ1IMJcXwBxYtHUa
v7L44RN+LwVrK1LraI7puUKuf0AqqLC14vMZFsoKKoxDzwPT1JhPLnQnS3sTV3YC
iUq3Nx0kEeJohgS+XxCk1AtGykAYWPtgGggp++D2ek27VthqPfP6WfcI1AumnH81
2D9PfIHVYFekz7uKwVQBOjEGCaxvf7G9zzI8sXIJAr5BBhGykdStmDYiMeLI301B
UGTKkHpurGXc7UaQE+z10MA5Cq3QwI75MlnOIEugMDrjEjeUGXX2H15LVG9TZ9vV
o76I1VZYvd2RGo+u/y4QtUjuU/2FisymaYHNrH+BmvHbb3rJlRo3HEbSw3jqr9r0
`protect END_PROTECTED
