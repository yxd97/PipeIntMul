`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ms/PxPrA+FvE7JRUwqaEImAvw/LGAzD0YvF08i+yF6mHu2C4+IHclWvlxchclTt
kkt1GQ1RYUYDrJxtns0h7FGlhOPKNfESc0i9hj4mHfLI84rNepK2M2HjEXyKKmdA
Y58fFD4h9Fw0PCyZ8OUgxkfS9nUiqPpWrGZqrds/c/u0Pv41Cdd3LV/Pq6zdTRM+
t9AUn76UHn7u0/aOHw6iwqEkDj8CDH29ilfXl8ht4QFWJsh9JrCtT/6nT8+J6GsT
pIKdyDfnCkIhtZC0jtJk6VcOJIIMEQM9iSvCopo9Lo8oqKtk5RwvIa66YkdyeoDQ
AxMnUvbpD8sIWwOLI6aD88gaKMjYu+hbtm7sPzjouq8wn3gkcgV/cm49JwUnwtoz
X/NdRr7niHZV3fop/SQ0f0kYv4BjmKOgkUWFon+R/JAwmZR4poePmL9+Lx9Hyhsj
tsdhQuWx2QDrS9pzNvr01I/U4UR+vNs7ZanxL9Ga78wSOlmRDs1Q9SgiCKX+YaGT
WJpDRWJXiqZhHXABsltlkjHW5q7pUyZ8yWLAi7gHM1VuLEZ8agHFyaNEskMFIwau
fN92Skn2tM45dkDW9/JeCo2h2vzJLQ0t6HcQPy5MoXg=
`protect END_PROTECTED
