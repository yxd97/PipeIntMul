`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cd1TEmSMRNx8an945O1fzOuoDk6cUgdxoYw51IjDXP9YPyAqMEsqkC82PNAgnYOz
9fzAV6jowOkKnOhX+EHZTl+Zh8AGQMJ1EhfYpOFr+ggh7ELtHlfBqtgVdXgBnjr9
uZ67lthRHlpQcBFm4Aj0KvNtQe+1MjeDLyr2dKC/LzJD08jOpUZqF12lGm/lrhal
qUc2syu80D6dStrQW8ye4m1CbuFS+dKExG7ihg6SNWXMqqCKJSEQ4PPLfvQxeGLh
dm29XchZ/wj1swypPeZU6NCPlmf7V735N/lTR9WokEd8iRwCoffaTOogbXE5Rse0
HOi58qV41UPBp8IUZfBxVBwRbndu/TT9d81KCgdzindezkI1tOkrVtFdyp+fSKyU
A49jdTwdl0KUXj+FrGJUA6OvGG32T79P3X4YprHMgz5+toUIQP5Ci9r+Irika1A2
za+ZIW3UTJLLQEAGvaFfYt8cAA+bncTYVBAYW0xkwFSqzdEBVKR5jYImwWRkEp0N
A4Qr+JC3W26ksIvIbpzZe/eOETO3UuZ8pcsjIun3bSyJZlViSpSFqU+W91umJePa
YOa7vl/UFSAyckBMYYyobg==
`protect END_PROTECTED
