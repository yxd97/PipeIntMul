`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxyCh++EKWFt1K2mfjNQyKVwx6XJOl3lsx+OB02CyYAU7k/g50fxgXootfrmEWOK
O2Mon5gJ+poqpavYcG4bzWJNg2/wyJpG88PzJmFARP1GisX/sOXuIpcKayIqRM4M
UTmGEoq260F0UVmnaEUfGuQ5QJpo867b3HaJtYahnNBYdg0adHHa7ABPmKykjc4b
W7Riw3GYiYbXRv7nA9RZS0vpAPw+I/4/oVnRPDnQGthHyycJQd2lgL7mxmlfFepy
sAgTGclfrbk2D9wv7r90OC2koeX0SDIin53SDVDRv0Z1XXEvBCY2lqu8cPb1NQ2N
yWVYn8cEVSlCviw1x5Mu7Zlkc40W3cZlyQOc3Kue6uVWoYiUIpk91ExW4xF7Iw0A
`protect END_PROTECTED
