`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yqea6D7QVJIJGJzzSlAbi1beHJw5Hd8/FgRCs+v92jhyTvEHWMI6YtAHeN88m1f5
DiUbpvmWPR11s9UvkItnpYDMitpUES6WVF9jajcuRmoHGA3JoTPClNAlCoGqdLrk
j2VkwPWOrYSJ2vz9UbLf83F5KThsdX974CI33bnLZTA1is+PxF1M4i40qJ3whyGL
YyyPTVbEUUjOPGXVO/9UoiBRh1gB+LI8Xq2kl3CgtOz58nakbyKj1ztYy1lzEB5K
+NXWkOmAqFcU9d5uKlJcaQ==
`protect END_PROTECTED
