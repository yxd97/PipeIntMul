`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cIP32v1P1O/DkL0iB6AyxnEYpZrttWUWKJneYKFTEzBcvHda/FGcHrD0UP20/H/R
DvxCzHozHAXaRanE+xnBFdE9yFRhzmNKI+dSOFuUZtB1Z2HXfogoNTIDr7DyRpVq
1g4Q6kPNIFaHge9xBlWCR91LUXzGPf9o0EEs0pSG7BiMALwz/1EZPNCJfG/WInVu
sgB82PQaFvLQ1mEO24VRqy2wLGo7PO6ZNy34jpRv6t2IVAu9IGVftFVHSNb0kbH6
1OMyZrzJuyV7chd/FJllXfto6xGN1kX/PgXbsXXiLsRYx29+moBIUM5Chl533eqf
OVxwlOpFfUZie+evHWWfHv9lscpsGH314y63OSEn/X9CWDuYMR36X/T3N0x5Z+vH
3gAchhDGrfAn37CnzJyB+3+518qqyEIBQdg2bi7+Rms+k19majy26ydEcMdETMu+
wewyLWjMy4PwrN+WbyLBHArj9jwG1F8JUIzadlX21daYPTt8i5v1pky1+jO8Le3B
H1dydIbXZogiSpPQeMFpoiwwbN6N/fVNSyU37VN0wjFjbkXZ2vcAAzo93vtD3QK/
V0BqS5FqpbT8saNpaNt+bOJ96XFe/l6Z/cZ8+z72ZOzfKYKkisBmHjebBikb8rpC
ChoxNhGdFLhYwcNo2G4ewsMR+mvFq5agbttBNz/fGeT+pJZU/6Psyugx1gki5peV
23ylFEcpQytP5IX7QG4fUarQbLjJcdNcTc1Y6wlNePe0Iq6phEtB8T2K3sW1MHEK
JPbb0csDXGNmwYgUJYNt6KDf/G09EXUYrFtMP79hGZZDEbmii/VPIr6eLAaYU8XZ
Uly+rLuk8xpFyfM7105Mja8cGw3HQJ0feXaKWbTAaLqRLWbv/fRkmFfSg06ToU6f
z6IjTrL7pzueNA9MzlXpWtU/IBsJocgO++3WHUbZedVIibei3HnBtFvt4MwY43oa
htfD+dLavkXSbx8YSNCCsEjAxxXVs6EFt5Mn28a4CCTNM0gUnNkhf2+O2xcLf9vF
gcwBY9HxltHUQXO/5d0B9x2/rJ7aWz1JIVdEANTK5UYRDVQmrub6cDdSjGvd/GgN
n96mrqYMhkQ9XUFvZDWwhl9KJGQ+0XJvVBEIBTyxtqzUQzk1KRBpFXEZIVs2lTdp
zrT8ZHWVRuhnqW0KKWi3UZk9v7yEkcr1SvL1TDnOziY7t9qDPGzU0r0VIV5nIC1C
sMZ3lTbeq1nuo4lYqHrgmyKnI5lIQrd1WdMGPe6ld0IG0t7EvA+lj3cDEX5IdWnV
Qp3Cun8vNslHq5xBIPU6r6G7RDlaFuva+QOEODXlakp9z8BjHJ1t8gAlymGIJGNj
AIIPO13UXgggHMoCQbMrV18MS7/OV2f+M6nbEi4KkanizHNr9UmjBLFdc3WQlfkY
ioAf6JOhSd6wyM5se1UeeRpiArFbaVyqXZyMLEm6mXl8H6UF3JoVNuB+7unHrV+/
50QxuZPAc5ER2gS170iHSGerqxQUaGQ0/NqSzGeRA/oVCyAVoGbuitsUQU55Tp7I
FdksPyN7fPiAQLMzR2D7Y5tN0IM34CNzwGrcQuZX/1bxthK10lGwUZ06MHAwuaw7
eK3XJKGKK3RI0LVffJvu3X8/dZzNaHhcNZWvcB8lDX9f5nDQr7YkDVTh5LtEr/rN
KksXXxP+HStTAIJfAuN6WO8CgC77Ae2JX83frBrE2Z+VdrgTzrArdEKp3pOteWLn
TpXAShtMkrDFoJ/f0dk1z78bo+NvFvWCFyIYxE6inzZ+1UvlNBXEzGzTkARLtici
oiFfbbfqNqM/+UYVkfQWU8WzwvnlvBfWiuKs3UCbTgMzeYxpVMlr1cu0b0OAAWFC
oTzKJ/1F3tU6/DDD7XyTlF3bLqwAf9/cdD6/DHdUjpr+BSFE9cc4evfNTXG2EHbi
1EdUNycpfXshqoJ7Kbyn1TWUMeAmJY2BO5HW+s3ZsOURCnvojeuCuSfrgJ7F98FN
4vflWeuA2HBnjRuIXUMBxlfJgJHU45N29Xxviq/jUygY1G3rbT8+r/Ias5QSMu5o
ob+L9UBVHV1drgTb8dlNZWJ3ZPGexesRju1f3bJM9YBs6Evs35euYaHTyg4KbO+Y
QAJwCBoHDEcu3BJ/ZfRcGmfNeOTgOVr8NXIJ8VCKdR8EwHSleq2chVEBP5dIc03M
5SYVvS3MZ8//oLii6q/PblXTTqjFTspBfVMTwZXg5K4YZHGWLhI1a57mT/F0cul1
6vPs+/u3ksEEXd+ntspbvQlz2rFJbtTpr9853+aEvnOG46dhPf0DxnJaOUBi1j7E
IZhllvHuA1diVVyRVHde16JK+LtpL+HqKTWPwBvrvtqRu0XnE0JnmrUjo3E78cKU
LxbwPOsZaB2M0y64yIXdU/3RAyTaOzvn4y4dQ5Hz/5DFI1wELJBFp6cVOLxrOMof
ES5YFKiAETaWR2YBbBY5xflGV7jCyqe1ms8afPAN8Tew7W0bZEU6EH6jtfn8McMk
J+tjKp6mnpr3oTL85vVqXFnjgeUmGSPh35cz8Bvz2HrhGtwyvfnAUafhA5gI4VpT
s1XYvv6fkYPOeSM71A7tIRlCcmMhUN0gicX9E/Kg8emVw55eosYeOcINFJRVGgYg
wRigFWYN1kKWIvektmsSdts0edpa973Bkuk0Y2hRR5l2FsFcBNUoIoneexVpwLyE
icgk0LEt+0IjBGkM6RAX2IeRS6UL8oStzKmettO2wa93XNz82H2rpdjC85tLvLzl
q42jtCKgvAWVqrDz+Xk0n2rt/qoBuCG/SSOZCRnO9FlX3BW5O1oG5s/0lqGEvf3L
vkVaViH8h9tCbU3tqjEZVQWcb00sYkCyOq1lQLZHiKj54q4FcjJi8jZ5eoWN5BOU
M6eA2UEaupEspVm9uNZtPoLXP+ZhYCGdqYTtobe1k7UriyQTJysXbBXFByBaXvQ1
Z1oW7YaOOTLMpW22HenLoohOiDTT6Auu3Ip7iWYGjcrzER+EqjE8jd5DofL4HBbw
lfK5w4v7EbkEfqwq3NtuHw2QMNDEPk1kYXUgKUryJJu6Gh5eBNdsspLrXs0gFZ4U
Yx+r2gCH3rf+yUECcK2GBq8VD3lZFxyi+ToP/DVWo7rivfA+Gd3nNVtRHP490ziT
JYh/pX9I92cz4QSVrC5lY6ExLe8Z5va8SYUoOPj7kvDVSCHWzwL8+nga3AgCucd6
Rgi4u4gvT6mDzgNlAiLuFiZkQj5c9/oj96ZVT/waYZRjCIaAmNMpLDTBU8jGJitl
ha8+4jJ6GKkcIwYFPKUoq3Yix9pCTDWArnOnr3ejwEQOtKIuBbeNhh5nwPbGXPCE
GvsyQsMa8wG6KmNGzabJ5uPd9BxcxkcphKThwo7uKh/74n/OOv0HLXxHgyP9jhi4
TGRqIwJDOTIuza+UjG9p25KbA0Ui0frIcicQft4+C8jw7+TeZoUqPPUaPnArmv4p
P8kstixHYDE+RR62aA5VFXjoPBRFyPfZuXtKX1c2T0gUQbe+N5CBfpdgLgjP7xTK
5/O8dHyrJjxw2qWtTOGXCeKrQPXQXIIMYoep30EZVRbcaNYxWy24hCrhSWwaIBX1
2pW38E5lLDut4b/SYLf/csB1YzCSFAn/I+bPVH+cc3Xy0z5xTp/zqlNxUnZ+BK7E
XgY5rIiflg+Yry6My8xNYL0dBVzP0dzmaO5xSY5ont76mw2nrW8k2k1LRhIaKlrw
nHHz0gm5HNeILUb2pm+GBJp9CJY6T1o18dqV53mqASawqjVRP0KxEM6LYu/wXnnW
WHV+6PRmqoXdg4vwJwoP6ua6UCV+4V7Q2/UeuvBJaCPnY5RA+ff9/AQu6lOTy21e
iVhvkAtQ4ZIkL5ECVPaskJJ7LGalRAXLsIVS2dL/AmcQo9NXFWeLn06T8QQLrw/i
7Tva+oZzgJUcYDK7KJ+zC82Y8Xnk1WuOdY+xXhWNWjZJbv3/gguK+jrJgHDJSbNe
8GuORigRCUGOBrT5vp55fHeLkHK8uQvvbir84ER0F6CbTTRQhZ94yagMAFNvsAtT
HA18qasn9JnjTLif8pPWCGdVs2pEAUx7D6ZMwKowT5NZX3qby6xH637SbXim+pnF
Bj9NKB6mvsfZxkRuBdZogzu7xVyeaTbiKeorOnflE74P9B1+ibNSzEYqtFARgUrB
TsftrHM7HzGWSXgxBSwqVVmz8h218Aub/LXqtCuJoYqD7sS6nVKDGDyCBDfed6Qt
dSPsG7wbj5amN9CNcvZsmstd4oln2CJlsIRM7MgFYWEi34hD5SrTkSvLSV3Oh9Y/
6QNWMPcycfL1O/onAZQMYjg+4dddBSEJnOMCnyfes/mAVwY0WKpeWS+WHRfnD0Er
LVKEMc1Umkjt+xfNL/16iXYdrUR+lSvNQIfomv5GcE+gfT0pJ9N9AQgukZ0XOCi/
a/Qt8p40sNXcdF7sUy1aBpTCMubJZHdiD9PxFbV8DNQ8oXh5RkSR8xY8Lfn4kkdA
CSoiUbdh06+M63L9TihkEslf1HI3VEeiLkI1BMTWvgLUn/To0xDxepLWD/4xZmHt
XYP5wv1vnz9pI8QNqovM6QDZXlW/nBHhXW/wmkNUgKPPWmHAtHKS/kaeUcXeiVKH
4VOIASj36V3HFG/1MXEBT+TDyVOsIRATMiX+xiuzrXKlABJXYaWysa+ev9MfI2XP
FVInnx1Fhx/MwLwmGB2KK9Z+I+dv0LG3HL430AbHJg9oUGWvXbl2VIEh9l/2l6FC
BM/kVIjchCiQmJUCX1rn2E8FE7c/2xFa3yQamWxp6LGsNQrFRcS/bJFCkGYwRTu9
09yxzIXptxOgiNe95MAAbP6hyimbMAZz2BFj0EGj2y66v/Ha+XST4p0ELjLBEmeU
gJqPj50sIAvbiZseWkrLpYVCqkBJI9og0anne1NWfV0c8JV8rMPcPpCbXW3F/7DI
jdqlfl7vl/yjnvunjOH9DHIgdr2fQ/6TOaKa8Y1fCXNm/tXAfmnsdvM0sRe6Rn50
zwaBZp0OZoKvWDugGkyzGtSp30MTIoIiQDzUAdzrzdHaiBidb8oKiJUNJRvlNWLt
phbDWbm9drbLilRcRu1/tNlW6JbNCSAhWoUQvi54qdwf0XqQgESonGeX2cDl2JtB
aubFxqXD/wpDQDSdh4Y14KFjiF+/+zdYK507jKhXaZY0/0ajVQp5dGDpFCQZQck7
g1T4ykMwjzl3LdHkY0ZNsyYtX47rdCafAz+rai8o78dD8teBXopQmWCIFqMs/vrL
fha5uUq4VadiGNGP8Tj/Ag9YmYAupoulhEHYmS4J4NzvXe8xJO85PBpSkdn+fKPO
hIgrENsd5JG07YmwLAUZgA3CNS8HSJ/TdYUSU/+KywL4Q/NFqFh+xKLCgZfITQfB
DB4Fxsm9cMKx76x8fMCIg6LXrvWVp5pR5ExtaeS47qvO571eP/SlcYoM3El5oOFn
YYPYENzI6zEXTAoDFmWUikv71b5jagGpXpeBRQmOFMdiA3DWkBBxX6dyhRlk2j8C
WGsii1S+FJv/zQZN8NSLmTGHQSQoguuh/oajf8cqzAfAbghRkW89yn//UrMxmvTL
k1+qhTovgcg7TBoEVnPczhATgjgZxqV59NTtC+as6UUfJWt0W1+m84WwsJNUxyAD
uIJQ/oyk1cFtMkpOSctyhpoNjNeuNH0Z0zWlOkjvDgU6cFIxhMamyZWwmUjmi21I
X8OuZhM0YRgG/ZcHqc/P1XlHvh5O1p/hqm/8Z74XNjmAN89OXD0Pm+f1jRl0n/Iz
6TSB9tRr+wR7eTWugGYOThYwrAmkn7Ecfitz5+r1n4+AjQ+WtWC3baSfgvOaS34X
C8+ys0LYyI9DrRkaz1ikf9P318e2M7reJPlKjWMw7mEwqLTRBzMekus09KIUH0+u
yJak4JgODFUn+uSYZPmGvXetVJIcKcl5RUNZnuVEj4z9V0VVrxbiDFSfgw769SdC
oCUsRwD0OBGosRqjZ24lBnTK/mmvAeZvDuFKMeHTFW/+atBZcxQBCMjm6FYp5wXH
CGfUF1PjZTSB456Lhupr36776QpYcmFWJ4stzCrRlBDh7z1JsQVn3hqqpCttmCRo
Idty5syZtLHspEtDCDoJgfnNCBjoBBgpJnV+4jA0QxaqqBD8EYQ0Yt7VSWAa2WBe
dgEquHNEj89Go8d2Ntbi3eKEre1FC0I+cC8tcwKPNLxxNMN368NgNkrHaAssE7k7
ILAHqsWTEr/hJzMULXGME1tfZC8jf4pgPdePzs2lTji5SoUGaVlv48xzUabUBhaG
b/I/vyfyxihvpW1hhLdYamfbWVlN0Dt4UWq3QBLeOZL08YTow/lhSa/B9w2FCDYv
e5uFGV3F5d0cQ/yCczU9nUlbsG6Rals9hVmo7XlH8CvAVEfTXkSycdHrkBw98eXs
qK1ClkadNsMr/ZtQnklyb7Oq04XUUC2cFOPRLuF8Y5mTz+6NX7X8UO94RAMqYDrS
duwtgALF8V80pYr+oYs2sR4fPMUBrcWi4sYbFaUgy0fljTJx3axRNnTFajh8Ao3u
fTTq19oGxG53yd4C06AE0Z6coULyeC+IAQczsz+srknkaKMx/d/BQj6E4p+aBDjM
0vJM2RpiweRGjaIyU0JBfL5tysg4uDiVD3/Gh8c/pu5uMfZ4/+BXiXQGAuTuKL78
gm+tssPzxoDrhulUaV7m9WBWaJNTrXbWFese2jjyBC0Df9qwcEufvAceyYYhgFQw
tmde2hhyYoliEr9L4QNSTLQZir3zTTToOxQ2x9GqZyMvbrSiqIkKHddpiSiZ0ANU
j8NfUaUY47tinHzOGAlLJQLLCJ0bbCVSvq0N7U9sm5PUE/EQQQnelWabSE3A02fe
v8U8SOjUGrlNaoWBJ9dBtMmSZQ38P7gZ0MZMASiBKSQwN/JzclJcn2qQ1q6vVbtQ
HQ6xBXBEbnKW2Qaudp7o0ttc41SsqFj9kawHfX+0dS3+WrcM0S57U+agTOc/kGiV
pTUrKfoiRAXIr0QbFst/pOaCSRw/P4ZJDEv239XzbzWAjYGm8EgihDBxQcZJGW0I
L1WDaHl4s6dzIB4yOBR8+yQNdAsTJT4G3cNEwd/zMvkODdcBEiN9hDIYJXGP+EGm
D/pV+KFr2aDNpCjR7cGk5W/levRqC+t4IeEhgzrXuf8LHIYC95UYlgUs0vr+Oywe
Qku6k7yBVdaeD0LZablk23mAfT1ybFSGUbv+R9OSQ/swiugUJuuTQ2tR7WGZJtE1
vAy3/IWBkAQJCAlHYjy3x10QuDG6dZYXzoWNp2XK9ms5piaF+4m/3HRHYtxt/sxy
ROBoKbX8OxM0ko4ip0vo9llOX6y5Ek+HfXtL6J7pC7WVH5FE+yroof907t03wekg
b5qVNqZ3FERaYV13GBCiipzi9sz8LqUR7esjkhGKvtL+pYvHKBXcyqPsbM39cr2H
reCdr0MrVkSX6l9yNBe73nXFM3OkheXfqgFq5M1RGZr/og8ivh7KG4wye/kdPvDX
Sqm5zZDiDHwXGM0kANR+8QZaooGmhW+CH27p5yzwNQaev5mrtsFNGfbI8g6E5D0D
pY5dnUbY8IQgJNzFa3j5rXPM1YrHyUTuV0VUhHEWZz7rcgVnGC8HZsecGBcgMQpx
87E1faX5L4HI5UVhSi4kswbTgzMB+fkiVKmjCH8HwKO+k0PvrV0awVu5sJ2mVl2L
Xhd9c6C7x0OXV+mAdsfafgzwNlMUYKBRfgA6cAnESYJrwznGtvCTp8hvo6K+JcGL
LIFPkeqTfPImQ/eHrIQ28/f3AlAcA+x8r812xLTFSyezsoLPJLZ11e0TPx+0PEfH
27AlSkmB6IoQh9KdPA1OVchDaU9c/SKbbHUX7ABUjog+FQN8gWABL7AgUtywoxHz
b5a0tWmM6wcHOJcZgIbgCGqlvXDaWngm/aGEggEVjs0C1tOGcJFXncGePZYEh0Ce
9VBPHDMdcDShjRT9/qK3N95KN1OYBFfZqPbt7nN14Vs3AhMPmUlyMBB0d11hIKRn
4rbQ8R5jMm9dWeJtueBdViW8BJs5YfAUmwM2ihP7rvQw+djmoE3UQmKYXCzqjZ7l
FV2tWO7rzJp6pav0LvN5nfpPI/z/R8LInxUE3RJFZSOn2Q7d2m3l+vFxSETLVQwo
Wrz5IhfBdlfeem+oGnlBFH/VTYV1er7nokoZzWmcYTiX5ITmesF8FSTl65b3h9sV
2d89riQpJhwT7fJGGP8qbxDvwvtJgUeO22CE+PCzXPvnFX0QC889pqg5RCND4IJi
ZRyuGWP+zlqFNisvSCPyiYm7NweSwUHxM/lz2OGpySJKbLoGNnccCNzqPQpuwx8p
wiZU9H3cWmlHT0VpHHFhnQUAIZcqR/X4TsQGO/iUVuLNqbQo/V4lZ7pwaMMYC4VW
noeMAv0qlG3hVrMheeh0lsHZZHB7UgCpCARm34PkoiBUcv6fOHvL8y3zgW4cbDbC
Yf+4hMaWxValLxt3Jv71hu3S1fTSb2IqKlH72yS9ggtMfVJKfE2SK45zwDgb/QQY
Lxkw1g1RQe/lPL2Y+2pviW2NBKaN38pZMweaK7KKpZyGZ0glpPJycSVFrxad5GLH
kfuzOrPf27cIBCfjTnAxZkuiD6ayE3eVPIN65ZrP2Wnrei8YnxB0hrk8QZf0u+Ed
8ef6VNlmLpVjlJ939TPOMlDkKHs9hgt+ACheMi138CO2it7BsoEIBePDUZRcZJnK
jnmN/T9pidR0X53Nfpu5fbbACA89FRDruqtay9IoIOBig3ew9JyJ5oW6RFrUKzdh
WtPp/tKxDkXN2pkrgIKDaGhaqY0a/KSOvRTKCp8YjLX0NTK3o1o2gigVKVYF+jMA
C48gx+PKkzarFUCBloy9iTf4P9sy1pziZ4AblLKCcGPS1gzIcwgV8Zd1uZaggeKI
TB9hiIgrEv8x7LwC3Vm1lP5NYX4i5ANRR0NunVROtdXf9/CW1RY2dQjzL4LMqkhD
oQ8/NR8GipUyAklpjFnWr2301yuM6u1qWN3EtaZMBGQNZWsSnzmBAeQz1EhISo1l
W6qOCTIW7ZxMrVl9F8RLnAUwPJXz9OUhak+gFA6o+Gaanzf1so0sLaoFacXBMXfH
cnQwtgV3aWWbtf3cncglLL0yF9lkwbF9VUG9SaOABB2GnZwx9WUugkhwYAGm2tv+
EgvsP2V1X1RiFUkE1l+yOK1nMlMSPZ8fEFqYNHBUaEIkk7xIXaRQWL4TStZMj76S
XhFu8vinn0qQ8Rq5/gDndYaePSwNQAhUu8KYIlgHF50RBWDxOFdatP50j1NXHWF2
c3+o2ok5Yf8QXcSaBhFhdNjsEjiM2x/MGlP2IlejoEW6+yDnJkJyu/4VkiP2R5l2
iE5ipe3yugZhK4fyHsSYN1WFFrKm0ndsiuMXQl90EVskl1NP8j/fGgxdkmLqqbvw
xf7rtUot0M1dgZDAJgdonGmkde85BGzcN6yKAShvu61KdCX6aNeQDqjD+n+pwmVJ
O7aFzRSXnapbWJtPb674MXE9nyZq/hdlwjDJKFTA4v2PT6CcPRYSUyh+pGQToXz0
1+dDPihJCNcLvmGmel2anJBBs+JnB/oCvP2jZ1xofIWsL3IfiyX46VcWDg+QzVqW
l5SlJCf6VHcWvJ1eoh7aZApCbvuFvzLIAX3UTZYU+kPs9QBx2gMhzuRBEIq3kq00
/wRvKR1ZbJ6Yfh02VcysEdFsWOw7LxWvbpbCJw58Fjr5zbuvFA4pQbNlhCGRM7h8
RQKjLlvn2391zzL7C+wcVmfeHMoCzokPgtCiHTQQTRF6+LFB9X9JF5yc/PhJnwgQ
H72lxRDlMtM59l4nnStTR8PqLa/PsnigYCmWSy0Bv+3p+ejemWVo+4eYlV2v0I2b
wnBwT/CQSK5jt5B4R6ivvH6NHaFAk0YHMJcGNWZutTXfiQHUBtnDXhcOmTdi6/80
0EhMsTjmGrow0BidxQD4OKIi1DYueACvSGGCapB0xYDu4WZWgcExzNJyGUkJxMdP
SXW+GJLIb0RgGyBABFvRe0Nj5AWWmcDWG7jARBVNFXVeMyTueQeUZxFMdAbZiKq/
g3iWpvqMlduYLslHhuEql26jakZedUMwv4Sl4XUERg73SkU4Fq76Detj05vnWg1P
44UnTx/t5D01ISsA3hs5NfmrskdZPX40zBIGJGD5ZtMa3SadgWdLyADV/Zwk0qwu
vME+SxPHPjT5IKvZ8NyHDa0LL7beju/vcLq40BZTQAgeAIzoKchlbSrLyAwo/pP9
mEo7U82YSbIdyhc5Qi0eD3H/VhhPqRrPCPqrkM+GY2/VHBbbSlYzgjYuPoXx/lPb
TsWufHycIH8R4UtyfPsM/e0euWZv9Fl1pmTMS5NOGOK/A1rxQgQ1vSfJiH3sM25g
ZKjv+74Z6KRyi72bLR6P+crX3YI7/ldtwu00OvjiLuXPxg5CXx+VLlETRbMA19uc
54Lpo2TtwTl3PPClif8H0cnjtmFKABTOnLDYi1+VQbmMGo7evi4ZJfp0W65vAJt6
TJR0s5AQ8oBpZpjJd401BtSgML7nA+52ROix6c9Asqa3qy16Vj04OII76ta39M70
47nRwgIvhA5DDLoYX6XyrgCxNDWUehYLcdM+/bCR787YxrR2N/+8MGNKza8sskWa
fXG9koEQsUF6eIMFzrEEAZR+X0Phv7cunTzjZJoYKQgwxJ584Ij7ZJvMTIi9mt8w
m8rwng0ulRTjdZfaiQVFZXan/f0KJ3ZOLM27wNRxoyrx1GO0dfPF9M2E+JqJ3GWW
8dcM70OzGOucZ7mUVHOTuhETrh+LdHn62CEmSO9Y7ZuPaIUcV9x/I3V62R75aNuJ
NaPQfuUEzgkw2uwP7h7OGamknVT3o288rOjw3soQ3KkFL4DjEysxEl8RsP3++Ok0
X0iGYiRpAtPMEWLGs21tT3UZcKy2q+H+EOM85wqZ7er34LlFE4IJQc2hEbj0HJ9l
QdmmXwlmVyhon+Jvw3Rn7LpVaRdr0RPu5biRAHPDzTDIqZKpM53GpYdE4q2KMmql
n8g7nIeM4wcW6bsBZj7RlquIUC8kggHKF+PqjtXyGNL5sGYHgC9Pk+AfKixajWbj
wNrlquO98qFDdNEIWi5GezNOeLEEq/XoEIFeld/NKto6yPTwU9DXhgEYLXDgiupr
IHmr7KxOBVPWvdAQtBEFJaNyhRMlAtiwI9HV15NAZLIJ20/Oy5rzbOT15h+nC6Lr
ADV91kPeW72SmnEwqER3QnoDBd+8GYX+d17F0ruxeyGPhKR9vXNSCYCKtEbDjS9w
Q1HjIRCvYZktvJWjP2f0oDhSsGvoCWh1J3dtx/nQBzhkmtXepiMzh6ugoYwKa1Jw
Rcpg8433YlHCrkRr7S/BUqYm1m2PmBCCc+Dn9v9KKTrjyG6Tu4rc/RQ9q0DTP70G
+SImVuIH19GT4QQ7m8AjjH5T5kjWW9hdv639z/pOrE+Z3QArdhduE1nE0aHQFn6/
Xvt4rt1QgTqcmBcjPES0FNkdCrrXny7O2oUbk9ofQv9u4MEuO8Yu0ohjBT/4BNOB
JrPzYFZPpwmzmf7tQopzpeBji796S6fy3yKGTnER28GXgvCMnFj5YizGyenncKdy
uwaXSvcKlnKGf4Jz0ADPgHxOMRWCmliO/UQAuEzGIIwwhyzVmUKuI5nddxizb7UC
DOFpjiVS9vLF/jbRS4suVLfjLWNmucp+0w6BsnCaYbHbb2TtZtOE0aYWR60O+r+x
04fh+JKoSiNzKutlPE9wczUjwWeMSEEPm71Xcgc8dRSI4/JWfZVqEtQRMbyNU8ME
YBkjw6jVoEAOVYhxxJxDJjovBZF3IycULf90lKxEizxdgZ5HGYWKx6uAbB4UlYfe
y5R32ShLv5qshno9gUdsGO4Jqz3Bn3Qxe0N34oiLyO2mLa6Z0bS/8Jzpw4btBx6z
iipP2ZdpwWUSYHP46Tz2fByfpQKmmiuEb4H8SjHAi806bj/Rvi6dHA6VarBPFzNm
swUN0wwMxM78x6hGbxrS41cFhpoN4kSxYaFAb+K4YjllyyDAV6GjYHc+zXBIBO0b
zuSA/wJ/PZCbT1T02cJHwGCp2uKIor4wCrgPJOfsblm2v8TRATs4NMgMhen2YmOs
NwO1XsCxAFnitnIoAIAYi8tTi0C2tkj/ahRjWfNBc5LzKeuLAV4R0Tm2hfb+q2Vr
RS4Boyv3EC8xj4JkW4hPK5ooQ+yDY8GkOE8zyQOsLl0P1omvXxjaYI9bWeWKqaSH
NU+sYsRrmEAeuS/XIJ37tECeXqu33wFfTJ0hzP4kFiUbEE8sz/mBFyZzNbnKCLsA
g6i1VltWYfzOtk8qNTiypzDASH/7hCfnXW42KEaudKA5xjSvgUnkbXWOmrH1fOxt
F+ohtNpkDPOUXmYp+P6yfnjbe5fjWFVNwVzF0pxukBPnru9wxg/Kfijd47zXfeK/
mhVeItOXUJIYhhupixFfgquvkNWUTgna0tZNyMMZBabIBkRMm4aUbvGhXOTpzOKF
b+cxA2gq6/muNgpgfKR+JRfBcnq/nizJfSVePLXpA/zlrJmF9+q5kktUimCToSEn
KNqvzoNBWlGDwUu+LVrqRNJ741ni6L6nwDjKhWNgeZjJLZdW7i5kBHL3BcqmK+qi
o2mu5miTb9pPe1YODewjhnpXhYd03ryB3pnwlXi6bHNv0LkxAxtLC+d5PpU9UBEP
6zoKzPHgwEHIZOPD5K1Mo3J6qR/heO9zXDa66CCSd1yEcFXr9FGzMbiBeGdmC90G
WQWaZVwFT5XzGvW8w4Jr+2LimH18B2XlXizOIyi31jwbivsEH2DWhIdtQXO8wJQZ
7vFroyuZj799zQJnbr8EzQ/Kc93UaJ+YF73GaCcDtLKRswRqZ3dHkKWrzYcMiBYx
pPp58OaLhv159AYq5+B7UrOp1Aobi/dFK4wxtVzjmBJxaKyXdEbqkJsEjrNOlpeG
spsjc7+c0aJJdiKDgl0cKH1aNfx0+J6I3ssdLEgH96KVi5XWxUeBUkqNe3FHMNiY
RvYYKA2EslDtOnyY+pK90r9JB+Yl7KvAZSEDgBMXPwbN4cSSmUwY033CAPmbEwPV
NZuEZCMv6xpSDKfYDb0+B04uYmgI59IXOfwHSt6QtW7h0Y09FiNnSx5/ODbMjdAF
6hU9fy+gXG1nChftLLwUtJ3XuSN/qWDFbkXtEuniL8u7xWSvqb8z85g53Ly/PELW
DuMo0o15FpCxdRJFwx1EXL50BfQIgy9A2Lj5eTL66C+YRKYXGWnFUc941TUQ5znh
xXCq5NY4vZHgzQBYnOu6SHGFtaJQWihrcC57PJFrH19M5GZUT5ByUFTqAEWJCAwf
1OQRurAHJD8xY51GiECczdo6ld8eXCz3kCKGVeTnJ+05JvIQDio5X+vrlHewho2m
yIaQ69ziXkgd9ieQeGQpVSSWBP54xomkn16sedeibrY/vZa21JfSlbaDFiotAj6m
2cmIMqoAyIu830fA1uzkQRoQlSOauC1/DEdiHnG4rnfYsQDeEOgwhnhEiioTfB3r
hHXaBCnFDTC4y1zPrDXnepSb1I2E39zF+hxZ3ChUZFUZ5DBdAUmK0QFNbjzUry28
zvipqOzh2MYiDkpoWNTwUcXdkzzpXtZUpV2ardtI2SA3UZ9PmPgOJdemOYzJeC3M
XV2V2/jZoSe3gRd8FpR+GZZDMwEL4WuF7c0jaGxm9uBfstRSVCOztNpRplKfae8o
pBBRLmpZZU3myGAUD+KORXeVQMfiBr2UcdVqNr9TeKpmXS+QDiPGWJDNUe1cSW6z
2DKMQYoBIiGESGW8/yE/kHK0MX5jbpFWTp2ceyz5ler2nfb4+KBS6sK8VrcnLW8R
r+3jjZDmvY/14OQO3+dxq+KwxjCNF6Hhcc+CdNNTVwPFsPmHVxpcY6iRNBkB4vdR
dH5SrhZBo6i50aQFbQA6HEGgt9pKDZKlPEYjY9Y0OpHba8nhR/0J6JUFSjoX8Bxi
IjYiWgJNziHUlL2CpboH4X7RvBU9MxJEVGC5euYUi0lxbBZeSIBRppZevWKr8/D4
/c1++NNj6ynbnXtKsN0O7FS5fvZGjvPhi7xRxfUAcJ/VPA38pHjXkv/EyFI4uJh7
ZZEqCRhWKs95xQkJ7uWPTFVl81Mol5qrwbtOdlPpM6tvgSXe6WbYgcV0mRZoaul0
Mfsa19FbWpxGzHZSjFozk++Hz0r/mCcfuWfJfvLl4iTvzpfpw/l8pZyTpmgtRP3C
VCcH2h6AI8hXRyfrgyDQAol0ahBkOlW9f/gLJmQYgtTUGwIOySQ2RiKHsHF+KjGn
61tK3uZ0B8BcQvwQ8+aj5q1u1rVB2iDkhAMk/hfnmDrsJHOf0kOLPQzuABDTS2Uk
vzyV74QcMMNOchEaPGCDJGSo8F6QbRMNW1cc4J2TrJwd/md8S4KSnXdf4DBj7zWg
GfUKWhhX7g45Gs66zUoF5edHzpXOF3Q0DEs9suYMGdMa3Gdgw819gQPuPUzhDXnX
j0/vgJrEz1uxJeEIgVp5mKWO+IK1GiZNA9XfFqsInhWy7p7chD0AADLcM6IrWt7D
AKsD4FHf8nfgVI0zC2PkXcvLD3XAsPjEKgE+feDggT84ZtMKIaqPIXdaO4WRNyhu
1IjySOowt73Ie0c4fLk5OLR/32JCgUEbtluClew6f2s4Yry/fgqOqzbL5ZLtw/WB
QyFpyLZ7zsWVVSYOgjkHHWZytAhnz+jJ4C4/e/1472uM4r9+xtbLV6GY/oOJJzeu
/ZiCUWpsa8UwLmCKv6j/tvXEEcV1z1aTxWuFJpiIRGccsydiUyS9IIppwmFTwlET
gZvfJUqWjTYfD1j0uO44MVByAyLc/dmVCGGo4jShFBVakdzkQOJLkwHA2doHngMJ
gTRH/0jAr/KD3mLVXZdo9H1aK3pV3hXJ62TISVbvftRot4su3vw6r2qsxvpVXHTz
43hrVzcwfwKC9YXYVti6UnDQBuOsQl1aqDkRpYrZiQm3+mgE3pLNnEhutulNgp9w
TyBnAKyBjuAYuq5W9sS3CIiSwc/755WzbuMZ159RGqAf+szJ4OmawIQSmfRIufk/
Sl1V6DOUMX1eXb2MBO0G47r2zPGVleRYzsNg0bNQ/OfHVN/3IJDdDQRfrfzVq5yu
Hq6J09r1OEX0S7Wf0q58xMOeJzm+4QCbKd/voMagK5YPkxbX6jlXe8USO8BD3j78
UYsHC2F2I4r8xtkL/Sjynd5+qAvFOPTm/diES9BZlal5mT6jVVqvxzzs41lF0qyM
RKHQ4Ti0nd9BQO6FbzirWTxpzvt4pqxs7/60BiKGtBPcSM+0kR4mEZhK2sQOrqLg
cSS/13UoM/FAzmDk9VyYzuM/a4C8vb5spOJvbBm9gNfFqCKc8Lk7XsB9/Odeli9Q
D/FCZM281bM3AwCNxRoNYsQwlEjtKrrPY8uyLcZGD1GlXztOB9LQe5QsNxFTaJQc
pLmQIWXZsKeuYmjzWo565ujGES0zhyeVMKF9uC0N/JbHrosbqpCGnFUZ4oRF3i9B
47gHA/mwByibWwgFL7AKVw3J9rGnCyPaNAjvIc9flSJSeNTGx6Nu5OLgkKOgyN3I
WOQtzq1imTLiDvysyAGiHGtQO0e9cLtyWnmPwH6rsH0s7Ai6QW+TVo0IqWAH/h/W
57+MKFDqcODzVugBH4TIDy0oNlqFlfImsPlA/f+RIjCDk0AasF0TuBDMAVWFV+jk
Q+SSnfIFapBEgtFA9/1KejTXWYDrVHxpJCNh/f+7JQuc1OTek0UaTdfbnXGQoopM
sLOpVtq46YdYbE6dyRPreU1r5mWtPLHpH5dMYIihw5Bi8+sxspuCDK/1ZbyvWuZp
+ad2amAdqTJ0IEDYyi67+ooEWT3CBb48riSo6CxK0pQCxQHjQa6cVJxrOuIJbACb
VNePGsIJZ29e6svrgX1YIwp/sNWhpy94LRnfAyzoiGwwQKRBOKFRG5NFsrpexidg
jup+9ioPoqU8ubWGCku7DFpEiwTmUotkuzjkrAHG3O7sYnXxbcn24P9qg2cRJOEr
o1Gjjkq2kHKuNc50QmrYdO18IZMuxBRiz5r7iuTRuU4sRgF2OtYNC3FSmRSsz7mR
fHjrHLBYQuoD8xkkcSDD3zKTQHd0tvtAyUpi8sXqDWy+vxnpLNkXmf2DbLHkzsb3
JJKvXtcjfVBiWk/PAXs3q1314vymP8Phu719kbx6ksntvz+lRBF6iS0RWVr0Y0+t
kNzzz2t8G89lguafr7bMXs8T63TDqDwVKIHsJqRdznvH9mjOKcKRiwb8hr5W+Erc
PcgBljPa8+LWvd9nei7veF7/+7TsuancxJpgYsFNa403uKOpl+Z4OdGLx4dsOe/Y
EJWmYtCN7JDfq6JGfoCTJCewj73CGYnyuWyoF/5RguGNfxrB7+vmDkAAL7F8UY90
L9dSKB35bBQMuykDsXadmzrh7hdT5Tnw8AFiC73LP5SfeX1SZFlqfd1c+a4hri2B
XXAu76m9Ving+Ve7gX7XIk3ShLSGpV5E8rwvFVDjQ9P4DFzmD4mBQkyMxdGuhs96
0HBEixeg2vnB73wwxwaCOQ+H3Iu3NIoFg613NFiRZ/vt/Qmc/spqeKHPLSS3WFBz
ju6pd2q5I5lskGOdG4tmilIbPi0jM8qCxaIXqNv1nigSTFpARguSe9nLKdpzOGT5
7ptjwAyG+EVi8tw3miACi9wRd+CAcebcwO90kn1Tjybr8PcIAQwbkT+sZoxKykdT
I2anJw56cxYLWb03xrCMPQWDEZ2Od4cdJlq7Xzp1n0cWffjkr8JHUGm+wn7v2ju3
RIVkACh1UfAq8qSbIRBHeeThy1cCQYja7/DHVMrqrRjNXMQeSMpVM/thHmNs4x0g
zbHi/hV2eyGEehK8oP0E9ROOrammUlgmRe1a9exxUkEL9vKYcNUsnCJHP805nqFM
WPwPxGXquxRdAGTE9REKO4YQo7Ne82LXh8gVxgbBNPuLdOux/ahONM6SGJ7+1fPt
wsONmOVz/ryC8Ha2K6AoiJl+DoNrweMh+jKaEEHZe2atUmIEKfiS95e6hKn0Tx6+
I9CCBx4yvzBfim5uRYE/NAtyz5XvCAVsLlDxAPWxxX/Bz950anaRob9Wda5edjaj
lQQvfKwDyU0jhNLG7kb9eS4uSakKb/5paix6orc0kLwHi/lRbO2WJFtVFP7mTHmM
NPnYAKU36O5D60VJyMQwJxB6Kt1MT2ADuNprv6Gic4zmxjI7NiITsg/ewdkFFKTv
RHDQclC/Hqs92qXp4WjPDg1KwIN5N8247vikosmcQCMHRbCs8ZqImYTNRbEimzwO
9vGhYs29/ITh+kFQWlmRB+jeaQlA28j0XqRyrnJ/r/+GUB04i771RrlxumlPUrgO
ZM1nHwvV7vvC4V9h2PiNJCI5G8H257fuTY/Zc3C22DBiFJh5kb5ebRadC99T38ex
aWOyDfJFqx5Yy7rbBLcQ2zWw2BYsOUA78BdbNn3E1h6HQCP/4D4vx+49U7zgVciR
Va0SnP8vESIYX6D+uZa571+9yPBiAJ//W1h3wMFndU/Lm9DhePyWZAJgDrjyB5IX
N7svMJvgja65DGRfKOchv2yf2Odl7XaMcMr5Okz1HHjR1ZTO3EdQ61M3kcPIzbb2
Q/lndG1kmCpQ6r8AIXMG/OGSLVgC3WFeHHocpgptp23VE11oi2F8ZHrHoRtA+SOh
TfpSeSRvjX/7zOHrl6giqOSCdfNSGAADvFn0oGLi18xKlJZEWtCRFhc5YbdoKpkF
NikirDcfvXuumtzZDfni7XgYSRYL2rNb+2pta9T013DXioeFNlrlEhDtEiFx7KOo
ov9r01qATdy9bdqKzzFIbGI8oeT/B9lFajtWBfPKFjLZLQ0j6KQT6TLvgiEDE1UJ
yL7zcAcrzdwWDv42V1GYofDuxw9d4KPYVQx5bLv7E5Z/yMUk7wSG2tTXS3k/Z0fB
7CqkD70T0QkEQCEw6hKK0vAy3x9t8qSiG6IsXUuXoNWmbeDRUEOs4j6goMmmPHcj
fQWsoczP9AGi4pbOD1jEX5ZR1hgnHsIHP1NS19dXE757pDqFasjABRJKRzH0eW9d
+J1Ds587io7G9UdfDkQZYK9/5ERVZs4mcfCjqSptCmJzs5UvvMni3brthy/tyw8W
qPGwvh1aFZGxH7iZtG8BCFXebArYlKURLGZ4OHZlL4bQbDTRjrAZjeWC7S9wkEY7
3oTuezyRYtLznYMCftsRMLS4aqWCMZPBlMUw5Cqh54V/B+t/LJtU30ivCfle+0OT
Ke5yJsBRCc22cPZkrdZCguH7fr+dxIEe35ioUwpRy25mIQjrIqX+BKO6b51mFIkf
ZKhFaks5alx+Ct6KHIU3lqcrjZlxOzVxcFS3JiqMkx/oPCkgE5BxvYyyTlEUdI31
UrK7FqQiXxQeD2bO+KzCGePD6lkAHg1hKl6EKuleq2hKYvXKNN31gNz4lN6sWynF
yKAov6cYwllLsn8GCMPfUgNR5CIbuz20Wuu+jRwkoGsfm0NWT1dqYvKPjyoV0uKE
ykYqinLlsHcNY39tK0zbGG1SbeTW7+L9dwZFHytq4y+1qGspvVptEDl34bPq0ugC
bmFjhy8ZuXUYTf8j9NVHyr45hm3YkQh0pm4Fc1IyGUIsVIl72KILtVZF0rdGjhed
JFIx3Cp8/n0Ke+W/CC5zeYq5I3WPpC9Yna+d5g3Eu0z3sT3kQ4bKfd8DJn8TzjmX
n1M6OFQMxuF8szULqq8UdMxRn4on75eHD4vzX9lHaR3dJNN/pM3d34yhHkGxRV4T
GiKXLsbvS4++f5DxIcoEZJcHshv9JbLBMM0RhAthC5cLbJZLrE6n/NNakMiWgxzv
QbeOiuOZW1br9d8PAI2bmWUFWm705krD1AoAudV/Rb5D+e0nSWb21wo5EsPfJB6j
IgJxXLCTVY4dYwZhrqMsHU20fZUIn+lCBhTPgcJeXXotvKMiFotfja/fz+rhQkJl
lMUcV8yO6cTOF65jcSVzm6NP+frdX93VOUnqLJhtFB60EFCSiU+89Nax+NOTr63P
PmwtyxKSCwUL1BDTiKJfe4RuM/OfNHsj+7j6rh8hcvmXIkdGDaSayt8/MRE/baG5
KdiupJNyWHyKkPNGkwVXcEA1TCnJxsrQdYKbY/2iu4gd0PSyqlXOnEVcLP6nlpgS
jFsQJGA8K7X1ZIInnBFYp/MPZeM28BYUw7i+vxoT29klHpctGUtvM9hI1z46Ec8U
MWSI337/hvfR4Hb08ryWf0IDyGwoh8zYbJ4UPyRkcHo1bTUsw9Y42N2B80BCvCSd
QdCLUU9Y1AGhbi2p4zSBuBBtA9QN3TKgP5imy8eo/cRPwKHgkFFtlTRuMfJVJ5dE
w+2MA+ImH+HONeZvCxAXIFokw43aQ3n+69SFtfT3TgS8pHk+iHKRysiVgVkNYwD1
0pmlJtNKIDd+gVFPyK3fU57kqsu/Xt2wrr8sZ9Xtgd5KBPTIrhUC2H8qZVVZifHg
V8/i1Su0L66XEAeypvAoskLcWLFUrczpbMe0U+bCraYd9bA3ULv2hHYQ67oIiB2c
od0FC8tHtnNdQEtAvldv4Pr4omLSg7hgExMHigZcefQFXyVhh8CavkhliXTG1BJz
IDvkwChGQ6ubuC6t7IVTyDHqCZ6Gqmx4vZ0nnL7wiY27IB4k0Btm7mFz3u0DzzKH
FL/WrXM/HmfjiUvonpCpOffwe5gEzZxTETCvkN/Nr4sntnBoZwHNEHyNn9kSPu0G
PEB+MTmcGV2sr3M8DcP8iTkAHIluv3iRTChaLNlnWzl1SBmLjYCWTSOJT2RbqC/L
PumoN697XNgtaia/M8vfrfm7eGb5DN7Cza6Aeh+6PVpTkUtTNloWvmQtF0ILSE3L
oXOqPjGBSpZWjku4MbmpihQ7EIS7BB9cDrOJ38zYYLjkAqMr8MYU8UF3YGUh5Syt
I1lbsnqs03QFqjeuGsy4kAqfR6Qdi36RGEIKjTy+SlPRMI1oxdQ4j/lCFm8Ev8dV
iPtFceRBoAVqXM9fToT5uBW/FUK8BfCKm+tPmJkSLtrqznvBCWjWpvDDYtOSq72Z
XhLG6yV/K/GM5je51LQQSbE3LgfJC71swYKSPyiRihGB/glup/2eupq5ww7oCqGb
21i9aeuMm1IF9sqjCdJ6kRXIYMnLiol9RL9MhBzTHspAJd0fcjiQLQ7QTivErJm4
cVj8NIiEqlT6ctv+xg/liJd2w7V7AO2yne9YagGJN3iHQ1jU4n5jNoDeGcMrd9Y0
NE1xDyV+dQiuA74N2AfUMzgRAYtOkicOvIRW7utVJZiz7W3Aaivb72pQNtaZEq9O
hWtfnfJllB+BInPUmxuHkXyWdVrdSoRHNvQnlf3bWHJ0ORrZE6Ao8ylkfuqXsJOA
pmE+kpJzI3pU8TbyLYazdJKMlBrMmyEau+urrDhrzwpkqDusnSAOIh8tiME/n4RQ
hKtCnLPL20N8jzHCXDutYWnsBLB/c9BvVkDEzXJ8i+HppRE02Drya6fTG115WiEf
ddxRB6FnOmuGxybugvq15Apq+/ukiAhsyj81ftHo8ez5kzdZfTTdoHhCEV2KhsBv
4oIaSX7JlBkKgUhM110VkqEWSJtU8f5BtBiRBK43qYo5I/BpPAYRCkY1dsiYWoPp
Arr7mEa7SRRiUpJWdO8A515XcULkE+f6AJGfx8Lls4OA3kf4K1XhCHxvtPvGpy+n
YGNWI1nr77KRoVZAGBASCdanpB4hozBz1bIP3HyJOjK1c9sX6he9M2LdSW7rE88m
d30LFs2vdnFUXcweM134PKqX6uke4kDVcLouZQiOmCa+6FCpiBgMD3VP9AvDgaFU
c9QzrwpWPS+tB7BUcjOYzbAP0t6dM22Qn6y5KXglIGupKVUMo2/R++WcltGzDWx/
/0Vbr3sYq+nmgzdPHy8UDAx3gZfplccge1p9JlGbaU+W7Nf6qHejkHqB/zglUnkV
A+EAahQGtg5JD0gK+H7L5AfUwRW55gWRwi3x7Tqr0UanEoCVTcvwdJ1+m4mEHa/r
fnNlhZ3xz64xnCnKpxkm7xfFCfOpx/LU/xPv1sQyF0K92Uictt+u2Xx02xOqGJ5h
ssJwok2mB9naXKNmkj0ozuAqIdphTgihKe9Rr531nKRnTJRT3mbxDpdRh1qUHeNT
iyNhLIHjQY1TQsdCHgoJ2fpjctpOUheN8RyAIg/8+yaQR7xEUNK8ldaP2C+NCSh1
DVEwZkKbpHZQ/2VOZd+JeqY0GrnAVuavj1cabG9iutEADjU6IQ7vD38kdJGLAcal
Eh9IoVri5WkQY0BmBbFgTwg1X+Q9vsYsR5VB/BvdwKoA8SIPVlTQmOKiN3Rzpob0
WzaOLA4Nbwh9y9RAXuqa4O6PvJ4/dMRjZ4CMbRV1pxeF64EbfIslgXa5YyrSLBqx
rsI49n2/c3zxPoPaVVjUY9v6qPGzOAlBv2vY17szL37j6ss5f1MAJHcIqsgzdt2d
yTG4oyU3zUfV7IR4fhnZWwrC5aCExG24LlxOSaTeIhAIX1nidOxcsyOto5gXGpPR
lARfgkTfoQEhqPrQ2SPI4mea6nPewnFrRlSEEjw//KmZT/97b6PHkOLtEuOfi/m0
l7228MGlOeKTWrjPWXWAeigMEvJ8gfJbxCxIgwlJMCioIMzEeevfOYo6271YeDnh
KWpw7W7bo3z/eGn5j7Qj8kXxFXGSIWgNGm5mHfGCC8kXTrMnIkdu8O6INlbJvrAF
/x/uYsLkzXg14NvjHczHLoCraBZb2IRbJIdesYpXmX4gxRTaysqfj3vMFVTx2cD6
sYCBMlOhdvJluzAl6idiNPOWfQA/dqUkJFobgC1wfRaOZzEzx7CTjJY0F1wkrToy
807IJ7n3SPGtRwaMS4kmwfKQCM6iiNT2peJlCVFZo3siQmxVUXsHVt+6DWkET07d
GS3gKcBkp72yNOmYjLy5BewlVgForleNKnxcw+yEH0rgZ1cy16XsA6qow2+yN+z6
0WvrvyNm5AXW8fRoRCR4FeU/bLVL06titsxp6Rb5yHvULfHP7YJvv2FxL1Ap0FL2
r/JsC4aGYRl24trOv2F2Dl9hHyirfgSbsmEiTykHKClJG6SEJ2HqRy8SYxNo70Ba
wquYszVooBrqB/f/r04n6sf0rm80jJ3DI4LEK2jspXg+E+Kr9rMAnfQb8gtKiHv4
2jTWMqpg+DG3PoSinf/Z0BBtlIwftucWROtSxgP5l+4aszz6oT7UivDHm+z+ak1t
aLM1NNatNlyj7n1ORIpAu5y0UNcJmMnIRlpPKEa35bPjYddsHlbieWMcfEi0gHX4
e1DeaKbThrbosWJ9E/CalETPHUSFms6u7BhTRmY7YDDVJbfcmvNNNKEZ1b+VK3kZ
Ofj0BiqRBq+nTj3x8tl0chjc64klz8TaCQz2Y9Mo5O/TJV36QeBtJKZ2RPZz8jdI
VzN8mAiFrOgd2RRsF04EuFQavOs1L19SLCDPv9D++dls1pxayyLegdGVUODG3KMH
f4DOEiRsSjpEMBNzkfGwJGsySI4xeQ05kQ9Itn76WR6FTHYAqaF67oXZg+N4+aqz
Vu2HC7OwseLm05ZwXZ7o7pu6xj7HXjjMoLHYmW/buTW3LtAkrpGDfSGjwOt8281B
j55RAH8YA+TBZVw+LhUIWr9drdqsbgWy2il7hVZxrGR0fD8j+szt3M5CQE2iWN6Z
k+WYMgVR6sF4X1OEJmRxZJ/pnXQID0mk8TIp+qZ8LfWDRzh38+Lqe7YwIdErFCGz
DjO7iP5kSIrad8zpQGHnJ7RbKc1c1v9eG6YtYQNX+P+S8GlhyOUdXzMPEeFsHDwY
zw6fV0EBFjf/+5mzIIhtgRgfWjcYD6BVtkZTb/8kTNLxVptwF8IsmFj3MOxxu+gj
41wDqsU/0keartzRB8aZUTAYYfnBj/dD1hucX0Zz6qydutNiBRkRCSFSkixCLR72
SmRa3M4+KFjbiI4sw+L5JmMafp68YrxAamLq8CHu6mCTgA+oztrrSOXkz04/7mhW
RSkGRm6KiTCNg3HcxIQgnPYFOQOQqPhvNpoIPfBfwMLMY09aEtpaTOHYQUhDRLfq
/I/GsO6KM4vtEyrNeB06eYs0MpLyj7PYGwD6Fad8LeQ21/3Lwvhi2BuO36ctSaF6
t88WW1SlMw05spGNjDPl6z+Mnb2ivUSWmyp+QrCCkepImz5/vNjQ08M4Y02llGuS
JUE7j2E+lE/3rvuadshj5xNu8Q/3t1WtVfA9smlpv0XEJIlAMGih2ZX2JyoExZdC
twF8PIm/FiwFUoDwbLZzeva8LDYWgpV041Cj7IKIQFyr6ACQgSd+ti9V4yjLcPqq
n17hw+eCkRHnZoHdXXkZ/t7GHXak4h8dtRf8PNNWeoBCEJBXi63OlGskiXmNIE5+
i6USppA1Cs0f1c7nBmRTPBXIZaq42amTYQLl7rqviHjxTb2T9BuaXWfgcMBH6BPJ
Dj6Y9HuKoy3W5gxjaWJdE4FrdMhsXgDOINPyOoqBEeIojrYffyh6w+n7jvDp04JK
d0kkAnn9Vx0OwDdpT41LOgzyXiz+tTAtpySQL0A+5b7942FBjWCxTiBcRi4BoGrm
uNTJZZSXGcHJOVPF4rSIdKt94hTzWWnXigFdSQPnJutxhxr1W/2Km+I2CLs0otfG
DpK1vgRg0vIHsXWxwPdBQJlTVtLXeWXsD3iFfltoRGoxrkMsGOK5wylIdjza0nIJ
Oq5Xa7z/k2zkO88AxYNWwr/PZxJWWhIj+aW5usvzMyQFD2fQK+jtW8GhUWfcc+52
ZBnq/8gxM+pLSwE5jYz2U7oBZQavbwvoxagm0OvaDSIVgBf/thT0dTGBc0Yq7D0N
lmUkNo1Jm/xO+KztgJ+kdtJkdd4va6sy4oZz7TTAM3qkgQgQrsHXhztt4RxMo5N4
MTEDdkuRb9YfmPK0Sk8iRZ0T1At6+l7RMqc37/3tlgrpsZ4ce0sxf34rLBnsEkEm
pxyyM4Ujjq0ISl88sVYaXdarnPdM9h1qXs25+uilDXt/ZxKWduojl5rSjOzayC83
d4EQmtXIesMXOxrutlciQz8gbOM2tIxx5p/7oBSiJmzaYlr4Nl1gRK1hy2+88oIY
7yRdzN8Mv7hEn2avqVbjIsR4eNWmloDU12MDOucgl3K0qeAdW4WiPxT1/WfkVbo6
vDYS8VahjrUMnQxA3cuk4kK3ZpXAU9f46Jl5WIVw/7ywj5xx2Y+tKOybZOPkv73/
shZULvhqUO3RJ59IdsGfMsx1TzSpJGeWIX3kgS964xY4FTat0AyEFovTVkTeqUzE
1+c5MEI3pq6eGN/16H6zSCoE1PzE6JBWDFZOIqfQjqopAoVwk/hnoKVRKPW3aXJw
/u4iFaDru+txh9KDlaOml1FZoWpBsGRU2fOWzKUxOyn4RDUq9G6+yPL88HZsECjC
BHDpRoW4nOHjNjwRvBW+4kw+4PifC+fof21T/bdS1Q/VPoFk1uOBFY1y+fUzJv1e
qAHED3sQVaPrIruBpiVa4gmXBKzSaagselTWABfbaq5COOoyYbMPTIr+4LkILWLP
haz/cgAGFCMIey9VpQ/0/u5uiaKiOM/ncO6Krhel1H8c+214uB7Tiow/EAN6MZSd
5fV7ughFtqRWpN9/qr9XnjdrJBhesOKGaRiIWpDvIZD0El47Oygndk+RrB/fP9Wi
cJfYk2nsL5Z3jv8Jldyx0ZEqdpf50XSC24h+9c5QPpe5wzYwN9KycHNBvx2dyjVs
rTUNMGsMCn1qcuaWJ6l4zCz8VzVM83SD0wNDUPvOuYQcfjZ0PFHff/WOHhCFPNlW
kHt1d6iXc3sLCxKfn052iZcV32UMBIY7hDSuW0Y1Ft9Lw7qCFvejElVL0od3HBP4
1tUgOYwa9e4B7r/s80k7ImXlZEanl6z1xlnGuxoilU8HYQ0RfrGgQ0W2taK6B9I/
2aWzjwFlr4a1jmJgoyPhKaIFmH2b8wFNBDRf69yOr/ZeJythlWvA9hfJOS2FOgWt
Helc4D7vlAnaMhCOYBUQsqI9FT7ixCMnYo4mq8sF8nZxDvtNxPog6po5yd7kl8/a
9N008hcjGYGhLq0ESjhGkWD4IPXz6ydHfZEEPo00mzkO0uLG3gBoS4sddHnLFtsl
oaU+rCUsz9bOMc6tQQy1GwglTlinmu0xgEk5d3ewgKpoN0iGUbPbAwe1ulni6p+s
61U1Z8EY1Plxma1dlO10syw0cBHDP4pw5+aD3nGKQ3tERasP+DaFvR7o8nm97rRQ
eweEXeP1JgPARblPvgJAe7EXc3N6Q10obtKr8iJGoJZ70DyHLlluevPePL/Hjx8g
sBOUQEtPMuqgSuVBDI4joY8oE8xpQRhm46XVviTK3yd0BapF5sTm26pqRPVYIWGm
dGq3kJnpER/XF01oDgMvQzYLgkOLCue/ioqzNuYwOpr/YAmvuOxntKzrP/5KObSA
iJyugMxj7mFCz9t6WshCX2M878plJm7kz+qVrhmLf6A13Gllb+gNy9cPB//q4fKS
xU8AhvWJxUO1LchI5ETCSjKHL8/TkLXa6cMqoWpPNCsUk8nrSmb831XD/Z2DOgcu
SPtwzeMYVfmSRp6epD4zoZqeqEQjVRTySncwwG4pgN4SU3DgI+TyfyoPUE2Dz8tN
aJE3I9KwNq0voHFiBYYsr6Jc0bBaQyFKcsEeiYJgo8ys0xDtfyrUb2T4YYabuFSO
xM+eYVipGhcKJ+zrl/v+h3HFXocCTfZrcSR1mq8Z/trPWubHFzrW9f0OssmNW8kR
OjVbW0qYGBgl4hlNlUJG1X+q65/rEwJgJvVKzRwM2nHAELZ9KP+Sr5L6vSLPvLHk
DMKGwOuNz1mLOZr1DaTtToGrnvA7Nud5jQVYq/UncbcVYEMhyOPYLrEVH8tVd7QL
aW74mV3LkjrBeO7cZprpdKG1AVIkdzayWIRAaFXDQTIgF3ZGm2c1EJKP1XcIsHP0
bvYLA5ihlPr3ZY99XpDd22kveLnF0BZtHdjp5CW54yyBRTqSKSnhak0IoA+pf2oy
P9v5c9iZUuf0fEohV7SYNrpKYhMVpV5XqxFsAL6ih63nhRZTCFa9Bx5hUkyPTIuZ
eJUtVbE0prO1qcdNLf6mu6VrudcGAB5kUz+txjAkzpQfhU+vzdtPT+ev2+/PHARy
bJPbFP8iHRGjwzTMJU4iO1FVv9oPuN+6iGmO3V8AbtSLq9ZcL0OKDeSLSBg+V4JA
ajVJAj0CjSx9eqkJ/kJ26rBDpli+nLaVdEeJeO9vXNn3HfU+884tQy5isJ/cx8/A
p5HjPRXY4u1FcwaNKlVR3qTZBOBW9OPOW4w4aPEn5Psat/sfdetd16CSdaRxGdD/
IXPagqYTPXNtvS+ZJMONYlbo25eGrUIig4bAtL21sgdUF6o6VqFb9qKRS/f/JiJ5
asI8y5SpN1a9j1mXtk+XzcyVvFWHfR19uaueFl/HnyDi7ZhJSYSBfpORKlsHLJII
Fxr57lfwvO+ZQVCcERz/3ZIk2qrCU4MBEdmC5UnJ0d1SuilsWrQleQk35XU3FZJF
eXQ0neYvVJ38BH8WbiKuwtU6winNfZKU+uz6u77zUsteQjyNflwuh6X5OVb+gg08
ZPfNj1A/zWwD6JYXvXvZE+1vphw3RNfFbbPCaqwunMRxMBmU+IXzHbL1WPMz3r7A
wE6t0Ed3wsfeSGOlrMwUUX5OOM+daWiWOEVhYedgFI6TXtrbQfJCYaKeHsmS2W6x
odyDe1EsnC9BUkZbUMcggYp0Qmlin8IuyD5tOH+8IGqpwpolAzBEoiqFYBhHuhN9
Gj1j2nvLe6NZ6FCmpHiXSNgAMUlRrxFd6jbDnDkceDnaB4G9L8l1SgDWl+trAwRO
f8eD+++TJSQJGh9D/IeIQhmNsyMSvg9pjwz0BpVghgkkgVi0WV3Qcc5NhY50qxPl
QUCOHte5W2trNccterEP64zAbWsnxWUfqQboRVQ2EeFGba4f67yguz0OdH73ydXk
J3jQvewGjHLxC0d46M9CW/oUmjk0BsVsJsVDtANYlgShZxo4vkcUztn7Qm68sXzM
7ek1Dw9jcWLhbGhcHnhmgfYI0hRVCRqdu6LGfEv0L0JxeB93Jp/qhQ57qIl12v3G
TS4JTKcerOGZdkJ6WA4V7NmUi9cHd7s1MiBIAHf6MHoRmYah0NTLQVEXpbFgosoy
YYPYVoFKuP6N8ZuUD30ZNHX2iMvAauIuOmLbJ0BpbXfLbRLoYzeVMNGY5cKkC8KV
Se55G/OZs47HKqNmQbbmEjHaTa0I/P99inF9dn4hJET8CT1sFkuXp/vUsOqCCBDz
yeT3f5HnzGoRyOcVw90IcSva1DNqdsufbhCwvc1GLXVUxX3wchmPn5A1Ur2cidT2
hXTZgmvl++DI0F1ytMQxbfv/KsAPmF9JgX7ayfxoKfHBvFvIRrjh4EfRN7zcJHqt
FKIa4PYc5y6oCGnuogdRcTf2zET2ZgtYNmbXwFQy44GfXPVc998IBqYUFhDaPj2b
FiEBrYkifXk0hQuKad+5P63JCbCF2pj5w4tSmwa4al9Q6EFZP5dU7hqkFldvtTR/
0rA43L9kfZJ+xNCeTXxrsAE49qThNJkgHWjQIpcYSV7q7ysVk+EbTGBrvNrfNVYd
t5cqDmJtCduSB5wAuNF/OFZL2D7K3fgRm3UIEsgyuXNWNlJNTXbx5uQy/cMzGTAJ
VI6Ir3JQSy8Za591nWGyEpnHoV7GW8oDuauZ8wYFxfa4u5q75MbfNKHVEWct2etV
0rcKeVKrtk6iRZet/NpMRnMt2G1DP+U1RdliF7vUuil+/kwT0BlhZJDJ9QCxMnr7
MChuN5iQpoXesgMMCqUTvYEvHIiFyeoqu+9/YTFSTIgCAKP0hvUq873zJRFJJTfm
qyUqrdTyB96SJ0JbK0huQnbPDQNllIAti30k0bf7qgx5Z6XRd9pFNrYJV0O1SbhY
x4/jtb3Ldzoz2ddQrnLSjZMUwyYps+KQU4sgEoWUwI9uTtkOIu69DUB1f3DUG6Vm
2uVhgRdB4ftH9BlJQVaLLwheHrb8bz1eofpc4bP/juIzIEdXbK7meqNALpyZEaEW
sfxgfUgbK51VkyT1+Bj4IcHIvFM/eyEDC7zBocYBL83A2AjYrIaRPHgjqddAgYRm
8gD9+ElmZOIOBvFEBrSvnvAqXrYeMzmkennn2ipE0EVe8qupsO99yRAiEXVSPWMA
VQmfye7le3k8PzurPFBV7cRsv+ct7Kbhr424G2wsFjX3qkR5lugqKX9RBaxPrUKb
cUsG1hpPnOmHKdx5bv7I4PHh1VmIAfCiycqN+AO8ZeElIPSW1sx8AZhNejZSYeD/
l8p67F1/QqQwhSvAGsl2a5CX3XSjvyo6W98xLcCZhMilCB5H6aTtOJk0j2n7tJWQ
4VnoHS9C9T6yNbYqmStkDEuuDCFORt5i2NuR4jaV3dXDrxP8ozhReWzWT/ruH1Yl
XWM/4OtRFdplnczGCUtFETwI5W+tnUvbx8JqAG3po5TIr3DBaZKz56Ofhq1xNOMH
6y4+2xY6VuhvzioCs5Hc8txuzIvdpSo0aWMPtN4DROeXr1iBrpOfrQh5tASqatRL
QNLmKtRMJ6MyF/9eAB6RAWFYZPbHbGbMCLTIKac2Z3md5hKo34B4b5yZCKBGbF0W
c9rvqtOe/I5p0ZIj+GNWeWXegKy7U0YwGS21eWd+A9U2MN2SWaLLYXQ5pt4kwxWg
DCG68iOMjxHd4eCP4eUL7tUwl4pV7EhrmuQqjmOEz7oCkCfyOFqxfwEBS4zxtLTU
rpx8q7mWti6eoVirfssEGL8SxF6dK3Jy2HCInh82LM/8l69Cf2UwA29EcEr0HVRX
ZKFoFturW+BvFpW+8UgbKgzghRMwd4hkIgf0ljGkrgdT5ACEG6FrxI7xPztJNZai
05VkK5lSqLeLds/q2ei/UtLNsfn2w4uhVF7efxSlzvd2H8wLdr8z0AS4pSdX6Z6s
nUp+KLwi6j3ZJy0w+f/yl/WLgFJXFB2v7jwQzXceux9aTCJmfoZjeV1dO1jwwYIO
hl+cx94i13HAS6/8OBMZiIhSznaqX/FyAo6PXCwNUCYrzpzECNppoCusSW+svEA3
/E5b66vcoFIPED7mcsD2kmf7WznBrgvl8eb/llk5unTD9q5aYkDq9cIwPzH+37ZF
TWACHA88d2bqabGeU4E+yAE5w8KFeU5Jp7Vgn3/54IyiEvLzi1zamjPNpmkD40M2
6saZTsYQt0bLqE+QCAYYay0a+WDT0Sgu88/w0w7l7JU6TAROjxTJdTbrh+GaAzkP
5fvj5LIyuC7rPM/WzcnEpBEfYbUv7R13GLAcJFwd8Demz2TgL/Yzuffm/MhD9TKL
GTO6AY45uuiYbHLn1T0a8Ns4f9bclD36E7C98QbjAZxd+tppC+DyiXFKAq33XrWX
QWvPozbXkhmjwX9lIfOd9v4H4K2RuPbEXVnftSUHneko3THefg/Onxp1j0D2rjtK
XM0QEBSVUkOPnlHhLWVwDoThcPpoQaQ60f0k4vyoYEydsEhbQ44oKYFnRZeuZzZk
tMPOd+Ei8z1DOJ1uG0+yIHScSkiFFxvrgQ5ecMk5jTyH0HZFlIfRvET1Ixd3EX/m
I5WlIcO4XYGd+Ly/+4wn+IFiGVxq1fRqcZE/Sum5RIjfyUPpyljR8RnmIT5r47fW
UU9FKbZ5/6LrFCFnAT4NWb/6y6jXNyxKD5yDiQ525dH8jfx92cfRtma5NWX1h09z
Pq/aCvfKba/nr8tzSqPCa2+Mxiix8X6e7x2WQmaWUM4ILNyU08LSSAH4wXW7Pw7x
Kj2QE6MTf0UBcvJ60vT+TFrOvKwmE7JOtC5kZKJcbUxXkqPOwU67Wc4rChBCV5HL
mtrJJNmSrNbfL0A/B15gAUuOuZj3vf2kg6YO981LLGG2sJ1RTxj2N72C8N8BuxOk
CkOW2DeLzSTgRSKp7LX5AUX/pXtj261NIGQBFccyXG8S2cBE/F2yg9POMYxEPBzb
n1KLLUBd2rWIdJwsQzP40jHW3gCKae4OwoUefSgNLUGmlDhFJiatT54aOchoxKgp
3/ibG8GD7BZ3DRCJJA4nIkHjIswtZUX4A0cXS5Hi731jmlIlXXbkL+W3LGcSuaN2
shT3sYJShCe/N/p/9bSnERHkke4YWLBVvy0v9YLE8Ne6iijEJ38jfKguM8LICLeC
uMSlS/9tmp2CeRrCl5mGlHSdlxdVAZsj5B2mhUK85rI+Jv1DMNO0lI2opBacS+kC
PYcCQA3lDF4R6m81B5srMjw9sSXs6PlQ42hRXfXHBnlbZR8i8oPyTHSaOEXewHI6
bYjiTwAHVThnMWjBU5WVcfAUs2/lM8q5rHeQymHTsum5bkBnWU3lmkb05FL1/aHc
rWqs+6Ba/avqXfY8sM9H74F2yOFgf1z/yFEv9rjRS8RrUhBY5XKR+dI2B90CLSid
wEMTarXAbcEbjTuArxvwhUjNfhIhcPUy+UsoarjOFFEs32YU+oEXcTOE15aUbH4E
eNOZUbItnDeWe8o7vY5kNoyogCbuYKt3O6B2asAnk647BHxi6hTTT1JGoAl3bwRw
SdJfM0HktQxuVonwmMOgPOiyUwsPuFa9KYoHAFzPSeNXaGYb7f6Brj/4pH5buTU7
RcYYg3ZlmU04gG74MynA+U/71svflAubddfILQes10jRs+k3x7CUcJnofkZNjvKn
v6fBpFs72NGkOk5K64bK0QlgDjifl+wYNwlw6CjBKzLAQ4BaXABnK4xmiE6Tv1Lp
L7GKmCr3nRsHqxv307f6WrWY++pHF5fWOpfIioeEew8S/P6j/Kct4GCWe0WEs9uv
qid0xkBFXExrrqsPvbWt/2VdhLluB9wf+00ubXJmFbPxWPjKQaKwJAyN8vuYbN60
3HuoOYo3zx72vEqPXPyggB3Q79h+RSQyiLhhPGLNh97Scx1uYjkRzedyl0vzNgjC
gGDuV4DHT4XqyWT+qbdAunq5DqDizh/ur38kJ1mkw8AcHsfx9Ve3xKn9xsqu2nyV
s/kfKDCRC203I0PzCRTgF/DVswDodqowiM9yaECT+iP6LI3c+N9zXvz1PVmigTiT
VtdKZ7KxQll0w1E0Jw3Z7CvcUAbd8PUx++0GTgytxPlwwVWcMBdE2O8X88/kDkjt
3H3qMVqREnb6BWM4Y14rrMpEHK6U7iWFA4EHqWXtoCpXO6xWlRkakrUadF1EDyfR
8tAo8QJ3J6IdKT3jf0EXM+FLXdSvU2nlQGXTjMpXhhSdUF08E2XkxK4h1RfXcDR7
YEEcTUEa7dBmR5vNJIdBTlMn69cTVgT8RnP1SasIXu6OdYovx4J02HeQYQOXw2Cb
k+7xrBOulNgxqvJZSyIvzDarrc8PPsCZn4G3q0vWwlWpvhmG3BhEmyVMS9csL6ac
zObSBQdFKnLJ+Jcg/7PZeFp6wyO2wXU57ML3EMl/EOqZWCL+mzuVcYWzLrdhPbSa
45XbWf7rgQydAh+nOTTfAyQxKYBCYWzLbuOEjCpwOWRt7P5ozSrhSQ7vpqwTG9UF
986t53QOH+X+XEVtOEqvPrUQgDC9UowV3wgrsVymA+UTUtM9eWn+kLBSz04W/Iym
jxPL2Tw092B+bS3ciMj1L3Hdi306lNNTSzd0iSNNK6uCCnuxJVQ5ZcflgSRLytaZ
SQEfDTUUuX/TMGKK0wfZfidY6am85Ow5i+GuGffr+3PDZ2FRqAfZ+3Jpm7pGiTiI
VfgYpLHxW4gjvTr8Fepld/uVTXuJ5143fzZnvzgAvUPCeisVe32oR/djcJHUYG3z
z09RfD1xMOxXc56EfFGD/QMQKJacOGhiCUk7MQnDJkAy86KCRiGUfVKHhckfelyd
2sZ1nTqBnMRMdW6/v532o99qBmvj6y81SdouFgpJVbkd4c8CYe39mz3wL85Q8EkH
vHVpYery12Z0pC69ZOHkeq1aX+wrtOSa/YKWC06B6e69XruPUhCeDoPeAU/owkNh
kN3zTvG6cWCeeHc9bn7B5daxBSw3pWOWeL7mURXcwtCTYVxQPfpQGt2b7tVTv8EZ
3nlpbO8wutW2cLq2NWrB29bGMfRXPNbJs/PKTG1SE7MOXKpAYDdjeSal13UlB8K+
5cKss9K6qcQX728eOEbKmVfhVVqZD1XF0TbJlC4ZmUNt47nuoExPa/ktmmZgMrMD
mTQqA8+JlzcxjL1QlL6xR17KrR7JnJ0Fxkw+IiF2lDQB40cbyV3KRY03Y016XVW8
HZlhn0bi07P2Gn6dskqWrGr5peu5wyJHRQssgW/8lPNJQvuDcRT8bTamE+yEqdrC
f+rfGT8JODNxs/KIRTY0Uqvfk+Duc1UlWXvWaZl9leeeAjICDw9dVrvcNaXJMZu5
5wZyQHzR2H0/opD/ubtTFMgywxn9Ch/pC1/PhbBt7O2yp24wyNUN2rFGRHwHfh8e
x1kozuAujGEkMHlDbaMEXpsVM+ZWxQDgNGfgJgCwg1H9iE83tLy7NZFcg3pLwAEZ
iuU0+djBCuADcbZKlYCSUqvQBkwdbEHY/PlBmK7HaC7YEq1kO2UEnfBzMviCXffL
58tXazBspJ4jhM9osQSXbWyBRvgdjStfDkqXRPUYBDaNcJ8IN4oYZtFPVjmCHS7Z
KP1p5I8kVGPLroJHcqWcgJO1lNQZmiEM03m2vzG/7XDE+TAEv4zl9ym3ThZnFIwJ
XcIffKPaRubWqWTpGKYFw90nEpI2X7s6PBzFw+c9eYkQgnZ4Xnpvb03xRho2wRaC
gy4q8albUtpzIkDeswgmpK+Ix3hrBMw58ZcEL0sxuBkckZ3PTf+fWHyHkhCrv4Yf
fQONSkoMrJmD0n7/22+4uswGWhPc1wPgaUkzMthsNqqBh9ZXVvvhQXG5BAz6sIgJ
xX6Pc4NruLxH1w/wGf2UxYBMVIBjEc3SzHoQgnHbH6PhLlqV5wIdYDVcSmirz+xY
B5pu0XMMQKQYdMbNaJjfzFUOZ/CjpHLl7RGSfySTeujSnLGRMq1XxW03vUBP7BVL
3xiFQ4Ejj+jVCIZAxVtz0EfI7gPwSRd2MgrBZ9ObrF3mipwJ827jPnHLFV6yyx/9
hcf1rzzOKr9yTpffxHlbvpQ154wEM4DA/GmNWirKLZPr188LjHaGMSUtqYySJjEy
Ct7V+2mZ98IkiaF0Ck954X2AIYBjAp2WlTwwamFENDX6MTFYJwlU77rwqOzyeHJG
HUS16vIEdMk2C68W0eTBMuFiaNQYb9Ki3WkJLw/eKU5knbI9JbKuUlRwz2QDdvGi
h+Ermykw9/akPX4XAOnzYfVX+8LaWgeWbK4Zvj9ozcJUsyX3mUd61MG3WZcCE5N/
l3KAlDIMtU5XNHv2PJ388CqKZQ4UmhLZenMC9U1W7f1gYbTOTum+6quLfrMBbMJF
JAoTELRSqurW45DBF1vvUWYcH0Bgf1MQOyKey+0Y3OUdC2c1aC5qHbJs4D3+ie2i
smSjj9HGNi3vkIN7ex9ckrYEgEyjNUQ7wWr/tWL8VFPNN/+I2k8es2jUNSzTgj45
MjHIFEqFd8KC5J0g/PEAbAK8E9MokMpjl3jHFaYgJRnDI6GhujaNuTGRR6mKek4a
l/A1MHLoV/vQgtct80Kjfnk4WP3y/vMkQ5oHXxuvRg1txb4vVTz7WP6VWrzVDPGM
f8llVcSc8ynDaqJFqdjqVcsGZGLue8u8ke7Ae+UFylPFItHcpUu5vaxR7hIQOiti
rHwZUCPb+VjBU9PxfV8sK2MIqzUqso8gU9njfbUiVRHv1ANOX54n4I2KKDlwdXeL
kwtnqPso1K5Td+qkDBoK2wc97L/giXu5sFz+ewS4nyCne2VQSgov81ZJRlG6ODV0
ybNIhUchptlp+iw/mSdoUwVd7frAiYzvOuR5zZjixZnj9EyMgw+WADMzIriTgRlT
DG2U30IDcEhToCmvlr4E7CS2YspZMZv24tW2vwV82ecDO6PB2JMQBw6Z3h9x/H3u
8etk7HeUl5hOOZXxgEbhUHp4TL84HHVHSvRcwDNtKMsGeg5zDgfhJMjy4rgpYDzC
vi444scEKQytQogPjJA+7ZftofiWpIFZzPnNvS8kjxuFdEugcQor2tvSk3P+569g
ICgq+c+FwUIr3EzmLacVfL6dzhUaFMRb65zHwnpEl/yOger50c4XQWHL86M4bLdb
Q79QWHASnOtMfPaV+KXUCwgsuiqqLbjLknrAP3efPHqTZL6SO18sN2H4y2Asey5v
tYYctz+7oPHNpMmo7FFeT2/RHfV7FmcQzfzSZJ3+fF2c9g3kvITc8eO27yzRqasx
/sWrv5ng150j3G4ywrvLlszZCARHL3EuEhySfdrXy351NkeN3PMng86XcvXg/pOz
e8qr6V5fTTqU4Qa0WP912VUs3CCfqp5CScdNUVsWDrtD3if3ZPboChMGnOW5bldx
bYIRmfNZJDiu/E+9Jv5yktfd2WagAB/TVB3TCOrJ2hZyO2wrJJXjX94+vNumj/zQ
F5ecFd4x2AVchitSFdUwEy10+234wvSHa8RroDNKD3P76dJWFXxrcxZkzjnd2y26
JU7G+ltuz/xCEae68U7M58dAP9ntAa6/CBCh9SH35ajCz+h7NzdFtMdA6oAj/02e
GqG5a+7ZdSRPzKjNRpEg8I4R8PLBNe8Tsb5Vg7PChLbQrsui/QIjkrHXKutbUi47
akiFqOYxU1zh/QHXH7/Ktehis3iVZRJphAS94Knoji7kM4uCovGdqzEO54Sx/66q
U5aIIV1o1WDd4+j4oxo4E3z0iI/4JD1X8mp8E1dK+FHBBC/XZIsvg7IYOG5HghbG
KR+8i2aJNEQNnqMWfl5qltgDbta7eS8qk1UAbZbit3pwJAHTSvD5vPYpdVAL1C7F
xs9d0C86R75Gmnwkcnm4eCKctJiL1I8U5LYuhloZxjjgMclTx6oIxyOrJAYn4nPC
sPIBbLDGq3BMHUOAr9I2bMF/YSERzJJDTvhQx+MXE5K62pakwJ85vJK3ItuIA5MR
AEkjmzDBJqkcctHJpTXIrGEV23pSp6OPBSiFZQS6MsQnZWAokoOS4oeFK7l02IdJ
qkrCssy7Ha0348tXRWnGjepB2Y4WLMTa03A6wLuzO8U+mFuzFq00Gf8PHlZxuAT+
IYG7kn5Q2ybCqKhx3VDzWeagyD+EioApdq5w241Nduc1k/vmoDDOn/5swxWEbip1
I/Ub0833xx38w4K8ot+IAkyYi+qHDG8DFocz3c8493kqA2qJJQz6tib1z6KZVVCH
uMl2RGAl5K8mzRxKVtr5IAYjIyC1463l2pN4T+v1nDK3LS8/KWx3nw1W/+ockOFl
LVhcm3set9zFN3BpoxJ4GoaocpxLPgSI6SmxPx+zFCjIymRLK9nAsNoGyBC69qih
rVEqT2VnffsY3QjOB7hwYBvISXi9mvw7G4fCzoREDb7pMSNjf3rG+yyL2/IyyMzw
qS2RzSBPFBi7X5kv9+DkB2UjxjQ0ymtalDt8Qz5LdCLBrXwZ1LEwxivdJsJZDUBQ
N9cmmKcaT0e3RC7geK4x4Xdz091E91s555TvqEKkNrx2tcAX9Ew/qOdRzRi8DBsv
qxeW/KiH1424j83q2FlljV2fbqFTSVXM88MxSpyMkiWH30nvzSf+JhbCbAJDvlfv
cjxphzaDOVdb1h6ZItGOHeTWugFG6wfB9JBmhLgwwTsb6mc+nORVOAYHhFSfRIs5
Wy1fW6LeKAX5iGMykyha/L8NHFnbITRo2RgHbDs3O+m+Y7AqZhb55hwTcIFjDdM3
G71JzOUlSylTs035zTS1RehspI8I7w7Wv+6v7iIPZstcrHrxrDehxmbDoMb+utJ8
jdLuyjHkTeAwuybQxPLHn/1X6DTyZ3u3pZR9FmpnKWwZyuEnptH2bnwTEgN19GxT
bxIclnLkGyrgwf5Z/RhcxIpvhX/9cnLCCwTJkbfdBY+98F4h5g00lF2xIsIxlIqR
mNHh4zNQ/ph+m/OKCaSoGo66L1uiOWdf+Xxd8wPsMVn6swZyefeoriUV/mdtJE8+
oKKKw7NxIK00C1/CQ0KY0bRQyuSgylm1VW2HkB8SD3MT0myC5n3NHXeqwCSflaEq
3b/dakSo0mKfALVi4pXvkm68F80p+KW8X/DtfKsABLa0srlHRSFCa0RJIOtNGPZa
gmhdnhMkl6xvenEphuQHK708TxMWROjg+GEeGJRcPp3gR0bGzleZ1JjoDZKkbPvh
n7vdImb5SOZ+NDbo+8znkRrhOTwhHctQ68jhVBqGi9xXZyIbd44ztEIBgl/X4JmM
mNr++wfHfcGKl5TnR8/Jm0M1JXgyWVKc3T3pxUYy4Z0+cC3nJQFpHkUcKLKMsmd+
g4DwOAjfu9MfEMWSGU2ywbpmtrRXgcJJlH3kbnXXPIsPemrDFKlTSK9X1Db7448U
NLtMUYMwy/nkMzrOvsD2XSodJcpyaotwsdfmaC7vZMbiCwuiFF0qsPGDHjK8bSOI
p8P4BvM9jzhgsbWt9cGPrPqaqckrdGC9oDkSeXfPG4BPHUbYXK/XwFsUABPTxEKH
+vVB/arqfpXaTh6Uxy1rySVkD3MYn1n1qRAHcx4OEbd1P4L3FV/Bm74JSzL7AJ1M
UooC9xLTHDWZKB6g+waDixViFd+4Wg56II8nNAwD29SsqThlGTUAisuHA9cc6opx
/6WS2B79Ye5lWDPS/DbUeFyDbhPdp9N/WlcFxkCSjxOqyH9QmI4ZW9kBPmhx82XR
DlrFmVYa35I42xoYdWNGiSh2zwDjr4ix6OUgyS/BKWK+WS3h5CxbtZDzBTgz5D3P
oe+Q7T4iQ3FUvQFcqAPPZcDlLpVS9FHwVWfArXx6V/+uIY3h3SZ95uU0LEKp0mkl
oUhenu+0VsV6zwVJhRX7mFNSA64etidPZL7UbwF+yM/gl2NTpWtrBMmPPKNtY4mA
GGNGe/PKpX6xPhakS3PX3w/hdIu2rdogVX4OjvC8vsX9Extg2cBEyuj7YzfrYHpi
emgUCWhAxAdDANRANsFoyyFQnx48n8eojKsTX90JTDWFQAUqcmWDm7iAQ5CHzk8n
mnoQNsLeV0nxwg/nyPzLZTKHS3GCXpB0sw+ExobgB0j3zgPquZqJwRwumawqzBBT
cVr80QFR2o1zRhQ8kocur2ZkBeek35eHCUkmZagSaC7hwdBfzsAHHLtRUgFNZIHX
9iofVag7ZAhoZ+2coPXItkM8Uqazj2w1wdkKnN4wpxw/GIy/G5+SYtJw/KLbxBGq
8rh3Z8w8MV6Pn5tb2a/8vTJgzRbcbGmHe0g992HRD9aOprtSOqk2KJMsS6L5O+IK
HYUikPJxdWv7omewpWyR6n/TvQ63L6at4/lQs5COV+Lir0Sg4nZLOS/cWj5grTaL
AK9FvlI7AAgCxELIsNhSGQjb6TfHgPuCasK1fvcEqdNrlXD5agfhneNTMn9hMOaP
IHuOMPl/dwGK812GOwpAS2YeCAOYWBCCM+dZobMMS5RqtG+4NseKx4dYQBHJOoTo
VqiHOR1NMCL0wwb9mcMcn1ZN9oDrwRmvAbpsFQfXidONyr07g/QTf+p6ld5mtmD4
B35GrURYeRYLCd5H5RBxtY4S3MTOINxE2AfzuEQXh912wJ/Iv7zdpjLNv8PDsS+5
LV9lwGggmGh50TxrIMvhuP2igGFoOTED+6gqrNv0Z+VXVCTwTljI8RhUBW5B8sVm
12TNfrdHGEPBJ0futzguZHs0Lt1G03Qrun8wvUaVWXE/uJLVQ1UCAWi0hjsja61B
bL4esZa5wfkM/GzkGJ1Aul1Y2CV74fuKlOlr3nuFS2QUQ9cpf2o0nwUMDodkykxM
F9KqrMpLeamHraDJchY20soI6Obxk3judBXEZTI6XLRjKZA5EntJR2jLQygcdL8n
ChIb3vFTrKg4Sk62twNMsBs+Pg+nQceF/UpY72LoeWPaEJANIV5gQzdVSFih4qDS
bwhvsnFTk9aswap3EXbU/6giR9CYuhgfmM61BJ6xmdHBphFPmZ1C2bL5Awfyf2dn
EISf2W2w7oO5QDfXjRVXf/yUMf34lX9nBbS3N27k24JvnkXF1HnzNnOp11ed9nwT
76rk+1UERbnacRMbVXuxPmOS0UakphcPSvByaossBGAI+v+2+8KCq/+hyO9q5jFn
/H8uLx442BgDORk80AJYP+u7AZCwLBUNsRCbYiTUyNsS+JNDCwkhkL8mklzfYUb5
zFsGeINLQ+kZkrg+AMmT+eeLKlTptitcWbKcXtmGEW4Z3Q5+ZV0qucVVOzc8RZpE
tsIhErTxhyEkcUsnOzlx1csXHZfGr+ywqyblgYs5dtY9OqhkSLJAI7kq/DlKvo60
ZD0YQHzqf7ZwF+mzSCzHuPt5gkYvz9Yf3HJlCFR1SqNKrJFOK5JRS9PYILHE1XyN
mo9xfkk56XR5jW3Juk8NzWSzpizTxfbQ0tTVgXssvPC+9tx3KvH58yAB3YhMk+Le
jAUICQZY2hWNB4ilKAiwgdv7QDY/hGmXgEFT2zcZ8vD+nrzNmKBtoY3L+v0g1Efo
mb4GvFgoT2h24WKUlcgs4ley44II7k82vtvT3kv3s2X+bTcC9kXL1Rlir9kv1APH
Sq0H0Cuq3WKRUDmdVBhn5kBwmLT2rsFpCuJMQA1QmD9oQ6tNnacWXIS9PJpfZBhe
/CkHd1pjs2cunXSOhxclNGncCJAS5DzMLsglbZorfpX3wtzo/RY0K7nTFbRmJY+d
0esveqbghuVNd7t4ii03kkDlKjA8Bjuc8N4WLjJ9FohP1ilG4Wh4huWZj8Vguw3g
c8FmLl8ZcchwGPnJiTujsttc8mt8HtsSUZfxVnLKZffeaW1j958GSqDBHHvJWTMv
vAP5jQM2hC+bx7oJon7c8lvG1fKq/Paq4X3rfFDQ+YuJoYwex5crW3VGieMfZs4/
dzHDQ8xrxJCysfv3FtuKpxo/qfPSAVyrrDO8kscfVNiDpLPcvgcT6ROO6GzVPTp2
S7EXGmkqmkY+ex4q8MN4iqaUvxrzf0ZsSDJceHM5y8VwxQxQQnidfPa4J1FpXstl
WEdnaf5YQJVV+CDtxPZc9nAe7uIjRPDqyihKXdF5P/F6tsZkzWp6nmyGd+3dHEHL
09eAi5LS4B/v/NW18Qp0jfFQb39IVyZeNB8VQbKTFzq/8cChfXl+v2oDVH746vus
JNONuo+/KLGfkw6L8d/qDJ3c4zgESgZxE48lCmdt8vbMd7xWXy5s49w+G2iIiQDc
4SF/0+NruswvL+Y/NfApKnesuxmITIXCwb+52p9X6xty/u0rqkkZavq3z2tc7aJo
mWAdp+uRtMSHk+T+btGy0MwVy9fP583XcWgOPUa8EJoOX2bAn02vcY7MNZuSqtWN
7n5+OTtwb0DnJtVk3e2rgvgx3sZoDMc8H1Qr+Ok1sPLxjlD5TfhG8Qii3mAs60m9
aRUijmYaAogYAY0tE4DkR9lwv93BofIukZAA3Ct2Yw/ilDpoigvqUhOZpXg72svk
mT7Ro+PuWM9I0ZYzbqNuBVZhgqyAJIxSTM5XR/sxfNB2faYSop0I+hj+7g5V7mum
luJftP2dAWUAIE0V7YxLWtgmXos+HFxtRFXnsPhhcmckBkZMJYL6eQ00Vnd9jtnh
3JVQHEplrCTUfOLM2OcTXSsz2hGVJwNfnSCcvY7iZAxSPFgTM1TJhPmBRhtJ5HxI
elbd85UldCsQSmsAVUOZiyKm+07bzz2Uydmbz+93Vi58vZw+iRSH/QJ2iunhOE0Z
w9r24AYfO7z4xRM0jilVDSCB/gqdQzKeEqt9ZCyvvY3KAqIdFkYVSrZlNR2xJiwH
+PKKTIvc+MJ9q59gQENlKLaG2+8Z+KLVgzhS/T3wfFr3wDHB4q8HQOK76Oivhc4n
J64fbCCr50RWOwjUsG8x4Ftnc2+DK/2/IsUOCElv8oMNmq0+6VrSbJS7BN72CoIy
sOLH0D4kOQZfZ68BU1Cgj+QcpeJB4ADI9fax72v8S40vE9mNUTriDcZfP2YTP+/m
6/s7WpsAb26gInNNNzPpiRTkT+rn50fOhSkDUyxIns1uh8MA8TRS9Ins/D6vrjPm
RBYJy+ZnZBB3cqRDefXm/VDyUHCpe9TfhBR8ArXUtoCEclPMCk9OQl9KFcuVHRVP
Rhdlbvx+ksA30BofIC4uIyq5qNVUYzM3jPxZCvsQixz+SgaEQhK6cHPHcVFfO7Di
0M/z2IY5nKHlXJLbGud8iRQ/jAJwJgl10znzZa5Ud1yCD9k2Dm7yW9GfgUjQWS3h
0Ukec7HU1eR6f2yDlJ2yHsInIQj6tKUhPsKsDxoDEZf1/ALeMSyEtcSM6kfs+x0S
P2BsZ2bCSW26UmVVNjSLhQ/LmBhXyjYd+zpxWrEajD9sJM0q5FRahhPFlPptJFMR
Py0WRHTwp1VTPokDAUL0qIzlYjd1UjiTLSbQ/vsBOtnjRpwGD8WE3P822KhbvQzU
Gsp+xFZjanF0pcbpZ5CFYAkMp5zxtFy2cSc9fhxwfjncIUwIhMjgCz92J4QnKkd8
1Re3K+PKBhzgVuQ5l+GvVXT+r33BxcqxCncnRXxmO/wn9jN1P06yGqzKQIsfVHTW
3078aAyjdqsyW2mmwp2k0l2ri6ZNye3w47d4n+DeAZB6uRNKyosZn9qOWIQ9T2CJ
nttQ4QmTb+WSXfyRCF2LySdxpcscKHLeqwgIG9O8i+AagoS7lsv0308P8Gzru2HJ
okd2Y2bZgHVa5Lm+vJddnY9v68qGzdnvQPaJRpypO1FeMWx7WgA8TbHEAv9Lm1Wo
xeCp4ixFEsCAPGbjpsg8IsGVDS70jwmA/MuzeXJtctAE348Svra5wjVAntLJkNTJ
tFrPDxeBmZZF8L6NDy9LB6GCirmSOACD0yfES/Jkm/pYs8ZldUCXhm/cwuJtJxLo
nqoHWE4Bo5czK0+BZyTQx/boF+JEHEP3VOolBq7A3vXWG7QmJPTa4nO21P5eKbT1
x96C1Mp/NMCUdRRQ7M5v2NMwGZ8N5PTO2b/YzkNOZfGZzKcpzTk3Prj/tp96Ub+g
qccN6kBl5snRvk2wo0o0fH5bBz/AwuNgQeeFirrtVbeTBdIXIH7lHx4rJdbxu9rA
6wqU+a63EexI1rE2BU/dUTRL8+m5QcLSkQ6TjqPIMu4ppv5FNlR3X6Xno5ue2EFt
YYsoufAvMuCSdP89KLgUbvsZjhExttLYIILrAdsPa1b87ilTvz9lwiAU+CFh2xv7
Ejh0/8tlR/tzq/dFgA4Nt0Gjw61YxVV5/PvESBCFkjLDXiFHKaoVNLM7thhCBC5o
WxeFYaK+L/eRs/UvHC0Ze08sEOwsndzSB0S0nx8etqukkBZZWDHtIqWauDRpfHhQ
l0JLUGjTnxjIwS0kU9M4GxXSacbkPMdfXBKXFgGywH38bTLP7jGFAEyhLx2ZAI5T
CwK/Wub3ca01TnyYAWNyXPYo4StdimeivazYEgZ9Ut7YcJy2FTZoQy6yt4cpdfWI
wEn2fmsvY//wjOFxibkgsLpuvxwC22x7NbHx7DbrzTkNLt2Q274JsnWlAEl+esMG
1rJJdukhVpdttle5ATRMMhXdZEfKUbg5GPHjIjWiw1hUVlmNWtB8uFQ2NvTmwROB
7goU6XgmI4dKT+r+kzhO7/dPv83FH/y2eLPMGGKmj1kUtmHET/vnfCh9Cu7LTVvQ
UjTghlEyv8GiKX0usgED2vwvodf7I+vCiyHvWkesYEq7qynUSaa1h43uN7OG9aj7
9S4g7niTFwSC909g3MZnsrZqTD64lwepp9LZ8pvfToB++PygBOE9rMsdl9l0KkQ0
wE10Pmg2f6n+Wz4O01ziIOR+/V+UMwNYTQpIQ22Ed5MTtXM8HSLEcNMfjRjBf2eV
wAX5067QQrkhRRy61bhNPdduz3vmPO5FB62KO+7v25VHZmYBVpg8YNL5nmK9auaU
XqvD09Bdusrwy7cNYNVqF+lnPtsoNjlD9VtuSwybdaMyDfrZeuiTRdGq+6DPfRM0
HPn6signooiXdo1M1esAjfX+KvoOAOnGQu49ewTK29BNHjLbZ+DQSZ3kVlq7nnbu
JheQLtNjTcdizfXFnxmCu+y5XiLXOA9ZnV66HbkpytztLIa7UWByw/yNa4r3NPe+
lmxb87ja6JgDewHJT4IDg5pi/CztBWu5mruhtjn6d9hkWDaiJxiHn1fNk2OLK4Pn
dClDys6TFO5rrma9NEURbbQNk2+jbteQXwRtFe3AHy4HCmbEeM88Jx8PqRPTgWhd
8aNu7Sgi0SEe/nGtTkhvYeJVvIVbL/Sv3P79H9erm4dTmAb1wCk841tkUAliI3th
TZ+g0WOSobjr6s0Vx/Em+92CJ8f5rHamTC+uDcR/dIiTx9bOR6mMzfA2jQOhz2iK
P+796twJZw0GtSmjsGtPtzZxg+W6dtKiANm4PWL1wf4ciEWQ8BZAEYqron83WvlV
bJ/3wcpSx5mAN8Hz5m5ZySk/OwyhBHPynVrdHXg60ml1lx/3c4CEXqwUMgve2OQD
WKGqIrAXZU5gaTTBB9B+PCrWFlsQo/5ouSlSTMGNFAyNM+z+0yGKrr/S0QqTMj2N
ndnFyHmT98cReztsgm/FUj0O2We3inEpTnI82fo7CIr/MR+evcINHQqf2F68m7NS
N/03Ves8YsAWBqC9+PtM7+MK1fgMDKk48eycoKyDpvXMeQAuKkUe5WZOS/kI5FFL
bh9M8JPc8Pl0jOW2GPj/sNyrxz1uws66iQYH+3TuIf9Z74lYIUngki2jC152d2SG
3AAtVKnYSbFJ2uUIP6RhARKWRl0pQgQ22ggFnQPngXGCf2/Er2SjkWQR/mNfXV9x
fML2SUOE01RVTUpJMoqYkgl/n7hJ9cnMe4PHLV3/fUJ5r5lMBb9EDxzDcTuJw+SY
aWxN2UkTRJW0zcMwTPQrwkgcon/ShXLqf9LF6RSDBFGrtSGO7n2iLX0d1XWW0xp+
2c6xT1udPkjEQfOnPPsTkCC4WCoFzJuc1W33cScsEM2/9MWV5a2ik9UcBT9J3TtE
tmXBCTt4Jg1/Pd6h9YWbAeJeoGVdAfG0R5JAMxnvGjnbC9TNeQtCUnKLXxTpqkdS
9d/SCESAQ2vwKBnXVjd61Is3rSHZV7mhFJV55Er2U38mlhf/7osDStawT9ZEWdeN
/Fseg8DAQELpKk6d14e2E9DNYX0ELxC17wzJEHUta4G0vDOC+/OVkvm3+nF41Sei
HwP9VJNdZcS4/R35S6Z8z016O+HJhZiNXCAZ0aNIxV7H3kQGq8FwZ5D3Z/3PdRXr
ZK7glZTNTuo9Vd8NqNcYfLFKEeFl67Z1Yyveux//TVL1qUtaYDbHopuIdugcqXYi
CCBMPhbLpE1qYqAFr8ipGQnuhTC9AApfoF+xnk2inEMzHjymteDB30w5wHAZARve
LYehPTjMR3nHeZyRjqOGeekKU/3sd7mm8xXyuJWbLPc9I77a+Fv6CbkwGXvBe8Sc
eVu7oRmCt6dIqWvSGERomtKgqC9Spm0A15PSAehDgJ5R8tlbxA9gX7P0DMrMdHbg
qUqcWhGiTfpY1rsxOgyWyLLTqiI/FpfLkJ4JBNcQE2F5LM+sy0pJiDFy8PtpGFbd
LJ61loJSIQnoLfCBIiBQlgJfZ6E+fQ3BLMw9dKMxpvO7hHS4/LfD/g0/yj7Tlt+5
QvcyJBjMtmu5EdsA60OtLv2+U/wTiQORrkdbMht+3jE4btWPOKOljeBIWrohLRE4
qpSkNQXFMqgxNLBQ/FVXU9EseNx6lSyfm71UqFUmoXuWH9gMQF7I7B9QvwGdOjTf
QrMSdOO1RWSGoTRISYqdKyGEH77Q0M+2DA48DSfJZySYltlWnFRbPbxSuILR5683
hXyk04RIESwWBl84NAVxJfntfDMrFbM6dTfrL4jnR9413jFtWR01aK7sNZyyW5Ss
AcZQCZnMrOC673KpNJeE0j4zK8UJr4gPtA6mLX4Qja8jXQVInA4m38WZRc+o/ZLV
bqMOySS/+Yluc5sKKxAFtWBJCIMnPcMQWQs310fbIgL2UuwQfI2yvJGkKVN4VAUw
GuMOjDwnbTvUZa3y8YfXT2dDJSPOjt2wdzrgIYE2U0gfpRCqqcW8ChcMmJzMX95v
rz4PNfJJ43ME6cj/TSEgDnAFMvo6uedwdKewcsVLY39mldrXMGKKb/Brz7wCfIXD
vvkeEG2nTyenBBTztGDy2ISe8Y0aU4xMEdiYnvel43BFypUIZtRybXXBLx/2hUJ8
kRa0puKVubMBD48yrJHZNiaLB8LNjEM28QO+SxajwvBBvu/Xg0KyNUiwxCSMpsMf
SupHm0uvedUonL/24g2cAIgE66yf6LsfXEhKUrTfBtmgXNEcIKvIEaE1qGa4aoSJ
2PkRWUFyftgGm6fRj3ypXU/dDlHv0Rl85sbcZvQwYt8zskaHnCbZ5wG7LWjhx2mB
wZ0nfBv9QHTvnNNAECioY8HNt026szLMPxurQZVE6x+bYO2AEXLDUH1Ab6dSGHG1
Tf4ZP0r+G/yXoWBIlxhm+ex7dC/wE56hli+AonJUUSyn23zBXnB9QPz1iWoxTgpp
3vKKzw+0ybVkDFHOnjCzlfy2iyByoYCSegvqIfV1OkTRk0AwciGqtpqo17+BbEL/
ViIVV5slkSNfrUwveRSkg0y3mrAhgOehafAUE/JOpLW0euL55hMAm0//BgSq/8+C
/tVqZpW38P162ypN3H/iLHiNGbYPf6a8f8Sve9YgUziwejTHuKwZg2Xt7eTJwzHq
xNFllGPGCqF1JHOum1y59bywLtJXyfOvB47wwAKj2S7PH7f90twTNCR3JDSuRehi
hgEUKYboPdNrB1Z2hGPBsxcENprNdjwUe6H02X6AqwyTnZWnPRBsPFJBlkGXukdp
hrhrCbAXWymqkPWqtEeze8WIPcqYTLrLVXPxFXLsdRpi/bNH87k1JGhZUC+B4R4I
wHbRE424svC5aPwT2PvaYhm5H0xI0OZI/2MYZu0CxACr/7zS0jTad9Uv/PCNnjCA
/aZX3MPXQLV39r2yd5ZqmcRQL7ibCCy/6vGS3ZYro8tw0yUrnCLGJJKsnJBTglMT
gehvWJn2olGPMEo6ZOT7A3JD5cH7CHxlhgowW6uMBo/+OVB8qahAxtOjgfV72WtO
WjoV+gphsEc22IiY2CEnHQ6TNBgQJrM8saYrc3QgszVv7NY8Cq+y3ATDt0shfQ6G
cfMpYdrXqnKf+vYayqjTmzVHiin8kndBftKoh95/89RWNg97pTyoBVpfPHqfYvpi
aZb7OuIguc3irz58Ln6yaoLK+D84IjnM+tV9VeMzqqm4FN8nNLxLHrkBd+9RMm5b
ASkBu0S/FF7ErTN9A7ZqctMG+5ZEjF0/7Uevm5/XN3RihIA5kYlJzaDOhmo8MBSn
jiRziK8mLSEickAU626MH2OJLhPhucm8W/+0JR906glJkG/8bmHVgy3LiggpasMM
FuaKRT/nCGDJQ9JPnt6wez9lR0RCcflr++kSV8elyUxsAhKvMLSdn2VJ15sCDhqr
nvVZA6A+3Wcr/ejrPVZkH6VTGMMN1qwEhg4PjCwZeUa2Lef9d1ZzEm8MxmGPPNEg
XXStPsFm1V1ymqY1Vvp8bE3pLwctrWjwt+NxK3kQfVv6k3VlVigsPZxGQ2YkurpW
qXqphY6TnW+aqd9MLEl/6jRlH/vCXbbAZH7qEuii52q7dVTtMhdRFu2IcbxZieYu
sd6ygxvi5lNGYhdcPUVzcB2IHHMPrWNMjVdWIrUXMVTEzXbQQCUihH7P1I8jd9Kw
9AuPawqMlwnRrQlfEaPH4TBSfF7oh4xHP5YMLvd0wFXQqGfrIUOwxs180TiVJMR+
rOsx/vD79Fpf6rA/y6V4g2jKBslmnftMX3A041SC+2S93IH3TvRlPTn0HasA3Q47
Uc4KyEn1IH7p4r7/IYzQngKYt2fgRq/KonfVq45TfqzEbYjOcTbxdAVbGZmG9a3r
hYY2jaqCMOahwg84UuWU+Q8hEHPFpDpimr7wtEaedU8zA+b3dAIo8B7gcR1Ln2tA
Rqg90XAcQh7h1XmX33tcUhjya3X3UIaVTiKaAz7iuPhpqiaiMDpfvX+Q080xHpY1
Q8CNANGzZwclYCD1mskID8blwWeSllfmN1ecAujXJsu3qBXejAn4cQgZ/CzYUdl2
DZ1+4uUT7qkaMN2ZFjC7Bx2GgSI4xzDK6sw5BYapCdSU7jim9g0ifyvbHarU7Zjf
dWpT/rbU6o6JUTfN5/Tx7S9MxHjW7uAwEVXvpCxVXHVzOPqf+BzGjAcl3vIdJU9D
CDtBgPDFd9TwAZoW/0u7JXv4jF9rmw+uiwGSourCAk61sc0oFJu/qso5qm6uHKT/
kdxrGYJsiDCMxEcxaXeLTLMqUZK9d9EZzilot1Bzlzft2CTJAy6nwEdTNWzfC7rz
B87EwJ06dvSUKJ2nUdJZM3i6Xhr5aTbEcBRJHQ44rhTvWJ9U4jiM99Cf4OHXIWpO
MaVReHdhd5ZbsZM0xV7+vC6dKn7AWoIm4b8PzHz4eDb8I4HANni4J+18DXPVKINk
focCjHSnfeUN6WwYQEGcjRzEzfabfVxTFMQbbgjJR3ozeSyDUUa2lIeAJKd4IfAq
7V6SIRUW99PKPVQil3ib8Jy6z6VMBHeFrSrfc3cX1mmd7s0gPKYjhiiiIHn365ce
pSMA4FWZ8XQDpu1dqtXWGScfqyMbfS1kBqgOtU6F/ERdLsvxYf+NKa00UsEcgnax
xW3SpbaytOGw6E6A5ztMChxg/GOAu3bhNmENKPYD0iItxAG73paT/VBGCqI0YhNK
hHclPx+/YWxClhBODcsxSi5bGkNqYXpgNVR9gVsLgSbabdu7KXduGZr0RWlg0y8h
zzFH4eXB26EW7dnOMOYnbPqp5+hEWVk4pZ1BWR0YFYiqjqsuObXN2umfDXR+kHTu
OgzZz/nWA7UdvRp5Oez5ycAjdEsLmlEqnpTk6lZuIKCXKMA3iWMuFTh5TU74Hmt1
rAbNcBPiZKo3twnQQeps1KX6cIyzdx+v1jy+mGLBaz0Z821Nu/BsvbQycu/F8MjC
d8vtMyXpOXyTnQKhk9Ee6DBHWacjf5rETK6AcTjkgGYBKPBM/zCOFgT1WDK/yL7h
kLaxlMI0K8fmXUU77dins8irv2hGsmNho4C+QDdSlqrA0PpddwMly0TBVKmFhbGt
Xnuy/Bs40dhstg7Ul3CvdIZ7z05DIPYo5ce/8Sr7zbH54QGoLvYBEEWkOR99Zcko
whjFY6qjSA/8Los3QmriS5cq9tzWQX0MtwvjRQ1Hc4uGDzbdKG38GG8DcwAyXEis
qaRyykM/nYV3pF2IhcHDCLsBWsOqaywJI5HYW6v2gPOUcdV8fmmKPYAaDp0uO2DP
g2aouSRYe8nAkhlOKcpgeXRCWsQGeYko3JYAT/q/cLUrPYyGUDFCV1Hv7aWEOzlO
S9fbRKI0NQoKDLVsFJWDe3lNIvr7rrfHLKcwOf51QSuhutC9FBIAoifnvvpb7Nos
BY8iC8A7Xc4mNjBDPyVbMV5b0C/Q4yXBUz0zKJ9Wc+XHLicbnDcojtvdGbACONuk
Cd3qPkdSRNKPJE+bsl39YiJTaSUJH2O4Wk4KYq2Z9FW/JIROMyZ+t5SWGU0gg4GX
EqLxpXE1PaJE8tRecjM4T5WxRxO6u/s0i4vAzmlsIHakrIwzqm5XhS5Jdg+rCFda
AZrz/BtjAytawWBReMiIqty7CE9Zpr2Nk6rqedYLPCznEjS9xAovd2QJKz60YxhZ
9Ye0YzIRojrqw6tUqEw+FKiD7Ae3G0rX+u2CSup7Nxk649kAictVOjIZdbee8k8i
KtCANHrU7Yi3QZHFxX70nkJv1mbzQW+Z/vkbtMPvi8sBa9bsuBQTISDZruO58vad
OsG79Gn0NbmEbKum8Po1g8XsxvAZdyRHL+WuY8gWdXfHeS56furq5id0QIjN+Buj
jC/z8770aJY+9wcbJpjy5jpuXaVVRLs5779AXiajIv0+lRRzP8O72Xb1fO3oJ10+
GAZdU2HGFuuKVeBSwW32YFE4e6lZHDzK6m3awFroJ6Iv9xFqvfRIaj3xsdH+mS2z
Hj53j2qLHRXL9Ozm/na+48+gvKn3PDCi7llya1U+/kotIFo+EpM2ulMO161a0pyd
DuhXqLox4D1mZWvQdPYaBTFzSsZXKwD6MOrCryM3ccjmJq99RiaxFA36lHlezvxC
xzahSQmFsyxeB5TsxKMH/C9kE9XHt/U6AF0xq9j3nagTQW90AN+3hyrSztTsvPUD
4Xv3xhn8t8NBb6qCfQivbQVm+amx1xPKBXKLKvE3CcHDBnww9bGwy8SVgNQ6fzqZ
4Mq8y/VFzs6IcYtruOCPAepKhEZyGV/T3Phr2+o+65crTw1DKL830Jeevh0CBeW2
U++IDFBQ69oLY6+eBUfAjBk9OUfLx4OxRhwgMdbCjFMNllq0i7WDtaHVwX09nwF6
cnB5ArWRGEBorUvzySKx3aRW8UrWx6ItE49vWszJ1kQ5Y7RTWcifVmIGhvJrWZ8l
md7zaq2EgiQWnmF3MKRkuQaLlbdcC6P9Z2PtEFTThuzxmEhJuSAkgxKm+6iYw5sF
NMg/JwSESOTATBJzzZ1baABnl11DB6QojvaLM6F6kjRildoPtVZIkdgalZzz6yc2
SyJk2/aMx3u2//wL9ODXMNPU50McHH3KitaWA531cmYb3//aa7kwd94PZ5uHkxRF
K3KKZp9qpd+I4ABe/3qLUttLt5P38dOMroFdHEiIXWZW3YAOV9O7Dpw/tkZZQ/8A
JWAMxbgjSVlsLhdObGSPdRYbgUpvXB7wXcROTu3H0JBZenz58RQfCaewrKgEKPbN
vVstvRzAN5kNAj7i9JjgZaHUG7q8brfv0fKwe0sgNeLDM9jFTu+6LXRrPrV+FNzS
wFE0xta6joaDKp8T+4H6eASWk7UeCbdAj0ZpHFXL6FKZX5kz8hCFQmPy1GSO9Osr
IiaviqbvVDI8MuII7H9RJbvtmyU9X3JEYDyIm+sbE0p6TYukGtm7XQ3Qb0ptpXgU
8ni0/mS6aocZLZbg6Lq+UOowf4G3Mfy+7uw6mkui0LM7UGyZRktoB7Y8h5KgFvzw
nvvEaLc/J1tIMTeAWGY6lAlYE8fMcC8LF5PDtcokSt96rxy8M2m5qvIDsMDZ7Hmu
xpvoRrUJQnTsoc2QYRpR7GzDplJ5/ezf/pPr4otuAmUUQcnrhXUJiIDZD0WwWn+b
WHud0jmB+yd79P9gmJuZGoMEShaAPb5oSDYnn9ah/TCMH5ho+qnBtjRO1TGWuia8
Q7moVlcVlMb44EbdXNZ6idy0MNxCh0gLn4fAXuLqx2kH+504Tw5qb5DXrpUhNs3m
dVWiY5qOw3dFL/KnEM6Bebpy020nKhKA1zR/W8qIoWLS0ANtdpnaLnPEJ273BKXB
z/152qI7THCqQCAOU2epXca7O4ppTl4EOPQkVFukpyeSZ1HMYI8Fn2ksWk+J5xXr
8EeIA2a2oWOuQlEgUGznkLxyjR0jiGUMGJTGoIZOKqs3ANyBdcY221OPA4UDDlsc
WPYtynKZ8sUe7njNAe0UJZVu98QBfNe2ZYTMHa4F6egH8qAsLqihLka0fVfAK8x4
fpgqW9aCBAcbkz7yQaTeVUukw2E5aU2v+JXWEk6GBdvGhPlVTySduF54vQxS0I8n
h53fMacKIO8xyHmYtPSPKkj735HbFy5MtW9EXZLqOAiFH+MkDOavrK/aeHlBffPr
exj6s/aT3ktrlZfBE8jfkxzr07xcy/4XftFEoCs1KGeGQxrOlwerbwcd8mnCIWYI
3supr4BiIRX+Kvf+ctOhSBkDaeTlV2vFDZqEHYFzHWx/5x5YebQvU6jOWdc8YjwH
a8jzCu/A2w9EjE8vcNSAQ8gx4XQHOI3GV5LOGAxKRPFtvO/BHOSfiYhDmD0naIA3
jAVXNhuzzNrm/gBOqQXj5Pky1d4gK1keESSchu6sARCVLvMnTmSOJI2FtMOgKq4f
D+lquHsHH6wa67yCBI9Zeg1DHK2kQROCLtBskGi5lsqOiNXz7QqMN7VACBgs02Jc
Ikma87Y1os4GgcDnAilriLvAha3kvev4eKCsRPHc30n9J2SkizazZj7UufowtTv2
dbvZMegt1vg+UXu200+NWqbOvEakRp3dUsXMmahF7uEND0/CXNl/ZoOFEC/uv7qQ
zTNrd7PHB34OJ4gwpU+p1UvX7qgRxm6IvBZ/V4E+dzoRhfVzwKq1BxpfNkN5T20n
JdC+Ohdkdw84Xnm8jqR3pga4P4hxRChA6G9qxI4MiindQ4nWE/u3PqDoItSViBfO
NnHpKZNCDGUt0gEOdOjl/YGuzDq9d4H8Emkz/3BdNCQ6AfDJBohDCi83HielcJyZ
hhTXT5kZ0KVU07+hbJKp4uaVm5SFlGzctqtlzeldSyS42nIShGImE3Soz6XqZqQd
YT2i0jW/wYJ81i9P9NWmrmOzWxKG4MOk9UdGAyiC6/51FU2DmbNUObJOIIrq9DtU
TnyuY4iJwfREPC8EQHSvooEHerLkMTHW+jcofbJU9Y359IZfp2Cq763oWPLG48yI
7A1s+M4abmWos4pwYMq1ZVkM+4sJgU3BBZ0SG8pdZIXmrtIV3TNRxp1VzFpnkm6f
M+v3lVZSaZuDVO1s6NT821VlGKO1lJNkjFxq1kizmeN954f2R8QdDQwQu5bRg/tN
qKCpTR/QAlG9orqCJIiuRF0ENFHqql5wEhWW57Qz/QyIMeDFLdaZ3ABVq+LLNY9G
wmLNsuEo8ATCnQY9xf9yjsrOFampGjQHt96PmcuBBmBxqOu9OyTwSDjPKfwVu6Nt
cA4jnzC6OFRCwHOzRCTEcTjT4u2wNxFzBSj5t32eGGi+sXEFPJuAZGrs5XNHHJII
2rf0+1JJdtzHmUPxMZoZUq32ST2Yd00/YCZ8aHO0mwEyfPiMZ6n+uyiLg22fQRBf
Yx0R9RzY6E5yj5snwQVyGtz/amtfiq9EfjVd8wR+oHg2+ChTjhoVQ43rRHX6SNdx
S8WQq5uLu5wOjQT6fTbHAJ5F4Uf8bNaxumpy18aP5IDg6Bud1tZBpaFVVvJ6FUmx
a6M5JdWDU2NDcz7OfhjVM/b+mLIWpk3+y802iYseB5Wg+5/gWO/FXHwpjPdzMmVH
rhYUZJLYuljKgJfx9GyHOycvlgF3JFhg19w+TOJYc96EYhc2UaI3elxDstOEAzyf
znnTlxe3T3nK0uAwfA37oDhIzo9LKiug8CBAUp7wnXtfziYKWpQeWkN3sWPJfnkb
DM3DcTiSqzuwHe7bPUX+q47iCYGyz2xP3GXyONixzmyKgRkF8bONW0BUhYCrp3iR
wCZ47f3DiY19FNwavbfXjHBxHgbXiIPzso9stS6vet4AyHW8UWARDZ8gZRVoE9/X
GlDBc6laq2Rk+a/Mqn8FF3CNe3uLvceqpSwAC1vmvbCROSayLLvEaYDn+yWjKEpC
Z0VqbKIMAjZmuOcAyPcPTeLGPxc9Q1ALFkScprcHi392IquYPlaLbA71vQdRbhq7
PmLEh8Paa4LkUHHgEHmvGkN/8EE38H8jpdlX9K33gpIsgrIgM6Ys2i8YakLuD+gj
qNuVKdUuF1o3DWdH9URC/vKFIM/cLQCo8q8YbetPFRjtaI0E9F+0vNqt9XTfyW1w
l8tGIvtmmK52NEUBGlCKPsn4/WO+Zn0qmQh7nxPv0tDI1rftumh6dH+nlcj9vCNb
DIiGShOJJ9BVMbYGyim7aR0GciOxEmED53z+6Udiio1eK8f6bLskuEkQ9W9Qa4ZV
JyLlaH66UagUbQop+CTNJb0uDIDzrkKAg+6PmL7n2TtRZScn47wrWKv/0u+gxuBE
rfNWGhmhN+pYyWYV1NvXuFQNI+1SVnPKLdBeJvEfc6dmGE1kl/VFHb17vD7tu6+g
HKvxf6AThVZjErW6aoIgJVA/+ghADA1tLDCS0HcMML044lTsH08ReVt50pNx89ha
0XGQkFTaJkBYce3iwAiUayUQK2CFXIIm73sWC5aFXkThU1QiHGXCxVNlTs4ouMUP
leviiJk+W8ZTA5q0/gWlorDyQeWF8cZximZWV6WfQqrTUgk90thrOz2snTJFZ2Vw
jc/dwbU21TTnrr+BckvYOrYDCGUeH1q9PQpdC6bio63XTjtpguqb1i41LWxDEdKN
hoz5GookiXwV0JJjhnOYLHa9dRzeo8SFoM0LaShY0ekrtOWkpFb210mLaX1r2K9/
8KUpTHvtgj3MEc623UJQZ+80yOBNlLdJ6965sZHKcIWEYprBKfvl/DtXn9vWYQb4
aEgpVOnlUQp+ovwJ/mfsMFa+C1a72wcCoajpD6UlrG1VBhq3jrISi8x4vKynwY9+
RBPr0+05R67meFzCY0QAyq0qm1UEfvT9rDm24yyZGudOw5PaG+OKpSyGM8GytAgg
dhzoboCV8sCp6pMau/f11s51cTMdUnXxPOz9pH1RpJl2CixvYdI8GAIvNs2giXiH
p1b7W18V0hdhjLJitpMXvoLGP/k5m81J9/1eUpdyPASJli6I/Hx9OHn3ab84fcqf
kg1U4QboMKUDvyON+4Io8qOZcItHIgfo3nn4EL2tlsk/6lwgZml3sC9JDr4ndw6u
pR5IpoMgyOnH9FtN/Kzodnj5cIPUqZB4EbHbGBWRB0Ak0raoywEsQvikXg247MXq
f2wF7NwxjlzwEUkXhyd8VzcFVrwAjI7L6v0MPJgnXqe6xsuPfnsxAR5a8xeg/Kim
QFklICGddZf4phmY0Jga0GUGRt2+Ap5TXC29cWSG45STPP7oMGTniHhuy0mAh/Pq
HnmQPbrK6ob9QhmJT5wpCK80IRNsF8PK0EFw0Tbm64Z6i3OaU7IB3QiQSx65Ftp2
IFTJubT5Wb4mV1Sc61y7xl9gaNNtLEFRHqaBF2bY08pWsrSrK4ebLtXApsMNgn0M
Ph8QaVV1l/6ugSgiL0XjHZ4cJzvUUdb17ouGJey2TLOuIHBUiKEhacxHYl7mnB+M
Mnk3gEz8VpzxOAOKF9RitMu0oigtIdfuB6bMexikDIRnvm68Xdl4pBwGDrerd30I
tueSFZ41jDLhbY3T8KTxlMU6klfNrTs/irR8PG97amjmddojMIIMDFKO3Vu/k+dX
Xst2K0MvuL7Kfls82RaOmj9gtxNUjoonMiCx24O/CjOIiheuXchMl/L7aE/cA7NK
Nz4cqHCA89gs5HXq0oC4M6pEadV4PhJ57Y7kf9ZPhjF+uCaG+KYV3cnG/N048sIy
pYTSyheIUGO56rJNyYQgGaZj9aahawFXeeUCJZflf6YLDLWPJs4CHDxWfWlrKPyg
T68u6kNwsKBCNmUBqWWcByJSULyOhd5zsaFXh2tmi29ILJrmvfpaKEVpOQY+SC/H
Xtc77HZwuwDhi0I76H3QpAZ/JV/ef0x3uasNbztC+4LhXNJi6Q86vclYyve4Q7R0
/q90UaYkCxwZ5E6a4bHzCFWqNUuqyPnRVxtvpt3VuAQx/gqL+EYVp6medrTAFocB
5KHko7sOcsdRo8VKIdH86k5srM+ZRX0qujDZ+uW/qVHhTzHeXJk7ya/cYM1iqtAM
G3acO4ObmxpsdWnPjo0R92stWQ8/iSx1GVou3UberqE08y1NHF27qfIl/x+Hnn1i
s5WiAh+BPXWqcu69bBgnx+GSFe082YmTLG3tl5PA4c9xAJJA6iNOS22nL0m4rPcT
a4C5tvXeTgToXxhsyxpWag7Ut/7ZH0oDKVGewriE+IsWteITmTTwPCxHLV3f7fsv
TeK2/r5Qd2hxYcZE8tGKTFKyu51oRrazRDfzj8fpHR7/RhSe2BG+gP/bHX/bwlwe
jOiCcQ0or9LnCuaDYIOCvfxd/AlqCf/8zytgkq0a1l0zXx/5zwO9X8OXra2z/9Gr
O8RPHdJgfyEOyfV8Vbbh4GJ4S/4H/lWweXiCv0ypM5obv/Z8RFa7dzf6WY+kj9EH
TKSLLBHkrkqJgtXpVZ+O1Qz+bVHvRE2mKTIxmTPL6JmRa0T2XsvqqlailAhdQRzz
/cJ4j8ApCbkFYGRzHbpygdkShfX7XgiGiN5fpcXKwWO7QeDRPyVoaV1LR2gPiuek
clLSPb+HewxRE2hQv+RXkold9hvOfT7lEInY7cGTOz7HBx6qKthuIAztLllD+ahs
J0XlwQMOZ+m7H+raXUiCdn4bpio4RjyLx7dhdbw7B1DP4/KMqcWLiVGjZ+uulMZD
GkJrFcJk3951rn4dpgrRiJroHnsqY4KEhjOtoSxynOOfrQnqoNbnE/83/qs0TbGP
A2LsgxUxXC2b3CcznRd42BDXOkP3YgR0dEeDUsJluZDWoi5DKsBgYBRFdn0cK6hA
+V52w+QdX64TW664Xdw4GNhnZo0n8NNlX9Dfa+THnRaOb2SFHWPkmz4ROtTOsZeK
aVVcDw/x+6i9NQ0gjHwB6mUhRSU8Uw5kkaM22FKDCgMBVH8Oo26mjM8rQovX6o5n
Z+xsutwppRzB7USb+a8QwGoq1Wg9U/0DnnnjVSS3JZKCHs0zOMFk2PfBihjsyyyU
65c+sNK56JmzhPt513sQ2vN7omB9libBOqJ85pO7KoLGH2TE2IaHzdClkEokJ6Lx
wVC3wTNmogDbeyhACPHK31BnlErj6y0B1EcM+71RBX+6mlqttqJQV2LkOFmX8dXk
a5vOKGr1hw6IjDn0LMwi5oM++cxHvpyv/rfP81WGi0sRUv+1JUeXbmffFF7PumPE
koZNjH8wKE5co5B8VA4zcWcpcSD+XOWrXzbhM1XniMGzLjihZX9FkvQvLt02V1w1
EhuWCSwOaXp0HhCBy0p8RDbqw3JLMGTwHo0yLUTSVr9l9CSfkyRbdY44jhSpXcoz
ouV0MN49/mRPq0oMzTDx5n7R7BY73heyP0thtNqgJb7EMi2qEzPyPX8rT1EgrqYf
8RlyBqcVF/oDqJ2bfypdVMMcCMJBgF++dLx22qf0nHgUSYsZ1hYQQd6vGS/GTrDy
rly5B0j6xzCmnFTk6X+DAEl0Sh/VU6YVU0S+JokwIQbVCbMgysRe84WPXylfHL8U
SutEbcgHTgGHNp9VISUBiEMwF9MDSpymkHZOtcKEgNfR7GUesCEyjo4h0bLLHrI7
AN5rrpYmWP2szgIfnbmpQmZYiPC1gMcncdNQtrpt1t99ihR3aZ2SchjMxIfCzLUx
6dm5MfjndeiLuD26TYQxpIZqZTZUQj/VLC+0KKSz5kiFYpP/6mF1mQVPyjMNdq5G
fvpMtGXUBjQytaHqXA2JUvET+XlLMTmgtcWOxJxV2IjZ+5V7e4uUa0Z9hUCtyE2t
j/gVyRdNz6FDdD+mC3q1NJnGeFbhkX0154UUvpRX0R9H5QA4GVkQSOwh1HwHEVPo
uuMkwRi9Kq7mZhAkM8bnjQnfoeG4/Ov9twYyoj9r/xyS2TBeWxYMVICT26cqp6wz
4Dofm27qwQ7C02SUppFZ/NqPzi6p7QrNtYvwPzL6+8z8x/7NB3Q3gR/4hEs4EB7y
mJcdJ+CfaGc15BlPXMZ/kINfGeuEgDqT6vikBchdxoEVUw4UU5hKVUbo/EfgMryQ
Z+RNIkmOKBPojECEpHEJywvnoBZWjrcQLvhz7pPempOSxmaYLlczRQkxQpdPf2RJ
tMkKFzI1RAmrJ5xdD0PaIllpf5oXWLiS1Re8DJuUhwFRC/cULmS9SC9CS2IeLYqy
KqO03B0odOUClONH90KwUHm9QjtjXM5ATmzzFSiaz1go9qLPXEUzvls+gpqRnJbh
L4o2XxS3Yd2c3s5X+S1eQZR7V2XTNffxJQHEae/w41ndUBhjwMybVCS/ofMq6Tdh
HuCyMUhPGj22bMxChuq49tgUDjtRo870IZqByKg2BDrqJnLVGTNQmbbXPU64gJ4d
dQuMbw7kqM/Nwv6LoVxR7RHRfksVnNxsiJJHcStSYaTvpJDR/hUJPQ7GjbZAMggl
d0fbzZ8GqUoLw4T6RA2mGwpatH4bpsLK6gvdgJkpsScqU3uTPIqVAVLiXIzG9/K5
qtkHYtq4WJ9DUhKZFE8Zmpxi87PC7yYb8uMRf+vFIum09q6eGRauIQ15LpxQRI/U
Q4/s65BngaZCVIfMRKIGjvW+Hv/zdVdWZjz+exzbXRPHqdtbjImqwx1UJtpFwA/4
C0xw6FBm/Lhv0v0KHSEL6Ghcn8qf62wmGpR7Yg8BWkh9jTisKRyF3r5fCRcm8ZaP
bFIHsnyslrwghxnvazSti5dtpLVr3SrblFxBvvcVtawN3rO0hoA0NyVHO2nLj/Ae
LUyLz0lwEYuO85hWKuVkFt5tJgzvLYZnDsmxxACc8FZ4S+IBnQQZ52Oi8OyUIaF5
hl6NvKA9HnQXEIMQU3tG2UDNv3yhE2Y0mRsUQGWqZBdg31T15I1hhAV8hlxcGKmZ
0M/KUXVYDl+ebFLykanWZHqWBLA0Rt3C7k8fRFFoaPESeCfQFA6BZlf4a25Meno3
pzdNuzsb8E6OWNREz2/CuS1vCEmVyHLLiBXlGLdugc7Nyzvl+Kb5y/dmOtWujnI/
KPJ6vKCh/7lH95k9sNvjA9STQO7Erf3kWJO9RNc8VIA6I+CzncOSUKxImd6iV/1B
JDxCFhvtpzQXFEPvSNbF1ulUJFpHEAQ58s8aKypZWBEg+Tpcbs+Te54Z03KsnaV0
utizyX2B8bc/pIw2t9IKAOItB9UOXvN8p9RQDkU4h7eX1kZuGlIXOSYaAJwrYwYW
JBXSEdya+G3RBUp7rBEyTsJJSIr+3BttLO+N4VjyoKomeGC65a/3j7bu7gM44xT/
NQH6Yzov9pau0v1wL5kW4PqkELEzUNHytSseReVLBvUliaV45GxXBlUajZoWe3to
lemZAlHhJ9IbBOLj6Zcoz8pVfOvlCUKBZfICKxKMsvDZTg7VhySPes/pQI3cO5d1
xH7kd1uScGD/LLdTD0ZUWmdcbqbaHmmEJEFtP8cpxajG2ddYR3hXXkYeJIWxQYIV
q+BkSYUdXak5a2Fyo7illAhE7Ob9obYNMBjxFiR4FDadwRsA/zeg4WPOy1iQ2QRs
74qImeC6YNPN3/FZodWqPWDdfYJTk11h4YLvN/Wm4EIEXVx4NRtzkZF8Uums/6yK
6q8dp/+AUi0olupMnX/IcDqEHJv5Iu1oh+uLTMY+MNSyDQkl3vstvP+8t/HvnN8Y
5vPRVGAJzQLlpywntgVMArhlvo9UziOU8/4vEG3zSOyWq/ZTQtMnhN1jwoTu6pmS
TQQudkWyc0BNU8ObsS8PwmmR+lbNpxBLfjrAPY2qX7KP2IckB/9awouniBsI15fo
IPgM4U47bnfJaBvAGKRQd+t/j504O64h5+gL/og8W+PEJheqM48BerNmZNpyk+kc
0T/hIcFvv3jcoGpmUoyviC4knUS80O8Crp71+wE+58GNbW0Ms6T/+QysXlxoCiYP
+REmQqjJjEHc4t5eVoWdLK8ZeyaMcd9f/Nr7vKs25ybE0L0jFlRwyKLY/UxYkezV
dsYh9l0/jPTiM2VTlZ17jcQu9lYAVajoTioGL7KC267kkw/g4P1NMEqPCeS5JO7w
2UefLQ75dRWbg8GL6hVoKUWC9gNhe0T5ywJNrrzgpDIIzN0WoTOaANMOTZgqDUuu
kIe5BHyODxeoXTOlG3UnoNKJNzp9dB2mC6euM6UpG6WfMvYk/tOWmr4D2w6xTB7v
Gdt8f1Vi4QGI7QjsTuZ4aDKoVytyywKi7aWB3At7PFyeWBNJZEU45CE6i+VyQ5uA
RcSUVzDUD3W1ZXud6JOprRCd//2K+pl49nhMxerIqm1W3QRkTANu+AxpR6EBds82
F/UN3sthdkZcZP3lE10LCBpCsYkhpBRIo17Eu9Dsry1KPRdtbMLdbsMiiUDblNU4
/mVgCmsYkB9nYC1o3dW+2+gqqWlXQHXZWku0Com+A3zgJ2m03JbOwKidZAPn9yVn
tiyPB2UYMSI9iN3ckXp++tj2Bh9Z9rlKPiLW/xpmxWzCy0TB22/C7Y+ZuyNumwMq
Sfyb3Vos4RQ3NeYfgQ9itS60DZrhDS3mK2hmiaB8lNlNz0kBTdLYdz3TZ35iRvXW
CAUvvmkWsHcNwdc80wNPQOL6gKhsC1DWv46Ts6iOyPSOv4UbrX93kJ+v9B6LcNlc
ANrPB4YQ2fDzH+XrOfxcrjFuvdEEoCqbOpvtqJikgWB6BA2jsK/aeZKhCkjAXosF
BzBzR97JDQWDmlu3bx196n+AgkYcasZ5UXcmSxzdQbtMwW/6j4bNYS5DZogOOyb7
NBeUEQp/GemhkjIIbZNEx4Teqsjk90lz8YZAVqQvSTbeGcP6Pjfx7lugP6A/aHEq
4QuzVNv4uhfB3LbDODxOXZnMD4I7+9r8XmWFGauzQSusANmsWf2wfrJH1GDNA04Q
rj0/KvaQKqh1CZQyynWGoZJ6seAiMW8UIC7JUtGHUeLpegAjPUplWEAbjp9DIcbv
J6ciZ2mGY307sTHsjkc/Zak0TqKyjPAa7NgwXL60XMjf6N//J5PNnc0d7uVRCtZz
WtwXQw+/6/l6E6Pd2hwH0IfXydoXKVUsV24C9kdLZOYcqfBo7Oly3TGxvd+US1CK
rrh08FpuZT/JFQjFWYmloQBEFyW7Z2y8LxY8IHSmvjA8WNh8mJB6ZJ8DZhzAV+6Q
+Av9Fp6pgPIZJou1b8jGwEkdifVgEoiEwaMmwN0hdRfjb5lUZqGzAWwJIHOLk0mS
Wsdj3yRH/fPeg5Yfvh0z1ZRRNgP/R3krGNeYNUWI6QhZpCd2t4Bx6bVdWzVAcZev
mhpcvJb+X85gH5eZKdzySAHZOibrtx11CinoeA1JDu0GMRgu35X/CnlRfS1tevdN
frdbv177LDqNnpboYuOlsKaV+Q3jyUxNo7Ly1tAANkL5KBbZo/jxd92b8VqI6bP7
HjDxRB7Ms9P9WZRTlAjVXSECFM8ogs1u+O+8oYURFbyfpg2rJr02wCqDH52Zbdld
9Og8/dQF8aHnAQ0w2Wi2T48P3J/B0fFFoo+IVYd4nZDDo7fR6gIDfp9rG14/7OI8
AEm14l7mi9UrILjkHgcM+qckL0c4Q4NWtXWQzzBafvSDZlgqhnGbTyraSONTaXnH
rpsUwNM2dNzuYjsNVrsE0w5znRINZxH+XX0G0k6H9pOVJVPpYrDwhmrucLUMvYb/
Xxgt9csLGhjjMnlOmzmVWFsPlwD2c0UqSIS68MT7bp8pingoXep5Em2XZObvvC3H
oxicsOf8XzcioHxdfX59Mj1TPOz38LCZ9+02W6nnsbcrPw//o206N4PNl/diBV3d
Sy8tDxp3BP86KwY2fM+xLruMJ1S+J2+0mdCwPhKjPbL6BRZHDqGBBpupp517VfaC
NcSC2dtji7kA4hatCxy7eNK0LIYoxa8vUuXyaLTzuD8TnO37WudaBr3fpylma9Ks
BJiNd4RWc2E+TzsxfdYa4GAdg20Sn62C+BP8bruKKVSP5BiDduBG5YcFcCUB0WZv
sKe6yq84XnFA/BZFnvzdsuP4AJJjW4xSn4Mx6YdMqulz0DdxCNJW35gPkNyGMq0a
e6/1fOC0sOpOjFWMSTO7g3Pige2YdrtRIj2QQTQmHMAdp2QuigMn6UJ+pQpjyCSy
lgUdq/3gfRWGRYbqvrmjQ3Am9oJ4S7n4p5N1U06HVczrWgx26piSltk/FMeuXVhz
2UL5b4PqVd4pGicWzQxLg11AjeAskuPa9frkJhWpZEKNRePAnZGU3L9U+jaWPBT0
QIbbLPvBpTNH+8LWuFKyOeXoCq+goWMjmKnSvmNpgk3oA32WQiL5PqM2chsvrccN
IlH6ZxKEjRc4WrR0WwSCXszcpLNv8aMNjmG1aivzsiVBiJ6v60NbYgi5FhvnIXLh
UtHy9JhLdXwTD7RkJyKd/8cOx0Qz1i4fmVIgEsI0yUSUxw3oDIHKecxp9LWULitW
CM+DtMKpzQGO39OSniEuo7Ub52a5+VWuSYdVz1Sf4d1cR4uQlA/eenmf6d++poFg
wH8q07ITcsVxxT428opiPL6GFwdSra939B0Cdv3IyL34vjq3KPSxMVYOt4TMkKmg
j9McqdCPGiEKIZ6kz2dY32zeivvyt0QfIphELolgz1RpTiCjslDer0pTufKSo1HI
ufSXfc3H3JR6o2a4c6f6+tA+X4TaPn1QiJ16+wGS6DoSggfOGcaL0zA7ilK5v885
vFyBS/eQoJnBYfDpyXTmiv/yO19nab16sj/X9cpLLYDeF0EYFyTdaC5ertCabehA
LpuP/j7c9FsTEn8vtZPpy6huJpPIov0kZB0xa5EZFf4A3yHtmtjMW6d4Zr9/YgFe
lgncqdxs8Nt5U6M1NvNpLPmpWl+dRF/lf8XN7U+w2mAq4CmMFekU4Wdz4COvJ3jv
dc1qlGwy4LMkUjstA09iaRPz4uvxS9H+UE8DblYq2OBAfiWEahu07oN8vUO3lw+d
znuXzBFiHbZwFwIKmudUKzLW8c9rrLlpEh8fKLSqhSiSOKMlUNU0AwEbMwhhQXVb
vAHJNC5g3cg7AXTwuwSdoJPtgtqohExd2s+VJ3TTL7RO33GoP15vRG98qGlqSXff
djpMOdU/ZNakbXDZWG99AWsK+ZWCPZ0fZ6Cbl+2T7R8eUxl+WIKcrsmRuWhZNvZc
gBeM1z32U2/78EQw5BJPQgZbQstnZjm46Q2AzzLR4ycGWK45DwsPdH1OV8yiJgJZ
Xhvvq6SI04k0vGsZQExfx9jVP128MvdZBc8wZ3pP616Q/xylXfGVTrBy59K3pTrL
rI0kJT/IqLWBy94RSREBcviR5oKovpc8K1gEgKOroGMWHCJZ8sYWp7z4yxmQDVDD
m5+pgEhDE1TWmV/VppUhtck6/ZSWwg1gNnqU3qw0ldIiCYB3dhK9JKYRFNpf7IX/
ZjjRBg3WGUs3cEYTAgw4Q38o77V4kEhlYNr3vn2PlpHxwIwE27YS0Js1kWvlLCON
bcuM49TpSR8mFG4Xl0J9eFwyXqztQBHRZiUnxm5l5QXFFP6pDn7946EGXy7aEo+M
dyOf4uwDIpvnH59MmQY1+ELE2Fpn41RJJ1xU3uih6S4I58x5pX9Fh22qrcaLk786
bCbQz+LSRu3wgwc/EPZ84rs/tc42h0IWuO6FI+ydgxXL1PLtKe7qjLNaPM4G0AB8
df+lQav23fCJGyuefmbAFpBQcNXytzn32ckJr6mHY8nqZfcENfudd0LQqtTVCNtp
3df9AbVhQnx+PdmLYcgHAqAhwK6LO7NO62joxR3VsSYvxdWC3YfrA3WBlMXBQYrw
WywwpO+Nh0ML3Gpy1HpkXxY6EOJEXtwRGss+4HxEigIwxa+GIRVg8l3jBMyqou+N
mRaODzNCTbkJyDTSRDMl5lMlc9fhfPGqhBBFg5HmLcm2v7ECNOlqI0y8yMkONsMJ
ketkkcZJn6/nDjq4E26ilF6YiPJ+w4+7fB+pneTyYc9TwmPBOdCwfel+cAzTdMjX
QDShaS+wNuOW7lY2o8iEb2eHRzyxN5xAZ8fSzALLYSUh2oJlWW0EgYiB6snauSKK
vTFdUKlCHGI97YUEn+qAyr4jXonG5wY7XbUX5TwLxOGxNjElLqrjOS927JPzzaAq
MUydRb/f/+FFpNiqxQ730DdGTjat41yegt9cdBktys0FzSJqRTPdIV2Blh6LISCj
9Bby7/yCfRRerdwY3a6VtrFM9Ncc4UKJFynnRrM5zhe3e0uX0rTkSC9zfhJTNumB
JsMYBCCXZBm0cseEvvtHEg21NAdaj7y05+KLyIzfpjCiVkd2i2erB/XMCAlupiKK
Y/oIzlIGb6B6u5G9rOqVTFzgrjGyhCCxabnupUpedPrZyfEni6ZGjsWpGVeWnacT
DJWhhHDuqMywzwO67Pp0H61ETcWc2pcFXFqFJRfB/pFvDaKm6ueI8C7yhJANFEUo
1mXvxMJQ7FGfuNZrz3v8mghyqrFnIxmF5ZlxF8dDitjNpaPoWaOoMeR08i7/CIKB
kMVfi6OboZBPgJmLKcvXSjATL6B3lCtSysPdGd+nf+lhAZLc4ZB+r5erbYLTk99X
FOmDnyNlYkEYsA52/u29RCZsgVxbpCJYcJi3RBRHdKa5Istgtjdyv03K3Fk/Z76a
H/+xCXfp6yxFb/Z8LraVZ0xI9x1ou3GmzAcXAT8jmH8wB6zPgVBcKGMZ4soAVJis
PjpdorrG33U+2/HGodjc8g+t7ysowefOBp+xnP+QLElEVyt9R91qVimV8LiAorAa
qbdGMgBW0tt9pwwlFHm6U+Jy4FkqvqKQMl0RuyX7OoJhVRu3kXRfuC6YMr31/q5G
svFABHKZOesYuLVFaFtDWKTR9mTGgGcnuzIO2q3QCymOunOaVNlTzk5IqzQN06Ly
oQwoxtQw35l0qs7z2UkkRslLI3q+y19iuaXNL6bD6I3xyrvl9fiSuSueoMSgqLvI
BYxeH31NnjKd8Xb+DU/dk97Gr1VU+x0USsp5bSIyPBn9fZ66PMvfjAa/NnKFmfcj
NbGXrYWudUt0b1Xg3qKgcUjw64A7giLFJ7DMNzN+mZucpKL85FZzXQXma3fInNQ5
nCgl4QfItZXvn4mEF5BpUGCBUl3VhFya6Oc97EYHKFzHoSqom3H6CprgTw3LXso5
RvfT2saXEui1xbrBXlh5802HGsYsln8tPBW/1hK53WoFlgNLQTsd5z9A75UnqCKM
FABAg0JhKLXBNAXKoipUw/Ea8EcnSlSZheLwdcpDEgSaPGC0psHI2IedJlhFw8Hg
PwgDj0ybRGb+P0jbJ2am2Tm9EO/59kVJYAMOFGml7l57R9pt13fppgH6h09o0G5V
VNjPCtpxVRoGdfnZ4M88pGLLpLpXDXpifaRgaspywO1/fRvIdpc91qJqD1e6qOM9
AErsKXloJa50wVlYh64TeW/KBGQWmpuBA56SnXsoxytXTUNWgR6QPF5G66L/4Dkj
Kv6qXbNsOKCEwOIjEmVmqu261WjEBVNMwp6cY7iDsfQ1PF2ixZatH3umrXSbehUx
3jJDUyJ+A6y/5SViG7omDq6sG+ZVRdw3vvXPjT4EYs6U1ughVUy+o0nXbYzFJ2Pq
Etxhl+R1bz9fnIHBfboeavBIgyPF3+MLOJKzNkfPxhXDcw3akehy8Jp9MotYHNGd
iWLaRXADDHwi+jqS0YRc9t46cd0FPZu7Mpx97Dl9befBp8BMRhQtyO5V5nX6RPRs
QsJdvqsB3pIz7c5Virbz4e9bEG0cDeFTOy3Ew6dscDlLJBAMC98d0F8czcyJhsQ0
vinzgHrifGPipc9WtnB68E3HaF15OkCCkZO9/BfOiuWD5Z3YTjZL+2D/3ZhEpIn+
cbeIttJ7wdqkfgqqk7BGYXa8uIv4VTwigGrXDu/MDRUQI1ZMH8IKwaMRQdgbsXPi
rU40NX3J8lvTqamAcM/OnVPVfw5syR7rPae8gDXKq28RqCXByCn21z7YLemBkar0
OUN9tLVUkcq46dwd+YM4dStgsxdsc69sEqH/p+k34YVrpoUUhP8mRMKv+pzOfs7m
AlTfoFpeHrj9G0H2adrom1jX8Kw2T5H0lDugABcbkWuHuGOSDT/EJ8yTiuo6BJdj
Wz1dwcn4JesY36QRkM/IK9m7QupIeB99xGvGziCUfWUmB/DENaxJsry6Npttjo4b
0tBiXexXfWO2+J1eQXm8ARqRgbNlOPpz8XEvYz/Dh3pq8wL2HBqu3QxU5nBoAsqM
9jydIiwLF6wva6uIsYu5zRNDLCPXOcWkSHkwrhwL442LqNI7KnwuTdtxn9g37q+8
JK3sf46F5YAaHFesZqCsPnxN5Xl5yGfb2sn0osdrEXKZMgYU/qlncyt5wvfrI9Vo
GjJ3IvsGHU/uNSZwKIyuJJkqfO3LQWb7vRBN5rhs6lCIqbaPzSdkdb0EdUBOiTJR
kZUYtmsUbmHCWRHLikmMUTzL8iyNurbJOGfWetyoyj76YUQAgmRzT5fnlMr6nlt7
N7yT+JXW+UGatw0CKkQ8oZoLbYTIVloveqrbKi9pZTw97IeKwPu/Ol62TeC5qgBH
Gj0E2CZXFyvxn4201sfC98KHG9p8QZSE4KTl5YD0fIw1auic5v1jflYabCqtE/0f
ZrwGZuIiRCQ0s+RtDF6C5VxoZFth9b0XyZns3QA2LD+0RSS+NR/2PnfQ2jtrf7t6
pmzL+m/Xx1Yfq+J0U1h7KPl9ngx1Ym+ZTGlgTbIlcpSGD1kLR9b1rmixNEGshTKH
UjgM2DxiIUrlGxbU60AtZaX0LLkoYSEF/cgalgKMq+p3YcHPG2Q1nSmo+v5+y0Gp
RwjAlIhM4A+qeXn4lbwOvHyr4OXqi98EWtedIHvbc0WU2OzLgCmqiUKt3ygaD4eY
EyLQrzAwMKD9iJ02lK0GQVhjzIIsUXsPzpZYIlLKwxHgtk24/97ulFzQu5FH7n3s
D897BksviHllOTi2ReCwpcyfID+A6xzsH8rZWwm8ciEsCRS4hbmwtDPsuNDS7WSQ
38OOJKo8Iyt3zmDvZhFn49I1BVyURHC6qZ/2sc8C8M1X6XxfYtjn8g5yXPOuuLTZ
7INf2xG031Qc7fGjJY/okNxIqJXWoklbeDvkCnOUssUpSE9TbQ5oJ+lWiPBRFKdd
03cSoF1ZRA+vBTubNPTxIYm+1nFnDoTQmQyBVDC08QyN8FV7g9aXQ3ERqEAE0ab2
ROMOYvxvxoe4wGkwOHA3j+VvEWddU97njAPxtIF9dCyEByeOj8UtSWIkijK7CVW1
CWO/fhLzmccLdoOasYg8SRQOGPG1oF8T08ebSW0C9X6O0v2miQ/ryI1kNDfqML6q
dcbbrKTVm35pfMq6lADFtGrB5lb7R1fWn+2Y+CKk2Kh8qbF3TEjrQ+SuQAwvHiMg
mTwRZYRQZCpsdeEMYeQ5eC+bRSZahgsGZxQjnx6jl0Jw2E8Sh3CGVNH98QYNToFu
nyTmhJbnFRBrXsn9OJTn+6Y2N/D38SGXN3j8/JELiFGj4ehKwyg4lpwWSHUBqsMg
RPwRfMNSrvp4yLsH1dm43e13kv9SMwFGxSWhMC14LIofYirpZmcJEIaCtu4s2Hzi
F8FNivewj18AOBp6bhv0oHxhvjNPWrW0ugc9UkrnYt56V/036mVk6HcJFtuyg9SW
Xav+3XVvbZ95lHJZUGIN/edJ2m7/rdARypTG1/NEWl16MNMQO26sVGNDKCtv2jKA
hL7yfGMYkwpRL/GS5ViA6vNoojUtqbVPy/1gq8KL1iJcNbY24pUYVHVmT4Li0Mcr
/yfvI3vSiDly/F20B0yX+OmbKmuEoeCEwBiywkdpf+1+63ysJRVOl4rqcynw3d6K
qFUtW1p98k8GaPU3gZ8HReKtOvp0B90/mA0huSh3jyhT/rZXi2pdWrtqmIGLlahl
gs+Vba0X9EY0+R3OYS04Z82AHqZe1gus3D5F+Le9nSzzXykGRq6MC6eEOofraDwU
EnBsjZtyQSPyNEhNJ0pJBapybpK/IC8O/ThL/x4urPVK/YJm+GoRJncBgzhkWlVF
Iu5IZKH4oomoYlXpDysQQaJqYJ2XW1w6Ii5SaIWG/7OrLDuPsvzqkaLaD0fABNAZ
hQMip2Hp6FTeZw2ZOHE5WsJI1F95gHZrdCinkLgq1VQuS7fAa8v1S1s3pOdTMxr6
Tt+IaUAOoBkoGWIOot9+Jgv9M+Qe8hJb3PgT4BfRNibwxnBZqbs8SAPdupns4Qis
QQBkeSZ07n4hiSC34gUzdgYun9QAUcARN9cBfAjTvvkZJn+cS0yNRfpcdJpOx3Iu
+YAovb+HT7TbDDIDwvZPKJ5B/hC2nfvdt3s/CmG8H/ZVr987Gec7tZCRvMQx8hwl
Qyvx6ecMwLjpfkul56TXBWoX+F3pkdxlSaoWKoesvJ4DNCh6NtYodjxdECvIw326
pfVuN3dYqLrnwYrP2wIxO1oOJMU1MBTOsPmEmpIFVXToifbW8yanwsfo3eXKR2Yt
b2ZGZUXptXr+0EnDZGBdCy1ikQabE1w7AbS1PULvIXJicHS2XxmcoK34/vW4UfMo
7ASM91UB2m/rdD0052j3yIyIT3FkdUkjbu1ZACj71lOWX6JvZTDOy8NHPVqSvyQt
mVV0vrqJy3PZzI00JG3j2mWMuhQxneiXqFlp/NerOOjCaRj0f7sb5mvJal7CnNPf
QZPymNLg5XOj7gdsPBw+s+Pnl8PKfT3AJPbzPVN3KeoG6IgXZYbKjwp4fUNZq1So
CnTXNhTyrlT0ea7giC3NGYYdukQr0+ZignQxeZWKoDwirVNjoAxxAs8mG0/RiTDT
76HQNxztg+c/GzRbaJyGoZ9GVsBfh3eyi9UzTCRzkMsQ+rWcHN6FMaSiK0sY+aD3
qhjLnkTt46humbhPYZ8CP2LHC3Er/fQHgmgK2aK4IsX0+bZxG80eMGCYsFk/txCW
jgxyf1thLd8ycSIiqJjZlpdLnLrxGpGCH8O5restlUaMbjNe8Oc0C57r3Y0tjjjf
pinvQAux7T9oRO2qlQi2O0/xm8x851zXpuCQ2meRwjtjKaKy3f+Da9AVCCrRTzXg
jUqgUkPLq1en5vz5YqHcG9ImCLXhG+gp0PQWshWURRF9mdKXnZOp6HmAe7hl/phb
KhmEFZj8bxDYXOFiatHqTD/aNGKhoypsgwPCi9ozgFwoF9yUIFYmA9pCRKwlL+UI
xlYihzb9qG04BExbHKn+Vl9txDWC25uzh1yrz76gXmPiTkZwwOI9PdPV3GzOWimn
erkeiXhcZFY424cv7FgBeJPsCKRBx7VUASaRDfPW94xisUCo9CBoaQOmm33kHVqV
tadYXFU419OriEgnMSuQeXNBfcMjcMReqvVm2BF61s8DW5ski7l5h24C56iwRWh+
XXXkb3i87C5is7qPMZ3AHh18ipZtItR5nKby51eoixo2tmhra8EDx+n5o+MiJHNU
IWszXfu156lBveoU4JRzARknfbYU13xKlvfQf49xa77DWQYKWgkxzCkWduxaNEBr
Sh2RsLlDKJOAmqgqZeaOpjkeQFULYJ+PbeZLXDwa+/v2377SMNKD/e67W9nXSkPd
OMTylcpGiFAUwrqdGHXW2KcaOh1YB+hrS8IwXZIl9Qc1HBgx6hCZzBk/cPej/AIa
SA8N5Bu2Ob9I4sa5sIqox3FLFi9rdXtvf+mN/GC25kfUrsPoE14Re0IQGhmbKBMS
DgZshUuxSlDKjS08jGKjYEfwHJ88alkkTNjUg7H2wcyu17MEVq6lfThPlIGilaKV
jyC/PFriE+1cIiW3OgE5T73+c8K9bLG2+f9YRjjnBMa9icyvH69UrtsUAuHJlHMv
WGHoO6UfgbFeBuZbC1xTUBybQ2u/S2YKH4O6mfnnR5pF/y54l+cbNIep/JnJRxF1
dPty6MBOJy2AKQR9Kc8j+CsePVRhbqOtJgVMNPK6GZ8BmRB0oVELjWTRoy6/85i4
0ipQrLprAYCEWVeAdoJFkFvV0Jpku25wsyVA9S/MVH+5eMGj7NSSoFE2PioeKWj4
gu44jCivj+n8180CmqZRH1b+7wc/Rrigp4l9eemw2BhcplTm90rMFLkaTbTOgbe7
o4VkZUDWgjfOB06+a4yLUD93VTts3F0smiE2mmh762NpQPVG9aQpydQ78M0nS3+2
vEKxMQcU27PxasqB19pTWXzm8mEYgnfqFWiIUxS4ZCflB3XZhz41ANl25PU5DWxG
1x6iP8w8cayDDATNUeR2JJQi59hF+t0TxF7W7pcHugbcxsOow86Oginw+UHdPGkn
m/WzKpLtJfZniUoO12611aiAedeoVOPD1QILL6WelrGR6D5lYgL6m9x/89ptOg2D
ZE9U8Xaxow9D6AAX/jqAgub6HTs7+IHVImjRD85LPwgEZDWlI4G38Jzt3F76Xy9+
6MMN+5mDUILODX7OLKsW+jU14Z5w6Wq/dODkUaiKFQwixHwuhFVUFcAmAP8s3+hq
bDOP5D7Ekt1olpomKs5Q43qSeA0UND3/K2A0UpYGFElOKCCl43X0lvD037ESLDjg
YW75olOjcaFWCOkY+ba4BU1Zh58k/uX7WHZcM/LYsnXopX+LbWCm1KrZnlqmCvyw
wIiEvoQYFsFLE8lklXq/1nS4piqmQfz0B6MFYGq77Za0UylLT54Sz0BdNSGpF4Ok
8+ZkAtgZvxUdVuu5a1EFy8ysykH1mDPKyFH+Gl/qv1/QpQHIFWRQwxomhkSZr59I
dJ1tZpBBTJrZFEGXHDooY+l7kfAtI4h4raHB7BdWvDsAb+edNnyxCg4cOqwPoV/0
rMT4NzdY8uHgUzOf5ANINTvssvqxm/HzM467lZ2G7kjQG6OXZG+Wb+J17PWPYEOV
taHEEHcmdOO5JH0SY/YlizrCuvjILQX9YdB1iARvOcunhmiAy16PExZ2F/ONFoiM
OTIi30mGqylT0o61TT/DdiXUZfnRW+WCPD+AgaaJG0ssq3gyVRM2HrsQbxpEaaB/
3CMLtfTHF40dxqhRzYxfzbPnNlxYqH+i8zZwPbAVYZk6mkDeQSK23Dk3ZXXfDtaA
vRb526y9fm8aqU8ZjliMZ1UIxFxPJKeNh7zcZwYe1J/zxbrlHukWV6FLL4jnr0GR
7V3Ulgpol8uflFJTX8T9/RyKsJFn+MPTzRgrvCbriFsBLvxoTZiRezTKPzKCiABb
vKSVqj+9CqSVyxsuYlxSXx20Gty0Nwm8Kz+DOoR+OGt/c2CKdwR3/oB5xx3P4lhy
4fRCJiccKLMo4kUopp7vQJBSt5IlJmdBEgF9eDIKGQ4KvakntgTeJVBz2ts3/5kY
Mv8NFjIJaaEsHHujXAUtYQ7cGd95kuuW1cF4fbmutqP6Bpnm6+IpaBJTdRlkNUwA
HdyZfGcUy9eBu2laLpLzurNXEgyX6xkRBhkMNaDqb9Rvu/dKq3WQr9aAdFh5L8em
n9qLH/mpwRIsxFQU0qgwu3Y9ITJeu3/BYEtmE1utvOc=
`protect END_PROTECTED
