`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0idY1XWGsbhVS2/FZbc0W3yhMqpx49StZkAFkL2uKZwjKYet8lAuRPO+T4+8aw88
edrFuHJFOPDcD4p6yD1i6BWCB0H+H4j4FqcPfnrh/uXkUvcBqMNiOrSilyQb9LgJ
fO7BVqT/nHywNFqVrIH62HurUS6cLqxNmQAmLQyKBNYc6YlpkvNQjM/GhcaqhzpB
FWirOWhgtx/RaX31QXTB9t8cLAMX0FREXWXsO2CpWXOHt1fiJUEvrtNMTJHPY57J
qP8+AjwDYVKigCJ+Q0dzvyVUhJNMkzKZOgx562HLgHycNX3Z2USy1nm0KphlzkjW
Wb9bnaopEhaYbMJBfaxqXYKmen3dcz+aQR5cLosx8m18OUvrVqjPWaemUrEAcUCD
uTfi47RgEZe2zHh546fmWuwsmFO0z3Tfe9FH86MyIgs=
`protect END_PROTECTED
