`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKrzPw/ZcQA+p/K7YxIWGEsU9lceIs5vBchscBGa20JJmCOJtVrt5Th2fu/bMt03
Bko7wj5PVTUbn+BPN49r0mih9sOaLd8e21YafjmfXhjsJFTf7iK3/ugmWtAFc/zJ
WtATGTSG9pAlTvJ+aitCHKu+tq+0qR76AKCRHkJBmQTvcfTRJt1crKvcp4cVgNFA
MTGd1tB7665Meungi9kPxv/SBGdoCqeZYoqTJpkxgA4aK1hV3cIkH9hguFXKAxUN
qUqXDEJm0GzW7yuzNhKQGCj9Na+DAKpGsQqaGYZGqnYHaQn3NdmhW3/EKpQxW0kk
tNq+LXgqxchE7OXaS0Ykt2arpKNPnx+nrv/tEy9F4ObYMRAXAJosx0Of4MR7SeIm
nDUXBaPxwAPPSk8KftCZ0w==
`protect END_PROTECTED
