`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T/6gAb9jqOr4eX7NtbgSkEzlIf46NeUQ5XChxOu0GvgRRHAlfkMN7MPe1lKRSKAO
8b8gTetj6csAOP3ZAEGFf0ClckrnRz8/uHdA4Wwj6tv7LbKGxm5wE6Lunv2rsAfa
Tr3E9k9Qs1prpJVawwAJkibe5JAj8r07w9pQNgBeA6SYgEN+I2dFb4pR+dzEVbxz
lyDtljthGpY5c/0DSh004/zI2B9AgmY9A8DXGrOQcSDv9Z0XKwZg3qgIbiU1JPc3
uIIoQO9yd9RFq+f4OOubN+xmnbEPt3SrUsIrj9HjBvorTXFXqsic9HNqCRN5YPZh
0vAO4jU1UgdymTZo9P+J7S7LpqmlEXakdsbCGourJhxbLDrUcaRX9hEzEcarfEje
li2u7NiAKEYckv5LZLTAvcW61EdfHClPt/1jEqE3hRKx2qgXtijt/PJZ6/MV1Nau
Sirg8UMuDXBxvsN7ISFeia5HOoR+VmZU2svK1cS5e2yOaS3yFNdP2xvPhYf3xD1z
rwnnZsgtmQOS9D6jh32g6XXs5phrxz9tvcLcxk8kuWRtDXFMz34Wo2xqo5Jqqhng
U3L5nGVXJUWOuVYvO07q93pXM2IEXMZcsNcCKVm0iNHlchVjUovHyU5BSuvEqU/0
oV+dCupeKJkgBtm4iH1ZNGlCCB6s/ggCcr+YnbpZFxgrMDv6pDi3kxYss+O/jThS
Aw8GYxSlcBS+Um+Mr43AUOtla9yrHRNiArWrS4u3mCTewa2DjPkqvMbCK6lm9hBW
ZuqZRWJw1sIPmzSBcKYmPMBNLq7XYkendV+mA/rU0ON7nVwY5Ht08CWrPmJkNb+x
9Ow+I4jPyaUnXDeTqfWwwDI8GheJykP1B89wbrX+gJHpwICjyImvgBjG17b+N/TE
1Ob2bRMDvFK4yYyzqPxgfiaAJ3BEIwLFMNYwz18FKS4amvZCJlZXcnWzGsYfKpuO
zCL1GxFGePNAzpHYcvbMpXWPXpzsL/IwVcgOmwSY+/Fb7r9joy1MvmPAXy4ZLgzk
qdoMpMYDy1xL7Fgllh7G8B9uBRPDcOlncej9SdMCg60YzpDU0BMlgElvjL3qbTsI
md2BCg0/+IOmmhns18SwXNpYyELJxcE3vtNTr29waDalkChXxn5rZf/hqhuR4dJs
X/dihoQNAsjft3VlEY75cAHeXhIktNkb0yI7oIg2huyFclSZuiQZAElq10oM7TET
mk90CmKDwo5ZmKQDKJhy6HzSNBZNcBshxBh1IJ3V7e6FHBsvCroYLnAhx4KqjHyb
tlV/i0d3AmicB0mwkHi2vJyT5CO0mgD2Nhfkbc7XWrKBXkG1oQ+fEGq6bc/rbBG3
bvF3xlbVqGKkXwcXnY+CW3D2MWWFLvZZk7W8bq3vBqlBO7Mp1MVcI2Oy1xhuqXz7
AH4yJZIr521QLhjd2deqPq58QA8jmVviTdIWdPxLIv9S7iQ7wRWS4LU0sOw/NNxb
iZ+RYpuprCgrsdD4qjr3se6CpprWdOvQ1TB5xLSs58A+wZLj6tniqYl8zxBPovzA
DHqH9S45zM1JAxsSLVRv1lqSdyEthQ5MP8pj6W4IB+kkhdV8K3dwPyoe/kAi5x9h
9JC+yz94EHubmxJPB8nNH7UaLyKFByBVnfPDif2vNOV5N16Kli88VAriOBGFLpKo
tcr3u8pOzvduDQaG/sROdoRWGz4G9QU5e8SDf6Pojr5fxi90MrCmEEUgnpcUeK2p
pYGQFZXJabaHbGQFuj1680LWFCje0KZkhx7cEoBnpxnZLNL+HCMqds3Q7ePwOZSt
+BZ1h6JmEKKFFW8lLWyuUZEHJ+8KwQhGYZyoin9NbZTeR0NsIeIrO2zA3jtrCjR7
J8JxRb1dVeEFpGI+wW3mvsyoplHHihFz48ZSKErWPkakbFDAmT2o5DlguPHaHMx1
1d1ltNlq/GAj5X6QlvFUMtjh35xE2f+SmfJ8OR+Gh1C2aNAvvOg3siL9k4SK6Kbt
Kjs9TuSOLjlEp1vClpvUeC2SRgbzIqrRm8kpzWqFmcOWlAWNBlOV3PIYgA7fHMxj
OcWdMBgqiElw57jHALuwJMdKsups5WzGFPAtI3SpcpynWAj7poYtYtPG48N8UaDT
jBcFL3XaeC3n9PJkRWUDT18hqI+7vpPb/uTfdm7qwmxQI2QLOt5bcgOOv/vgkd5K
Ror1nejrVENOM2vHVjFctLUy5lPIJT+ZNN+hKRPuFqda6ZyIMrevegSU84gQu0K5
gAb8Em+p91I54gSlOOVdh8s18oRf7c+ivPyOVhbN2x30Ez2b+blH5YURs/AkVFk0
YZN5aSbMKfKS9xvDB4TuQ0zU3vgWr0eewqzCJQyHo3JHJ1AgAP/kq8xhItjfOJk7
X3bUcTTBraZHrtitFk9+JPyixhpPSyA3fb/n4paV3fk4Dazcep7//kPW2KDssCin
y9HpOZwVt+kR3GCkyM97hgzfedy4qOupLR+8qzDejcSkeru6Qfld3wXSnSinv5NO
wezk3PSwDrhY5p/yo3/5OtabdQkiqDYjAnQhrCQ5FNceGLnvpQ9D0nVVhBU8qhlY
P5I3keBwkCdGwPRYb434yFBMxmNu9dKKRVwrBVwKEVJLd9t+0H/Zr4hcJEeL1v+y
AnrETRnfjp7Z9lDvYsOHVHLfgjq7Omg2YrCvWWq4lxGlZnK2o+jgIL/jLsvBmQly
uagFmOkgC7CJvmTnUiCt60KFEe0vZ1BOYsnhUWtDlhl+AhYQLr1LZWRGVqZtFMcY
8rBcDPXewyKI+u3efpTJ5YPq5Cbq/h04NT1f4hJwgmrR8f2F2V6EHtw2bHm9+Zr3
OF00CO0awrPvO4nQTUmdJUSFDc7ehLEWzOPUyqki3sNDG5DWwE0EvQKGZQQ44SSd
p7y4BvCLw4XV6omEfkVskAJiaNsyjkxGHYk+cqAANHf/LB5/CBSIzHpSNdp5KO/T
4yaAZgQ86PZQuVcEBrMruRl+V2kTBVcBe3Unt5eXg7AwdI/NYHlJ0JqkN/Vqhhp5
p2a3pAJl3kY759p1YdBa5iGwpMqYVlqhewPlmeDPgL2VbzRdQXxmP22IBBpOI/qU
dv3Hh4RnfXtqiaIvsa8PLw==
`protect END_PROTECTED
