`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGajYkETg5m47FRXYPUyfxfeAh3qtEvoBiaIjKe7XieOeNBpNuWlzSpfTGAzKCRE
nBKTz0Etdjdr8R6b2egO4lVWv8qO3F7qjGnIcWwBZ4ILpwSx/6tN3UuLwcnCebXl
3HfYM3HZIR9BuJvBIPUqqMDDC0NdME4SMd0uiI4hpy0/MFrCeC1WKsPkfcEIuKYo
ZtATg8/VsFFAR/j70Li8RCdKqnpFkkOmpG/BT7tijALM3nV+lr1urUe/S/4C5zo8
RXHH4cjnmDYuZIWDw73SyWY4+NzWY3rvmupluV+RpfqwhLHXad6C/lYNOghu0Vn6
bmvB6705sWiRL8/4n+xyPAuC6o0EPcQ+zaI8MnBPnb5KDZh20opsC4MMMLpPeYmk
OXBcUToewQG24/u6wUV7Ei9kgrbOc7EklySrEHHu99EV1i0hasYc33UXru76Ma3w
7a0xzItvPorcQcWpB6r8hdKkQ4i4JslEYgjJjUkWCOVmySOuvUL7Q59+7kBA6hg1
r/WDxqvuWXTcgwafaS/hPg3lz+v3loLhhj5iniNbaTwgmODzoB6OYCCPeqMeSH0m
r7AhZY2LN85lXwBdsV4Wr40J0O8jPVFIePmNhrI0q+VbmEOvDEF1M+e9avngYdQ/
1jxdOwU2P2VaD6KKcxjUmvtvTLD+N9dmAJfK4K7lNmBWqkMZaYzd+TRPfi8U+02m
KysMMEpOcvGkLjIRglTO1HEau5hCVxkZkmBGgPXATfUXWEm9U7NWqKU43w01xTpW
pyBTmuAVbSBMVhAxlLRV2AR+l21BPW1G9ed+NdragVwX25XwGXx4eUQ2bePEnBpF
4tKjNInNaD5YcKkNA3LHHdE9AdGMwq9d/V9BHDLY85rh6YTxxyI+SfWR+MoeIYtB
fqpCpODVWkQpq1Zvdtkt8Oq+VCj28KEmGHaNaYJljGByh3ytGdy42JD4JCa2x6+L
YNMNkAX7KvahOKXizOMHx1QypjTjzEg8rF9qmJ/39YI99f1CAoViyOCCd+8+X+qG
k+MogrRdNyztoCTU5i2HLWuRK44Bc2EtBMslM107iNJv+PEaZ3cj6wqDsdPCLPtR
QYdt7BovrPuyXNBdI3XLTSi2b9r/pHKzWXtPtp34yHsGURLIWb0tdGxRjmzI/CCN
rF+vrMCTr3Kiwd1txJEb0VDknYv6y2Baa1DP1pBNcOQOqVDFri6vnRvpP1qtJE4h
fT7G7H5DF8rZ7KvlDh8aa41oZ4H/NoNZVSf/2oy/7oLt+Fi2rUDKPu8vEPCvIrqO
8DK4c3bXRpsca+7mTL3P+c1MtnA+PB6KVZIZOEltF7g5LQxV1H2A3yx3+uyCdSJ9
+fH+MzXwb1jo2Zw+m7OOfR4xSInnh0ypR60qfve9iFSZrLWKhPXpncqzVN13+4Qu
tYICauANA5dWRcG8pDUS+d7nMrKZZQ+eQ+FVfGf3TafayWPrFvp9e+uVCNRG3O0g
q8ZZwFVBJErgw1V7eatX+1mLvYQujBk5TojeWV+szQOhVLWinIpoGUzDxUivYTY2
p3tSK6D+uuBRxIx7QwI3IcNbl4obiCDQw9vK1AI9WZJ6KZC6QuPwiPVInC5hCbmO
LSbA2egboIYiBSgBxCHsBLsE6Bv/RZcSrVt0aV8KTb5l/ITHB79PxOw9pvp4sjmR
52g+733xWiWkVwwDbUHsYpPW5UaTm+M/k33Vp94ZWH8AWE4U0drzWB/cWRnBrnrO
NuSWObmPYtFgwnWO6CDw8mJ+iSyRGIY4oBrNIzkszZZzv2IwnjIzuY45apQd6x9/
tSFIcCaUzq7HXkeXMrpAQ1kF+P2UjImSoX+1Pra3+PrAembeHakV2ETRLV8jXmmu
iVlV2X7VdSW5GSOe8tHIByIrlhXxJU/vEWB9nEnDtrTupxcN5of4KIHaHhK5LoPR
dJREO3n5YZdU8e9gTTAQsgP5J1F/42lW+5GA9+JewGP+CHAplIYBry1ktdrbOpw4
DF9ndhMnW4UYnO0rthHnrLZ7KYCJtr88r44FtqhA943FgFLFKI5xxHqUZVOxFNkF
OVjK/ILR1Ktnt9XVkRKeGQQliuEznq+0M/E2XB15pzaWM6tcx+ct80T7gbMkp/M0
RAqsNJry6QyptUtP7sCVqJOIxHGO0q2RNN7XLZT/np1OmFHcwtYJkAsN/Gca3+bf
e15XFOrHD4CPDQUV82zLPox3juyCA+9We3LkgKAIcWn2/QHCRuwhdBDX/YX8ljoc
31x00RODCx7uiQfvU8X9eCovWDoQxR4XoWnspxrbSXggaJr0XnQNSanaKjgR3eIK
0hDGUtCM8pUE8aPtUE2tdhjGKFQgAnqztdVI/WOL5jheLRrhuuUEJpEl7lqA6pJQ
eQVaQxkYzpSBoOl1vAsHCXQm0ytC8Dzh2M6DqXTXECX7abzPDzQdf5u9j7oRI4QJ
i4j/4A7sr0y7X6cvnylUK+NNdZtpVxA3aM75o0gU2bkXr7OzPpYmaj3wMF7BmgKP
a6YUUE11Tax/zHhMEEKkf5wqpLeBv1YFefEFNg5EeJVvVvGOAj13StykU6arkbt2
qYajkA/waGO7P5Uo4rO1sb3xLKfEBW21nS+r/7zncmnmq6TuMM5i3TJldfB2AtDB
aWmfmaaQWOXeV0CTwd+aGt095MoKugYWNIgQy8CmXSyFePzgNcI1B6XRLZn0BOV8
41wHufMYf+i7zinNxOOeYO3WsRvJzOTtw8VVsE36FSZJccyw4oP8DaB5DO1MI3WT
6Re27+HvD3FOg+OE593i11HpZfh3CRoQd+QlYFDk+JjsDacK1mxbdx6plPRqtviq
wgBOGH5a0gDaCTjVOKXHn+D69Wxx7WsuTRHpcEgGLtm6XNsOXMnUFqYwPVmmpjAo
`protect END_PROTECTED
