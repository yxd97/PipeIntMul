`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
en6gdPJixWpnIlQMhlSudP82LYaOXUGumSOilktbm9GnZ/pE/TFbMpkq2Ul2Wk1J
/ve0FWBQIcjkSnzoAvRkKC/BNrpH1f93vFu+ddTpFdrconaEe0uxfO+4eVGrYe3h
FQvN8eE06+EbV0kVswEAVmmk8nWF8NM6CKdQOQ+Y5kYv/fBwh74Fnua6Dkt/k4fA
VAX0exjl43fsmbUDJ+7r40ypr63jOeqQah9VxSBN9FkFB7t5k1f1yEp0IDZg1PYu
MwEL8m6uQk9cBGrn/Hr4/f2Y3igJbQ26/luF6CjMWPumzKzFMihzHM9499EF7qbn
LPbbC4CLZ2Qzt+MHU2aipljxXGqHq8U/xyCT2SAAnykO3QkW16SzD8GJmN3BCfWf
5vkw1pxVPznoL2BQs2WpjM/RLwFAo/erQGLdXO4IGKU=
`protect END_PROTECTED
