`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZqqCwBvFCCQMFhns5Lo2Uu/yE8axWDR5K31VCZjmbiN1LDNbnAw+uQ8lqP8s5AW
ChRtmo4k6M8jM4sOVafSgBt0+4HtecmgtnHEV54/MraCvnu3qoBKFYhAJDdUCYka
YteSDKaRdlXUSpaVLtV5zf+vBY5gUezZNlgFFtByH7ZUNqg8DLEx+xSlsxBSRy16
ckDPK7teaLfWS3IcipGpqSCx3SeFWIj9BlIK3E3TFz0GpoioIvN8+ZgFZKN4mwj0
mnDcRF7dtjgcy7WXkvrmuPDlV6Ud8Xe//CdF9/MFYFMi+brl2QNBbfGWJubKqP5t
ZSD67jDA2CbUI9m1AQ3r+6hTcq66w7ZJqG9eaPJ+0BLFpQfx21lNuB6uldukJZC7
`protect END_PROTECTED
