`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdPYUVhHAQ3cV3KcJrL13bhsMZh55lDsFwEd3JD2ktJ+R1Pwt3JDgHjpr1A0U1EQ
P4qvy6Q98vBH90jhu9eV11gTv9FlmWPiAPzR5jZWLijCJanWjcaZahNVXQhaw84J
KwYZqoo3ky4YV041O/MpFQyftJAxdxyihxVBZ9r51ZpNbXAUxbMuwwbRYyo49Vlu
dZDIsJntNM9WcJZU7tbzEabu0Q0GfYCY8a67GtC1Qn5uG8aHZx0ntm+xac8IsFdJ
FHaNH+qV3j1CSi7W9qbXRDC/fWB+7u7UfdlfYKHOlICNrDCyuKN0DVEGXrV5eGev
2Kr1Xrs7V0fDiqGijyJ1mHHJniXIe418LuWlT6S9rft0+8aQGZtf/R3WGC1X3mI7
anAAqqVi9v1cm0i35w1OCEWDmJJ0czXXINrdfHaAG1o0J34YtBHqV5DfTyJjZWif
cKcwi89XJCScXV7qUWzHc0F2Ao1f8+2ZQHDGrHRzxdZTjbO6wPPYXUyuDJUUYjrN
JL216yi9lmWmO8HZ/6ijoLJNjdIdMC+WrmRgl6NbHnEhJeVOjv8YcX1JBA7gNzEK
6BWaYiSchKPd514ePrgagLbDbVmBDDsrs3CyjFTHENa9Wu5opdGjbftB+4nW1/N1
vwy1Nf8NZBwacf8LmC3r7kLp1WymzbuF70Eb/Xycbf/rFRjmdk3Dx059IgClziRw
LslsTStRVn/A5ykHq1oOE9BOe7BLN8L0tyGEtq+MkKupkepv4GpciL9/dvXh0qpQ
+T6FSdbxjqBl0ef5O8dCNtzB/9a1KbZmDRLvlkDcDoLBhyUeG9F6MvizCwPmoZ7d
eNOwT6d6TaS3/pDg2hE5upiD86RO8C4QCUziSmSW0PSSKoY/fp51nnE8OSu5Fzgy
QyLW6reBCzY5l27eB//Iq4OJhorIgms1IdB0JKVxRO5dUl2OwMj0CU20J3QD39s9
XE5q58TM0UW4s7bJXCOhnHTCwFH2nVoSkM4TigdcdYP9z8LI9C7MYlcMObg6Zo/k
XGtGFBP/Af65B1OHpsA7f3AQf3HG4isn93LcNhBpUyRLXxV09IpCRLEzNYCAW4no
305IDNVdyXXHvhzDFH6iVq/AxbwruinoAAPAosRpTfuZjKVFK9uYDQo6hP3w934y
BZPSUmTGlq+F9QxaT7kclWxgzaSibq+E8ydoV6iRxZG/9dDhq5Y1nyAnPcy5aNo0
OnszVfITtwfoYNNU8SdH6sJ2dteYHtN44MPaVq8Ib4Lqz6+Sv/P1d0WqUZWNYFoU
hUxSJWbCR65p7EFQPo1eXTxyOOQTX1otu1aXuAenKBwOSwftuc8gv3urOWuGVkqu
CnRsNaGy989kHNAbgxS6uc5XczW0hNLgWOGGf3mQgY4OlSJxfz09J5xXu6dQgHOr
8LOTkzPNN+bfRqCVYrl7M6eXAy42iwaqpdLK0LXWa4UB+1APJk/xsXh9QnZmHkk4
emBUjNnAqMi3DN7nnx01EyZOMvyv7gUxzZfMilZV5batSSMKxXnN3HArlcBj+uzj
8dC5LZin0ISsIkO3l1JNl0bjzlsnQZUGOHd6BWEflMI57rl1IaZ31cKp1t5fKzNd
NNy1DPqtmRqtwbXH6N6c7xxszy8C4EoS8qUwkJu9Muu52MmbhRNSS478tPnG9B1f
XvUCA0LupV96IE6OymK544ANqd10VXfZ1lP/f7plaMwXh2FUjcBRkP2mf0zuOq1Y
whcmv0i1DjRCa9M04et6A160iTrGbCnNCcOMjZ6QUkPGd9iyQ//WYz8Y3WL+TXRA
7RyCoTMYteiS0DXffm+TQ6mnSk0lvjHLrvdXnjI1Y3MYdPzzkOM6JWS5f1kvP7zM
r5fIuHEzKnv98nwuVRb+dQ==
`protect END_PROTECTED
