`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0cGvn6OblPEnLi6UTV+8n688AfoXSOWXbpaJ1odxoF91Rmwo91N9Js7ZrMJg4QLg
PkKFSU5Kv3fyRKjEjEaAOBmPemosjDIwLpL7fG3tjinYybYmkqCJ88/PYYcwCSNN
aRvQxb4Ju4Pp5kLutf9IqtGBsIf2ojj98JU7ZVwMSIn3ltfi7JxFbxQOAscLd94a
ahDA0dR/JQABVY2IJN5MIQsAbBfkNKglusAPKsDvQqNfqsW4vKINz+72S3KZ1Nlu
JeZyXu2lHSyjPyb1/czt/FvJa9B8W0eP5Tu2gif2FEvHgvMk4UcmaP6EETD01SEl
nLbbOz6xJ/cgZDnh11HOlHMO8Bn+dQ6SDFtimjlrPUDBhAOf7qPMPVLadN82+LAA
HEBdqahCl13gTcBrA4AuiqokVP4n0SiQNvyRy4G2Asg=
`protect END_PROTECTED
