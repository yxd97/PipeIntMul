`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e42kTrCXQ87ewFTt182p18+905ikhguy6sQgVFU1eaT9bHvId9GsBFV8s0GHls7n
zzfzeh7CcLLgJB0P6KMmGCr4jMiMGxsbl/YeH+PX354RsW12UogAmM48pJP+Ihet
mm//wNgYqv3rCMyuzlMEaEoeQzvH4aNrUy4oW2R9HDRLcvUOZRwzeDAltPT1sRc9
enWJrI/BQ+5eXjCmZtB3K8EnlaVhZLBfJJlXQ6SrVADoBt3DcaOWBkNsqV6Or5BJ
llHjCHJhQlFfb7nl5bTAaA==
`protect END_PROTECTED
