`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3RXdtjE8NxRFp1gqdy8cceNxX74L8dwXvSdcOqtaTM5YLEU72uQvPzHIJwSAYLVN
XvCvCQfkMZVI6d5vph0w1xvHklyekYq6Jcs63t++BDpWU+W/EOkfhQEsARiIwKJI
CZrRWzh+PzG6yWnylv76B7oRZ+2sZsKnPNg8M7XjuRGYpPvXfRp16xqVexXraM31
0KnQeaXRTYOmmZZu+DkEghF2X9/AJkx9bmHb2jUfYCqfrL6r8jHoT4QbC7TSwunw
ZLXgrh5dASQauyzhU1/UfaC1Q65idT2GWtORJItufrU=
`protect END_PROTECTED
