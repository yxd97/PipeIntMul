`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+8cV6kVzUWMcUc/hyI/bPg5r8oBKrA3rxgng8S8DDLNFLJBcRZ0bKmXzxB0DPTa
AMxy9wfAn/WzUq/+hU+xIEuzokDS+Ysc8eWOweWSzYnUjvcczVriNuHYv5f//WsD
CUbXs4KuNjPpMYigvt7utkSQRppdO0vtIBISQp+jedXaGssRzjkRa4cOhkE3amPD
vzYWfYIIZcwW+SsfBstPzRfoRUtI9y4gFHT5v4iEUhRE7Mdw2CteaGYaWLM6lXXG
sMUCQUp3WeZF79QNvOjfDpJCOHdUDmpaucYA8GXbpDrA6IzdhYFmgEAcCuAXtexf
LFjltu8ySogQxNN/pwretZPSTLUuRRz3aYvg7DcHc6lWmDPhzA+XHu99PQqkzlcr
Fn9RDHLvPNZvn2KVt/khX6iOg5iVK5hwOdqPp3l24kLsX95l5WaFuQU3ZiDAFidm
meTReKBXUMLD9udeSEFA9yOg6k+jG0ZHVc4dXjZuJVQQEd5HQg730f7zAru/8OJ3
72ZOEVgbTgeZJvdK6eY51CrXQPfZ5xW73Ds+7kN5hCU6vNjStK9kIAS7nd+6bQqq
CReAEr4zd1u+T9wojHPASwu1bmoO4gbkUUUNAQWtRhWeVgUKNQFLAbWsRofGEA8b
YkYdfX8b9ycW9ZffGFK20ehI2+Y02TWNH1+1X9H3ddiYyndyqku/+ZWXfXLy42RY
eo/4vYuQDi4aF/aRDo4eHrAmWNhSZPmYc2VMBqebUa0/ctDRxJmh0J5UnXYE/ViR
NxqSlP27F6NFPsZAJxTQ7ncNONLBTQ6pzJjZF6jtte84B4t8ein7IY7CFUUeOrG+
flmdVDjrtJv44juhSIhEH2ohzpWDD10Q/NR03rytFhD3mzMPqdzXYw/rjF5a8dDT
CIo2dHH9Ih0gCLOtuoTMGA==
`protect END_PROTECTED
