`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6+9zFNCQ6kFwugPp19r7NWBixjWVbgJFjelGtv4riI1BX5UMwqq4//WVufpdQ2x
7mQ4R53y7ULz5sSBHq5GUyQbLnlku580RCL23IH/eoTn7lR1gz0UhVxV+T2XmZ9d
nwRVfGYct7acMUnwvVGFHktOs8IKSvcs0Wykf7UKtmA/prcMf9GJnqSbebMZo/Pq
Ew4Db1w3Bgqhr66ZzQhctHp3i0N72O+CpeGnGozW+CjmrlmiMnBf7Iqz0S15Utjw
1mACyGAFxqGjMGJo1TrvQ5H+BUsdxczG2mEsJRwZYzWutmllMAEM/jU22qUaF1Ta
JhytCue+NgwN8rdIfk0CIPI/9ZKuJwFs/K48pqiYhAzKxBmvq3HblkwvtSmHrfYH
czhTBiwo2tqPyryKQvw8G9lmZk4qK/Pc7gtrthYSC99Y0/sYMQfjzXXcR9RUn7/r
a0p997LIuo5GiLqR91iDfe7t+po4idatRIugp5t5CkjarTmfvI/tbcHPf+Duk7Bq
lXCiTRa+O+rlF7EugnEDZK45cvwPU+nX1Dwl8Daueubim/bISkq9fALKsewCWnma
NDJ1MptYxnsp7BNrbfuYq2/beDkxS1dcSflE8/sicQWOwPg3G/HhU8VGjhD7bKZQ
cYCJCOs2Qd1n+D2+rNOK/qLkYeqsvRGowExx6uIWk3aivY/6j9l6RF/xF9HSNLf1
YDhQrj9yT3Yhy8zsOj9epOc/Qit/LXhTHrASwTlkDbFreGX5ErrnQwAg3B9c4Sq7
NMtSTQCP4nDsubjqaEnbuog/5b1+CNZJAZN4loVSiiYCi4LHmOX9eDhrInrfhK2h
kjlB8nraGCPc3pcFZJf/EsdDX6JnAirUFX2+xAWuNOQg97q4Eli5SSUdya8uStcL
R2arKnIpzaQOOcQ+UIFMdEhUopodrQrz834r9QXVjnQ4Zrg1RXLu9IiyLM6edbyw
u4Vj2lSYwOIAC+DKdV2lPJvw10IRxJSm1cXKBnUSPITC58iut8k3wEfZ2ODDWr+8
SZNjgSpadBZ679L80JS3WFSqo1zLw/91JyLs1Mhj3930XdYzkMLQX5AUAept9sOU
cMkhtqS6zOuF77MHS8wxb/m37fI0iL2f2zfDAk0kV5hOGpC7F+UAJABaJ8svPZ3p
+nmdX9e9PzAXX3uP3q48Guwaa/m7BIiuMNfe/REbdE+Qw/o5YC6YSKnlW2hilhpn
UyMAq2wrBsfCIhYbwKn5NgT0TcnVX/cBqwJKQnDnZXZR3yp2PI4svbrQuFExowpH
clOXwQ1mX00YBuAiK3ySWVV1XAVMeOFnncrhRyw4s0d6v5gvwsHBiWi76qHPjyGP
j/ya7A3qEp3xpUWQUHauNJLLGaBdpHNCYHvJVgppkBCl0ouhXgeOGnBNNryi2pge
4V948T6pqtTB8V3sOjiTvOEHupcreHMMsqSZuRO2DeedjdwsPemJplOD458Nzcj1
i4tSwFw5oPncsj6b8TAcl5Lebo35LY3UjENRx0XUm8qcaH/hPSP0+Qlb9xMY1CU5
f+qC57JQS13ksMIbts+/G6qOf6ZwFunMLJn39846u44rRrdAsSuci9Kzobx8YR9h
uIVE3LaViRxqsL6fTRTfK+Tr9UBwYVZv/XvQNQtNmTP0dDdnaQ50JfeiAM4Skm8+
gvXeCUf3i6Dn3/NGTcrcVjd6KiLkiCH00o9BjEEZO8gzt/NDqlcnQwtSyR+y+cjc
gPMRROKWhZLaPuSQgDGfUHnRDA7NxSy0MDMKECidFYAeIuC1VtlcHONPtLaOlCls
8++WaoCwQLe76V/EJiwnUcWBsKmkKduiwO/AbPDwoyrm09Wquaz+Wpmv9QW6nmko
QIrzpn8cgYkEkfbHWYpU8jk2uo8cQH4JmeRf4IJNr3mBQpRB12cZPHD3WcKX6I22
NdSp4CmZhwngj6/kxDBbDqQ9qioV/ALpOOfw46SPiKpJbvr3y1dl/L5RA8gaC5tx
uIBTiUWzvU9rB6L35wVMOhsNBhl+EKkDaLNWA9Bz9EHDxShrc3VH5WXQOFMPVe19
g5c4F9PjZwx1BXa0veKx8WjwLJsGI0DeKle7SwdMmvUhfVYXcPXrFhAsL3ORUEeu
8vocoMjJAfQI+EGx1w4cx4m7tDTa9Fa8JZtDVhnjJkimxHPDtT16VyI0jIqGq4/r
WrB00sbXw9xjVYrsHnctULtuu8GD5SKax8xesI+lKSP+PPlpLo8OFO182n0ZoiAf
`protect END_PROTECTED
