`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWUe9QwR46guglv5/ZRcfcS1bcK1KunX2mY9Q4PkQJ1WhIB+GDo2A6W7hzVl4KHp
DPWDMLN6Q2JPpTZpBPB6ydo5z1Dk5xbcuzImLC1Sc8v+Rx8FCLMK2IRyIwmDpVhb
vm/PKTv6+sBPppSP9xVtDsufhJhS9Ywell6dcw8TPC6XmonL7Ttgh7ioKkG37kLm
mRdCiF4JXxp3EPrpWkJiQdxUuhr3K8WKrDzHf7pL2xAix/8+7KB448duSwGbha3R
FgR9jBOENPXOJ8Or5w6bcnn0hInGU6p/hYeJGP4WPMTFor4xIcgrIszBl8ttTQEZ
MvHzI59wZ2XHIZqr6zeC3lG30kR2cErYLqE0MsPGwEo+FQUs3jAH4iNYCXhVYVwQ
6rpv2nst1WhvIf3SA+vcUbowtJGN/rzBlNV0CUtyXl4/chhlyAzItypbMc37AKIB
p6gurb3UG0jvaJM8ovNJ6gCukEN+o7gMu9frv4zEBcvC/nr76Yoo+SpYLKa1zCGX
vdXkOW64OgGEuKUrpgTj+aWGRYqGVnaJKOnNmAUtz7bWyEm4A6fvRyjvbBfLQrVf
PW2SFI5M0GYQpZe8TkxEl7Mi0O248HboffXF5B5sFlt2KTq7aoGpBPFYbV0gV9KP
1lLGCIiBaGIinPM/Gh/kal+3pn5zYnltJfoVZ6uiCy9J0Qm/gVKfRce1WTqfRK9/
8Oj7vIRhZijvf+KRvs++dTZjizozEaAm9pe5OlfXEU8=
`protect END_PROTECTED
