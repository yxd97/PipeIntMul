`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T8dpt/BfRl1NufG90iucFp/lF7utzO6Zy99XQBGltGZQM5GVZw7fUXgwS+/gyjVn
F9RdgJmSXoyPLeM4++IGnDrTsxX92ZBECELaYHyUzzTLFiXE8/FCE6OVJd5rZbNw
h5Gcds8Pj0fpZjoFOXrZ7R2EPNL0GzfEXq13yfNqp60nxE9RRSBFE4IzyIw9k5WT
o56ne225PgRjO6/wKDjIZIOIvr91XEWyQfSoPpdn7sFaw3IYlgzLFN1u4k0nlFQB
ziUNhPwo87ZCncjL8scMl1JbXjxwFahTlf+l3lk/drWXpbIzPjcbXjDiDyy5rAKg
q1F0osfjVIyd0FZTjEa2plomomlQ9rmrWVbpwLpdnD5gfNezHn3BqTn4xAMB2tir
ArxoAhw2vhJZMJG19caq+Cy/4tkjA0gGCfxqwK2nv8y9WM2vJiuQExKIjbE7Ie2D
3P3IzhwH5NXuE5f4CeWTroFk3c/kgIY0ddot3SAuPcrJH3Fttz9EAXbvNSOJ7O1B
13PEapj86tRx3rUIdwZ2g1pDNnmOPdyAIAJCRiwcYmRfGtTA12Yg5WpH/sFRp1SF
foVvC9hYujlaum/dp7hH/CYINJ+bhubgnlbScJ2olZQsB4Q6V7p8g2hIwjFsgEuk
YujlGRC3gIXs8q7OuEp0koLOqKyxHRA/horiITBXtGRqnvxSjNUcFRkFVfoeNqqC
1ybBTrzjOls1BNMgM4UJenx/OZTzBLODu+mBAQziW8B6TkfNkrZAlIM0R5j7IdBH
0Ba0fIO48RxXEosxCQeRSe+84ziDZsbbX1gnvDuxYhz3B58ZzVDII3YnpX/9pTrv
yMGZxIVJeHRmHI8M6I1U8neybQl2AgmY3vl3JBk+rnOlhen6I7hDej+90SCT6dZ6
nYjkRN6p3h3h41T5tV0RXWNfEnkk2kJ863tUx1LJVHMnrLEL2ucnA7I4td5uW4OR
QRV/Jy8s7yjp/JHw+Y6BUAuh8qm/lRXZZTwb2iJD8E07b2k46ia486CLC9mAPTFr
W9Y+zdWWdNKYBx/9NiOVdNpRv/8tEOu5JUTlmoLAhEA8vubn2rPjvML0kzHbh+En
AonKQKeiE3TXEZ7/caTYIPiw/ufeH7ciBiNyTTubY2DfJfNZ+BhbUWn+nVWOF5UA
M8RF1vg94/C+/D2TxRQ3WG85duWU3XpeCB60vICaEQ9N4QyylyJUR6aWJ8Ar3oES
Yq2SIIQzXwZNPiCYFZUTV0HGXFaWu5GjxMZV1bUIcLqp9qgByCF/ScYZU3/MC5it
J20Jrhy1C7YdMBwRXgjm+goBD3dLlPX+U7sEZKGSmG/fqoqYABfwlYgTn5ht3Bw0
FGpRbGgLvWmSmB7ZHC3VB1TEvcaRLRgJjPMgS/ORX5v7Q7vO3sikW0xLzXMS+WVK
JKPSeVyWHI1stskww7t1z/ta3KG8M2UseekiN+UVI83oM7OaAZwtbnsggLR3eOq7
Ol9ZsUjXgn5ORtSAoMsL9yRffrYz1vc8biXztuG1QAygL9AIm1tWizBQBVNGAbEb
oCzHFi2Ob6wMCGpwzOy3Kac0+0XQBRjDwaCHvCoNrom4hEXuZkch6+UTVKRb/GLH
2OG503hLApv+/pwdUHKPxGkKKAvLfoIm0FWrK+7XLBGqM3zB2ffMPJW4vidObJuh
vgDcw8i19aOJsu/ptgXxBSxvsOttNdcHrDJfnm4+Qn3OuRyTT/N6C2ZaOSO0F3wb
fa8fqBmeQwzik9R35e9tn6bG3K+cfe1bBGxNvLNX6tGLb49IwHUx/+NqyihoP31w
ka5WmNtXJF7yzDiTIosDCfXKZ8qR/wMuSgwI8cMeK6AcBOmp7ePuXCja2hbPVr+V
19zR62BbDICc7IiWaAgCmsRuy7JF6f7b8DLAvW/dLuitk1wVkZ+VDWpcSOdqvRH+
2T80oHxw7R1TpoOdbQ3Nbpe6E+wnol37Ki1nMmV9y2buknnRRePTmJaSMx5NlTsL
+JxhWfoSXXqSoyKKlsYQlGEPVfzF18VsLjTXOpV8earVhAKdqklU8M99VE/42dMt
N6dp+tgiQKu1EEL32/NuOQvSuTB1073491J6YVyPf9Jr+vqopBakqmMzeaiHc9eg
4Zpip1STHzfWvKrieNYdxa0cC2RUP/oZRAvMorsYiAl3nXMVlg0PlFISh1ANWQsB
Cq85XhXpp4ImBwsdR27m5z8ie1oOXXMn8l+Cy8KvAiYd6bjiz4Fu1dG5hQ62Looj
/4ynD0mYfu8eSmmlZacgHcviACYJ+sp62yUpuv9kcmUyoDcqw1xdXBbXtJYtzelN
0bYMNdnrp5DYL+jf/eU6KCtiLehaV/c6rLhQL+YLdlJ74scaGPs8IAOJJBa/ljp+
d2uxHpW49GE007BkrMLfb8tcimfJy5QhYtE4UiSSySHJp5wnivf5rA6btrpbSlDz
PhE9WRVcWiUo/WDSD8BoDx/cuUe3JFMOp7a5qV9W4j/4bMo6UjewweBbaR2bFC+U
iQ2SugP2pqUOtTizhkFPk70dJJRHICOshPKQi4d7NcYGF8yoDK9lG7rbYHwaS0Ae
2GtR7LLx2dJGxMrljGgf2f/ukrgPyL/2G3OjF5uupo9HB2JUeusIHhP3+a+Yddwh
1ik7jj6fbSYEhcGrE6S6cuUkgoC2vn7ZP2nep0Wk3/jPRCrjGMF3x9oRnDsr/+mT
Z+Z4Gokn6ZmXH38z7edw3OiNDmDLxRlqdCeffl8iX4vNWQX/O9hb17CrOVJQibMJ
T/dH1guV9N4SxCx5JNE/r+BM5w5yvdQQY+E2sQrAd2IzfbrOen5lOpjfBRe+A7fS
60GJRSRwZirL5ws9Ue7HhCFnNL2+D5VhOEyzjDxUslN8AatDre/JsIHhsd4tveGy
ByhO5UDgHEVrf3UY+ZII0BceNOwX/wHYSIv0W1XHR8gA5Cvd60DNa4Pq1t0JQnYN
bgyVwEEpaQ2dyI/imOe9iJ5UBg18fihvMLb86cf5AobIqpQzLJa87y46Dip0IpfX
xWQbz+KkKJ0os6qmgmBaCYpRc5qihBk44weEFTvjrb5Z5F6xTJ6P3CqXr/5t3nSj
0Tr0e//+Cq1YXk4Rz7G0dzgSKqqeE5USQAQZnRX6cQg5vQZDPrNENbx7ILB01YAI
+GDntUwaoc4oTpmUOZRPrOQiFgSRu3/PkjIp1RzHXBemGlArI1ROWsTx2y2JWIrH
o8at3D01/Z/olALpczfzeMyPmilBWTAkS4l1+xje8CQWjJjwSPMOZ0+X8dByfHid
bFhkpYGeH1ls7mnnc/wjkLdNh2iiABmvnPnZWEhEkecZ4w/idztNf1xHUlvuUfAx
SIkwluaimwGKTlCMEPGFjsWj4mFmv+AAScp9aWx+CxNUqPdAFZstETQ3TVSp+ojv
kYBuIIDKGen+17I1Cluv1j4YrZ/n6KGLPcZvrGPgeMvBnDWkXm3ayLoC1IrPH3dF
3Moot3VRptqfQWOjmLTJEk4xNGUpQo6u/o6nLF3iK9/gtr4LF3skyuoixcx3iQS1
cbqQRo3JNRi/kPTVtGGxzgfpMNirzEvWPKrtTIzKkEhEpcIDq/bpg7jOq4kPA0cw
LT0kjB/Y0HQxinxwZZtTJXI2AO5hlFK2yOumqS6oKzSUoKg65tsVH94T+HjyP5n8
51PiSUVGP30cf2U9FOF34KD4ae7l1iPLqMumt9no0yiIK3HQWegE+xYDdnhFN+3U
hJuuzScatou9VxsZtG4X2wzl74bxQQCc69En3kaM+VkleFSrS4aO+hb1hPteJC/7
JzkfyKaeBE1GbtNyByLkajad9pDw4xD/uUm86PprO7nkrJB6ZDmXwM55lFi9psX0
4DfcvP/S8lJpMW4mcjDuLDOqzJNA4wfDXkZVec7Luat/1dTbNQJyx4U0aN0Ek/Yw
gcXIX25Ely3F4R5/j3pyDMVdGcdwrdv4mhHHfoCpsFXrB+uIUAvX8RdpTi1ZJvcx
bpOuhx0icLDpe6pHyMFWGc0FFwz4ctqj6aHtR0gELeES36iT4MycjzrdzB1YXKG/
eKLYAaX9rLPIHOE04OhwEAET99vCD5tUCX1qG79O/6xwxYFVvIGlX92QWRmJFtsv
ySksFxNYPdBsGbzjigLzYJEYIDs0duShPc8zdLiwutLjoyziIOT/JLZPLXlZlyoj
F/0LGq6GelhSSjI8QUWp2+dZtvP3mLiDi+6vQ45JOUoVu9uNpAkNOC/0T4M7NcNn
TKYXD4Vw5pSq/EHg+/NL4m1RCK2auknP4J1StYyCIiZcfxhaRBU+m5B7TRqZ9FsQ
wbKdAhbHPxBYp0Sqr9+6UX3unN9hkGLWP5CkZkEz8nVAzqB8NmX+K3Az1K5h1rWA
H3EF0O4h6oJLC5WYtD/HUY3b0kXq7Y5fQejWge4XZmvmjy0pcgnsGlfcIobJnABh
nYoO77YJUsuTiZIn0lEgGhDUNnfS9N++uZMyy/jpZ++2i2OLb65OBPunhrEsRhPG
gl+rEkdmCwtv83iNRK8MHVLqokkNVmYYrzCkoocWAhzh++1PsBZCjXOH0ZgE5W0i
caP4AegYOQhU6wL/G+mLV7qIya7KJkKvQ1xPB+vsxB3I5IiSkVoiTYYtZpbn1NAQ
QH++vN7vEUW/Z7pPiFoj439Qgp1ToUT7QkWmy+6fCSqW566/7g0mlLiHzS6DYF0S
146EgV+uOJusM0qklw8cc3pk320uzYYTGpLyNY8NUoRnvPqUhJZy0jlwc49ypWhK
J5zqcnEiI8J+EIE7RieYZ8EXnJvQlQuGp6GHviC6Eli1AXlGzD4NYf9Q6YUX5XTo
5I/sfs8RO+azoQiy4ntfyZhh0EBgdfrZtdQHll0PabnfhAKZLSzJoZijQRTkjftz
/WqGaHamTTasTeEYYav/CBm7fo11mcVl+G64Hrd5VJL09k616uTXDIwQqhw3Gqt3
DRcrIF0HCbkzKYfTxxUxajgId0J8PlAes28aOS/58OGOeunPl6QpkLQpsyBwzzgo
+0tXRpoc7QxifKWoZ8gtmwlTlg2EXFwhlJ0Sw/jWfM9gtN//Jd1RqtX4LGxXF/nv
dGioslDQXcfxBDb2UmiZxf3Pp1LgqZxi9fMnR8LuExwX1OUD5gQsC4m21QxZpB8D
EkISDnnM3qbmaiQYbWAE30342iDQPeGgZ1ZY9vhOS1w1ZQ1JL3pwOEHydW0xoJ57
8e64L9SK2agIEui5GhLhRRR78h3z+yxhsNLcXFV8IlCgE3W1xLMK9pNkqmDb1ZBT
jeU09wGUwRxuSwjEK9Q9/9Ga+vS+p4wpjxLCeaF7yWli3RFKgEk44QKto7ThP0Ck
VzpgTh+b2T+7XX2Yu92xNzHk3SfFROqGFJQvUzfrsNcLqLrpnsUtT+snWTnW9+1s
bNqHFAyW4YP93vc4HM/707Mbtc758PODUWKFVb7egxcwW7NsINiQAV2jR0YhD1eX
T+FC+fyRNNv8wUQ2TbFk9M/UfWtc6E0bARl1y+hFsf0sDtYEsilygIXBbnpRPOQu
QwaI8cmUUCRHY12cAialwZNs0lsjutu2gyMVpV8mOiga7VWJCnEF/ObAt2UmQeJI
rseFpLIBqFbd6p2yBGGYLqseSX4q1AOFN/orx/l+2vAhrGdsbmqsTl8GNhiGOHPT
Xjrs4LLZwOw9uC5f//x7S+wXn/tu9R7jCu9HaxohIYjwKN5C/MmDcoBiHHH7z0Rx
BvrTUeXfBAVFgJYA5OushDwfkvLI9382dQ68QZc2sE2iXpKWzexLDKRXQp7w0SUR
5+GuDLM74hOTZIy2wtT9k5PVaRdIZt5UbFi2F+nxsQvdn9lAWkCUxg3dTmzTBwwq
enk+W5zus3FkcBAA2A67jUAFeEYACiSkq9HxDD1fXjnwG0ffZQqs0H4lyDkCHH52
2HA5/Czn6osZuPHZ56TR21edqsRrbRw4U9SZ5cOIC7T4iRy07RdjZMkSTCVo4oBE
qJREielhRXZuuNO1JCvF5VOfKaE+I4V5uxTv0V+k3BK8i4RNZLBpqRgwwoPC9hfC
VRUCdILmNWpYn6LdioLCe4ZDhy/LbORj+ihqkY7Men7x9BIuLj5iFUygX4NokG6D
0XKPYzdQ675w5EhpwYuEppT+K2JY9eQV37i+iUVtavYhx10QkGi8sSQKxytzvYEp
2d5s/DUTRHie3V9vGKWKnHBiHMXNZB5zoJnIFlI/E2KQKdE/FiD+oyVI6JTySmi9
9WwwUJw5geVHZDcW4vbyQFjnj/6mgtJ0nxtUOmvjc6Bj8JKTlJ/sb/oxgpxTwkZW
XQJ9hMECmLo44P4FpWFDjP5Nx3oJhzvXcfAjCRpgx6vDWk2c+MvAA+pQFb+dik2X
MSuW6P/+PCE6TJU9ah3m+C2+rfmkAIOcpprJzbCueX69JVlF9KRUMBm2GvIYqqUQ
hBIcAmVkTFGsRtFqx7d8hf3Gp7I4x3YG72bj3HHXpqNn8Ux2lxFi5T+CntotyEIn
3xYXxEBa+9kVyH+U5dWb4ieBvxPq+LjUHwz6cJaf926ahmGOjHTFXkOoMN6ViMWN
pVi62ug9ub5YDpduyCF16+F6g1SNzPLGsR+2mpdEsvC3L/KSeCOBhSLmp5wRMlxL
3BNCXXx7Y3i9qdfBPOt/5EOwWlecLSF3Td08RNIdA+y5UqTNP00uYX/xcZYzvRDy
f9+kUALzcXaaL6alD7zHSdQrj7j5TvehbVCRudfcysloyLqEY1js0V53q+bdns5m
f+W8i5082nndM+Ywi5apSd38mTQQi3iCmZqpS5OMxAtQk9NYGAXLw76W2tDG4stZ
vj7vSNeU5jW4/IEt3cK54hL9cTaLhUlOgNe1LBbUl7odU7sliBf8sBlh622nz1jI
x4Vn6UAHmDPkjX+Usw0JdHUkuHn1b4a9fU1XXK5xzglUuTQxBwJGwkBm8YI0A90f
7sZ08HYb87J3/06hbzrQtiyg1WRpMCYeBJM8xivrrQRVGY0Vp7DDdxQarTKGxeQ6
qLwaLk7cjsumy5LH/tjOZWo3rv1Ybjc4RR/6s4GHZWvK0HrBa1A4std0UxnsfDMQ
tpZWmA+ftN2SSynfD5FUwDfT57WuMnwK6OVvkDT3GRdzLGXCFhCQqrwbHdPBg4mc
4ISW2XaJL3+VCUyhIJcy1fASfYz/TfLUPWw1/i6xms2McE+qwcbJncAAphFDEVMi
pOb3Lc6lBDWy2+FI1Lx0K7Nl0QdXh/vYOGXLSVJzEGsVp6ETXz/BpEQUJ9rwCCWM
P+6H/PjjX+iAYwDnZrcfljLidFlqKtLkOmv8Nloj0RVUAUgpgTGoVJHHnTY7/Mks
Tje7OzWiQr/r+UyH3Ol61XI0Tgk12uu4q6t3ECEsfZwbloAtPWKcdAGP999DFcAR
L9t5zMlRgTR+L+x9/SIz8liIm2T2jamhvkIgfPmZxYnHlfXZ3tADdch2cc9IDtFZ
MwVAciog0piB/CEVWsgTDtIAPIQbrxw9sncwwaeDqpeEAjXPJmRsmdwNOxMnRxRw
Oc4XbsEqYrP9zuAG5SWoK8HplMb+2Y5ZQ0YH+K5FdGTZF5K1bZDQgDNso4xlarba
K+6GDZTajMOpXd0CGu0E4HsO3dLXdudWcivEEK0Lt3a8vTevuX4bOaFDw9xqMKRO
q60UD0rzsZMBYfVuV4p7qpoEDL1ldecXmGmXJ2bQUquxclfmKBc3iPG2fGv2SQOg
2LfW+mUHdSKdF5fCNlY78eS7WmhVZxayl8JKrDMhRrMXaqAuRr+81gtVxGi9TQtI
l6phY/F7OOCmYDp0tImJstCeuw3Fr4wJA7JUiQ43V1XgSr1KWt1Fn90WXMtVpYmY
IKvtacLkENckjQlgIyrhIG2ysAHxG2x2KPIUyKg/IDVw1AXDpPC5QvHJxYtme5HQ
x2u6NZ5PUuWlLs1hHi03lO3WbEp9xmqzQvdAV3Yov3l+X0RMIJTxBVcKbhMK8EjX
nSDfPxXkLzKf0ac8aEoDoKoymRubk4nFjNSqOAIw0ziTmMt21uyEJv1KYX72bzxR
G0pAhagdo4wX7AF3ieiJLnfwLpAb5+qNxViy15nOkP11RYiuPpA2QMRmRZw0rf/4
hj7vTF0L4A0hGWzHMRbNVz1s5QRVh7RDPTqpsfVTboM0xYuTzdd+OsVL6hHD8jyz
BMaQZER7SmB39UTJUFJF5vwNLkJE9IBlaYCMqqoS4h6wejyHQd9m88ybAB1WzXLp
UE+WX98HPv6VCVD35o3g0ZCO4k2T/07Ge8VpaefY6HxGMIUylRmH6gcFVfGA7y5r
RUsEVIXUxX1c9g1+eGGe7BNZIJ0MDJF0XTGy1tyx94foOk57xeo+gSZ6XIVfcj6L
1jX2AIkYi8Pepy12WwFUrFqHAsJRUQLa9ATyfZPv4J4NneUx7Anh+C0IIGPsuCJm
rrmsI+4J+OopdHqdC/kpIojEkT/SXqGWrctyKWYSyKag0X5gYZ1RL7xpiWDJLY1U
GQEIIL7W/wJKSvw4sfDD8HF9AZBZFekGW2rF7Vqu7Ed6JZkV3neVqLTr+uyFVbPY
jRF7FIZ7F1lm1kaCLirIMDh0lu+lkYTVeuonRFXLqD67JlwbQYR8dxmzHAFv63wG
D1iMDA5SXOe6XIQOSgiyR0s9rXHf7OWzEf1kPPmtKm30tOivgd90orXZ1pCdkD4N
cEgpjoVDaYW0W4Ln1G5DGd+nbhrd1vcEET0JXILHXjjH1/pm62YvohNhrKWezcET
TK3SHFiO9ybwqB3fwk1D/+mrkffD6drENxV7FtL22GWiCRgZ9EqYZgi/mCg9k364
qccda38ouJY2JJvUpaa0Y1A9adsL4afYaL2W3UK49b+wX1oXBwDazCFhkKRWaeNm
YfoMtFD7xVqpL2fuq6YT2JP6gPCMCn3Lc5wepYSOJYNB/1/K5x4qXJQeD6r/rgLA
38MBAvd0Q2QY/Nnvg4Qp+as9ZReEVsTom2gBnVHwvnW400fs/Mczhm+wrJmxWwnk
5wPorHQbqd94D2ndSkQYDer/8I/UJYU3OJSh59TI2ygL3Qqb8NmCuHgcYdOny1H5
OeF/win4fdH4kDQn43HgB+yQJLV2nOdsor1jDv8LUAubNzZn2NZNcZ1lqZP8wS1f
5U2IUX1AkuPcrYZG99DNPBoj3MMvq/+uj3lbK1365/7i/SZ5FJqHlFoJMcHjtyUu
rjx9Kcou8JzydV+NdFlTyWsFizjfL7YLfKlmqOg8ypmC+t8P+6VWyNRYk1H+P02F
SqlUO08TzzLfkYq4nSXExemauuDZq+nuzgTf42fKkZQQOfSn+W/1VxJVqTC3cODd
gqlL7h11O7d1gQBUqXx6qdEEzW6kHBjqs2QD+aYxb4GorsjM/HPNcWF68hTa3ntv
A5qTldouzxLrBBk3lhpLcGdk9KFeK/fnlOTOMJ0DzGPtaiyqsnGVaRpQWo2q9MDI
O/wbrYiiLMeW0gUpnvfhF3DR3d6Cr/7h3b1aFRcfpJkci3UfNq83m6iQ5minxIvj
bCzrNDO7yimPTJdJcPqgXua8PZYNd4Rx51f9tgc8qM3+N/cS6eEbhAT+wQ/72TJB
IU+cP9dSK/NVFOUzDikT9qXs+DGCqEgEI4mhepGsSBwdpwGO4c/v7sVesBqzS8CE
QBSiMbcejV8OsypGkbhjPw1c0/1Q+MGT6DZsZwHOl0TopzOQqsWGOWHthbpgur2V
UNi8MtthAX+QMyP7C57IyiL9DV99iiiM+rZiJENv9+ExWnTsG0IFKW7N/x84GrVV
rPdSvE3kY2fk26wTFWOruZkGdohQeBPW9O1+OvlsxVLUFh4LIGgStBWUiRkgVQpw
ewvQRas7GkVPLYQ6OuWRXoICB4+KCrPfKwtjdnhIAQeGah97MOC0U6etCojN1irM
6RuhhSA7Z8HfVttkO+kEeWYNHuW9Iid4KySUNAWaUG/aBS4HHR/7V7ANHlefT8xx
u4YqK5yyJsKzTXdpkTlIPkV47xhXaKsp5UNGCuNrJfmEpeidzC1rrZcZb/egq6S4
+DzpxsvMwaC+MLz+/ecGRq+c6xv4xyuNtvV32en5FMLOoyNHBhauoVE2XAS5ZTsK
2vlXuggoIsbmzBCnTCqid+Iy53kD5stAkZ9DRh2kKHh4g6z42a6BeZoC39CzskhG
6cLxuwrBMpWT0ILdzPS55S8P1r2x7NPFiT7/z24s/RUjcbVwfSC1kDeuen8eW8V1
21tlk2to7i9FtD3PaoHXl4CjgsrEmuXwryLuKFgMJEvsqIYJ7hKh6rvcFiOxHZ50
fR2OmA1hKOjzNbvMLIHtzC7bwKXDIqTcPBWrydlIG2PWSgThv+PdI5KntJQoTXuI
JzsHZKR3I+S17D6Aglh0oDd6DuqvTkSC82/ChuS6NQJYR76/04EvsXl/eXN5sqNu
6p7zdl5FGGgBQK+MCsnrisFpOfkpI2Yc5ML5Y4+vO6SZ3zl+VjetgpcP5Ln30JkI
Zhx9yyll86COBk+K35UwAGOCl6qwLPNdsY07XWYV4sEGiD1WWgs4eH+po4/Ml8JR
jSdxspXTBTan/QDqP6uKHbKPMHsqTq7bh9XqpNEw1iAgVl0uLtXbklbtCTWTlOTo
qclw6tJ2JX3qus32ywxqGAekI3DTeZf3T84ILhLpHgTCjZ0/gnZDBZ+cRrBsreas
yN6kZqW4aE7W5GgZ1Lo9r8oe6Xmsj0spSqANQ6pAF1IQG/PQ/iPnHjrmUj5/Awzi
ZKYKXhPnQgwPCn9garc+3qjQLoL/U3uz+ZkzsNSiZcWp0SQJkWqq2hMi9u/mx7FR
/Iak1rI6RvexPSW9AN/YHkzxdEFPWWXVLE9j+zbS9YsssDYgIkW6QpLIXigyFp+h
pL0cvQ5rTGOs+iEUfOPe+s4ync9R87+EKLrgsKdsJrKMmotDDgQZXZfPrmPxHbiB
S1OObirtFUEf/WloWO21gNbLYXr8hWNKFnTdVzAx/wE55LZRLQlcrxogOe2oN/PC
oWeqoFkTvnRszOsRXt0fKNFIyHl8OPCA4YcZfPzX97oy/cGi9uV8QelOx+Llv5Ng
6l+kBukpRnk9VDcfdLz+iEOjOCwwDcSNXI935PoWnGILOX0hal/RGyYEzhd1xdJi
w1/AV2/bCVjhhy8nVP8/Llkt2HmfZawElflG29dVlcaYDzV0jzQ7Gx40Cl8AC2DC
Nwh/wyMo+2aqzvL7EzZDlyRlPVErlMYq3SbmavDTA94LW7ogl/H5/7zf2xpNTNNr
YP6bLjNVq4x/onLz3Y2B2jAvqhZadcnl4nbvHaBKAPqzafzwqr8vHTkTfrgHNnPA
kRQXG02QvaUBNDDILuwQ2luFa5disNhi8Iw+cx6egAMID5xgW0LGgsvxVrkLlooZ
vaQT0Gq2DPms+M12YIHJxQxnhBmrJeWeECO+QftSlLCdIpuKSEiiHOUESY2G/DsQ
AkEmi3DzPYaWofF9eayhDlQ2z32fdmgA5zAH5vtApF2YECqskXZ8H+EQQsW9qAaE
tf1V6feHrKM2491KTp+Lcv3rebtTkQjdxQ36DRImIq8PCEStaeJzbCgl8EbpjeFA
vnS4sRuYM/yUHDeTX9W1BIW6ohSIYj9VRgL9ysoMkQYx7uYPPQ9BDSP9Zov64oVE
L0OjnTXqW9+5bXtwDS3B2MFGVnVm8cbYkAWy8fiq5UP5yVM1J5V6+fgCMBP4s7+A
AaeixHBBPwhaEZEAfnaADVP34tupuAq9kPF1Tr07CqVmFSJdZNDWTHYtgSgjScIy
zeZarWA5btvcLhEE24y3BnY0g9S1AEHDUgqjuwrCw9YVXk0utawxISO4HpZfq7+u
ApCJwHjrmKHcvhDE6xIIsykw0wBSYC6wZH1ueFSCr3IrfEphojgDXIpXGsWJ9App
UXF/GLLvOkkDGPJHQXHX8dRvKJJSD7dRYdmSVj0QttncdR7L8y/81pvrcRl+RZ/C
p6iVo6w/TydQU+BLfqCdFdkxuyrxqqcAK2KV95VEHAmsHitbb+MeDKTVPNYFdUxy
5As0PJVRFB5hNQN9ulNexWiAqWjQg3i2yjielqGRWYp6+nI9lH8mhDgeswBfDf78
BdkLXxEm/1Nwe0RVOMD3GvzJo3o6jr3gIdycOq+EBLpMRgnNrDL85h9YLQP7uZQQ
XstosElBtIjMv/w+xcetViqmI4ca4v2XNk5h6Ndeg4jUqukXmN0aV5qdOSnH33Z5
BQ2Hc5l+CqtYQv9frP+uNPbCPoUonMdXYnBtDhZuEGb05ndj5kkNsKUAUh2HpZ7s
+EIZLJiKZV2UKoUJWHeHYea0+63RbT/KDh/84LFIqefChX2jWODkEpWzXQqj1BvX
GVFqV//xliY2XALTGQlVoDzEcG620zPaPJ1JfIF96cwAiku+xSCOp4zklK//uPOu
+5z5UQ8udpAQ+Xngt5Ly4kMv+LIUTVAbpl8SB5z3V7GkLodxBbc5l/sUjujoImwZ
vIOGXYOJREXGD6L8pksxEZw98v4VR6jBPNsVn3nEliojxZwzIr6muhyuooRJQBSz
dm3EFoBE2A3kh3xHvltCNIf9sFo91U5Ujoo/oiNpgSl5491wOPnjzqEY80Km/FnZ
WqvJwRSB/5eW7LWHIvMIkywub+YmAzWOw3824Pqbj84XcUO3fq9DrklgENl1EmMV
gMTo/ibKldnsiO0rF3W5zeDrsj+z+GjHx91zW7vcseJ6Z2t2EVwsxGRNzeUJPdMI
omMQCCnF7HiVm217jbp4SctNvD1Yk1MXesKBhZh6S52fqKMOI+HCHLSCtKnE8rhV
kiI9V1dtiA1k8lb95vNdQqJiklbJT32es8ZDyO5CM9Lghaws45sdQnu2GKKEvzkV
GYljjt+874DNhZZnjghg9rGftjfujHv0rzSE1fdGQVm4p4b4xHrfuGNrykf8CVJn
0J6YUz7E0rHJBYTogq/x8yqOWVf8dOc8sNNZfjurtuatgVAmAzoNdA4h/quKFwvl
0wEEFVO/Glxx4Qf3BV9Msd9g8iP/0aazAp1hgSjxMofiuToJh64Hn4+ePFeezDxi
eEY1inFJnrIaRADIHaUAYOnckRnk1wcMRQ6f3kZ0nLIaFb2CL3Q6mPYzziB1H2lc
2/6agNI/dwpHezJUr0+2nL0MondvI7bMBeU0H/L/sTIi1WtpAHvwoa5e8UygulBm
WwM6vKEtZ2mKfFfmxXiD3yiPSHj40TT8qCm2cb/NoNtwuv9hhCQQ4AKvOb0WeRWP
ugrJh1RcFNOJPkB4JxWbnktEoLArrmkbFRg8wj7xIfgwc5lkY4VzLcjqXTH2nQvy
V5bN3euZBL1iiQj18ndlSBWSLnn6n798oVg33G1+1Tp5HACse0NGcZ3fNa/EERqi
xM8wxguik6ZUvCxtrpLXL90w4LsyJbGUMinF7YYDQlHM1SSyIlp6XggT7vpVBoFN
/d3Bl8HJv0uoX06zWQRYkKT9O4VX+CaZOYCJESn6btcurHzQdttXYvKcAD0TrYTJ
hpOmZmEKaupHEYGsO5pcGPMOmchT3bXSuZxNDqzhZA1p54L6/xElMOUV/7Aq7dIU
+P2gj+oIczPKbvqEpDdzi7wDlVzA7PYVoxyE4cNQ4/vm4fVqeS2fhQ867oif+NKu
YxFmXSRWvcqybxnOWj1rzyH6pWhSkNHO38nNDyhJw1Si2+5d9qjwtBBUuycVp7vl
NSkAcUCi2PHE+1GiVlLJXP3LHGjizndG1BncQJGSffxDEO8qqnENpDokxNnMlQEk
sl0A2w9Mzn1+XV4Ruva1pRXuST63mYTGAEIkTeniNm8QpcaVpi7AP4mIWAw7tH6f
2hYpghQPc4v7apvoEyV63yloJkpEQ/y6/tynjHbsKz13GinqXkDPNvA7NAQpivb4
4Sm/1SvvbdKaMIYKEM4iHh59YreV/z+PE6AYTFn1Mnwx8ZLB+cqEBwfkWkDgpm3e
msTBMQak0CNymSKzG/99w2Zma9FoSuFISKV9n3BWTjfo960MRRkEi6+nxngBn0gA
NDkmjQR/ixZqVjz9yqiuP/lcAm33bxQssda558UVi1wJTwW1XpXe6N73XUeRLSjx
jQn1gg87LDakn17hy5lSO0YJTZ5ZBqY2w1w7BjZp3vXD6IztcpiKhAqW87Mj7w09
FUQwmK3Blhl5PJZI3iGyNsWTBQU09rEPi8p0+fn+2rhjO9bfd7nWtf1uB61FcBve
D1+5HH2F9U9N44jSExQqjcoYT8hZlh5KDVtWTez2OZ7hgCeqM6HTzzsROm/Rf5jh
vbZGZ39j4TWCh7DLcMS8gy1MlJYV5lhexiOTijQ/Fzg/ycf/LSymqYG23QABUpkK
25KfCqr9MMgdIT+WBlsXXS8XOM4yKf5eG6ApFluo33fg+XnDC5Xn5o5L0M4FA+ug
t4MXadYlcfK92qL88qqeOQJFz7s5JgqE+G26/AKxEruAGtOtBSUuwCrCpb8Gfy0K
6a7ldQ5Lr2aALZ6N1d9OijNIriUUtVdSZnZsF0sZYld+r+7R1a9t4mYthxfWjcAc
fq0CrVfGZSlmciNJ7I5kWo4hmo84Xcs0v4f1BsrKD/dvy5VyRWKMg7x6hRXR76YH
da5UYgmDbt4HtVZ2JySTGH34ZfHPaWUqUubtXaZGtWCk4GP1Rws3sZVwoa9Brb+2
tEJelnkXfuEPZvmBJCQtclQOcrXavEfwwAuK6MMVf4E51gBNBZS/fUaDlN1NMSna
G3gZZmbAtLPycpVGNJ4DRi+WTEvl3q74sjCYQDYJVmVK3kQ9j7rl3n9uU+9JGBVx
Sep40X3tmPRP38jORtMyikUiQatvMnWWW9qFR6TPB7zKe0wuav4LA/ZAINb3Wnft
wDW1tnSt/3oy/fkHJT84vUTvOgsC0CMmxRCTcZAHGF4hi9ySjuePAn2mjpp1It6g
UJeHL7c+h1z6ez4ZkN4GlG631Ln/puaz8BOTXYmSAinlkxZfuYt2ldGc4w+BQgWA
lxGH/0UQF/7y8KCFEOIMEDznOpGYcDytcLV+DkFSE1XuqijPax4mA2tpv5Bz+93R
j1Geutz4O0/ou7Rm5SVKf04VWJ69RI+OK5wDRraZrFOrCqcGhH19FILPVrLSUAv+
/0ukrbK2icDC0M+k8BJX/pWqa8p4nFKRDHiOTxrOnTQXrxz8xzz9ff0C3qR6z8Y2
9vSnPpBKz+ISH/KvGS0yDz/iGTITEHY+N6jOHwtiWV4JeI7Ykt9/daL4ZDYYMbqL
bJsoHYUAuaXL1ReiQlA68y2TaTMZ5NzgCFIzR3cBd7cnjej2cYigT6g1E7l6OjfE
rAlSVo2P1AVgXRaHsmBgu+HQMTjVj63WWySQ8eSWGNi21N6YjER77/YZEL4Inrjc
74ne2taq0cjZWjR4y7YrJdTf1HTvWIQ6IDMByWgIDnYY4pQavPURxLujrwXIfsz8
IYP3/c+g345y0ERe7p2V2Xw73VaW3+vfwF1Fn0oBhL7aJtqm0U2s8B2vDNkRw4fw
2bQFpaJ9+hmV7yPbHBfTJZEcnUbSSL5wzdf/glc3IngxbUluR/8PPxXIlhbkd3Lf
KGdV+2HFCF4tbLY4ncUwApMbc1oORFj4mEgyNjWV/FeCBzNX0DKFYWju8zaP40gq
Q/PjWVI/RzNhDVgjpm4n3iydlBGcjg9+leQV9FYgYsvryYMTvH3uXfhoRD18EWHL
S7KPCBdWq6zYVg5HCTxlfJ+opG3mLta8Ll+Zq174XAjZ9g+eLZZB3rdDqELzwM8G
N7LCf3GE6rAHQwmdvzE0X6hF999p6GsmCD59WW7K28AbLQBoaRgNnndAuFgqp7EA
DyMMG1mOE9EeCQXsP5dbNbyO3RVucTepOO+Vdd9+WvqmWuhj6ZpNmL5p5lKoqEJW
DuE40GCEHMDxaN1mD5+P6flDBcbL89IgEsT2S5BsH9emVjcBcrQ9wrshtx5BFCzr
G+ci6O8B5vkB1PMUnrk4Q9hSH/uChkBxEhvY+C5gLK+oxavUXxHwkzpF3ELnjsTz
0qs+BJvrlXkK+/J4bERmjrEoNlt4B0fNOX8qBp8ZxTXrAb6Nb4yVTrYnQ1EmEq3X
pTssbOi8tdgwQ5n9y3BKTvZcsB9K2r1uvuOBRPgLiLPlWW/ibct7YvTMsoEDp7qt
XU0298aYpYcKaZOKW39WbC81lhrByS8dPpkMPaqi2LlbF9OA2ADb9bEvkK6BQvMB
W8xQit/6YzONVA8qNXXh4IoFXVCgDlfwa1+Lv7umGaNLgXLxXJ9Shq8Fr9REMJfQ
ENQ5HNXO1F4UeYYf3CWevFmfY1d5+3uL08RcN00l3My8Icmg08Z0K6j7McuYPDks
pme6W+K8dmmIZ894Ps9XGw78wrRMKgreVPUUVrj4fGVYCWy0GRmQ2gMCVUHmZGDv
IovsabcN9mw1TjyNdHrbCBLfbe7KLnCm+YtjAbjtkUUjhSoATIgvPNKRw8+V3QYN
//ygM0F93DNuvIXMnJuQ5o6FE9luVeysto+Oz76aDTRwxl7IHqauDp0fJhXNSEZz
Sg15jSez/COAa6rkGxZ8ivXlEw51zws41wA/LjdpQwHEJN6IsqOXWEvLWNyUsjEF
HDk7uSlEzixeLAyKYIsVxiC+Tx10rFVyAkewEblBVGJZw3UMbvX8pOXZ0ArUDqZc
K2QOP5MePdMzKQ3huMYezCtiBZhq+uXeaFP466/8GOp7CHaQwZR1o2Oe4Q1bEhtE
9GOkD76MV9Np6uidrZsUGzRCBHrOxhk+idsaQfxTQZNN9JzRVdsazI7RFaJdf4Nk
CKn1HkGpaxuFwgURzsaEpQExcTQ4z1oN3vliljYIGlQVcM0CTJ9wboxnqMv+r4jD
vwZL5oeuI8eab8YeT88xlg8U5NfIIxl0JoNQj5SIXYygLfNjKK/a3hRRyDWwPpFd
xWMLXxpVY8m/+XuEgCbliyjoaoQGdTbN9gHP4yhUE6KXUfdOVMNeilVnsi4zfl9Z
Mu+z7PKkRX4QhHPVg0ve2Yh2gBjtTtGFp8K/Wm5yQzN7s7p1+d2/oqZh/HMzfleW
5mhL4cE6h89zlQ08OT2Ifx94GxoSyKO0PgzZ4hNtAcSEYx99HSpwG9v8EDIDJnHa
AGvzEOERz7JudBugr9Hj17V755YVHZ8XoDlXavixs/vhqab92ApxrivpEhomBDeA
oeehaMji4//Ns+sUU4wixppy10ls/pQ/Selajw424J57jJ4gw1uM6WJz1OfI3tQw
OwII9YiiveU70kqYP9Wpmi77dObqsk5cXRRpCHq3wkGUgnQDf6dSajleqnzdh/rb
JrVH+8Oae0//94gqd4lSD2KO7w91zDXrTx9rqjb7/acFAMZlmgWCMtR8bXxFURX3
fyzsfbiDBsJR4lUGy2kfyAnWVcx3d+/E1fv8+deJiGIGjTp3ldZwUQHRS03LTjZm
++0WNagzyc/NYREeB51NrIixsBIOOxRA0/S9GlDMWHOY4HJp7Pgr5oVYFL8Ld3o5
gqUAxbOqglq8F9ajmMIu7DXQM4KPxntmqSo/Jhu9rJHvJ2lLDVeVJwV0wQt2kqep
fcWzK5Oj0ReabMQi3Wvt91zfpK+iILHNh+w276lXyxo+e9Fe5K1UDpbzWn7DttAQ
kPBIBFmR48sllMjEolKZn1JhtyGEpxCqQuPEndE1YcpTFy6cxaPJW9+CIYwYJ4xD
aN00xy0U80+U/h6KGb3aVjS7bWNJK4p8zRsep9IFhXFrDET+bad6TZ8mGf3B7TNB
0BmTuvSlGRIfgsFPAQtoBH3g3ipYDZqByCLbfoWMcu2JSzaVdbavSxGS4+tV2KwM
XagNt53zlgjQ9zahxLpFrNrtofsr+wXW0QkCet8yfg/2qH3twc8avSZ3gdDhsPuB
LOorfQAGld3+Dx0EuFF6pgenpnbNpy6+M9HuhNR8qT8CY/S+x6D40nM4q3TmOtx9
iZbWPCFNHa6kciJlmyucPfPwSmg9R2u3ZC+l1m5HfZMNirZ6wr/MbmgLf/hK7RS+
BOycaF9XcXlC4eVR060y4HSNKyikAJHPKfg/dBP7op5d8a/ArA59vxlEsKNcSFWI
85ehxcLqgUQgn7lXcZIcib5TWg4+MGNSOp8K2+Bq0VhojyXQS5bBY2L9b+uk7qWW
XGgS8jOvLt74wzMBHPlEpezSu1vEvczISIr0JXB/uJewR8PAQXH4927DE7trg3q5
w8VpvNP617LWSFd6QPXmsFVip8WGeKcDuQnlhVNOYBChqzKYWdoJna+H1bzHEkXx
FAeXx2MPAESCz/m3whm7RoBQiMY4Fmy71ykfr0dZewsrhNHKCiZSPBUKSI99kkkA
JMpTZXL5LSWLHC14/oc2PA51m1T+c7n/no4lhhDJa+Ga3DNg1kAnpw78dguN0jna
GWh1ybfVGLzc38EEekydIeFM6oP5jMUBtDYQ0WpGf3Ddu+KfJGsQpqFfMmGvwD+y
7G2jUSwLJosGiuWtFFkrDFa15OsdVWL8BmRqmUDL+jaM0eeY6FCAXsg7hQef3n+F
RjtQN/ReOV5rVG1dKEayj8f06CEnjKyG/gG/ton5zX3XCoZmmpPlDSURUAXLGwU8
FLSoM/XhKzv36cyglPNCky8Kd2Hxn1npbQcU+1nS92rZWN8xeAPs3FqtsLQMVkAC
6VBxB2E+Z+AHg5olOI5DH+Qw2ZMublQI9kK7T8B1Sp/7/8oxDBC7kIVRz6DukHGV
mJYO+TISMr/w1mynqxFFkXtIrZcqLZGLi+mIaboBnllHT9hl1hOnGuMSNt1uQdmh
Rh9d8ITmZePQICGPqsY5boUAwPxNqeD2Xd3ETvRlCZCxioV0wpTVqEp4kv0T+E4U
2UdVrFNGSdj/TAoHQLnIiA9PCpJXB2cnc08y0Heb+Dlc/IbROlaGtkpw9BDdjW4B
8nc7UUhauFluQNIOL+wjAkJzLukf4f4CqMUVi/QBbk+YzLzBfwlvh4e7GtVcp/9X
Jt5vivseCi9GmkvRxdbfLZ8xSQLRatAvBTmVTjU4eAR3hLT3T+1uY+LmRJlCKqzg
ubjzdTFUHJPdqc2lvYQGNX6JKwLe6m94UXuldq0kE2WO8pI6gZ+1TJy4gZr651kX
oA8V87FntwC6ap+v0YIPoq9AyizDuA4cRA/dTTxB382mND7qKc35dm4L1fA6jlTp
lLjl96yagRsobQy3EqTx7N71DO0YacfVSjHoOOq/Ms8bAOmyjgr9W9+9nKfG+hZD
PCPinah1kRfDjyolPYOZrtlvA9GXUib+13ZeMSFmSrwTrPZHxyyEWhE9atSQvZQJ
vgBtUV8fgixcfysv74opP6g60+NxRYN/enPXbPvto1QKSqHojjYWSGFMAq6xprGq
gZs8CmQXGDyxxGcIzIRvlPuSfg70rpJefZmlKDDwZ8VdhBk/ueJigzPhCJJSeGdb
gsDmKZvvXdOlxLLWmCFOJ5lu0+XEUxr4nIX/a6IgZOd197rEAVHrRtb1kcO4TM/p
4Ji6YFWdIcEnDqUVOFIP5MlC7UyxFioNf3lIO/bOgVQ7KpiC+eSDlOCmUChrNioe
3HHp6GzE6wWPwe9CrRoNk+tkEe2JIwa7FuIES3P9/v7CYwXxqDtH8VxMKCPsvrFU
n5z5ofz++k6fJfOXfeqaOCFLTWJrJxWpzhFlzTj38I2Nfwb5I0+QgMbfPuGtxtp8
7l0pBUEdAuB3689PbMkqbW77ep1/953/bfOTpcmH6N89E8YMHQD4Nl9Pj3wsEyjz
LeWO9rI+jADEoF2lBE00ek0jy8wxH4sG0T7kqovJHs+JO4HDZqY6u0kQTIGiHj3K
LurKxfC6TMtItAPOwq06ByJJ3+f7YFy8QAYoOBMsQXgeVIZ5sMiLVHnw0nAbJQHg
MFKUlk3Aiauk6jZQU2cI4IlFVo1y3I1LZaFPE4nI0sQ+yTnQnBD4/HGR+HRjYWPC
9QhJ863EkGzvNXiYln7pW1HUtko8n5h/Y4dwanN8ipe4ln8enN07Rkz+o25Jepcf
vIar1hX1owMMpVMHipr0GPKFDYWLrPf7q5pgzMaP6u/8MOPxkNkgMiY6LItuy87b
jy+vLbxn4Dcvi7qD/IEq+IN3RmG3Y7Niz9zoQzmJD+fc1ZrZZ8hsn5t9zVbJ3ooa
44z/yeKulQH/5bkyOGCdgJlbHol/JzMbH3C3sVvB8L4pQkhvD7x1DS1MSSp5TsLH
tcDZbU3SG022cs5jHrd5PPADMTAGROorSNsUf9C2b8rkgvmgGp52Sqsy21FJ27Eu
YUJuSO10Sbkor8rJrjiLzm+DuEi0anCZMBoSLRyy7n5++LKpO8AI+x73B+L/9VV8
qQ/joO3XS5+INEc+Z+XwZHlwCAqs56D5WTTb7yR/txRUPShS8IYB3kXwVQTxi6Oo
ZwELfZKtbPr9DDGgKC0H6sBjJrapXUr0KWvrnxLktTUJivpprQ04Q9NAXEuTYTy+
g9YtfIFCixeaHiJyO4Yu3Vi7J6nNis9mQIRkdlkMxUdDRchQ7xWiGMowdFuCCY94
bwWmJ7k+yqT9yhFXYj07EG9fA0Z/lTZOE46NTmuyjyGfYN9FpTjO3PMbr0+ZLVlU
Lmfh3GpFL10BHp9/ZbLNk1ccYZ2qLYPTZEq5qIZZ124iPTe5S2BlCCjksloBxwOG
95qjLeKW82e3F06uHSsuBZJ3XeCgZWBXFuz44MYSBawZVnGf5sDVtZX/7lOAWzpC
iRGjVKe30rlmAw+u0yDS7KbEOZYm+6Iz9+nha26PsCT4adXWZHCb1G36CrbqvfoY
ozPFMlBF6eUWresyYguks8tRvbvsgiqHMdLYAWMTq7UM9M3lEK8bPWuN9cNT1fws
I+N04r61ynr6qYqVEXxgXHnUOWvdoBJdlubM+c5299bykVvIdDoFSYr3GDUAgw47
yYYVVcbq8SVwOD/GF914BtoQ7kXuo+J7c1c18BfOxlJwqO2n/6mqsAT8jhw4UNi/
SAq4aQhMv/LKSXb0p/wQgeasiWzzl8be8ENI1NZZeWrbq5qrPaFSTQy9Up15Y/HM
TlRhWzutfP037+wIFBazK4pwYaiArCjpPaYJqQvWlDO+jTNyAKuJsLQej2oEaop3
duy4f5WLf4vY4VLxZXyURQ/JdeewH6eovDzhNnPiqz5Pp8Yc4BWJ7h4IhrFvHiSp
nJIH1G/ftR6W+DAWGQpYEiykm+vk+owrunHdKp/JAR6bjPjnbGalrw/h3tVMs5Z0
PgEHhQ3T6yZpnOoZeHsBSrJw5zyYE+O8+JzwY+C/oCO7RK5GaPQl6vqVvYbKSs0J
BhIgTKodY2yHHX/11wnRnteSa5Ki00ZSfKuTHMf8Ta/RxTZUNGpduNXUBPJtaEpn
+JVy9R7K1HmGrq3r6BmyD+VquykS/6beFaM3MgkPbQYt9l5fgoKvwWc5mdo/vw7X
NUA25PQrXROGmNXOxrzrVeOsWNbrrlI8tQ/uCwdBjgQLUx3GoS5gUD02DyTY5O+5
46olYAMi6Tx0dmPHDHU611qGSQKPh2frchqinnFURsMs18Bpj9ttATVKMTt2PbZM
jagtEe1ux7nhC5dEt9ffs/AiDK8CiHwDe0BcYfOQLV4xHSAjSbshZi1NybvtrbiJ
aK/Q5suoZNyD1Y6aKQSUnRnJcFS5QLIaOCEytbYETeF3WAk8B++ZOCNoWzsIdSA9
fGbIpfGWmxhr7RHH9pLqgaaBSxUPqBaoVLG/zRdoAJ4P4kagjlONneaMtD7y//TU
30O2NQPPLuhvL3NBurgwunjKxf4D+SjN2+wwFvUTfnybitq34s2lmaoEZcku8ya1
qoWwtQVk3p3+7OEoDKYxquwarOQRXZWEP34NdOweXtsHJaHwZGgLM45LXgzhANvh
D36pWjgv9LF6fPnRHxaT+TVY/iZCQdldAMXfO/DZkRzyR32lC/s5yODacZymQY6Z
2BE7p7IPS5YpSN6BK7EhCY8NX0yjDjhZWDYTJM9NEVrxxZIuZjNNP97d+ZEwEInW
h0kcph9MqBoE5xkSgmyjNiQXztRgwwZOa8OqmXsns5/N7XH9OeGV8mXlss1J+TB7
Szw6/b6VQr1zOb5edHcJSO9O7oQJ97s8BTpRbdXFd8a3IYxMKiAlTlbr7agfNvK1
VLElg2FJfnJ2trRaJN0q9tlOd/T9i5qhw1lhjAA3Vi3kbBN8Xaow2wg6jF38bRHQ
Hx1WaMrVFzG3Y2ffFUW8KrmIYBQ+CN94lT4jbD2iZcXowT8P158WrUjUwrK1Jltt
Hxlp6vLQUT4JUsWdCjhmgBVI/yd0VvfUF4v1/ohhAL9Z7+8WM3dqgstPkvr6bQip
J+T4//vvCz5ernfZ4V24qHEDr2kv9YCCK0fbYWOeEr2utphbHwWh2RVdqhhDdzio
LO7xX+xXKknAiwlXb0DOzDwXkUYu5yHiFPQ/7UYGw53oCZefPZOtJeKS+HiPsCnU
6ngU2fb76wpcL2anoJJQkFq9qTiC505CTfM8AIyCmfmwWny9EISfEsOwrY48tA0G
3ZGenhBdzMSDj60T5QmFkgSkqQH/NCuiGA5Hy5byxK6YfN6HlnUmpbqd1b9jZN5/
PlT3uHzW+Yb7EqYC+cNkIvIRll9hNlaKUZNHgEHWIaUpqgaKQd9Qk4UKKb5HkUaZ
Adi+uja01eEoQPi5cfqnlW6awXk1TB0t+4wwxI6PrKfYQAhWHPvJ5/EFo0e/liMB
TZLZ+ZOJ2rR0XzSu4RPh3DTPhMzi8Pe7mXLWVc9pfHGhGl+p15p95fKLrvXpbTPq
y2YdpRKN0nLBwnjarsbuedYKG26kV7nmb4sJ/BiwAuKyovIcBy7yffETapj/AME4
9HcpzCtSundkTD71GDV7C4dPkzuOQqLk1LWd8rOk8JdPrUtGPHnG+JQnmuYExDHl
c7e9Pt9GSgY1a58/0JEGOT6qdGMpTYDgjjt1FUKB4frcr/Ydxiy5QZ/qkX55LSG8
WunHlJY5GqiQX957kEVuAx2XRPGkckPcsmDpC9wD27fZtALApK/iMfylFPv7YWhY
KGc04IdWq8zK0DYIlXx3anR8SxSmV33WGbtjtBMyELs9i0h2nohLOaaCdmcNd00a
WF+YILu9CtF4GUsMf+r3J0RlRhhwWU6oei13u+/Pgq66ZaFZI8pF4ZqOQj4JRogE
nRhGoTH62cCqiz1S/WgaetMg20ZmgzJP+jPFi71QIvwNvsuw+vSk9GtXLr7Tck6O
/AkRH84pj15aUfxzIIQWQKNHPY/pvCnB6O2Rfk5BlyehXe/NTboW9VGs/ZIGRAGV
pBcypaFqDYd9lwCqggLF93ImrDvHsjUaUGDeIJ9NoVVkoTDNvFE83GsAKfm2BAxB
MLxK2cnhgJogDai7HVG2VnbTR/PvtaVIL2fkzBQyLHmfLEQaYmhg5SsZuGECuzaK
PadNMGFWW8poctjm4Zz0YO05cU82m+4FayMChhG6akAQEfyTYnHfDulNgYIwlp6p
OBse4EG49B83iKWEqgv3eEX3JoJR317McEsbHUOUwzZxD9ZEUg4mxrsWMeXfAA/M
ayMdR0h2DTHtQPvFL1F8QboRC5NNz4htHaH5hqdTPmG+Cwcgl2exSNlIdSWY16e2
PIv0SflMg1p61Ipp3cJ8wF0GK+qpoUkugMtGmJJUjDo/yZZkT4ld3GmCcvM0PHQr
LyOIPx5bzYTMmdq2yzqsQwcXNkUjTurC7RSLO9kPVows6e+0IA+ewVlzso+9O7cD
ipRaqAXkPR0iQJuMdj9VoBoR1t3au4P/YqlLpHCIZ2pzBLPrvSkRzb4zEBzOE2Cs
VQh88D0Wk2bOw/0KQI/4LvEcMYI0MB4Gc8tSGXIAyM7HXAwnO1E/g6glSH7klb+g
PWqXO/zUNZtUCdeBqBC/hUENv22PyEnY71rg3RzahG+FnxuY6rgvJ9mCbQMYBax3
20MTlpRJii7azphhF+nVioPhlr34RX6jEhoiMZQowPIBC0DHoQK31PANVNhxnTMZ
bypCfkw3aVqjn7j75xbJFq+FsWEH61goIHqs6hZkzi6QT+ZL9r0ZakCSUJ/U3emh
nWBitutoH84GPVpmQQg1cxjp2XyqLw+VJjtONBjq2nVp+U/npsywhiYG9D51DQLP
zitW59su5N5wcIYE1j7+NixdwQ1+i2pYjaYztEYSX1tVtowscyRPOo+T3wu6crzU
Dg/K2G3LsCZY4soTfsAVXHfFEHuT3dgEoOwqfpk9zjQKyfhFLU5OLNE/oNYTFKpz
CbbhAxzB3fE4RQzeKzKSNvdZoP5CiF4rEu8+IHUJEonDmNQT07KcRhnbprXRwu1H
ykbMlWqRgTN6fzB2Ttq9I9ppmg9VnnpE8tyPiLJgJSkLZ6ZsJNqMTYSSYZ/TXQHH
11Cy+MUrtqoiWzTAHck635kGoIdGAffF8xKl+5dJZZqE2OeHCLpzpQthLpY817xI
8417RfjugxmB0MNulJnYrsmkOVgizoZdA5Ud8PjPf7OxUyvl/cGeUY5UBsa9qcbu
m65TpkKAr1jM1xG3roZgaMpF292IL9KYqzcyAyzavNmEYi+qy9BVKR8H0i6MzbrA
cc0owk67qbTHzmQDCL2IzJGuR5rgMqLgP5k6nJDqD9m7zUphF6FbwID8y8t1Cr1t
bwtqQaNgUP1hx4oWcbNzb2j0evVQIFrHtX2Vtnn/ni5HU12uH4Pf6cpT/eu0CwRs
Az2dB3JYJKWQeaya6QfgBuU1gsC3StJfxGB5b8vl1n9QqU2qlZHjm1LKR9/DW6LD
zL2C+/yViP2nc6g5pc00ZmKioegl9Oi9fSSozhu7NEhDK0e+1kAleDT2H7xpTe2S
sWl0AOq4kcOFNQRODDLZwxIWTGzl5la8dcbAMkgJPdyk0kFwgMO1mFmPZdQ9C20d
yuy0wpikmbWSc3U0Z+gbYM3jSPmyc9U7EGnR1RKT4GIfWX2+IGG3tkgv+7CScJ7Y
96vyVbJ6EfwGYJRWrw6hF7gFnIA70hasafz1pUgKnsSfP1MjwAYgcUBWpVbeXo7Q
UdgHyBdo0rxuGgWVdC8de6pBdRBw6yOHtFfHwPgMbp6zIvgRHfE6gkmGl9llAYLa
3vNxTb2iYDedKl9zF7r0MKIiPEHfdP0fT1Axwy2jHygdR4xWhEoI7IObcnO5U9SO
+6A7hHmqLbjauv3w49l+Gm4q8mVVgSDkaxW5teRj5mMvzm8O++RxEFFrBneurLmO
lQJIGZq9jIwNMpcr1OE158cukMb/Om6EYOG/wubj0YKAifr5RWEOFxYN67tbiMv8
Fbc5Rj2zsjHwS/cBvD6KQ3FeSxGhx25CH5AI7ZowNZ0k1+HjoJbKLdCZuY89NfMZ
xHKFjN4Yn7w+pEnpVjS7UtEsJmVh1McaXSEvzISZZB/TlYEcSjYGqYIm2m5q1Dk+
7X8um01OySiiOqCU7h0en+aDWQ4cqvwAJbZFj7jfbFM3rdJr6Ut+XSpv5fX6W+KW
Lq/zJB2iBbKrwffQKGlgT1apGEd3NM5XcjNKX4UNd9DQYWhDqfxgma47NPr2c9Vh
WbXSYn3m2PVnBdBbHDQpxN5CsKHJIgWJ1bApGX2VUHjejZvhFXNzzmgx0VHe5AXv
1mpVqh6ZI1P00416vN/FCD4zRMD3DqV/NazBCPlcYvR9B55ahX9XBhWE1u5GKFf2
ZFKi3e9KXVHk7EJppiwqh6zmcCLMQwYc33bcoY6a6LDf1r1fEmO2WfcPPzK5wQZV
Oy6Go/GbmiV4uBPrkk0NvbK1O2lkOdVwsDIWL/ecXfz0vfMB8pAfRC90s5g1iinD
kPIhwWbSignW9ouYP3GWcqmlUDwg/n/sUp6xf/ZovD547/OghcjWYwQCqwajVOEm
o04x1xAXr9cPbZgZQLzQ2jFOTwkmkRBkcMlJV2SddgVYpeiW/QjCDFEzNMKtQ/Hl
TUEyUt/Nd1A+wwR6b7aBeqBoPvR749nFwe6AdWMtA2wM/XZNThki5RCDSFx2K9gm
f4dq/YSW24aPC2lGi1N24UybqN+hqAid9hxym2/q3Ea2yCNfmcQELvEPe3hsaxn2
8uxKfbByoWm/hOXU27AG8hzMRZ27zfIUntNyEvvZBTLPtDGL5rvdet75E+o040GJ
9PYo3zFqfJ+X9Q9ejTUXNSTpceWe7Nnzs83LDEHdSSxLusSELPxRtyM268hm6ZaX
CfgaSyapniCNOOA6XS3iUkE4SFSx+C53oYhKdjtIcFpm4i8g70SDE+f3vccJUW67
jpUPxDw/peEJ8UHYbymm76wZuXL6NqyKxSF3fYunoiPI3b3Uy1C8iyFdzdD2ZbFt
s8ENBQg9GK2sX9BJgCphD3htxf5aBptW1O6e2HmMAxLaY24A4tDZ4SwkHaFo5lWD
IOD8xYsQnHv7zZ5p63s/GO8EzonjiY32xnXEbVxThL3b0DsuccD4PBXsDLWf5wll
VUjl8nkHnKoxK+eM918wcrVwfQJd53P3hLiwUj+iHedn7zA5+lMeUNbCkKxA496q
WgFs0D5qKvaILAFF4iracAn80e89g7ACWpsk4C1FQB26UpitoMqRSJcD3iDNpBJ2
O/F+lmI6WvQdPWpAChHgcit/AwEsBBAx1k5ganwMfEY17vM4GKpshFR4Db9RlxoZ
GDGaXoq3bPVfw5tIOHpzigfZJQXUhljezUod56++zKMK1nEKfdZPD0/6K39aT1le
E8507OKXZ/JxmH84/2sENBxVFPG6xEZO7GB8OVdxaDQSdC0c40rqtBMiJ/w3xkx3
OaKpnYiyKFd3HNdYEOP1F3Y1N5ALdFMIBtsHDeDy5jLFwAGSbDks8entT1bMpalF
VW8bstb1sAC1BZOmcMxczDh9lkJiX/h/Bu9w33hMVaCiuhN4dE74brT1cuvf0uh7
orguOLpPGCInfjbN+l+EMCsPQFaE9uryIvecnRuYTzV4hEHA0OhvKV7DxEYkMsck
I99sydy2lY5O2s4wAZnPZTLeDvQPgNtjocuiANdbR1DWHyMo8BTjp1MXb3RlmSx/
okugrvZrOQWiJ4js9a4LvuFKVtlKwCk6sKO+6crHk08XRd4/QOjzLkotZuFsXWfS
mTaU4TEG1xyKl9f9h38WSbachuE50sHXdd33oK5opIIVvkx7yT2UXmjf/FwNW5x/
nXNiabSjxo43qHFIFTsZ+oRZHQit0141hOAagQt2AifvujVzg4eJ/fNkEOZCnLku
OWaMQ9DDS07KIgsSXdCbELq6mAAkM7NQ6lf+l/6z+CZJuvoROoZNRMmlo12CyceF
Ir2m0loo37qFpgaF/0I4XzHVKPSV0rrxtnMmAKfq4Vc/IdqWGtpSSARtblnP1YJm
Di6mogYE6mwBleMUq/ImO22oqpb157mz7UvPypH8/PXkGpVgFr1+hdx7HnJfdeR2
UUolbW0MDJEclGFaLWWrIkTFlFvEmxHm5Jg3QvmlzlzE/EPH/HEaRfHsjeBK4Rle
6lYAuPqy0G/ehRDP3XMKSQii/UyuVqBZRLZn5VhLTU7AP/IrHN+oYW3Ob+AjrYYN
Vu5SEQVIfKQUv+84JiqD0PCo64XoyOAc4s5EMwWoL7uuPUQbsBoZZDjLZwD32pcK
o0bVczcY+bWwn4kZWN0OlZMR+UyhtFl+CqyFyMUptYZbFOiZDSGCexpCsvE5x9lb
KD+eIWwpVGFNXt8IIyBJq+3m8TyyiN0CSRtinnlhMoa5xuq50z7yrC513ivXetJL
Cjf3ckvGjW1MvYYUOCwVj2C+mVBr2zpj/2PuMXcVT7rXgMLNs1lssLymsEEtnGk3
9ElZ/pjHZl/+jzMQ9YHUK2QNVEqPpgUYydclzAMLH+ckAlbfLLBrv8zblpGsMGZg
BEmA9uhgeCyIZz1mW5G/PgHWpjziOw+p8KwZZ3W3f9Pu9cFI9maRpPOySkcE6gYG
vzayhuEloOhDBYVIDHrLJ388jBY5JnL/nIgVkyjX9eWyLMTsb+y1prG8jFnuoyGH
uJWaFIMWAq9bCGgUQckGN0EyY5cx2MSbXLHJIJk1pjKPhv/sE72T9TJAetpRhwOj
oCLyI6YK690lx22bKkvqnw4ofW82IhgAdwj3Z3NvuH7Goze+BKW/ftVEV4KXxL/Z
wJMFWfsSHz7+jTYAPBOZxGdWe6YDK1QDeC3zHWUh6oJAL64jpIROj7pHFZuankNe
io+pn57SuD0r9FwXVAHXT/EkGfkbDJzvjLfYtlk0j6wHdYFncEXLw6oHqjWgfc2y
kcvmu16xKVJI1SUwgluD0OFV1ufJYTLsK4FemsLldZ2EuADpq1uF6Q6EydEj/LMK
JDEX8JkLmkxo8xK8YMBU5JvpgbuwcZgtxyuqMvr9+TgYwY5rjiU3Gv2u4kJTuriw
xnA3rOrynngTeAt1jbzTYWmY/AYk0HY78Lp8Vc3qI/XMudc8b5UXcLdkngnShkwg
1lTBoXnK4nr8uf2ga14hv+6y+vp3Pi/PsU50VeXsDHzqRwmHlC+7AxqFFQSslJNK
SJ4D/D7CuDmMbNa2WoMFGx2by1dlrT+g6K3il8Jn3exxUuVwjdRYiOCo2EyYdBuM
CH5MOkvcrf0tfjd9V/mhfz7sKx1heqB3XhJpyT0Y8z47wmtFmnAEK8CSenqn/Jf1
KWDg7ByiijigYFnqAz4gxcR/4yPrhj7CqXvsBYuUs64ilRtXU5phcnvHVfom+yg2
rstydwaXmQVqTWraSzglu26nMUNW3omgpXrzTGJx7TiH9MbwX/oqZNmsEqDktlU+
NHWk4ARg/BOWCcfMHRgg0iLpwBWQ5udwtboW1X0dmcQNR9cVycULZedA8CKvIdf4
lAF452EENWMh73uNkn2zyH45vpH4R53ctvjIGoDpfFAszDHQyCZtr7Z5lqiZB0cd
wBFFgLZ3CltfUjWW7ApuWD6eCABXO9uYo/ATiHMuyM5LLOCxz/2paIO/3XP+c139
jF8Q6Ix8HdwHKqPfGjfjomLFmaxdano9BOiImrbR5oOAf1PP6tQuAPHv++maZmHl
OJXCCifgsQI+vjC2ccvsrI3OORJeev5GWM2feBbBAg8EWp9+hoPqyTYkgClarqDO
jpzGb2sbqVYuCCwSqOiByW8LBxO3LFL/bUOV4XCZ8nwTXOMo/8pm24PUs7bwFxj2
c8MbCIoWaMTOzzKxQkUdEOiYjerYBpHoGnxc6/bJStEihYiArHyjK4Lthti4hpMs
jO1xt7WLFpowS1HPbKLqKVNoOka9nF/NB+IhwnkBG9m1H8B86AsW2f7zObvOkEDx
EdyXkX02UMXL4VWLz7TN07DhV/dqjingUraZVJjfzJIVI44/JCKIAYx5onrOrPCi
05gWdeT1sJS2E977LiClmEluJgtkPNyjJCzPGVfQJ6A7hD6WdT6oRwKFMdmbiCgW
Tma/leUowXILUB7SyMqc29KToLQnVMQ0HanU4tAryIxi5eKLOlRISya4vD6z1cBY
OFQS/e4hRgvDaI9ox/IwGOH4JepJ7A8gXuyG0/vJp/lzE6zakGhrVJuUn0Ks9HJx
RMPIbbMAgYCHUrg9uivPrxYSIUkmWtiwENuldqRMNfr2CiProycJVuCaNHdq4fU+
SaftvVaw2CvuiAAYyG/F7DL/twDn78FZnvqh1UYtgMK+Kq3pNhSprJVK02L6Hpcp
ehy4V7H9WQxWqMLkRjilGJrRdsxOkiKSUDMbNM1Y117/5UtrcvUmB6rpFR+XouYo
kzHsO2zwHv3pl3zg8eAKmslqvPN9Bpo53hT8wEwwu/ANccOzFCLAjECd/5EbUkmI
srSFPyw+cIatJzG8TtePtycFzgRvVlaA5LYXvP/gPjkYhhXBstJ9iPCR0oF3lPWG
AzS7o8CNldCpFSboh1/Iv8N22IossBZJeDkOIB7v9RzoLIPUz3rQ/7cBMV21ynZH
QkT5291prVL//TvUF2Vt3st3M5b1RwS0E6m0BO/xmSjjq198FCxZarkJ0XrJKnc8
ozgp/bEj8mUOD1RK1/EIT+wit5YfPuUiPFACLvKsT8hnOeB7SEuHzYaCPnsCcLxH
asXq+TEHTsLSuyfiL7M3GHPFKjEVGWWQudhu5OJ2ulU2rQPejSnjT4EVxATI7wCV
LXzuZZB2uIypFl1Sus6AmQ0WS50crFueay7Jcd3erxw0qIbg3sqvGxl1XV13G3gy
rUgWEiX66gOGwYgxh2LyRDBObjiw1Dn+yr3swghxWKI+kuyi/D4J24V5LxacpBgt
MUw/FwnnLgHnVghsMP+BzXcZGIFgjVQGTwZDB4bu1wkK6ZXyp3EGNIMDHaw3oPxW
AP1grpW5bn2t6Tur0P2YEOEvQHMb1AX1K2SfGSb//IjQnCQY6auKomXCpFxM24sS
N7XkainerXF6fCx2xW2kZC41HxLrSpZ2IOkEF0PplASgEq6wjeSmM2n7CcVjBLfO
ih3k0Cx5o7S9CTGkGjT6TERbSSx596DfuTyPRIb3SMt9MDTVNGSvHvEy46mWa3Zv
ybjSRGFC9cLCsUOasjVvcpw5jTxsLwRKQYCkUKmPfxa1hQLQflPrvlvoRvWXSB+v
wXNvxr4lahTo3bSrz+tz7Ujt05weO40Uvf1N/lL3m24KLOM6FF61eEVAloci/NLj
zIFjOfO+XBRCyAmVc/WgxFF7GHOQavzieqgz3y4B/4eaQ7ty5m9e32zMnU3ve1jd
oUj/jP2sj1EkmZ3WU4CwroRtjQtRJ53ZsJdjlfiESNSD+cS2r50P5ZTR32aMPsDM
Y5X8ExUajAwrCMVsYEoDcrTfftbBY4lGcRLdDAW/ghsrM/WGGclZUIW46AU2Z1Pa
yroVxgUWbF6C6esniaWIws0NjvcGbVu1S4UbsI1V9vfk6Ep8bolkOCj7v9b7aock
fwyg6MGE4H/TiRc2UysJr/7P9yiRj8Dekcx5YUjz7J8gh+pw5VoXbPkEtNLCbK3I
NYrQPj7JDH6Bvhx/nG55euamYojtKaL3SOuAM94ljSpOZUJghQET2xD9XQVBvFtm
d0Azkc2w5r21i4kmOOnm/LyPSF5n5l/I2iIN49azrN3gpJCCiKobAiCh8EgdZ9zu
habPhys4ZpOJE/6Y/tw50zjgJvgFN7T+9FXbzKjm6PNZnj2myWnHREIbikg4JJMi
BE89s6jhJKTgTNHd5ilb9kJiCu2qVONSuKXRVsQnNSTMuetNPdAd6lTKtJxowTD5
I01O0v/qR2Oe6yK/x+3Pu7jiXQa6YYMpB7HDCXVsBHxYYYNo0teQ6BLtQkasn4o+
lWVyahrF+4Iq87da0wDTzyzDraWm0LZDjDD9pv3P8MZ6Cr3ETnNPeqW8Cyic4uBN
1fZ24MIX/YasX5sfHdfr3g+VKkfsClOCpt/HIqZayxHhGgZKnzOIMXJXewKiK6Jy
fRRnpdHq3ccgc1japetSKGfFWjTUM43WO8oeB28F3IrqU2UQCBSxRVXV9jSbkIMP
lSByu7ypeEWprlyB4bldECSCK4ApQOgU6NP92SGg8DS7bDJHGV2aEJ9XvRfe7RWB
lZ+IOyiU5cGiWJEC21afV4VuiaVIsE/QqaXxhCyZcCVo4kkQUSIWMBtfDtQNk2nF
4o6aAt//Wk2wKmlZCBbEKoBPW4Rh6zEDHNZEIxLpLaNK2gmsgf9EnWoP3yshNGs8
ttbPuKNDh1rqFE1g1I7xJj6gQbmTWLNylPPwEJP0A2tEQWl+fCMLSwiu6ROXVc8N
1Gq0j1yZfByhnAOjepEtJT+xWQqrCBmQ/7lAtOZRTIHXP6jQp9MsSeAt4w/6liSL
be10p1HGKD6b/bnbOKK+sYoth3+jZAngcKCn9bfUAScVPiXmxV/AhEgeTCTq2Ix3
zO2rEgrJ6ARt3MMRbB+J5t+dRjY0dULldota9nh27NF87/FY+OX1stvAGWuq5L6A
09wgJuONomg4Z9QjgLif5oa762WwV6N+U1M2QzBcz+rBmEm0b864c9CYr53JGhMH
f5kWNTkQ31q/+ga0vCoX4JQqlMBO8rdj5MYj0p8QB3t0ylMZGskw+zPSCldn9RWK
bM2QF1uy8D6hB880113boZB6m2UfaknzX7/oyRJk+ygYtGOefAkSEcgynziU99kS
m0t9IGOX2GcRCnbhkEZVmUGmZg2C+GZP1mwTWx4P1ozmi6/jpJDSKb9YH07D5wyt
DH4e2spRc+AUFYuakiGIdO8V43ptuHmY8XjFmgxigG/ZbRxSe5COPy8zoEZGalx+
P7ug8LhQGX788cAs69gTYCzCFpBqc/sgO6isr9n3118DBss1mrBiDiHEnzMgXwIH
ILhl1L9Mr88QS3mW//7hnr5Q1RkFtydtl6y7FGtQ+xoDdFEIo0axcbGjAWzAqX3f
HTo7yZOycZ0ZB2ijgCke1LrkyT1qhg856GtJX19retykfY5FTiqHTcaNEJHBBF5T
OgQUzyowzORM4xI6a6OorXKmLIGHC65zwh3fCig4+CVcsxyQnk9MZwDy8644w77D
WBI1liUSQ+22vR4zisvNVaEzhwryEsh3aOTZtedVbblUEYCDob7SMAzNNAsiQLCM
tThnxgYmlhyaGIBzvUylZ1f4nMxnQAm+e2gwaDM1d9ssU/ZEYw4MIOL9uhNinEKz
UFeLuyKVw9TZIndmByWy1t9/860fiZb1aQHY8eRh2dF2FChtKqR7/LwKKbEsRuq6
IIfo3Hy6ZYbyXWQYV7RIF8U4vn7hhNW9vhc7GFb78xQX7bqJ6GmBDTI4P1dVA1EO
nKdIdR6ymgQr+cuik+Zm6laqtG4wW8EVlQuRQy9/GUA6JV6xMHmvTuGcfkaFsstb
SPIr716oJJwOtl/CTXVWBq3ivpJLoWOUODE7jhsfV+UMH9zfsAa76nk772pGBXHq
zQI4zvj0v7bz6zs11d8o2dc8cpKlgrbTfDZAyXqxXqISvZsTxWqTu6CiEIjQthu6
AXHMvvWWBPGWDblH+5u0QrX+9ef+/IFt+unTCAr7rH1/2M7hagTlaEi8CWmeAgt+
CanQShcYnBypU6cCnm9fSIM+7eDPTLh1mFyweaDb9tGxhdsusygr4WIUQJ5Nisow
sJXy3XKcQctklKWX4emxf0q/nHpxF78Bmp7UiAjDVfptSGnuXtkmn5KBM5trpFaF
V73zGIXT5XdNA07YJ35OQBTdwqqwiI0Q5GgQurWWq0sX2eZAfpCrIjvxTLG37EYI
+KgEdjy+NsBFtNInSWtdITMBjDeL5Lasfq6npSI3mks+4TRO7Ivd1uph1oISpjr0
V7trMSnBfjMHZMYNzbWq88i/YORGMi12hn6rFur1sg8gj+loBdFTMgVn5Xq4GN8Q
o7uSJWUd9DawLyo8UkACzbXPA7wXB5uMDrNKkMKVPUtGHw/SwQ1YPza6Jrc2mQ4D
BeHweC3/aneNFHKIM8gzcEBz5wo3sS+eXpnoeKNwG7DTZDORvt6k6irr8fyYZfrN
hcY3xWN/LxqXOd1N9JkDSZ6uvqnlFaqimc2czQuCqv5tRBW8yTN5wcJUaRnKl1nK
gYSDPEfiHnfBmdwBsqVZunYOa+2cw5sdPCVO8e/CbPz9JlIpHEplcLCvY9mXqBaZ
lqDsmfMyxLdcW0mQWXWJdw/EhutXj0Yig1OtRjZb6wFMoa5voo5ecnWvayn92h95
oinwzKM+QHShYd9S7VedGGGW/QredJ6BOB0A4EftE9TmUCSN9oWmUIUjawK4bMMT
AQQxjrH3dpM7Iymw9eu2kpCeNvH359FvDDWIvJKkd9c37+zzqD9tTak3GS8CQIxB
oQMxI+z4j+a0vHsKtKDY4K5lSmN/fr+ep81gkZeLZZiW/httB1RtZAojhsMc1B8n
6g88SrOQaN+pDFVzukGSf05HDXAddvYnBJDlYut//hSDF7rCns+BKjtnnrJmymru
PL0gIX8OONaCqynMBWqs9MFJh+JCQifS9Lap6ABRehuhnjy7i1d/dJoUpMbGSYEt
EQx8A95zAyhgAb4R/L5vkDHVM/0AVVHFqSNhz1xaemTA4Bzras9oJcsxmSmzXlNk
iEJfCWL7kAGvZMFcb8+noMbQ8W1s/YPt7u7mOvtboSmAZsw7zMiWX31FHoAuTZcm
U3RmFTgtlG/3ZDX650KyStj4+xkO0BHKRvtnnkKnGjsXXae7YULfJg43RxvZ+8qU
HYwOGn8SC6/CoYa4X4gIpgATQm9MccDKoPkt7/iPfSeDjrOkZhFFaGUVkqNw2UZF
d7D8iQHwcZkJH+CZtbDsLEn+/JKTVk7Dn4ozcC9RvNbOx4gWbvlwVxhtjHOZ2DJc
XpQDMOvlVUPPE1JfBSt0xOzA/5M97EmuMoKOLclwJHC9pPLS6LQGuQYOoZEb49qo
Mi4iM2/vX4zEeXxtAgQZfOnmwBgF9Pj+ZFRbPDTAY0DpdtQ08pGtIMCq2nr5s9ns
04bAOqVolfCo7+lNBaY/F/8pkbYtNyAxaGpw/fa3nflW04jYh+whC6Fjjz+8RuvC
pIkY8dIsVXai44u3+6jkOzRWqKCkzqRzHoZF3Ly0n31x1UJKAZyHAsVv4G0cSj/s
twhO3o2+9yDwm8+VRahUlkJ8zdGiHohbw0YOJcu9s9UuK39JBKZYT3llfi4OwsWS
BEO9ojBXGBClxdmbtR8a51cIg5qp5HX/Vg66KPiqgUp+o+GBdJGgcwpVSV+WCU8Z
oQyWmeuWVtm/OzeR14c+2HkkAC6JzGBpO3Kus4miD3+AxoKP/HdGNoCTVf4elWrb
o1KfH9T3+iaQhvwkFxT9I7UnZc1EBi8j0EVAEO3hZPy8z1uE/qr+LKQYyKUKoII5
VsQYAgvBY3QoltzMplYFxWwyju6CVynrQ+26Ey9hpdHO+mKIGLA/RwiCNM+8lJBs
Dd6cgXHpm6EdHox8pobxMKwh2ZFBJUQZg+rjBzlPf89cDwQ8ro4hfO64dBBTac2D
DwyEPOBCbk5Bwz5GA/DqS5QvzXYINOiHGmAhtUpkvtHY+U4a+8P8U+bM0XBHPs4p
yyMbLDSN5vJqeNQGgvchZ/cBiOiNIFACS0Le2rSYPrdNQiW3sVCm/G4+Mqp3QcSA
vlkfcmVWh1gLRIOGoKbqZAon7jUa1I71Wm62kIabu0Eb5ZyzbvrsvZBVh9chvHk3
uuE8obib7ADajw4wCXWasi+kyp2wtY7D3QqUgdYa32/dnkO/MLyshlO0Dr48G9G8
Hj3cmEw+W97GRbho/mcCTUD30TcJ1bYLhFiyxYH+nlO4tVZurF9O6ZUA4sRdJqpw
NnD8TLGMM8fZKEZ7nfHf8L2E06bDBQ/mZ13amG8QexYcssFxBDBg/yRmiWpJ1eB4
AZ8jXTmzo1RoL9Mar7BzPkEY70rnL1iGxhhp4GnJohp+GCoPi+COISvnQizEge62
5Y5ebtfh0XbmRPMU1H+POkMwTYBIDb35p0RIzBBts9qLuaXGna7v7cdscu0n0Dvh
K8EdrGeiIKlmpbRJsEb+rQKUj2cnA/+fJZfXR8Py3L9T7Cdf6V7PbrW5fNf1sH5r
4/mPKV7WZmdFjQYaNow/josD6Xk8nCC8vGXTBj5BpbLRvIID4Ud8jHzbySOrvMDd
Kz2z6tMbdzWga4NEOLsqKpf2joLMKR1zEdheByL+mJf38sDXqs1U5M/jb9iu0uwG
qBTrOgoJEyKqSZMefnkU2SnFanLE4musuzGMEoAqbWgAyb/2vDl030770g8SdOte
vDR0PWhG3s4RQRObgKEhgwGAoIIu1xO3pFHvF3+IksSNjJjXKaB2KrPiI0kuVktq
M0OWyXh9EsIfHICEmeUZ8KQOBpzH5n11YRB7MDU9MxGPlCKx35vwqTnreHxZfdCg
ueIQa6njQ6JftdhKScOivaEoP5UW27gY47s2vKLj/dD88lZ2oo947Uc/R7Vt4ir6
EdRuppPDX4DzrAnHMkj+X9VPG6u0DO/clnEuFIZLaWN0QRh3bCR7db/GJHfwG0cm
A8rCPjHIhxSIZWjiDECpkf6QO43sQFAVpWQm26J56V5ytUsPrOBrXooQ86Crk7XK
SuveRLoMAeiFfX/rnEekxhVwmV12EzuiSx+K5dqeSFhWu9aM/v+4jFkiL1/5q/xD
ZegLdkW6J7LkWalhJrgC7QvJIKHKWykBPe3WtBNcGwWRGNf1RZFyifYD/YVt6KEo
OZPwtUnaiezUsP1uuyjrlqJxTfwmk/kXcZJzsuorZElYEs27kuS9GDMDPAI3vTZj
bCA3gXdgzeKqP/ixdjzKzq/WiyUE3kiHeSev6+863eh9I3Z9Bcd32FgduAo2KkZw
KMdlV4zyKHA/G3FYY1mGyPVdAHWj+d5eJcJ14ZwxiCTPuSjxlDR61OYkgRtPkERW
Nfvm1ApDqltmUcl4gabo2SdrcBMt95y5WcHtANkfzlXJuBzL5nm8EdBUvcBLtb8Y
6wCV7GijZHKZkRqBgB5If0c5BuZehDFj/rRLE8ywJxtVXSQYffBsR+ivcY0F94o8
oQ2ZQUiQxsWYUrLcAK576mpA13GKDVwlJtCGgD38S2bBtMbWJYxk3KRQhFsmbwXC
gwHBJ8fh0fPTIg/C3pPpN8k2AToUs17OJJYCPJ2nxKiZNIFKGcgc7kjyFfGwIsvT
0R2HdqKr9mrskEFAJshnGEqeFfL+whdLgRxn+q5xL+dLomP9hEx61dCIaWpNdnTQ
cAO3mt47pJCiEVOdylj7/+oMnmiL4ZiM8lvcr5Ih4DjFi2uDzSx/sqVq56yodzav
W/oIQC2ikeB4Hvz7NIyZxaacGvy3Erc3THx1fMZmJLZyYM4UiUcKp5A3v/WcERBR
+GHJgfN+nCFJ61osoNW+xDORseqSezB0cGkf9xjTvoCr0BIdgeEEidwAAntxPNZ7
6jJRAwUmrkImsaWq33EiHMb3U/poH7J1nMsLy0b2PoRjTKmes4BOjWX1goSGJoPn
tHpDDCVYkDfbPL9mK4Id3PE/TGTmFrq/o2BNHC83VXDFLSG+LYJNirdl4qHYUqcT
/NczyBnUhkITYHOkWbsLYlpG1rCiYLnztDygD67V9Kw3PwLh6g2/TgpGj9fNrJK3
7wAiGCIWEeJKhnKFfDBdcPOAj+gDW0HMaUIaFVunNXjLWmG+f+Kc+Jd9Kfazn0oZ
r79YgC3eI4AdR0XEOGZEfF9e44PYZQTBTsgtqDKWotisedFVca/1kxmYVFtjxcNQ
4VFVPdXJijCmgcD0N5krqmapvZPxHU8M0+pmyeoZJpVcHKk/Y4xHxG5cRFGCEQ/1
Gp9iVIgXUYMQnn9pc1fVgPRx5ZxDyZwi68oKDinn3FULTg3y7fJGkfuzRcSlm5kM
1Auru+abaPo5616l/5q84wGkb0jUa5yTSwXbvY7Ik8VXKvDHzO3fjR7zrNCi+K7F
iARp2nynUreDrVPJNlc/tOSb0Z5KEE7EjiZcEGyY3h7B0n5yZ0Tu+e7v+vRqaVwI
DsdtspzQtFJuTbQb9A9Mt1K2xUU4kCYtkI5VH6sZiwLSPVY2hMOX+IdCyJIYz7gc
RjRzvxjiT5S1doUkJhte2+lTAKftbXpLUO6wt++k5OyDVjk3am5h5meVeqLHO07h
pUSJYYpBVYK6qUkLcfjX+rXtHJ9wFBTtEJZgK7m75SyIKYNlVSe+3aKs0Ndab6pb
qJzkfONx9UITl9RNCkQlWtIlflFoO4gkTzGh4wGsQ6mXyvu15JSZnAvUFb7EL7oV
cOHTAB/xa/J/1HxoI3NUt0reAHF/2xfxaTzYIaWtwqIYJD7z33M5XZsoA4hEX8KL
X9nWu9OUwTeTkOTJylSiIV/dbHgb8enm/XrDm7LsMf7BBwnJdeudIr2R9Hbvx6P9
+0KdL7PmcvEVPi1km1TxmzQf6uhEHG9RVBkZL/QkMxayqTsUEKAPwSlIfY4V/NbZ
rpzceQvdspN0QnuMsUW9nWeizHlAGJN2+pyp+qSWLLlnqGaI5pnBwntBmnRGqqFU
kUl4rbehpW8DRt477nc18H7177oOJvGOyxP0W+caA6jZSaSNLrzja5JN0RSJt26B
vf+tE07/EV99mY4/Vs0V4tstAJARhqwc5BitT4XdJdNSISjHDUjhraFo0nPFFXlL
m8diBWliiTkTaFGlaUkA9lyoauIRmEDAOFXnCUUCsCoINW5Z+MsTzzoOfEL2H+2y
kQsLWVvnr+a370fSEOcRaE9UWr/5Un7st0axT2TuMz3QSHXf56l4cSz3z+a2Czc1
kyPOck0MagS70CW7fnvuJBP5Uu5i+uu9A5OMBUjNt737v+hXFV+g00MG5N4/ikbA
oKDwm/ZuNpomeLiTWuGF5HXobsGGrcMS4eRcfX/gM5RQOc1YRC//yJlUBhJewign
vXqVWOcyNSjQi23GDwvjmoIOKrDJmg05YPWOHi8YfqVwrLp3rPe2anDEzoktcF3K
5Hpi8UOeaE9C+m4weewcMyGxfiTMexV217ipLO/8Kk4KmvGYLiQJMVhmDVDKnNoe
1Cv+lhImRxPma0tVn+wZdDGRGjkTXt7CanPLNIpLrktCleqm/MqL9iC2+LgxDwV/
LlBeLgE/kD+34tmgp5h7ZLb1H7UnEMPXMn19t9ZbdScS8SBbe/Ityt8qn0pMxZcx
6GnxjOZFC2aIqJFF1MKF5jtIK5OcPmJ5ra6yXxi1X3STiuOBwuZmvnAELbsiCYCz
YTMD1VHDBYpaHA+WASQ+frJsnPB8wiEttkCIzlEc7lahbR1K12ofCXBInx1l1hIQ
u0tL0rGpytyvtvi8SWlu0ML7KVat3jcg64UB57SB9u8cTBFW2RqO+M2k8SwuBY5q
yVH2s9cO8rkzhRTuFsz/vUQ4cV1QG/VD6H2dADzNbA8t8ZniD3wAYuxzmGxGCMEU
ZIRsqDF6hgZ8SIoegukdhLTBUB7fGozBZHDxAKxosjgqT8ncw7fninyuEpotspfV
tOdeL3268Ounl02DURr/MlnDlihlQb3OdfP+bjeA6VBTHr1DHKx57kDDrKmYjJJi
vdFR/WQBmCTIXkn7fabuTqKrl1ub7g2IVJnzJlInuzu30UE8LIyhDAAlKnIrznB/
stVwrLCyCY6ch3FxDhWausr/JVg6WizPzR+22UatG2XBWyqyOIB5+250pQpXTujk
G3MolpYdCoaRSt/cRGpsBZ1aF9okBQw3OsL44V2KX1KGvXrOLep0d/9nUGnrwgC1
CbWPkKsgli7BWrtYS7blqdveQGyQDq8aS0kG/4gMk12mqStuNdjnVZ0pnDfd2zw7
CbD20DG4w2hZqraL9uCJ7W936rttt0ij3pWbDdohrN1BRk/oZsnmbl2vxk7EupGA
DFK8z0VlbohGwhuw6mb6N11VBmuSBcuV6lLEGEEdXJOZgtV5H0g+eZYVAuTXvP4b
8S9GQxppIQxyQsz+HjCUYCms4G7V4d2X9MeckauZ+iR+aaCjpoxRjfeevjNcFTDi
rDKyuN/+MZJrHX4SZQ8ii/IQdbbulYQzdNFx4LpRZES1SOkxuBIJ9i/5vC59tZ/H
fdU9cS3bpsOpJvNjRjcBpY5sgYbn2jlsFQdrAsnZWbFWWDeHLBSsxih8bZ7GmF8E
er+Orzfz3K3q/jhBfqWQo7HCpCSD1n4Lxh2jOx2ubZ49IncOG4cW9mYmFHyfDdxe
EtkEko3ZE+TpucGJOLdpCKzs9sqHZknTenBhjTqoFnziuE/kLYHjZqsBX1jZg0fU
PtX6EmkWTraS8wOr1Xo0ypiAQXZNZ+Hzs5pPthOsS7h20MBa70tvZhLE+/KV5Ogd
KiVPYlYiJMRbXWaqp/kyDFzLJwsKpj2y52Pc8I4zrO+H4DuJHCz8SIXhAU9kYPAj
1uUs4Q4lKY5grSXIm+cljdxvaP0/gIR3JqRQkkcx5AedWDgIHP23V9VuAwU8bjxK
BvZfegpy3G1Xsiepx1i0couH9t+i1fDZ5RvsouPx8UJ3yJEiBOjj5z3Et5ynr58L
fzVvlsrtyL28tRAYFWYZtYbJnTSUwHUTzaXgloVV3FGvBIWhZ3wyq6S53w+0iH57
j0FvwCM+QTSCgI1LbYkS+wSj1d3edxNmG3mjuvyIfVXnD28a6Ri90D850fKWh58p
4TqvTvqBqFSYqg0uHFyfsBlasFlhmx5P3jWPqmPFglHh1SRFh18MU6TVCZxSm+71
i0mScOo2bDDNMnjMqabNNb9wHnLhcrVpyHGWvdYq1rG2ZoTMvV8/tmTqmRjCpIlS
qn0WMBGPhZYTzLvroLLqtb6ZokaQ2AYMe1qGmNQUi/t0Syf0LpAysYXcMvetF3ol
olJQPIMFSmuVqD1Gy3RaIbGbZM+bIEIC3toXrnxPVz/glfyXW1en6+xPhC9RMz63
L3OUD4CKX113XKt3xqrBdGK3oxXL/R75Dzr+8DMfL/vGdoMkCaf9bUtvk09oCDYT
2axy6Kux7IyM/tg5XNo38hLN+0ONwbTfgmqVb67MQbeiyAa5GOlD2nym6Ai36NWE
O/W8kICtp1YIHU7I1km9dO3TR5z5ItKRDumk5FC4Ey2OjaqZyyE9vwH+RrM93qPp
cKsg1SARPoinDkmScY9y/mGlwLt1RTRp64CeJwr/soKQKImYGJ9xeW6LB3N5GRPT
1Rf7r9UCzM4FbH4xg5rIUUTamjOZhIeG26Yy6bi8lbd3K6TfFww91BRcR1azeuYQ
0G0jmoQk32IUMIC1zDmjgebx9F74JqHXAxYcPfNdv4YOmNnj1WosJFXDNflc9MBY
x1rxPo0jAaYzeHbTP1hqT2JLUXTtfT0vKA10OeqldND/mfbQhVN+yNuULHdI7GfI
AxWZq4W8d3i+k4qcN2kE3dr9RgfTjmNNyUZ1nmam/cWKDFkOMgxqFzBmhZ6Tm2Sf
ZS/RyaculJZmCAsuXTFUFr8MJl7tZwPeyYKBYspap/JNKqeY4rYnZXmmDOoJTQgf
Ao9IREXotc3NhiMtiZCYPNuj76ZYTCzgodtEgRgMwrhsHJqOGeHnwr/mKFZJTU1z
gWNKqOiWRlezLevdu4t4L5siAuP2a/jzYy4Y1OBqmgkROdu+6BlUM/Nq8U+zfl+s
FzHl1Jl7bZjRXE/cXz/5JMg5LN65nmOu1L4dAk4kEiQdznYumjpYgL1hyqGfTGMK
iAjEWCPcM55gYpn2AckfqkHU8OggZlGzAgjJOp3z/PbXnLVDBVGyFkCt57Qx7pej
pmjfQSZ0RYPIneqpGSrp//AWdoMTBIUX424GQgrcyoat47eCYBIBED1S791OobXN
+4cad2AO3UFSU+0Nl9PaUk+OTF1lJukI+1wjBxhH3mAgxlgxFPo0lQ0/ncTQnOUL
hxgcvh61u68ISB4RVNYBy8rKl33rLnIOUhJpzJbV5IXwyIOiIJ1EO2km0zH/sMZC
cCPSIyfr+AlkwslvGUEWv8no11WaENCpYA4DSIKUvYGBOkHf//HSKSGoAxyVHJsr
XhZCdN6mrDI8WBJYOUlxtvYiLgiLZjfMWwrrlh8sgl+39EyuBgMBTU1Q4a+hdaK7
NZTA0X0RfyklxjakqWRYtfXekAKixVIOdk6QgX+Rjj1f7c/P5SeQA2RP2hDgbM1S
iBNi0zqZCcui97ZHRktEhQjBVz8oPZqZsgKonBqdRQWjEL4H1uHkh4tSE8DX8mk/
jNAxmJA4IH8W5tzx1TswYekLhI9ehNgdpDujxmp1IIxzT7A46SheLry2EYG7ss5J
YuGzAjzuUWU50MqR03bGegVakex7fLfNjn2oA8LifZf5ObnrnnlJIiDbESf/HOI0
iRUS7IeA/B0wgDfpzMrpt270mqDSBTpbiyt09IM6qxbUN72xppjVUqS+vUwhPTSf
VfytS+YhzBr8JYx0SfHKPK9I9Q9XJ1py/+ZMrGT+7QX+/o3bhZIJQbzRrDOaAmMg
cy8UNFVhU+0ny3DvGO3g7Ox/clwAJFKl8m7jM/O95+QMp+mg1nTma/0k407pJxs7
XmspWCT/puR1xEStwCZL5m+G6pe9Lm8beOuYRJJeoPFYqLGDzN5osoC+Vb0RReds
9LZ/RPZbKKIcTVS3BDYa47HUByjCetyxhMfMY08ki/YDKHAxknXq0Rq6bJct3y/N
IABPYNRSn5qv8sf9H0LuB4dvUH9ylQVqZNZ63e+dlAcdg66vGwOml84tV0z3oMJl
3SEuQLYs6uGGDsRWKVksl3pf1UEV3qIQ+GUAekWhKt4huC3y2eG4inCs5u4Iks+2
p1OdpYZm7OkilvwQyT+nKr3ZQE7/FUBtV+jDgZp5t93yTPIA3zccaPdK9gha4vra
onQJHjsWkzYEA2PbxDWGKs9LGA162lV/6UtZBkVf5AyWRIcW4p2jfcc5mtqx8o3y
efe5zKyWErshk/lEkUjjJkPRg34HvlRIFkHRRGL1HcN13LzZUzQTbn8A8bL197MW
L6KXFZIluD4ZtfFGvK3Se2EuGtSqTHj5IJmIw35Gs5jlRD3AztzPf9UdDMCBFRYe
wP9vvAo56342h/rU/cRbHaOj19Jxi3DqAENsjafoaErd4q4w/7fOiidhh/zj7MIR
U6+9Exud3nU4Ou12BaNpih3Blst9KD7KNAQAwTsXVqKAHAL0mtQ5tMfxHbyVU1pG
7uRBapKXS2ehWHJU/ZbFFwtag/4zR/otiTJBLIqR+2JI8Ar3D4mk/3AleowCTPgB
Bn8+EJFioovqldm4pqciNw5xAKSr9Ng7j+iCvvoEw+ROmzOmc9uKHJYUdEPElUjc
zcIbRUcJ0KWZrsYrraiGDi1OHGwZ7Z7lkVvhBeV0dVnGPsLDkF+QBqOPJzISeIqP
i93DWxaPHCpCPs3x4J7pjC6hUeWumjDBlumhUwF/FS9Zc14w3jmYNvcLiBhrg2ap
kIg3KbB7uqGxUSiycViBbgyBNHUwmA/eNpeTTj1zv7WJ6iFy2tVsec8DMSERWOzR
DE0nhE/kDRuD+PLFWwTLcSz6JYrmv9Lhi5v52W/Xp0v73bxQJNOMqiLBpm2UqSv1
JdDqiJOzQnXLRu6WUAEBw+XDV1IcexsXMEKGGzmW1RnwSJjHnFpyEHNLA84myGko
IhDhz8D8je14L0si2MIkU6NlMh2W0WAoijmO/FmWreMlGoXGWXH3tiBhUDtUwasV
lmirtL0W4+GfaI8MPmiakjDz04HoOHFv5vvFW1fz6NUJDuVa7tv6oPamsdNRKc96
L287C27gj5yhGL7tcToazgiuk/4ZY8hZ0Xz/a9rCDqMmR2jTLvBJADJzri4i3emo
XHNzDkhJXVohpHm8In9RiFtfIWpbiHWgdXDc0EmUb4LkHXZvnnb32n+URGWq0WNv
UMhFsiPuWkDOkNNTt67x0jjz5siLIC4aOEePLUAOpfNEbr+Evf322Td51pNlDVD7
EwCm93sQW45nvQvraPCWww59Rt9xl06crRgjmmzhEu3+oVo2K75ICT7GE927EV6I
xRmrWkYr2az+/oiV/tGP9g1FumA/BUNiNZwOQDivpv0Q/UGgXe9LPf5B7O+YAdWZ
Ol7YFbbO00vR0GAnQNKdI2obRUiPblP0FfwTtCqj4DJ/hJJEeFKbtaW/kDSNcaMV
xqb28XIJ040Cgfc+WT9MF/fnMQplFTOX8qbLjL0PbgY7vYkrgZwgZtDl8532bFAP
3z2+xt80oWrsi8cuTksy+v9wTGKtPct7WH6vN9wmDzew6BU7nQCFTLbxQbi1K7RU
+ySUcYuwwCIquCjC5cz/5PAWznJCNB34b5Yz9F2a18i8l+X4B6w3qkd3qwAPwvp5
RNnZDezvSGqdunLnMXsYD352Iszj2NZKXcxsyAPuulX+9K5cOyBPYosX4qHwl2J+
t+EzXYkE9p6p7D9nvDpM58XFqqYUSx0Vuyf2IZJBW6gWXnWddVlHxnLdoNB60JBG
5O+6bKMK37fUqkjz5lkgOoKZMAbMZ5O+cegxWgxfhIT1uIM0nobYVzsibpX0sW6K
xJGDXaSu3WuRIAyKyQVSJThq6jraHXRCdQ0IOWz7Yhz2l9upgDdmIMMesnza87Ws
IDNibqjL0FfZHIcVBUu/UPBvXJ8Q2Ei9mCb3Y6FhjCeBWzpQgKBCYT8y4PbiRuNQ
IHBJfpHCvzIWX9ledRT9a+82hpY6mzfvdf5DhCRT8VmkzoeCB6oAS3GVfNIzCJYY
+4H9gFHNMnIwmfoGX+wlf6/NLo++pYI5QVzCRrqJrKJox3NWaw8bnCeufEaDK641
Aik7lthmAMDzKJ9zjygeGvLAQ5JKkcnWmfDXN8HZ6Zqh/jw1TrO7yzBLn4ykaBYi
OF3mGeeVhFTkhSn//Mq1wwkoyjSok4piHZhtV8sdJLORnckKyBpZP2JmPqImWExv
3r/M77CmbRwnKPENKz7umrG0EaBT/faDRUTOBePnpHF1Bqp9HQKE2gYs9ph4ZDTy
KC8ukOKCmnsDYEL72qV+1Z1uM82QMZfsgzqJor46VMP3baONuWWRIKHuZl+zEbJz
T5UrtKKmLvDMWRyticU1Qch2nICEbKJfeJJc10ouIUGJdvC5OIPrq3yu/YHzO4no
VChqnMUIhR8M6W6vvAEMaYOB3l0KijvZFcDZ3HFiB8LrehbiYm8EjArCZDESmFBs
pTSdfhPb+X2daE8SDucE75m4MmR10OQhCv0L6RihOPHDpFlt89HOl48OAOAzy8Nq
57o1eVo4jrBUa/a6USilF21dQ4xOPBJgmtY2HsVmLgwzsnWvP7VgBZOS8crqxAi/
0uZZyImcGjmTwd4kk/JgXEWM2/B77M9DRNlWzufRTeX4G32e94ICS/dFJzL2tO71
wkuo1SNTIRiJ6aGH9iCKb1AlKI5XEIUQOyYfpsBa5dBxws5/4+IrHBC5uqAd/4yv
K4ogypKwuJ3H9Mk782rMYUOb/PtsfV5IpNATx5Qa6llrjb1C4K3teae5YZ9s6mHd
yDnG2KRzW8XP57mrAgdptm6AdJwo1Pq7A9xy1uI6ULPVQ6BUadyiAp3DyD7iqK9M
UzsWQYavnViD6mXoRl52k1CyitZmAv4Tl9+Ff04g29z2oAxOy9EWQuzyuAQaSNTx
NwUX7rn/sVGCUF8IDnHgzmZya9hq6v+OB0Toez3QC5juAUQQAf0itqhZN8ThaBIQ
eO8ysjLtihUHYzQNrRYUu/Sq02Jr4CwCsNBXFgf2sq2t3jJ0Vo5WpPWhpZuGr4ot
bn5LeyYI5DF1HTPLCu6PtOlG1/Upewgj0uaKZFhdsDgGKoAh1SYpBV0axI7Jg0bH
Aq3Q2n1qTBdKQ19xC7lgloJhLeUTOU6nfQctw8v1SiSdrydcP/B1nNvchn12lvLv
bUZgShobpfUPqIB02fCEQifPNGJ4uURvXtgs9gb33TDDiCgf1igVH7WyeRhSYF9O
Lc6cF5YbeTp2zQ6o0isNRWcKerUGrzaIBz4fxQYGbuN0GSiD7scqYPbjRzr4IJZU
EgIUz8BhgQiSwnXnYn+ZKmyLTvNjCfhBwAwiarvUdzWdDBm6MtRssWDIAic1z8u+
vwjGgg0aNB9ITNfS4yoqVHAomWKCZqDmW0dMuTIyQv79MR1T4yc1lBJK9abUCfNm
uBoIsccLKOlP1/m7ATmTZauVQwP5quv8xbP6cY7rbbbUCIGpqlc7/kusJrgSHHd6
/6xz9sg1ZqNMau+c8+73YSZQKrnss3Y1xG7Zsb0Ducqk+ZiMwRf4QrrDatGmdPRk
ayvYT73+fvb4anbnMyKgTTvyf3NEBkyZPxu66UIznEYCSpCHUBtNRipAJoHEEV0S
jWaXg6VvbeLHhh5jQkIh57hGFnq9ChAWSMHcPlYYLe9+wD8knHIw1QxW4P3iy64R
49Jy9RykjCtlN3R2UxYr1X76J7gWmR/nofVXZ8qZBvDyTyLGFAEBTNr8+LVsT1hV
oph1vAn6cDlRX4qMQBIDajss1dqCyhRu0CS4y4fO/11VHO+eFVsXq5BbOmjPR9Iy
zMtcfGYuHMjtZ79yQNxhCeOwUd06gxiUfZevYw3sz2tQHMoCVa5Tgw9W6pBANQBN
C0ZU36tA4na6OgLSrIaLKEZbn0el/gg0bKiwCetMiwTnRgCytqggghjVsCa2SMfw
laB3M/4EfKDhqPDHFOf8pbaaWSdUyxgD4EkflK2SpNKakt0nZi+ONjfm21Q76xOn
iXslkQB1lUwuQPFv0kYltFQVc19frfwpOPPBxPjaq59yFuD6pCqc1lBwNbij1d3m
3WcvNMRPnAwjP15WMaCNY4l2nq9HuUYtHY0tpmtdSpte+I3faVP8Kf9bmVe4yz4n
EYaSpGEbu9acFbNxXvg5CyyS7v+opBe19J2aFjFvDpZOhjECV0rV1lj01bGNZfPt
zqcjgIKAJYo7SxOmAagwlX7Yjt9FrjLdbhrmJjq4ZIZtvKBsaP4OYzVJhMKSM6NA
oJz8t8Kt2kGZ9pu9LErEUP2eAmiLglXv6vDKj0MPyzarhAJAb8UF4JEB52NvZnTe
Hez/URdBBl8+XbWMDAHZjvKI+vOln9Rfl+Km+zzw2onrP8DWmHsjf1eRvDkdnxMu
1j2PvM1eR2v42HYZoKAIIPtQVe8cTQ+aaN2PO4nmsYaeTrtZEtvZqrMw7M9bEvrF
xzljCRpCclVIgub9P+/BK3vfOSdVY0EfFo1BEKT7ojadN2kFanDFs9T3M1+unl2d
CxxIyvMdfezEiN0Jk2GvZFSF4Fmxw90O6JsbqY4ABPeQ7pXfCdP4SBg7ZLphnwFP
t1LSrPyM5sGvzz8twdUS4wHjO9ox9V6fSdB6AuqjOJqm2BKOsvyKAFj8LbnUQ8+c
UhArR8VnjmoqNH9LCQZbHxgWUywR64kgRg6IXhta1JLpPoYvT9BJHJnyORgh1DsL
+b0ofEBBkVM60xKEVb536xU+xyLdd7/u5TVWeBrKH/zpU1Qy1MrrhzXWxGRUtXz0
wCVskZA4I5cykcqZS69q2FmaBsLsv41M7T+q4MWpArCYJvOyarKh6ZdImEMv8gHE
SI5Mut7y2Q4wVzGxODaAq99tf1CH3OiwNn3ymzqhRmZJ65EaY7AB9Fzd6JKK2cDm
C/kjsdbaWgRwv265ARdK/+G5tQn/Be2YgxWdBvjaJIPzvK5iVA1KCLHl4fwW7UPn
ZMQTEuxmD4S/Lvi/8Q6OvStrYPC6XeP2pb89bAZm3/6soYR4WjernBua6Z2ymR3b
SH8h1xslNIYbH8/ZHQT75AjJFD43nLUtv01j8J3/1y85pksJsR657f7e9jmd23w7
XGqoPHTcxugoZUv+e/VUMKbamB0EvdZ72cSKvfohgVvD2160jngfDWuShx3FLcXF
UNuftPrkCegNpNSHD8dUxxabgJPWgpcDpqc4+1znGOqFirbx3rm7hIhvpepB8uZc
j1s/9wYcDf0IyofI8L9dcgx7NtySi/+XfiQeadeOst3847ygOib38kzsidgtTwS8
/s3kXLtbgYxbboLLYf8YJcgWLovgkrKMSIaYNL2IpibLwke3gtJMFbtg/I6f6VnR
T0R8fYFt8BawSHXc15jYBjyIzgJA+ASa7TRVjj6xeSh2d3+NVDQtx1Z2Mfe0v3IW
+yvC7N3rN/nF2Aw43+JOLy3ovlZGsLtLRmIhhSX5pc46pvFDT7J2KMS2SHUZS4kd
5qL5/ySjAFaw/lF8onkjp/XtdhYxqgpsaeyPMU2TFp3QrBZFnWMjMsrqt9f4cD6O
9+KTtekaa2JrZkTjpOoHWeYpPc5pqitZsGuBVc72vKSt3fcad5/hrUr/F4H/jkvM
ZWxOZEjHcVx4RVgjLCGBJ1mL2IXL0I3ojRoOziMSr8LtTeRUJNU9Q4dK/Kr2KEyx
tCxYvE9pgko36H1X1YAHjdZ4xpmSzTi9kQ8UigCNbOm1g1/oqfEew1k7kldT1iYC
eVwmcbvfpqRs7o4nUN9BTdUEDpPgGrZO6f2K9pq2atN2+SixnnxDxfLjN6XMQ836
KaMQFJOL9mCOiA/jX/Gk05pIcopzUTzIS6Rk7YA73wj0Cio1GUikMTDfSTPj1KQm
UizNRCIC2xzg6djMVcGaR69cdsRIZafJf9h2lEZuY8FoO/WAEfotTlbhzzqo/3Bk
LMj9PnC+oRmhLCSNBoUyj+vS3lEC6UTM3J9lFdL7ol+x9qWHKPHyXtlyfPJFxuFg
rgbZnwf3HH1EgIw6o2No1NgIz7po9UYouVvvM3j7kcWBcEOjY3rOjDSJz5CC7hk0
DH4zP6fm+d+WgO/VEMr+7vc8xE63J10RkmUDIsgARlUuxdfM3olonJdp75vneRwq
G3F6OAT1IytErG4n//Lbn5fnBsnq2rWGkawpqTwM7fnMs+gPbKxuVqXavzDc5Vre
zL+nOyeRIR/veEaOnIm+RdDbUbINleHpN18lQHGAZJtZi8paevG6vsSIVkRHkwtO
35Cn/CK0tNfn8OHhdX7cGoAgGBQEfaZ+XlN7LvD7cS/GOMpeP5h9hQpF1AE20mrL
fxnuu6LUqqvOjkDutYy10RSYu8VwVXnXQd/j1nNT+raTqaCISZmG9erSqoVxuSWj
YDdMltaVq/0CnyZ+xaJsFdunPThcxx2uNrU2YKrbEa1uMi4+TcDy4yXe9VwHxUMd
f7F+ikFSZhnKQOZYKq9x56ZgvcBohTVPLeHJLDXi4h82+S6zwRkUlKf2QODO4fUr
dM5XyKGlAfhKHcBvDoIFovOwwLsAjToN+U0oYvjnOHs2PFV8jfBqMv2eNaShWisw
E+EPb7kTcj7pZHfjgvNDmQfRMbhX+uOGyINPnLk72NEEURS3NIGqPyAsZQEGGenO
QBqUFKu8m18NeqJZ1lgEMhH6InYZ9IcydxQAMI5IV6JdKBg7sNY2ed32gEV4u2V3
f+21sJJVJgvwbN29zbvCopghRsOkoTdJNECiVtFYRhy/hEZ/Tkhsok2uUrCdQ8wJ
+U+ub91aDzag0u9IhK1Tu5pIE2NuWfdmuPqjZIyGH4IgC2gvRYISScaOci358Kko
8wgwtmK6v6DfmMPj+Q76j0LE6UHEpoPBn8FDktUvAe7l+VVXmMRjz5yub3CNXgWz
wHjviM7BfhwM2wk3ZLgezaKVQpx3+Swc7w4dHZN3xivgVs/+4851wuQ07FlcF1dK
TjYg1QBmdwWd2VZgykFuKZOsDtdcvAnDOaASuI5whbcuVp637vk1xJxZoD2wENiX
Ht9Tz9YNiLgSy5hZVapfMabBaQsbM7qeQxZn/VH+FAMkJ6DEFaczgtfcdukFa+5W
bI99+ldEuEacHkhqlxDpo6dSfn90NvZfHCE9see6NQRdM1xhGJwl6xVxRj8bR6wV
beVrKl17D01QRb7OO30twEvzK4ag7jXSKJl6Cap1EmwcyiOKAy7wiFOrbk0RXpgp
NDmZex8K9f1SPcnMK/ckFch0nVLD2XzAkNEV742jR4oljp6auW6e8Ni+QeTW0952
XCtosf7N01G7q7GPJzyuQD08a/KckGHKuFUHohuWnvhfQo+4zlENr/3HPd0EpE8n
6XOYR9AebDaemBFwGU2MqkOtcnLMfUpvoKNH8Nsz1eR8erhKA/4LVsM5Vh/wSRGV
LLmcJt9Rh05prWrv4ISJFjtg6KNfOT9n2hJ6sOEW9s4VkPryJn+EIWI05I6h5sm8
CFfgTWfZpKYIfxa8Gyxf0fydqHXaxv9WI5oqaIq44fLNPtNH9i+ch1lUzP94B7r/
VnOKZC9ICPrK9l0z0q1TwV+cj25c0m9pbku00gVFojqa0xSBFcybXTA+fraYZNL4
Vg3z/3Op6g70rF+yfH5lYOoq7ZJ2jhoaSes06Olu7JMKjMuH2BgbW5mGXE1ey9ma
amL6ZM/OlHBC34l+FWWq24IOjS5cDdGujMkH4W+b3ea+50HQskfozibCg3UGO4qi
onQxq4AFtvnSsQZBjzN6qCA+laJkuDSQ7ZAtvjbYmK6ytaSowTHYOL0ZBzZFyYSf
7ISLdWZwQZWeGJgjwUulNM1Oer0lhhfsFG6LrOjrrBFY/XvLT2d1sdsVteA1pW85
GbZNs6hfCqD8YzXQztJqzAeTw3GFF5qVsIf4x49iEL0TBD12czYttFj9IcxIpy+G
dlLdq5BJMCgcvUQz2GTYfHwGe0rcTqwcYpnPmcmD2hguEl55zA74w1PFgfClKRFy
RYAgPHA2rITPma48iCNfO8blo/r5vSV9nyzU1ADc8P7k/HS1ItH73fG86xTF26gv
34Ze4SlWlyIyGHyn0xeGZ/8CNGIMzQk3MrtAUoDhgvqbBsULp/1bsWAKcd0qSP3i
cL0QlXqncJfe60PvE1Y697C9+LiNFi5umJdd3cTT0+0s/9oC84aOP1ujMr1Ts1CT
vlN3m8tgtiq2DykLnBkHwi04qi0XN5ukR+wAeH3W1In9H5J16p6mJfWZIxXQKyZa
wy+NdTjgHSj4v6rD/iWmQSYprXKxl/y8JXZYImC+i/Y2nEE1jGKVbWHSyHu8ngXL
ttBcerW3ADsMYSgkiteLISmWzVkvCuNrcpCv53j7K20NBU2bM/jzAVy4dwAun3/B
YrK8YVW046QTeczlW+8CDUEy5ShkWqHcPfoQ8NjUDRod/wy1qfxa0gNn/6821K44
Os68CWqc1IEtzN3InqzxYasKfhTmoIXVTBz3MQagRNBwgbR/tl+KG4XE9/Nh00XL
hOgvAQYqzHct+V1A7kcMQESX7+YXGdSTUYgy6udhcuC0OVHElyBmLOB4RATFyykI
ujMw3mQ+pOmMGsmiov3I/YezwlftKOk0npRo5KqvprBCC7wQu3+qEtcFmYfG1WV/
T5R4r42gDv4blDRVH1Ni2EEpg9P2WF4d7CvTWrK+D/drMFppasHzC1C3ygork7Wk
KgEpJrCQhm+LyPxa5b0rGEmgwUuIqg0AnXx59AA3K21vIaQkrXhE2r7q3s00knTb
1X5XjJAPL9kTiUVifso3ncnzjnFFMciT3SoGqCsLGdTspFo7eThh42JCrqIizvwr
5lbG/ZhsHIh84R5jy3Af8PxxVR+36D34X+hIPNWWW445xQdFZM+/0hA01ZQvx5q+
D84qOqcwig4lZnIEuxMxRiKuSEWxCPeJMiXM6igbQoEyLrZvIDqzJXVIduWRAb+q
oGeyIRG1unO9EKalpoqwwi/vAhKLnkRxXjh3m6RKkYXn+ruY0U8g7F48DiR9DfdZ
p/xFpK3elRBwOxg3R+dJPHk4S1PsVCtsEyWxI0Pciy3pG/qzFa0bSDPXVQjxRpBd
AqHzA0iNmjWhhPZdqfD8H84NT203Zo0ulbu31+OmUi52jyWRX65bJ2Y2vBbi0WpM
b+aDamIfo1vQeu0KBO932iRUahbwMw4Bls2HFBEWsrfV/NxceDXsr0eECyI3fwmG
BNtqZetuzJ5DCrz7GFaT2TSMl3siBSUupy92q82+lAYE2NocUqwTLoJ+U6bWtx6n
e2kEWb5DlLBIBtZEOo5WUI6nnxZE+J1uEqbc6h1kzmpZpDTuhKFiTx+1gxgBURet
g+4FTLgjM50HM7fRZGD0wO72lTJ1mnpO4jVzwGvpUn0E1z+KoBxgis6Utl8dbhQL
RpI/oFMYeG0nDw/3LkyswMT44XiBuEHhsazw2X7GU9zelAG9IIJ1j84lHXycTXMq
dkYy7zImmZTNKv8nqJAF7l0sfVa8Ot8S5E7ZGSZ65X1jfF8+/+nGMWqzE1i14O1z
nCTJ+Jcv9CxewfU+7ho4WZMgy7IcXDikW9BvawuG9oGPJjpaa42MVUN2U+HsS886
ucSEMCnvSBt2riC7xa7s9wUQdF/iXuSehG6jqahxsY9uXTHWn/kifF57/1dGBIEG
oLr56Q4I7rMc5NRss4hqa6lJeMP0OC+fiYW/zkZdeDIqWhGy21yWwFkCVxk5sMCG
PU7K9cwavku5ieMExHhE4aEl3CFi0W0/fXimXDugf2EzCJD4bxbANi4N39x9R8a9
gcMfw/vB6YDtnTLtHVxV4S6Dr7sO7aALPv9yTR8NJdhKOe4SjcoCHHXz/hyDuKS1
EVBDgWerD1b0IQqGosYIEp/lrGQWI0xz+ejlHTqYndJSFu7BylL52sidJZpw4U3Y
mTUUEyWncEhy/dwbw3KzL1yMQC7yV482H0eFWmKivOtgO52FssSgKOpI4GmDJ7Tt
HsLHg2PleQUg9uPjeZ5W0DpPqH2BTKgjl4GoW5dKryRVHMnT74oxN/KupynSH6+z
Vzs9ZhiaM6zt040Xp/UMbjErhDFR5PNy+zALk4e/EYir8wfr7lSwXjJrB6yTFWEt
oq6l/i1McXHT4bEo0JEVlXmxT+PE3t5jsH1U7M9NkU1bZkqE3DoifP/GTr/bYo50
dB0imzJX0DqiL5nQCUJlnCFIKmpQDwC8TsCYunZyhB0Qbgbt/jNETw+WGTPXCnRv
nOWP4dAvaPPFxY562bjlNLyPz6SfCrGD+bS+LUUvuJDUYRndfxAtZjGvioHTFcVv
h1Xg8HQWCOaj7w3K7bles94n9Q4QFrqzSMv2SOoZ8yL3/l3x9HDvNbvmTddt7Qp9
XYaT7Ra4e3psz6lDhIXcQhV9FSTWDhOFfC0jfYh9EYQtnJOTQa5K6+PUyqH76G32
5UcNEDm1QDyiVkiAHo2MgBH9NXk4x38H+r3+j/ESG6323/+L/b2BYGpghe9wXwfu
hQm5hiO7pHkbORN4PC9v6297dM7P9307CifkkiPvrTr+4GZqBEYv1Pl2BItxj8Tf
eDtMU/W5pgC9qbQzYLZC6EK3UyWslURoJoDPByklJJnvy86G+IRCVz1t8lIDYE8K
xVyFO3pd/MayDaVrr/2NMllwH4IiGas16nptaLNbUB6PCAb2/3ZSRGX17d2uqQHS
8X7GGzJ27vr7PZLu4W4aqw4pDkPWjlBRp4gSsVK74d0y5WsyJlTI1EC9M5y8umqZ
Nsds167IE3HLbpgzfo7Y1lO9cxLMAlE0sMpGnvqfKSPKyrDNV/iUia5t3J01vn6D
xHd3dKEcP7yUzllFQaont6nabKG5KPznJdMhHSUPybAkFPuI1gjLbjgsKMJ/0kKp
6JOFo5959zPkH2RWOAGWBGI//iq2RzOKHIjrOyx9CuUG5h7KZRwN4I4gRdRft1Dz
hYy4ISJpXx9rSnMwcVM9LYZIZLS8ZSaSgEN5orWvy1F7KDW4D0LBrteWp8LJciJG
CVuJmtwA8XqmHwMQVrCM9LfzY3LDRjP2QiFCh0Jz6D4sw5+3sinq+OPOGPTRZQ8k
oxcoNkObWtp72zT/SrRVNFMvAaKXte5xqaTBf+YenvqH107V5mC5GQAg4Df30JuA
RO4oQjRcM5aqzc4q/GqoRp8jVnrcf73EyXUDyqbdJqKsCX8yq0SsbVH3rXsUboMO
ctNyGTTGTryL85q3VH7Lz4K2df/MVDLNMCuvfRYzItunks7eSaa3rr+KZM4jeExn
8BWpF+C4DH8ne/GajQNe9ZzusPJEeKjooSXFL4WtPD5OD3Jz5JIXKuTeYfcLpmdC
E7ba0oyMBdPLzNUMunn/qnfvgS2OdcH+xfKHlFUjtaCKGLTfr8gfiXE3O0UNLFFW
JR01EqjZCjE8/QgWocZ16jw3UU3oKT1gWMn4PJ0HFTlCkL1huPhm/ackzpQ2ra4P
E69gJMYFx8CgfXYP+soYC05QQOLq+gRRjCmqaYimWhgh8K0wtyaQ8wWAiId0djD7
6BpTi+52lvS46iIFwNQPFVo/KV7Ieuiuxz+qz5CZ7cJyM2qyQplHMMjahx0eRTdg
PuI4VKxCAKs0XmEV0Oa0picQ5gW+YwbZrRH5YRJPGkY0Ed9y86KZN3frWeD0YlmW
VTAExEqvJUb2arhlkxLzIz0n1R5aeql5683wjKXi6/3ilOS3es5emMbwa4p/o8IB
hiWysRn+j1Ikge3KZv17KSQae0bv9o658+046Lsfu+wiNmoYt5BcpghH8I4wIDIk
JH3jgZXwvUeZQYjJMQoYzqbRU21AtXVoZD8U+ja+BK4L3h6u6VEFn3opwK+V6FNr
lEGMKegmkgojCxMcgeAUdb+s2rCAotiBASCcAowW0e2qyNQc4AocoMmY3IpCcO+z
PFfQCDRlt/eFxYS+PlFfZpIlJgUHlfTh+NZjdg2vUmjSAgerltZGzdFqjoL9rUH8
aShbtCZXO5rAPBgjhSFKh2Y/jI1H9zoIB1d+4pLcLnfb5HfDnkPsH7uRMA20iIAk
sePYtdWZcNnk9xoZdacLr665qDwlalYJ4vsuA7ZmgOAPHSMCOQlcsm1HCX66cL/x
FnGM+Cbqu0Zut7UwzAMCNCB058vFhzMTxvDq+ng5tZF5SgEd0zH1k9x2WVbL1XQW
raaxkoSAiLQ9nmF/3hzymatavrFp19n1PC//uyGyZnttiwigzOFsgDZ8/scJhFyw
bM/20Z034wQGJpgOma5j9bwSN4wuD57AirWT7w4hqVJ0sOlLm3SsphYc5i2+Gvlq
yh8wuRSEhtNzoBPuxdkd3BUOU0YGAB+eutg4rCEMUhqBxKkEIm1IMqInkHgYs8Kw
Z090PZUA39SvpxMrmYgHcFEFd1KWawk2/E4cFLLSbOkfzZLflXwx55tf9AKZq/q7
g1ol4IO9Hl4Jh4e0fKUOrzsSMBIdHrlkTGZ3qzNJYIpRYBPPCGHYhSAB8B3FTWXR
DvC4/xn1s6YXjQ8SXXZKjtBMrKwYkoee/at2LQuLhQ5Lu/mcU0MUzeIBPlRkz8j8
lr1RxlcyWTtn9WhPTUYfdi6Eyhz2xQH0A/AERKySySTZab7p2RyzD5crmAzfYfUo
7+vg6tbzyaS/ad8fIChhDhrnO742SGgbtqnxhx9XPftMkonO7DHZnyZL1Put83+Y
xUDzwIngIYW9IJH02XOGsDTCQA0UWornsr1wilpI6XldN89Mx+kDuFmeREkVPW/w
vbqi/UQwlvQ9q9atG+YoupNjqSjciRtzgLD9fr9J+0JG+3q2Y9MjZRRtvIPmllxS
FaxoHhE5dwmE4+da1cyH37evlzphZxG/MDdyRk/KxwhUNyS0vccfkZn9aP568+8B
eA1NKjP0LRB+TbKALL2qkHyfX/vRWk6C6dSsEotgN/Yzu+ILUgeEeJtIRKtRSfje
v7I7UXP9NFSu7LJmd0t0hqZPxufIBXz0HvqxUb8aSne1fJjPczh9IbWgekICWLIu
F+Ogd01okDb4aY2+kZmX5I8cJId3gFAM1D6EDTIS1Mc7wgnXs9FDR9BdFsZgRvJa
Ps2l/zd51LdJ2ge+YpASe5I4dLC2juLPgrgwEssW7l3floYB5F5nWn3ZV42QzPpk
8uAzlSswdPWd0FQYC2s9cPa4nNonaVBmbPoTzlHXAkeobY3VRA4VGpsZxarO3Orj
HCNXln2Jsfi19CP7kf58btqq14AOpkO6oz9+d7Ln198hBC6Yge1i0hFnbz/vW01/
XQJBAAWxYoZVpY9YpZfzQvA7zm9ZV1eYNo2CwBRGgaElSXYhzCRvYSoPpT6PIMfm
1vY+a10jJ3ADxm5/W2ggPiJELWPpXxqGWqoGbEb6tI6ALN9lvxckpu+nycXABk1M
wvyScDvbn+0e7zN3dzMFTHsyQ5bul3HiHLeC0vpGI9Fj8LsoD3jbeyvUbXdYJgG+
0ZgjxX8KsfOj2vQP1SvD4g7tFTaMOV4MLr/QXB2E62IQWMHtPlFe9Bz4WrqIvRu3
Vo0Z1CTEvNTP+dqlOt0+VpfXEDbieUmNQ+iof9xCkET+2MZWU0k6JW7lmG+acdqR
zIm4hh0fGOKoKdeEQpd3brA1Eu+4N4lQfEsEKZvVcFfC16K8g4Ks/9EFNp9+uBmM
lBXewSYMZtqZbs6zanEtlvCbKsuJc4XCPPw4AZtuQYI01mdzhY7RAWUtFPVF6c9L
9u06WszV/6e4OMK7qXrzTQ6IqOMitvltLqmVSMvQGt0YjF3GUr+ozBDFIfswrjfK
rVwFCMsx3Y+w8JiRL0zXY7SSjMjooeO7mUEgXpvXnhrTelRSAn39RYigro2TTB3F
xkKMJlYyBlc4FnGp5HijNJcdlUS3n+0HFSFXRvZuh9UVbQ6z4sP85kAnVej+UVEU
GHGCoeuTq7P1CtqrHP3UdqVx+v9JAbtpmVWeZTBVQw7YlPy/dsXlpNnULlIwAQ4k
GRNPKWpFAmIyg+btd99B47eiBQUdIW7y1Tzd/44+uKIKLMecUxdyJu3tAXQnFmIo
88r3m+aPxPdKG/29K22MWWfCpagydrayqm6/dQUYC4tUHDilY801L+yMjYwPL7zO
CyZU3mP7Ql1YUmP1NmMyzot9LwzHV4MIEH957iykDbylOyql5/LoTojJQx2IHVUf
Z1+eFWGjghUFDB7bQ7OYHCKkcVueLr5S/QKqdLTGaGHFOlMzybrRWa9uMwK8+v+1
zw4vzlnFtEkTVMQAAbo18PCARjYAr9ZWuao4F54zlKiTw7hftHiFUNQScE4Wku3e
Zcdse91xmQmFuD3aUuHloztikd7q9YVelVxfmHfJ71hNqxSwC/4IfMoSqMuo+m0G
Ko9fPyzUboECoO73LS9jjgxFOSVcBy01ZXqpzjUVWgH+BqiClaT7SD9qbM+xC/U+
oBsbm8enn92oBfWWymfpQjkc/0kz0oGod9KPatpmkF6u+iOzT4kcwnKi0RySXwwa
Tnl1h2XD/DDTsZbFiZqxlEJWZ8+xPY4P1ys2CNg8qajgbzmBtyXfI6GzDanq1F+c
E2VnCvIurobTUrpWCefUXdzl+XUUiZKoH2fRVgytFXMEIqLALsefy+vCqGkPgg3s
Iq6i21wbRHyJzKIjhf7eq7L6lhszTxWYHQk/syPLtxFY3A8VSa9ODsnMs4LjHwCA
+/BriktrYVYGCsRNKh5rF4tTw6NO5oFlRkFpTTsiKp6rcnUxNcXkH0u9yzUert28
k1gxoZfWmzUQu3RrLhiB7MIkwGORO20wAhX5FKZpluVVnOt2K920B4Car7iCnZIu
MluoblA9YmQNkc7ZqIO37YnUEw8BI1MGHpyguQAKm5wvCxG5dHgRJ/Gbs2UBL+Li
FGvDAiHV/nx2ITQOdhSH5aQHYyZqiOvG/VTAvs+aJNCh+T1cNv/o3n6LBoQGIPpx
TmQqsQYesdLp4jUVBhyDcNlPSm2+s3NyR8JBKt9Ew+emVmO701jaenPDjUUdCNSr
U6TUjO02DDIZerexv5bgSotYdg9yGwWooAGaaT1W8LPhE+p02sVfC0KkohO8smZ0
xuS1qrlmjclaDrGVZulCtgF/a5uS9r/YTjOzjSWHCYX1hcEuO98zpdk9jClCeScW
Cug7+dGGFAyCTUNmC1rP/eP5H1jmJyA6SqfIvOPXinE3/ldNnaejqWseDoX6Ny4C
WCocoJJ/bTGkGhJeIpOzI5oltoJh44iBUc5CRcDczmcDLIj0dAAx8AX3PttxDFXH
5TqPBM/B6o7vLy3P9zEKKTnYX0A44g3Y4JRb6GmvTe0LBV3xAeJOiCREk1jDPDEk
YcgoSiNe0IvOM/da3oFhDO/GAtoP+BIAT6UpgEulWZjeVoMZc5x2kRUDddDYvHI5
Ovtods/jN/Egc9qaxnUPtnmgDPqRi0MgFIVZsYscb80trN2wX3W71/OMy8846NRS
wxX2q1R7WNbtICcowlhabTA6bRgRRxgcsZVNFELRp1AiiwDsUaMkzfi/N6xvi4sc
foTurLB6bSUrydJiyE7rULGFfsBmoWb2XjPWptRBn0IsrGvGUrI9n/dvKoUBWN0/
5shdruHdNkoDJpUzvx57159qbrXGjAN3qTU0QtG5zWDYrFeot127vDBQGwpCeDNc
fEmqNgLE2UvSemNyUOyzlmenHBzj/NdC3f/EWgwyFYMt2el++sdlIehDJNViI/mW
GUAawJC1AOcIeljsQa5oQqP+IzSndZUqwsCQGjzqZebzydtEcTmKqeZXHhnMJXDY
+he7CK8AW2TXUG0UD3jWiA7YNVcKdzlfPPSbsJ/nw6ffR0T087NevZ48uqsF4XPZ
ws/vbxLysOJePTg8yOr7LaV2bTY2bRSQSR/4hmb8BdouiObwK8TB8Oxo0AzBNmdq
OuRO09+pRmpnu7TI9eabu+9gyIzB3vfeM99/xe7d+af8mcsO3L26F5l51kLTuG9E
X5wHYaOUOY6WbAeZLlwjW3BMpHs61/M2MEGM4sjiXl/ExVfh1YbWd0LAz9wjOsuM
q+cO7cH/DPeoz1OiP+FzyYomutg3yGniSp/thOX4eZnWXME3icN3xMa8Vtr+3CIo
+0LOfCgHNWCl+K5I300V9+Pk7Em4qVLFoVmDnOiOLNupnuyNTTsCn+XUcdbbrZUn
2JZ1e4S84v2I3D6yB4E9q6g1mq5ll6bpzT2WIJf/MX5RLKhuVOvcxRXq1uXu0PIg
RtNUHfvykv/7QYavtJoaDko8qRgtE0SML7aOyPGAgmLj1eBMNL6B9jjGTvKoS7PA
+v4HF7skEQq6M7yCT3F9hkP1+RZ/5sbc7SN6pfSMyA4GianSl3Pqiaez21/kgbLV
LVoeDGGPT1aiLYehmFOLpfjrSMLyQ8Nn9A2Psav76ILakUdudAsbSCHGppEia6Ja
92xPvVOMcFAf4ZYMuJ2Xqsd8fHJWwKFdSgM9myytwF0IfiFyBOVQg+HZIgNHubUO
tzfgwfDl8t09FultYWd1EPq2C7CcGeZMvgWVP76VdY6tfu7UrtMZ1SpdMGaomXJp
mCUmN22LtQxtcdtPKoYQS0Xv/BlHoKh3ytDvVupVySwdE5w9lb3cA54sQRbcrSl+
cL9riryCnY3vHQbLLcHV6wIzMWuajQUiL3GYNOlp19jd20J4pG20IyxQqBeWwcuL
qHB0m/bMjwOBES3Iyh3wlHDMHbmt9fxeXMG40oLzkFX6nmmHhCZXpzq3hb6CJCDQ
DRR38iT+W3nS3fb6AvslPIPC9gD6YGG3p9HZ1nv/sfwjuUucKM5+/Z1UYU+irVKE
gXBf+ZBOVWoM/ALvmRFOjvXxBrrL1IjQnsFZFLaMx70f4aJxj/AsC+8xpX6gAP+J
9z30lT1z9fpMTq04mt+cHgMvpdQd27xLwhDVw92Z8zpPmc7B0k3O2oW78TLoF32m
rBNjatcbesjqceGzurwvLpfxuKcNuS7q7rUNH79VT4XkiVaYtW4VRwiZ2JBwyeyG
B2sFrKuWyYX9iUirA2oahD6DbZ4jKdCb9uqwAkEgzVOxSDHjNf/E/9luyCnpRNlp
nR4q8nfC0za3gV3DvMd45XkghYwFccc9RIZOAXpXyJc4xOAFCZe7krhHZiZ24qa3
2h+QbNakCbCvcP1TkvDpMJK7jQFO/0im1DwbqgYkO/R/O+fu2jB90CqO17mWVEqh
gbNlelLWDKTUzZuk55GJyKhYlAe4jvjOKeVwiVU4PoKy4HsqxMSRDOEgxps3PUh0
4C1MB/oEDgq51W1ZUpMkIpuOz/dWTYHwjpML3awnLjo5OvcXGfIknPkZzpr0wyqM
5XmfeSOMt9N/h1JudkMJF2dgZsf1+7nvcr5bAwPi8OnTzsp38UFRUqteL+Mt6pRL
wTOQGSKRn95Rm9dpVRT0p4KXaTijptIwKg6Juvy6oj7hQsIm7VVLKTC/4TAFwQo0
heiXLSzAT+MRgr4lwGo/UtWkMac/HPrVulbH5TVsxTCF/jCqYtULOyjQ0Mgmox7f
Jw/ZMrJQPT48feZQwIUmbFQb7ZBn4TTiuoYiOLygTdEJ+Gtx9TTcCTKRRg5XQsnb
3kMAA/+yDrf+gQwGXbvUV+XmdlWxlBJsdA5Igy0lM+ueYwDp30cUbFjQWEbUtrOQ
+r7w0VYLfh1QqSQ8jATJWvGgE93BK8C14DHeYvlWuuDTy2PJC0KR1TT31X7hW53o
uOKJd4vSTRHrFJuYeSr62/2K4ROQOHDz/Ium6DxMX27QvVLZQPtWVxMart6k9apa
tsP4tZWo3euG1ehD64nX3WhTfGA522DkL1l8N+Gst1aj7L0ZM4UuihGeic+F/3M7
Ehw/HMICpZ/+k2KZ0hokWcPOhw0KonOJoA29F/7yvmp7ens+AnJQV2jdLuwd5ma3
Grc1F+4TmxeNe8wMDGefzQnnqPD9FiHgmwi35MmytQcPsmKm02hcZ7miSOCg03yl
gtcFd/rQUfbBVzW7D6VfPxQUfG9S40+jK/whEtufpsk8SoPn65TSkUrP9wSmFiVU
cyzNBO5mPwALaBdU7X+A1NeJhSrVLpL1SuyZbcXhnqABcsREBvub+6bOZsck6c3G
voxjGqu1VivU3hKo4edeKZBc9r2UmzZZfN/MRuTbcd96Y7lb0Nn8q4wnhXZcWQ1p
IMsx7JkUzt0VMvB5ANHv69KK+UXHzQAxwIyESaq/pzRvAdzg80x1BOgivmE8DKqG
qDezbfsN1rvuGv+VsEa9QEAGJMKgnT7YYTrFkYdqkZcP4q7CbHXiYfPsZkZYBidA
4EsD2h4jPtUqd4Nz4ODkZBrmrIcIlNrHLgNmSQV2IMzykeSflnXZr/TkbAXt+2PN
iTgIo7ESFKkR18+rlNXL5BRVpXARheFOQKcNRYh0nwcL7hBMG0Mx+eHBB/utK8Dw
bIkOtKvvn4lrewK1eSIZhTGZGlFaxi/URJ2clj32vXuxU98XRnncf89k+g9pggmV
H6QaelPyepkAG4m7JxQLJLr2vtFNBSFQLjKsidyvyxrqps43QfzlTNDPX8xsuKUG
a8hYyUUbGp30UWd0TFDfn7ATFLp5YEJKX+T/Z7L5XZekCFS+5u4XyAkgVoMB63oW
L8AQymkAduF5zLqQhtfsr4gfliYUIWrB/N1hEmbLFWNUZ52zlWIbRd7XqqgK7qqO
U0KGeyNwOJxyLubhjBTYNVuqzW0YTODXJnboCeXmHEnb4VG8fHFOmeSLznqB78Zu
kcwR3YaGHh2A9UoezWXAtTMjxCkxYn03ssxeRqPU1WLN93DsE25HEEatDE9OWSrT
lOmvFtjaHGJ9/mTtHbR244etjjtbDNynOzDYbB+VbHvp2rauxHxweQyA9XfWj/d/
ZIP3gcs7Q3Cr3+76dw373Ae3FYTROPs+YPfAxPLQtDE8wBy7+ddToc0lNic65jCx
NgXPSUCyDiPMmR2CBRprDro+iPftmGVsNS3preLPYKPl5PjwEA3ZJocnxcSy4xFz
k+EWE5VTJz3NzbckG8zHHYgdUsZMEhXtKe2i4Jic4CA+UDrd8w/U7H4bWJlWkpXW
Ls/kP4fA6CTspHTgVCqpvn5Kq5dE9Rpu9ddX9juKEs89omfNdieozD/3dbsFdH+u
vqpOv6wHPalGyqHYvd7fnQdBBTAWCQQv4VppQyF/scH7k4EzZ71n0/wkr/45GoGz
YFCZCh47MzPw0UMzG/5wz7lnqiIMUstPUIlPUHly7aA+Q+CHg1jXw94xRVj9Bq2D
bsbfPgCGBHDKwpj/zvzfMCiLECI5oVJs8MPS1+iRkgfpsML2xv5gef6N/oeZdesr
uC7u2xS+4+zlmh3WUVZnG9m6+tqVcwxXn7ckbvNm1Bdfv0Zu04HfknxagP2HNVNN
iYJmFjnDfpQIqxiwTQdfUOJ35HtPQjlg4VnhPHbXz24CC3rUCaIEi1DtBEHEKbGj
k5pCyF8uENn8KF0YR3vB0rWTaSfPT8OQVvseCU8UP02bDMHiE0isOA1Us3FnBXY6
zobKoW59Q8coVgNR+8acdyNuIR2pOxd4Zpe2GNmfeDjYtdgTq+0p+4sIoN4pj8Ht
U2i1FnePdb8WGXM6uL8wetpQAemFBkgWyN8nzDvLB6WJ+3AhbUW2qH74FelWbGn3
pTzQv+9B6dVBEF+eYpVizlrDBVVLl2Hjvpjzms5uXc741d0Q6VO7to1c1+Xwf9yg
B4dspn47tK0RIMDo4a5mrr2VBfFeyWSbHqdb4U/lYH7N3TxidZtwoYAclJAYfL8P
UWWm+C2KVG5dNrffFRimQNr0K1umKV9rUATOvntUNxEQ2P5ZWsgWyi+ezSAfs2c+
H+z4UA4uXD1YEPEZupD5NNT+7yZ6KOKFO5y/ofeIYxpC9TlnTgfLZ6q0K4JGoDd3
xbTDs4n7XhoQJNkgm/SNbITdo9d2EcEquFCHpmMqt/1+U9FyCiAZmIUHdjSxqARj
asjbXdFPZHuR06naPGFbRH66toxbgIPkYCT0VULgXQyGSCLiIPs8pQyJFhPfZIaN
aco4n93Lwrxyxkiylz0XXnA4QSPtErBmrKBYPsE0+VmzNQRFLApGzT3fYFVR3W/b
YoFUAJoxWkiRwIJiBEUgJR3qlSRGE2FVrka2gUtLS5CgnlXLmVMeQg5zNRPWTFna
OF0GQ/EHznTX51vFTkNAAZ8owRDtZuX1jAIZOJ0qBH81VfCP0k6yUHlmOyZHF0Ul
bm4qMy18bkZpHzABD6OLZBORiU0kKVcu+FAMWoD8AFa4Diuv2bz4ko+BxdajeOgl
/NYTqTYXwjN2g/J3gaOFkXLPNo4odQTJ1rdi5GmUIyW5i9DUbSNkWC46DzyDzvz9
fA+aXxeYP7tVo9gix2b6jyq1266+QrAtejxiUDQXErxjwDC9Ej/T3ap4+qEsDfKh
j35Vyc6HQPml7ttM4Qdyh4Gsi2C3YHDlFzybT38Jb0tv+XkJ8NDnv4WX+AtYqgYv
/DK9logNO2Xb8ZYzyfPNcH/PsUxhroudKlxZhHZijhpMgmtldGweiG+a0KC+mykU
D8FDPawnYjkKuvpZ1S+BUMaNhKz3CyOr7iJZ5UTGOyPWPq7/GxcsTKh1ghXEIwV3
+k4M/F3xnlBRtZYWVeVXuSWf9OJNrZZB8+WWnfBq30jqJ6hBmYuxLSHkLvGXagDo
Y2Ievqj7HOtxWk3b7ugPvasJdzhxFkSCEfOC0Ti5LtZyvNMnmRG7/yUerCDTQR1E
kIOlmAE+Fkk9fZjaentPk+F2WGnDOlKTtvha9lFffPPaJQK76RQBjufuKxQc2F8H
lDE+7cNTt2c0uTwIIGy94Fne17jbGYgDMW+8ComBXJ1Z8kdUfrWkq9jIV9isNfgW
a7kSqqH5PN5anyn0TMUpJnRdV5wJBzJJpcCBghy2p83QxvrqQV3igJh7/wRvUENn
2Cyafn9/RjUKrCRh2h94hyun9BvgNiI4Y3Jq3q8gsQ2xzi6iVaKf7S2ORGHzJrlc
eUnjk/pFuLFCf90U8Rxj6OnxC2VkqsTBiiE13BClWN+E80dchX7IAOtLIj62YwyK
/NccXKUjFxML7ZmHXSA8aDD0+rx3kETFGJQgYtcpUVfa8cyhMV7qWPckUBQ3l0Aa
SBpoR8iZK9v5LkPUqWABmehJW1wxGAZKxgMucfRAAHxIbQFi2v4+bCzYeYXzMUKV
T70XqUlcSldZvAOcstwwsJFH6HVpDTpEPoNxpeE7P/zPJ34WpkuI8ryWI4671+L7
iWfprA6o3/BlQp+ihTduHR/uukqTq6tdmw4HSAW3YC2hfuLx29ffBRTz87V2XLFK
JkjJO9eYqvSCBAc3/hmMv+0GAwgG5zss+c6646+p02UNFbN6KF4HJEHUsUQXuP7o
B47mIJblJNPoFUChy+MX8H4vwXQd38vZBPuC5YNwRo8c/9tnhUQKdSB9mlkrGY6A
wtkYykoY2755TCSbTgQ22YDZixb3ypcGqunGT382PAG4CKq+yStHH/EhfK8exuIZ
eqz5O+NlTS7sj5lRzd9t3lYxOXBRc9vhoxlGN/nUImFgzzK1VqgbbWprDW3uM9UA
Qlp6OHkQYpW3Q+NljY9Si/ZzufNopVrN76Ym+8Ez1GF72/OM3PEo7BGcp7wBx4fG
jhzNgTTSLoR3/uNzmFYCvSL4iYZo/dN2/9QpjqH7OHdWhQZGJV/sdzTjYWr7YtHb
Jo1or6XAKMrQYQ22ltZk0RqSExj/ShzHpdVCdlc5AaQDz+mthAQLj7nR4j2UiZth
UqRi3N5RY+l91h0Ee0I+uHL+R1LX3wuml89C35HdijEVnqm2PSGClMhknK/nlora
0EqEd48WtamX8f3HfzYx2NSK4bp96/T4Vv8QNBuSjmXYWublMp/Qht9/uPMlctYf
h/Rbr0sQgXlf1cd2N1B/c3y0GF9E1wY9zQ4sH0s3pugz4BeReD4HdCAjudn9K5V4
GYqGmeQTt7h4Y14Gu8HE4e0yQHbMBIQNcxAdYqUWApNZWB8zQPSz1rBG6mZt0182
WniWp7DSW/3C4v7Cfx6YMcXpiXy7bEJUNLdLYdcFyWp/9WiGvMeluarj4BkI6i2q
nC2wDG2eeRDdwhHkMtDFUSPR9jsoPxFQEKZnP89/okgEPHE5wHgZ4kuMewlpj7i9
RBQuGuyNq9zEML19An5P6xZdLe548itwCzimdxKTxI5YDq0U2/kKY5nWRqF5bnfd
ZDV/qu6qfWDXEPtrRSV1UbHrX5hArTQ47xAY+ymZRu34EYApL1bfNULfo/KtnM1f
q2pNdqnvBAXk+D23uNTyxBMyjUrrpyWl3ylt3/sYRccHnWhXd4cuFLgKO7xTyFTu
Bv74Y8WgWN0HbN0dPGb/IqVRYRHW9FTzij4PhwxrV5ros94iZt+XfTasY2dBpsfO
e+HoMh53ewEZE7c9dBqOrwWpZK8PV6uZa5lKQvc7mikNt8qy72ycrlJyrbkmvhn7
Zdr0r4cSftgGdWl/vIKIlaQjvc7Vm6xl/725JgDgnk2kLNAN9HhgZiIPxsAvt3dG
7LYUrqJ5SCyxZjPuYs3yPVgXuQ5p1Y8wnFfawgpWG7q+vOEU0r8JL5QTIywwqrUx
drKGNeLej0xmMzk9TdbqpHMKb9rRem6d1qCTjFwcQ2R+IoiY//bViLwHi+yIWjI3
m5Mg4Ft4qflKiZq02o6V2+XnD+Q4SPa8efFa9a7pvTusEPis9lzCUxHWPcNbdlKk
X058cvaqbP9KEs/JdjeQzBUNPoTaT08FlWDNK6WjUtqoJMAJJt7lPVs9mJatN11R
S2lGlwtvfaBUVZNaS6Jrf7XnmqRAUQ0U8JuK2lTfiv/TGqLm7j8QA9Om2nXyYbMe
lrMoI57ltmtFdCtwOcZZvOhke6690fSkN+dAsFRIlLmNjRpRTfbbmf44uPXzcaLE
IMQbfLNRNn3VzITB5ze/RDDR30FCWDroH3gMgj3D/AE1rLelJqxGbA2mELm0ah6+
ZgDXLkzpeV63KJZNXTkmyKw4rGmjfuqJ9r6qnpltVYx1WxRlAYGIMKTF9AeYhPlq
CWWnqh/bAEHbPmM4u9tbhq2Oxn8Yvysuw4AHRhh0BnKKeI1v0L2vjytFut51WT8s
e0kojCWrkfo+ViNyQ63EWtgxd7PNi09aNbdEnDqTErdLz24SPGEBz4K27Z7lb7xC
IDutNgtQCDq4/2em1mvI+M14y4YJuExqcGUrl9ZrMuMkQrtFiKkvh60PPqKXeCQd
H1ZdkxVjOyQIWw66AggqqzagIftrEI8S7xHEr+yCl+55XPxBzX7BaQad7jm2vChl
X8ZxhIFyh8VHYFhXt4Gl0g6Np07PxnLab1839ira0HoLwsd+AbMu23OABx+vs8Lc
GNPLbfwSZYaB892yEg3By3fGHqiZNbhIxd2dwWXbllnzST2XH/PNXHbnS76grbe5
juuHBNin91pxbccG09dc06IVogKCo84Dklxy70Utm/TDr+1EOs/MY+8EPi2a7gi6
46I4QBzHU1CzXrhkdOud7CpHywpaEKT4XxVUtscGU+d52hy6iv9zYH1c9vi9Hx75
En24HTBCRz83yuMWyP2yCxVAnyfwzPoeCqIbofI3rTbcUv96iR9pMFGrTzRzYdvN
mhEidL0Ofo+X2gouMpNoWFZ/oPySBcgSrJQmYyQ592esLVKvR+CWacaOqtcW8UDG
mhdS0J3Vr1twD5BcB2D/sFDGzjUwc9SpOrariPPI5RQshI9gIfVwhhUoyTFmIVV5
siR3BeV5AWm1W3sIOBLhzDuafQ5rdsJSK8E7HnOp3hLC0naRe5tMdp8uqGGVXuWk
FZ5CxRKDE4rald437adnoIqZvYwXBDiSKbCfq2/ZZLih1uLSt8Hm63zipK5Eiezx
7ptCwAN7Crj3Ux3OcEpSOWZ63ROrN6d57CDqsbLxPmRJWbzE8aXykLURIlYv5nbT
zNWLvDnwkaM55NJq+CWrTW3T0ZuDr7k/x2gw9YhTiFOlIvVGMhyF7j2QJ5E+CFJH
5tM4DnoU5S4DYttvoK+vJhCKqDHyUTpEqRZojr0m/uEVo3kwB7KydP1WvBOhSKT8
1MLaZimWzpvd9QN86dE6DGIbqaQbDOG7ddS9KkyNaKJGfh7pvaF7QnPblpFYCNVm
xGcQWZvhEqKQrc54ifnlNxC7OHCPzYOCHagyAxPxQvnVsuzBbDH/+t6zNqLoVGLc
jnppHObmxEU9HlquKPlq3YXoCcNoO8DZQqtfxtAfxPtZiVZjrxHZwXEKvY/2UVvt
XoKttO4cYY2KVf7HAfQFUu/GdbiFmvrIO1Sce+k4e1xiwYDCBnb9xUeiTMkRF4/E
FTKmhkTVXFncGSbOnm4cV2D3kb1XA1EOD00NYQACFCn0BooTk7ulj4RFj0hT5Zuh
ULoJkS7WgQGx0wypGlTj1cKCUiWK0gSeyF+6IBv18qBhYTqt41DotZq10tjNT706
uC+1E1WFQIVoFMCEmUANAgFIvbODpqCG6IIhvKcPw/OlVzNKiHCHESyeTZVxpVmW
k9fCAfmLOaYx5EAhbFgZhnx0Rr8oN3BGKZB3iSDygvsKbaaOXgZkAkHXM9elwMne
Z4AAMsi6ZOZHq0G74k7Et9AEAk/D7JVwXuCV9MVfMpKMAu5aZIOcCAKylOI1OpUE
tyWJR11RpD9IoTCKhEBH0mLKjJz77yCTm2YbQ2oIzTIuQ/Z62eyjCDyxx+fvoFEE
iwjxl8rphOJvDr2m+qFHiLoF5PaWIbwvbDfLd2LPAuH8PcJejBCY5PTpBvDg/TAz
peQNWFjTh08DYMEnBN0vgY/bz7ePp9ynxoBjkG1KwKFt0XS8VaiTQSpttw96/Uho
5inwAj17f6MoRnxs6kO2e6AHm1WsaXP3gnz51a4Wnex7MfVJKnKc4eNukBS/7HHE
3lkcvytk1wXEnLkirShLICxEoSOFJPXDSl5otvhWKeNQnwk/qt4f/FjMLW+AsPJG
gKe0qPS6rTsQnOFxTNY2XCqfD3BC0U/ZwmnY1VgMZfltmRxHP/aYzeYJL3eZnVRZ
qjvvKdZLCkTy/8K6G7vO+D8/uR/ATTvATtr5OUDlyBfnQni5q0JyDgpfBX8HL8wW
ioFA+KD675YcvMqkvBJRSxRsvh15JHl/KxqI3ud7crcaPY62tK2ODnKr8vzFWd8C
TTqOqh39XHT8uW5TAqKIJg5pnSGxrZU5LZzLbOqROXFJHQ4nXsPep6N3g2E+oLsQ
4n2b6O9bnPcnCmTUPuq9NNr1/Bwg3WEeNWiV8OeKeoFhBhzJ/LJUo4dl8EQfSaYh
iLj2qpA3qieXQ0zab9dinK5tA3AoMwMSE/DRTmaQjpa7mFLQAAXkl5/NWzOyqyUj
vLBCqP7Cx8wuvMyYlDIMUsJIlKAbmA3Q4ZtDNpAgHucK1uhdCijVuMYilD1wrMwK
hW8TAQCBsFiRYN/HpxsU/sesCPLd0nq9p0+j+7qSYHZvTUhPCIzkv+6tP5MyColh
p9TPEbpfebYMYED4wjjYG5v45Q1k3P+BbDmQ/E9DG5ZkfiCiMA1hZkfIw9obu9XE
PtnDNUxJwpKLy5QcV9AC4k5czknsJMzvM1e9fVsuIPom/J8LA2+w2Oe5IsQj4qmc
3CYHkmjNvpDV8yzrfQp48taEjJA3ZnqqXEY1nKZftq+7a+/RnwCCfb/BzXDMDWkf
RSpfIT2MCFBnP7qitBj19jmk0T9dpEFkwDdU/vZTigS2/932NnyAHWWh3Th5AEtO
SzElwb+5/1EuCcrPe2nsjzE2+7xBEtjWqoXMYnHuHOVkQN1wYd8pTISUo+GSw54k
gGK4Ub4hYKAmab3Swy7+J3+IG+PdsLvUYlbrGI62/t8AhvIie2T3tjoGbEzDTB5E
tiNYIXwi9beh6642e2fzP2aFbaBRPfGuyKLCTo0VPqWOpcUbNoeftl6B3cCtUghW
BE2VPFCfKKLZtrnldBaGzfD2M4Q1pW/YZeDZDrJvdgCzFahHMzfiRNUldloVrJh/
eflFAVouk3g0PhM/+Z3U3OjNxysaxXMnhWPzadF88WsbLv7XRJj39AizJdkmJTEg
NjlSsTjUGAr0VVPlqgcS4NlFLaWUJk7Fp6VcSXMNCzH1SLHHQGVSkcxtSBxBa9TW
ZsZ4T8Qf8PXAf6W4NsnCG0snqA7T08a8cTN7aT5Qpef4h/fK9Gmms8O7+mQioczv
h7Q0paTBlzIbnfiYCt2VQ0OZKWc1gYJ4D4tKecZehtNORMc2SZ0fs8+ZrECrveNZ
iYv/5FUA7XsPCY2oVRkme5M0g5d8fToTWmBDhefjWLDnclDwy5qgmCZmEfqfu7Io
XJ7jtyHLHQj2AwlYVTXkgueIUqKd9kvxqmbKspCXc509Z3jha0bxKoMkZHS5Du33
/mACvZ1XuoPNpTcN7Tsczl8lLYWBr/hch8lPcA0ing0ArLm0H1Nl7pmMisHCa4Hr
nWsFHgOI6rpc6HxyI33pud5Z9fgzIky2sY8G8BqyHWyDbdjddQrxSLIpSjUP0YdP
90FC+sz9I1lilpHqS64jlfb3yBYUm7FXv4yxZOqCDG3ut3jT8m23L0HCx6181ScR
tN5TGvCF7N09/zZJOraRGzKGD/bYsymdJUPawhhrhveU+5JotN2hG+plGe6coSkD
4ITmtWd+AP560iTZGD1Rlt3MYDZ94VAlTkou2b3edj9XjXGXDnO5YnjwRB/AQ9x/
aDJGJ1jKNdBABx/kcPJAhcYPDA0Mh7HJUNugJ50zKy8=
`protect END_PROTECTED
