`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lANckj5WAAWb0uu+sYP5mxHNTY4yXKrf7oIhCzTDWS420YiFAu7yWrt0fsrMIka7
+wNpZYggkMYKBrnXM/daw9BF2efeWbUC8Rdm0kArZW2ieDvbxoEv2Gl3MdgD2fWc
8JqfFBZ48lMEJKMg3zFgJ9Zr4XY+zUK+ApCeEor+iStVOI/4yXpJdPITMF9GZHqE
4aoSfFhk+dTqGdQePoQ8LhMNSrsgbVcPd/phyzzPpZMBOoNUEfyaqLvv1TvAaw8s
mu+JlblQmXdBrLw43VAhXYKd94u8Hog1UORVAV6K9PZglTQmCnRoqcR+VDyYrUWJ
LbfyPro6SKvj4DOmMS5IBAOd4hVCQ0LmbfFQkQjFi5B3WzqLkf5oSBHzdf2YHyLd
+WZndVUKZqaoY5QESNH1mVJnaJKsKwWf8agsMmggUekIaSD626vwaTktbDvRNmfB
Yx7cLXqCpMMn+DoEYmVfiOVI/o+PIbvvkZJ4Or/X9WrWFEgHwVrZqmdCihCqYwaS
VnYmAlxhbd2PsSbYIr5OeksG1n5fDQDLPsG8EEbIyfPafa9U6eyOD/NPKAm+2JT2
q0ESk2xY2Equx0JfWHpZF/DWXoWzq2fOVltDjeDCoF4DuucSIkxKjWXTF+0pf/mE
52k6d2S5lrdZOMkG9NsQrU3YaK6QIECLwJQ6aYiCVweSXwRTW3/FAgvkJYw+p4fd
`protect END_PROTECTED
