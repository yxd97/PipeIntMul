`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/U2Sl5pUEW4s5E7ExLCgGytNC+ZE4JbSvKBA+ZI2PtUSl70lXyaRtN41Nrg/Xpa
FpvVkbvuYlibl09sFqUeYMn5hOH9klSew4mQtzhdrVmWekaOfNDYrXTmC9tjQ2kq
btBhok9y32nP64I593XJhVvYfZHg7CftdQjy5+pHhbcWyZTacer4y2pxjYQCPL/w
uSpSYQdqWreGBK6REuhlB+S8ZH67Yr6GveSLs05sS2RdoLxhtEgqikuaTvYQJLwk
uchXCu5u+UjyLp1T7vwhIbq1hbAGo359UpHeydRsLHMU/By7BBJtL1j30vi0cx6A
mTTQ8S4j3Y6EMc89BZPYtR4jNUw7Rd8l9dJKiC5ZXMccZyb7klffp0RzARYoOctE
TMpjDBh9+7Ez1Dnmv/NNScbTg7TG2GI4iGj6Xzmv7twNM3FxQ/+ivK0QSYBrvtP+
8IltxNOrnvGFegnp4T7EyTAcHSFFtb+q8IEtA1Kuk33Q/Vy9EKWIPpnmDfPgrZn7
wYxQ5dsfDL0iRNowfuBnJNVYfn9qe9ZwaSFofhKqdaqdpIWq79kSX6QDvXflkxp2
yABvsWJIdFyE6xSXQ020y8wJbGyL5HCU8ZLxsKuiRMflHosuax71spNVsFj0R0A3
Q2oN8+FZFILFFAKGCmH78grntflRSpj0N8IRYsqHOS2A1crHxQQsk07a1tbFAvsZ
5/47Q7N03YqTH1Dg+lDXYiSWTmuSjX2ldkVWTrfAZeexGuy71nj0XWzZk3mzrn7O
x6U+Pj8dVtbS5qOSuUp6UxKZ3iZ9FxzBg1OwOXCvPXTpERfrg1TOMVb5+lGrXBar
GyPOX7Jqf2cdorQjp2qlE33eyAEYZWSKtpVK6+gNkx2UxCOvA1zYtUbVR4SKVxQd
CanpK4gcsoF+Ic01Drt1xE2lOq5k1DDmit1M3I8fDT4R+2b6C4vHKbizbJG3kLgS
9MCVprFTXNpvAdMvBDu8VD0T9NxNw/oORxRMjj6058enxio1H82pJB2U1gHIvTeq
1Hq8LCfcwVBRAcSWJHdjVqIcmDOnk7g/qkZD/PGjFD2khB75hPHdKiLL2aEcLDQz
cYGnTD6onTrzVufkd1qxq54ulr9kHJYOfLj3H1sfLC/aTAJJaHsAXkVF3tF0ozaS
1Nkkv/IwNu3hjpXdtI9zO52cZE+CIo8YGHCIexalqbKEeeRtogNySukfhApJJ18l
JfhpsW0mo4Jk8x8oucHPs6GshgjrwrN3epVi4Ynk9W9nZgJOmnVSQth/qWVxuzwH
y3+hpjCQfsCNBGoasLJD7xbaJupF8mqOmpEpo4Bb52lG7e71AqlZMbntIbUQV4tN
K4R7LJzXCrWNy/fBRACohAX2BePHmDglFkGIgNWEoi2bUsAxnvHYCmC31WcvHYeL
EhGZnFinbfviiiMGrZGiDTfTu0SMkd/l2v1zA83NuA9aBpAymtSGMtuOdCS5gZSu
GslQS6+uPy/ThAcofQIccHYbnLRDTV9ole9FHblqbYBXg+dP/rWzl9mBNWGv4qQ3
AwHwIt6NcjGhY9IOCFOLYQbpt/mXzIi9U1ZWy89VingQG/ewFCSLv4D/DrEvG+BS
SbjdosPNVoBGEeD0dI+qIa+viySmyQ584D+QKeOe7xdZF5zRkUZOHd3vy1/JTxUU
qSPx1U8HppBqa33XmsgMe4R1R+Jq4/Lb+F6BRwdqbsv6L3VUAb1/axbWdkEzENeA
wD1Y4cuFHTDF8ETuc23TLs9RSyHRkasii9uQv7CFRyIJiD3NrKDCkVJeJfPMzTWz
fIabPRJKQ2+LObYFd8CWtsLPsXVAQJR+YaopQTBFSm4AUgYfer4mo+XAMbPu03sg
fbiHDMjltfpw04wMDI4CcbAeI0TSjj4Yj0XP7zlB0sxO/JoYnpUVER3VLu446gTX
wE7DmsD/Dsem4PRkFpebwYGEnZMDF0C3RBOzWuVAbK6Gz/0RiNlgoDE4UZGQji6o
M9bTQqGe+7CqGDUs2feisuUs/X6nPQtQiJL6HkLvWs7hILWjdvm2aDRAF1ACwvkh
UJCHjwS/41yKnX9/ClQti464e5CihFh4xfdU+jdtJlU+pYu7ZyG5S90kY5dX3sb1
xajV0cxCoOjhn/Vmc4rSEgRxv2rEaIJCuhEqP4OdBUOHyKcvpbla9DvNruM2LKTR
xDnOwLX9udvE2c0gyBGcSTuAN/rweQexp+uW6pV54D4Q9/WmPbuKrCMmEfn/ir8W
X+9fcK4zrKjSwjA9wH/ziVoncOoj5L01B0kW0B8U6TJ2ZFUSnwPApd8NIsngIZ/v
DW4Io/nNNYD4t96ZwK2C8tLKQG3phlbpgxAb0+0eIGXOnfohMYbUL3RIVlMmxwvr
J3uVs19+ko/WKsMO7j30bi3XIXptkA7Ay+0dnnhTc1DRRxD6p5Ec6aO5Jdw7wXfF
4htzRUEg4DFUEYRJR80rgaj9HLMGU++uzFUQvp039EsGMX858Rq54Vo1iezo3Exm
dbZr+XNRZ7J8XuT9wg0kB18NZLFc3sBcXYG6LFoV4ADrorkPlGoT59N9Ek3JcQcO
TV5+ecwJcXJy8YP4zvOnm/LIFpWlR8TvIYPQgbTBzmCTuGWJiO9zV1X+2G9U5dfb
AI0aBFPSZPCzp79H9OVV5b5MK2bPtFxommtJIQ3Pgbf42aVIlYpiic7KZ9rnyV0y
FSOW0BhDzqoxUvT3ec9C9FC7s7qWJpKR/a2N9RMY7FENwKobVuc4HLUclFR6VZKF
Aon0OoPiaQtLxE8ekSBmnGglvquSYErVMtrGst1ydtTXnhh+osIV6v3ENggAgdzA
YAU/ryxzvSTZDWBsTBMnIkyBvXezOUHVS+4JCafUtHRxkeuDbDEDD33YNl9ALJGU
Cd8lL1OFlk9LjwnH6oCMz9340tLAxeDS8qbkW2TecU481cKpBZr/Nby9CWB0ny2L
XsXD5g5YE84uAya1jQaMJ3rOgrf0rP3ptvJwFsUx2nMW2jT2+KRYfrAPoJONrITx
0ZzY/3F55HvLXPE+JkY05ehBbM5X9USijTIqh4vK0wpXcu7ujjzPD0taQUWdZTdj
Tus3RjqyTMfyc8Qb/tIKxuIZNNPmzkUmeNNgb6hzJq/R6DXBJRgJDis5Up3z0VnD
MDItcFu4Z7VZCBl/5AaJsgFI4gt5iWc2QFcs38jBwKHXRpFDCE0dWCMnYL+3II2S
VMnq2MB8fhw2SULM8Ieel4AA8Ksig0j+WC+zEYFjwWzWtXwiIMDtBv2SZDifF8f9
DX3bYHtaLcUGARMNzEhqdVjDlvZWw3JjWO6/FJk8J1ATd2h6jTAvtQUlDetKs821
E5aBj6W4I4QMLUypxSKG+z7aQTJnkGoGdOns3qcPYvNj2kfOQPQYXtPlmiyPFAV7
IUs8vGq/UfswYKB4dmXJsZ5fIAtNByQU4TTu5WzIyo0beclWNujRR7DwuOsotZto
NsP4ffr+QmIEgu8DFue8NUb/fmbI3WFq04DfhnRjf7M7Q3I9YZWIstc/pF3wwUpa
tK7J21yGnqQBE7dx9Pt1nWI99ajhgwm+iyE4y+MlXN8=
`protect END_PROTECTED
