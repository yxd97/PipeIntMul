`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+oUVCeX8fblfRLqG+e3sNMj+Bvi/v0Mh0JUcdeBYAx8/2qtCx8RwovhkiiaCmTd
UCDuAfLI4abdpa63s+lWjux2hixONnu1lrd0G1JqqW4I1WcRPt60/xsBFbCt7/Kd
amYDk3hjho6LV3gCp+I6F20NSFCTpNAkmncJ1o95O1w04EA5aqCD31UucsjrlUyL
gnHuSx64Aiqavr2OXVFp0L8t3zCaXuUfudCdPO4+yVZyPSTMD5u7t0dS24PqbOWe
o8rrmsWUNKgVNW/Q3YSGqTwWAWOnxIkpvNjvGiWxOEdbCSfqgtZ0wGkmI05PKHZE
OudzedEdczpU4DHek6DRpGv8Zx8tykc0lVxToiwrzfSTrqBH1jy96kNeSf0DmzgB
gebCfSq0NFShao8H5E4zQ2JcaLlJHgfDjXZjY0VXJKtk7tDvJddbCXtRbujJzOuT
pjUKmsbNFkL2USvwrqvwNFxcs5GJaor1b6NNaysQMZPpV1u0zj5i9mAeIC/UlOAa
sXNQ2qixXuQwwwNIIolBfKcPyG+vO4TRYI43wTTB1OdPEruqCHZyecJ2wGerdX1u
uwDSE4XhFO8dEYoO0OJu/klISzUoL2SY1aC1JTIFjYoYMUp89dWQBBa5OAw2IMun
J2+FleeX8hEke0BKZOw6og==
`protect END_PROTECTED
