`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6xIhQjejqDxh4D+xCpGCsSVy2JGExONJvgRLj314neZ2AR+3B0GKRwbLhJNNP8R
670UO77fsuEATmSJ7b5pvDtBSDHQSoBO+OGG2LncrVJS+0Hifi1yF83cfpBRZW7f
SZ8LYPQuwDX9d0Mtdo0NEi0VxUpc4Mypt+RoC4QgCRjLuAJ0v0spWCIL27mXNYn0
zdyXkxFfZWfTDjwDdVrd6jRjMQoQOecRwwejUh4vRAlgq6srthmobcZ9PMSa0FWm
cKW0W6Wlz3nAARtp6gQEoguOlgl8KKTfSyR6A6GjW5vTLJdHZqF2CRWt9KXQmrmJ
4j4SXdCQqynKVLQIulZPyLVlTaM/FosEPIp7FBi+m3pPL3xX1nwKuNqW4EfJX26m
YPKOawWyFexTI3dy9H15yxq/3CbBArGpSdi6cBLsO7N4qP2b3JTp2bUs/Zk/PZfQ
B6SqY4bq9RgDpG65dlH5Dbw5uQC7fG0oTn6ELyaLRxYD9QRGYOBtxf0XRw0k288w
n3PxoGnLV34Ps+p/VIINQ0Ci4JIDTO/fzJiMtxZpYJNiFBtdCLstFAlvfNvpEtaJ
LiVItTSMgTyTe8Skj609pGWcpMChVEd3yafEeZCc9z7Pd+gRpCmi4hR0NpvvqRfg
vDhCcHsHfCV26IjnZ8AnYHgwIsT5wT/cnZNIH3Xu5N9WQ1MzpqoCziymZnCQRTgP
PiJzgqNNvIKDm/hHGyBuL6uG6CC/3zqyC0/tiuD3ZD3NSHbBEXq/gb1owVkwN4zF
F0+/+PgK16ElTMN/BpsmAA==
`protect END_PROTECTED
