`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LoVx9en9fAelxKBIzlHg9fJGPt4vUKiuMjjgtH3Zo2p0Vc1z7DnGzY3nSJtR6yQ7
eITbA7z8SwyoNF3HEZp5pVuWLfJEUKxb3PYrEnxFMLa3d/PjzobajJDjLPqsGO4a
jhsVKUsRubJnmz5BCKEMZKiEfI+d+Muvldm74NCjnBZkBUQoJqOCcs6Kk6+9K2T3
HC3NcF3j1R1XM3NnJQJMq+jYXF9W5kxJyh/XfZUc+dLXdBtPzfvvfgkTQglFQyKV
JRyimbhNjyt25RUT4cIRt2kM0nc4urVy1cta6YysjLJsoHar0FOAiixwDh9pYZ6K
yBpunlN+Y8dB/5FyF1PC+lyGR0aOj2527EuQxHnt/99uEMRGeOSIGzLo/KzdgcMM
Z2Eem0pkmKrxGyMHxLKlIKlLoAHJayJriXOJmHz1hXg4eLyZnwy2rJnIIQXrW3pu
uuumWxIyBBUZOUmdh7kbDvCPPZphLvQGewvLgrcsulw/moHZNqjQi16TCX3KSSNO
Q+G+74y46Qi2RtxVjyICbSrrNNqvuT+G3sMNEVBVuEzF3/YM1PhJwsM6Pjvo3Ap8
pe+35byobfqxyUepn6lIAXZ6qoiPtedC6Nv+4+dphYqZHmmciUMVLPO2xnL5GWzm
EQLa3cUNT5B+lTKBx7yNE/8Xz2z70Q1iDDLw6EOLTGNIPFM3qGXL8+KHf6Ttm2Gi
l99/PcO+RWH7CuNFnoe0mzHR2TlUYuWRM71jqSN/QwzHCXLHaF65gfStRoOpxngM
X510nOHT07Qwne2IRC3ZjZtS1HJDO78IiEi2lJCfUcjKxcnWKVc5qxVgYOUfa6MD
Z6u88PyiCDtbI245l5Ivg/qD7yrjHsyeXrS9FAFteSFdDRYYnCB3YJ82aElzudj8
UKwRFoSjhjQSgK90Bs0vkM6KoeSnQ+Kxr67Ry2FPFtw=
`protect END_PROTECTED
