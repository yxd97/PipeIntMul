`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QN+9O9k4k4fIMArmAWbIe+yaF3g3CVM8dGgAMQM2sjGIxIYXcISPMqhJ1D/LZeg3
aN77+1fmATVg3Dlg9KelcMR2dGFOx3mZSBfsXNm5ioKLoEXmFdeQKHB9KMSVXdli
sQyVD5SAYSTqiCl76bUcZiAo/54XPpMExJg/9g5U0nw0kGda6s9eveSf7WBCyosE
vY+dWEAcflXmNA3xrgBCTUtaV2Ct5sVWPcPc7d24XVNBeklthqpTuNq5B3aIJT63
fFaQ+5A1uGGh2PZsX29UAO89qDsXx2AwA2z1L2UJuWcMxNp9pSS8ACc3pTXGZplc
q+W6RzgSQBNMJVusHm1+Au4IGxFYhzxEy5ZcpywyZwk2uYLg9ZyqOShjHlSDdMjx
UinsjpHsMv2xK7nSflvg/2zUHgliL8ivPlFNSFxxY1TtB6s0y1XL/w+XEdfNUhSg
+XqNn9K4ohLNlShrBY6c3ehzrRvofyrQqw8lHVfU+NtF5659hcIXn/+IGHbQvOGg
BA8KYIr8NREJByCMAgp91Q/UATf4uD+tjb0W6IRttNeUyusSgYAo/YalqlXDEWmj
LG+1f5tMFV2Icl7RTGX/xw+4s/oOCjvmISy3VaGJpEJ1oh/MHhl8H6tJuNvufTrF
N7DAD3F0ra9+A0lMSE9bNPZl6ZMMuWPOCX2cmtY7yme4JDBLSqxxDqIY1SYz2fkg
42zv0fFIam51dsmI9mlme9r2BIRoAZPxAbm2tcsGXik=
`protect END_PROTECTED
