`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3yBaAhNCyHXUohnbDN5b7EzxTBB7Hl9fgCxa6tEn4wNILbrQTeRP6D22HXsWF7X
IO4+0O+tfehXs6VQtw8ZrXsfWJdU5EzABc8et2Ouk24w74HKazGPBSzNjUpt2gcI
pMO7pTYlEU4qdmjMQyVrV2F2Z3mZb1a5FVzFAQM1D1/ihMIqQKVKou/IFK405aLW
Ih2ijP72JaYTbJCNTpDOb5nkQpNLOI0sWTqUoh/+/lP+XSDVK+9krY0LceOlh7dG
YyAA8irda9j59C+zHiblpmA0yiYWuOZf5fv/dwLtSRPJ3W9fNmpJpnHR6sBgjFho
A8sqmFDso52ai4xfgFPp7db3MiVxpEKvA6NxsSjeB0vvSIBe0G62DZWXS7hUXJCV
lWyLJTeFonWlXX2ltgFIj0lDOktyCk4YG/NnWNX3O4XYTMP2XYKEOieuRBP0yZh4
hMdnJHYgU8iKZ8R50649Lik95vgUaDW93dE5WOLLViXz8RqyarsrXs2lpLc6UuOt
oPUxT2Xs7yII13DdgNiUvA==
`protect END_PROTECTED
