`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VqBIojD/O2bcMRsGWbH9+Wf4eeTba2BoXsUKxWxyZXmveMjZOX6stvil7yZ0sjIt
mf7BvXTSzmbKjfXxfKubjDIQJbaS3CdgndKNtCJfCPbyfrguJCOWMQZY9E1p56zu
XCUrDAb8hZ4KuTKjxDZqQ4hXWyxtbgsIXWMH9QI7oF4fmmBKDCh7VNWkI6m88Sne
/MVJ4YX+zkqfxs+4tbMd4WyEYh6VE30srrtRFN9+yIyRSEry0XGigFaAhUf6kQvr
MCZjvt5U6NeC7BiGvmxtzjJhR71kARmfELnQCe3z+7xgl7ryqcfscrMlljw1CweH
bIRlm005TX0QPVH7eHlF0Fw5/MrXNPH58uiIxXZGPmLRzjC1xF1dcOtUiSHSm5cU
ZJGigC68OJLZxZL5NmdqLbzrPtiQ6ngpf74xDB7UiOZoteG1LjtlxYcT9Ax/gPN1
g7hz5S3TELpHPcK4D6af/2g2icmK7Et+wuv3otZ9aGbIUOWN36yUXFy1Aq/NRySP
T3wya8WFwCRcMnlVFsmJH0+vh6ULfVZQVGKVC6XxDO1jSOpngBu0RqIl01o7MYsw
r3yas0qpjbHre66LwutHZEoXpQCb4D7cy7aSZ0TH3jD+/PYL3kdbHvVG2DJwelI/
8jyhcsN8I+JcI38/byb6wBFA1A5pd9uW+EoMdHe+Y6kMTMfKlSZV+0WNvRMgOkYq
kG3hBZ2HHxfw7DC24GpDdJ71uG0XXBsoLPsclJ9fnB8XDrste298ypS4AMU2e489
JdBLW+Kwqc7XcParWaG/Xg==
`protect END_PROTECTED
