`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1oShjq8tR416c0ToZYX1KF7w/3NFFz6rklWVk6FJiLbY6asGDh0j9CxMeEBXqLWH
nmcJKnxLkldOkdSAD7bzfGQU38ahYDuPII64++M4p683XuzocHh7PXv3MKXzwQqe
suWLjm6kh9q4uW4iJt0NYyGCiVNLXf/EoC7am4fpyvNHqzsxdmDkZeGzCMTf8THI
jTD9GzJ7sDcbb+m1CBqMOnu0+ll0ivjYIChZ/0gz9me14nFeeO6KsMvGDO/Bmb/L
RkQZ8r1poJvbfSTDquPFJ71/i+BSZ0+vtvKJXG1POKN99jCl38hopFLf3pA2zWQE
7T0iwv0sIvfWa75mpVTbesLTerC8QybpxoRz/l//VEWIXpxn/1ximQI3h6PV3ncD
4iEQpviDZ2QEeqvt/I0ETe/6UoYUi+h3cBP8H/eWt9vpnTHaRO00/iIga0Rk/aFN
gh88gtq1MzXIpDdeAAnHD0hHrioycz5YjWmGRX0G9H/ecCrNRGVQwvvQp0GwiJNN
77CsqVbU7G3KgqOteyWW/lkH3jpxJM/+zen8ytgFCIXW1cY7fQ2O649yrrVgnL7c
X237L50H6JGoWr0S6Lwy5X46C/mZTigjXieiWjzle8DVYqw3PmkbAEIHDLIuskI+
IzgsYaAF38S4OKGXZlqYgRF7icIqjbGcU12KjJsqOTXwnC+izEzA6Le4k11r+Pzv
4n4Npjxko9RzokkLfUs+6OINImQWSjf3RQzA0tneD0grAKgsUuTwqb4C94AXz42R
HG2X/kqSzp7QrUIHY6LzKyg/2LhfNelGDHl/COlhTucdNGg6J2fPYgbUeZukQdo3
`protect END_PROTECTED
