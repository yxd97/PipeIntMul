`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6M8cP3heHwjvLNATvKXMX5ywam+bOwHNzkKgwBBhM5o5UWI/wH0/Y0C6NUIWi2Y
pi1wYATVW1RhNAdpXSYUFSt3t+OHPpBJiWdgC28fUShmK8b8UlG9cuX7fbhGJsH9
Mc4TqU4M5ITagOQ67A6kTwzLppMidHHzK8jv2y49HJl7FaoM1YTVnMXV004P9B8N
8fjCJz5KLyT9iFqkaSnV6ccy/RocpzP5isbqvnDr99gezpmH1CsW9e4O6+97ZcpW
auxp6f7Gx5Lb4aHGnm+B5QgoA6uDfHMKA9YSbBY/RIGylrJNRzpMomRYP5Z6D7Ni
rkuztRLAflvUbxglNc/qbtizH1bmvR6dbyTAtbz9XusNlGforxhCL/LjTo5ktiBb
vR6FEqv0JMY8HhTN7XjCp2aD1gykN242aGe0i5pEOUbOk0zLn/1VDNziYA329Kdu
UORQ8TihAfrYb71rFPhHA10f4eiwQvoOQAb4bpCtBHH+7rTfZssz5iMeQxWOgayK
pKFj3s4rXsSEBf6DpWO9GNBDSga2x5wp3BJJgri9YXafJW3SfchxpZTExT/ChvbR
`protect END_PROTECTED
