`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHuTwxivBUo3nNdox46jh0iT51o1qFzHRC/bhh5MSP+vdY6Lmz2lkT/VuY5iJm5a
8x1bnn9n5Osn70bQZwk0yfkf0od+bNRPKbh7wz3tDosZlRhuC4J+5xBb+gHimxF5
vqtA1JESvE3y9djytuaepX7fxMT87ynz4iJrot8q0vJxsvQR9VA59epArgUAUs28
kRNPwjRJyM5KYG8wjt36v2S5hPxvXjJzc3pKqE0mBDdKTx7Ig1AkD3KPT74EgbTL
ImS1WD3EpHXVmnJ7/akzPETL5Df8bh97STOD6aR5+u4F7RRG2luhVPbGPlsvNKYl
bVE3zkRvlx8rYxFNoeAayi6ME7I5EdD4mlGlTWmySDLc4SkPo667yl5gaL9ihobn
pDVJ07Cyx4P7Dn29Zh6aXEvZ1waMz+vpvxD5YgV6LnJAy73SZqx+7Iz8Q3bV7ree
xqaexvj+7fyIiwojWrs7+1Ypa2re6PdBOwQt20d49J5JvKzL6foJ+CuGd3vF+w3X
ISBjV5Dp0hmkiqmnHjGdG1HF4TL00vLPrynVkyyMDTGhsAWofhtciK+4QCJApWLf
UwYQ2KY54SnqddForK5mYWuTd2arUepnK0TGtdv03EBRKzn7jN8HR8yVs5k7CkUx
nyfhWtRBWbbE35L6PqEIvAv/ZoklTjyx59xRKBR1gzPvkWHhnXol5UyCuDhPVJ9x
OuiemRH/hbFG3lRJHT/umamHS/BqiF9hk6OozHJzDNm46j2vSFIIxyCY6YBjVHBT
AkBsB7m4uCtnmaAIBLgkKHIpBCFzLUG7J85zoEGQtWnEvCqrZuR/HSecoaw5TlrK
JsnOd/BzMjCUwKMiRwJMBSJum5dbmvHmbJniwu1DRCD75TlNItAzoRul6rNBQVjO
rSXjTuAEVDRZT/b7JYEd3hWHKkERhfU4IM3qiUqiQm0vDUrwnDHmLixMlA8L5g83
QktSpFyGK2ksPXx9oBzKz6kEbOLB1wPwuMlypYCPPY2K5Zmz4JmqxssH79Ro2jrk
ECNOlVWYaBAa8gnDz4mheH/KYkbhM8R5kdtN9ZhxeW+I++bD/lPeUoeWq8qhIPGv
PV3WhsUeJouTihpWie+LD6yHlO6XuQQ8oTkWq9n+uledmtHF9S4FJf8ZkW3rBA9J
/xgH2cRuwGqmDcCygMCURFpn/hxgLfLyRrQzaUocaC2NJLZIGVXa1+VsvUG39X/1
HF1ajt8WsKCSzapNpdV9YQ1/271wxhrXzvmIqB4nJVhHTpgxAdKcuHXi1k6SrFzr
XDdsEP4nOu/ni3aQ2cBdgFeGU4S2/m9XI1fLTudN7fpIQQcS0JR/xc0jGOeQzXXR
syH7xjgQbgpzcsXneLCyVpaaKfCFLa/4f0semFych8xG+Iw/xSl0j+zM3nW8Pb3q
azVxvo3DhagyVUM+Sf4Do37X7qaglZY+zuHrUVVlsPqrgPwkw9+JK9Rz3YLTqknq
Jxv9Yk43/RN/5HYwjajuUoVL6cf/QoV71pcUptN/7ObHbSn9U0Lhs2dskv7tE4GO
YVnKwD4CuJts2DnNc89kOc9VJ6vcTjA6wu6CwCjl7sbt5F5fZsLQqqm0mtOpBpvu
qKjBLqojtOg/f3dQ8Yp5hmMRMACipDKkFAL49aBOHSB5AVId9sCvlA2JOhiGancJ
B4EkLY0qo11eGsCIShLmxuJqFal7RHJgrr5NmX2KP/BaRF9p7QA7/R8Soec96TSa
RdlLZ5/Kh5RPmTDhshAABBSEAMqs4bAWGez7BsGCj5b/baIsjRSunHnH9nvXLsZs
fOckf60l5IqS/FAwxXBPmL4BFn0NpNy0CBeCLMGaSBtRJBB3se8QRs4LaYrtR8wz
gtiBgh0pJG9vLrmS3eCr/W18GgkbAlBNhfveZD+zrhCxkKmAmBsIHOnjwXHwQKRG
A2iiCn2GeaR64cXwvHRq4JggxkVhF1jgm9OkG2nGwDr65AJ7AaV2n6aR60qA/Buj
7CISqdP7UxxaaHu6jLUe96TTZ4LOmCkaGpunG4n0ihjUouDc4fRCYKjzpIaRhCaD
ZRsyG1IV46fV2OzM0H+iO2COcHpDdcYbJBg4F2cVA4Qs5Bep2FE78bvua9iW2PF6
iJb+lJ506o3HQWrzauXkWIJbkOoLcTrzEJ5HkJQ3u8AO9fsdDLj/21J36G35XgnY
0OhMgLBkisXgvu6V2qFy0Lb3qrICT3CncNP776aol4Y62b4qMSabPVcbq0YHGI3E
xH/8Cgq7aBdT1B2swB11pZtuKkcxviVM9qXYR3X34l59oLNICocqNwTrDMUlo8hN
hwfmzZRQCcEXqYhVK7H7KwPv2A8Ywp2WVVbrZkl1GKeUngcZDp7lRVoYjn8sQsi/
KjfRsr4uABjGeyk52CHia1+ql+RrwETsyI8eU65JkardsDM46XpGaKH8XBmymHpG
QaUMKMYji02LZmIv2GIY6DgvI3rUKIf7+fdY8WhY3JtZRyhqjWss+yOqJWRPlIQP
GmZSbAREOn7HfPf/BuJ+/chaSMMFK8QV2AjTy53gl6Qt2AySkV8tqlLzS+zkVjOk
nen33QRTGxFeg8LWOVRwM3NKklGWBMeDHhI5uq+RzvziTT4R4WP24Vw4EjfbV5gp
F6zuTMX2xNR+lSlIYVA7SgGIsFItrAJ4hpH1DrnLZjvMltmXFFVU3O9AhyzfNxEG
KlxHNxwtO//qWG/JWQcLf9vBfxd0CAaORFac87xxCJx93gUnV8Toblw97h7CftI3
MuLMqG187aOOJB4AtROFOAE1yCFvq0Pbiskqa+HsQ/67gzRgfl8SU6CvuZJApo/Y
qurFwuEEPN3ciwfF9XGyAnTEoBtcLpTzHSzASlV8X7DTyaDDluqWZ6xyUSTRnePH
s+0vPmPTafDwljbXGEDNajeKErALfFcoA4vpEi52Jm34vC2ONjb0BUe5UUsZ1JCU
l1jEvhs4gsd0Y6YeOFkVq4IZrRfcEf/uA/yU96RkL8wDf0Q3nzMWH9ALVVdqTrUU
dCLiObHFoi0HaSeONqmhpefUWXYyGDb6sFLZiMcXFZjpp9/jGJbCvHkbLyb2tOC3
yQMIgUrKXjXuz+E2+CV7g1Kr5h3kwTI0tZa8E3lTHK/XWZlAjk/7zhz/XEN32p0p
7UvNnSSi51cb6uTapWk+EnL0LgUXb3xJELzKNiStm87El7T3KedhnvE7gnR7HXXv
naIQG+p8Z8lBnXF3DIxDOq7xaPi87LQXfbAZ6u4p/eNUy5Cqv5lYh4PXYYgrVBse
FxM6WW8Q8VvmmgooroYgdtuT4MBJFYbmY4BvDgm3iDESk5r0Zws5N/c3gM/8ofC4
sB0bYDRn2FPkJS48fX/17iR0IYP8Acp3GgGQFWlx3piDRR6Ev720ZQloSmGcjdfO
9TyifS10+DCdhw+euwl/ft1W7++4zAcpGSXokvyfNGOCH2U41yKHGGDOMzx7plm3
yUXEMCRuVFl0Q8HgtBsn3SwCQT5qWFjBk85d5lCEOyrMhLTCvgt022ZAoQ2cojqn
8U6fqp5dqCwvmUlENidXXEK4i2aVJHqNfAeYN3mZSBBNmtYeb4g87DrAAkrJDpSR
C1RJh+ZWAAe1gBreLdzjCo9gm8chCr5zu6J5IuecqZU1C14OMjo62tqoi+lXBbtp
ISxXE9Od7Z+ymjL8lK/pve0NbYt4NWe6aAXd2Gf5b0kOctR8TeLnmbU3Mrm9g73G
Ufn4qJQwmnzWPRyrSgcHx67/iO0LvoDyaN/aFge6dsggrsKi0h40f+57cIku72sn
QekcOo7Lt9rTuakA6n9SHYrpbBKw0sE7tvMENtLWlS4EibIar3eFfVX3nE9Edq5v
7laSSc6RQbclnyfeEB1524xaYge4lfAC/lWjPhT/H6c=
`protect END_PROTECTED
