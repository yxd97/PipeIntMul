`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFzmYuL72aDluMnKj93bvspeQW7dZPvqwrddHZTZCrY92WxUSxMBbbF2B3lDDrgK
gt2Xryty5il52ZjjIVUvOpt5IdF/Zq1qGg7tuNwKbVkavik0PYuic8wpEtYMW4yw
lvnEPOXPG9j6R/Eak5F+D+m7czBwL1DDwKkyDe59v5taNCgCe458IdtJGleU4auq
DySdIxnq32jOWMghgrOjgwnyf17Me+K7smF535Wcv/xIr8YG1/Qm4v3+fGdtaHCj
im/R4iJa12/uzG5zpATYuOUg81pJF7V2wEOX0NotGRkWb7MVqX0M5MRJ/s5n/lMR
garUahhJYxIVFdLT0FkO4iEv/+sCFnASdZM1ZENKV2/Sk6LrTOZhr9YUo7uBrX7L
7gdcGYtlz+KEAQSVI4vknA==
`protect END_PROTECTED
