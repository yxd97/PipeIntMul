`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZH3QwJgafeVfJ8MpMR6YdlLr2/GYFWeSQVPICNwHhnNmy0rP35+gqi3BmcCLtgTz
BQXltoOGMgDkuMpC86uNOb23NZrZPEitF3KO52iUEIpucgdSz5s2heDtdXlH8DpX
6I6vf+PQBxkJ6+I/59XTdKqZyl9vGu4UlnCX4T2JzQ0s2n8LeWFbTPm1moWPzaAY
KxtroNaSPOlM0iryUv9+m6RyB4sYtaWvTqdoO6+WqEO+86Fpu2Ax5fECrz+9IUw8
b4Xc2bYB5gopafdOduOxegTFvHsWUAtG3AYNsKpFRu6Dtq0MVdYkFnL/PmClcRw+
zsZLhwL+jUeDWGkzjcYa1UGnF4wtfofNI+EoAun45hy9fiWsIbdR95fmdv9BiiTr
nPDHaVRwx6W3YgsutpGAhrBfJUVpUnqqgkdhJmMO3iYWatzuXydRucPCcuG8n8hH
sn8GArjwIckz2xR26OiHMKAyzsCXHuKwBpoZUIyfxGwmHQITUjkhm895nw9OtjXQ
DJWlatG9rxOZScN+HzgZ+tRQYswYRr0KtDMvGiV82O79UoqYJj2g430wflkgXYyj
cty3cxeybw9lx2MzHYAjQm5m9iuwgqJOPmR7rWQGPrM2O0SRNfGE7UxgwaPUF6in
qlihbfH6ZtivXHpYwlxfzw68GW67EzYeOdcTZavWHFg+DhlEIKkYA2FYwdPaIo3f
xo9KYPvrNCvV3j8wQOFLJjWKpkuS4waNzzSXbM8ZoMgzwWzAlGJRn5IpncF1/Dg6
tMSRcoC1W5ZoJ4BBiOQDuFb3DCHPFiClWb0DhXwiyH1l9wHcpl6VEo84ebEOHMas
WO3vtur1Bu6s9l5X5hhB0+9uPC0bgAPoE1eqTJ0L/38HI02l35SnOKT1S0bOjund
j5936WsnOCfH6TS/MyBPvrm/jjJTVdFe8BPYFhYMAD9sEJWAze/9pdSewI1EqLrc
P8Pj8YqZVBuBfL1oVWaSSAYZvShr8Mis5oPphcksNjpfNKovnl8THA+FprV8tX4T
oDpzIimmD4L+acxRHX0pHKu4goqnaSMcQXISEIBLjfFu6z0nGkWZmEy9Lm2cDtj6
0l4wRnrpQX/CoFygdKKZliVXhMNuj1y2AMCKeNMsO2son3KBfgfuh519WZTi1oh/
/4HGqgPcGmGTJhzi9DKp3Iz7vICa1f+mOwFmHlvBEAvcVNuEaq4Rsk3bpToVmiw+
MAM/+5NXLY1t7YZAc/mJagKr6FGdx0YlXVUdvOUAxR2yw88lvIVYPM7p3ImxYaLX
ZCE75/jN3d7hg8zrsw9NLT3EBDH/QPzM0NMgqriucztVq4Q5adMf51cG2BKc2Gza
eE/E23ybsZOqPFeYuNWAtYKBSOBX/rxGuIh1N+sEvoG9d9QLi+6DY04y4WBWYegv
GD36+IxP1hyrWG9meNe88Icm4Xb0DCAQ1GaPbvTq+1Hwe9zMdbrPnzCO1woXDn8v
ePVdF+7apoDnCz3KMzZuclbQlfx9vuQ+ufSPU1x3swCUNSI3J/55O0qh4g9kxaWU
oIC5zVxOTK2P2SENOEkH+dm1PDV1Jqg1VBMT108U+stZQ1ZdtFzxQWCmmoJ2YYM1
w0t2wNB9sU/A1pyF48sSffhlJP2ojXKpW8oPcI0BSuZ+eXQfuW00/c8np4ISSQYu
SHCpCaeZwPHSnEVp1nquHlefXaU/iY/jZTOnOEiDOt8qd93OSv9s947DzCaz4MTf
pqWj9GgkDcMB6X/n7cTVObtSIQWqf5JY4oeIkyHChNx/ww9SScZfNjn/6/tlkdUZ
1JAB88lgPTJ7uQcarUlY19MmNkanNaF1zsoLd/kcXat7YXoPYKzdxzZJNaANQIN5
324eWiYG1XYq6FjjfhNKlgOubuv7VCwDfCRPMFO1xV4zlNFNzb7nLL0xDn5PTBpZ
/adZXIRq/sLtdHVqWJlvFM/qs+/7jDvSd2HGVsQTCyhSnEygFMbF7/QSDh2e0uLk
lX8P9gonds+Wn8QQkUamtr5EiZArIWMxG7jRKJMmcXv047PfmtKmgnBqD+qURwRy
Ug0FY84CtKn8p8jGa+8x+8xS3YNANs0OsvR4vgHN2fvwfgFrF7o8Z0mCZG7L3Lyb
z6o10z137l3Hlvyh9bFGLj9E1n8SutMpy+6gMX7eWBVSQ82Sqd2i2bw+NR3u4PVe
g+n1MKwoIvdCmCJ9asu1vbsVhQ76TQVqqHV7cNUrnC/9uMJiVrXT3i1QvzoyfsUw
Gi7sI8QbWg0nxzZGqUW/1SmzSxQLdJzPnOhQISbHVph94gaIEr5ODzAgFXkmP8F5
Y1ykU5wYPTEsl6aWykA+S/mbf9LobBSGpDLdmmWrX5hK7CJV9XpAw3dz9lPz78Ro
Ki+xscOOqyen+Kzw0yH/vnJGJtcj2QH74hvburRIlNKExuEt9YfMchmY0j1WJSow
YLnkXZ40Y+s7AxVVMG5giQbtZQr2rWMgYVcp3icZiHS2SJq8y6X8zeR3y80Mk20u
EFBB4Csfy70yKTtMU9BnNmHEJaoEUoz9ots3SxJw1ulmKZTdCieq886Ej4QT3dPt
1QQPI9oAlgd3hvnAaTENGO6iPu0gXxFVQix062LIyrFo1VMf/1J6nei+J8n7E7QK
bUS3GZFZshRCLfR9887H6+6mv/3qV8nbqRo3v7fxc8IvnxtB076hMb75Ik27MWyX
fGTeneTDhL3TJUGoEBR9588W+nfWHrlF9vyw4fCa5rHgNQMYmhyL36pT38KefhMj
+6pIT3o3fwj2hNwr+mGMwy9QxxfqVG7gnlaEUN0Hd1WiWmxVDADjQKkYRuVcdGDZ
YKjsYehFtNvlS96xZ6XZTBWUtpsf/xQc+UNRuPdGKVUkgvZ1rTFQbFjPY/UJUFPM
mq9TCVXYabXUl2cpgoP/V3tveR/M5iE1FGMh/6fBIeFuQFdUErhpdvJTVKK4ddNT
B8NOHvsjAZU7vFZLtTqqqucWWbtAVoDSZCUcyZAXDMXYK1vAt3HX9rhOfqGTSTsK
4AYVXHmw4gDPF18ohIM4Aw2yELGPLD4vMxurzvksaF3i3cNS4btc24/neO2F62fI
q1rPQrZFVT4d1HIxUzCf8MoWa/mJuojsAON364FAtliyi+1+fylXt/cb37RTTbo5
bpVUCOTOMg0eeCl03yH95gJKcbWDmXz/JuSX/BFmWH7TV5YZIkX2mNqVB4yv3s8K
qp9YE9uqAADIDhbWK6wiFfaP7PsHh8fTG4ty9qQnT6awrL9FD8uQVTnl2qzJ3fU/
dNRIUeX4VyaK6s56x/9LhnigYnOIiU2XqZoXQ2MbA+LoGmZiBKjSo7Xi+uqqD8Hr
pZkKfM1bTWDnR2x36Zzoi69kd+ed/UwqdhG2q5X95Dh6vKRswGMZcTOrROxfDq9K
udXSAWzS9CzXqGXtfW7sH4AvR1hCmgMVIakYHn1Nftd9JKiSBvJ7QeJU7bwDEw3J
B8lBtsZ9/aMPROLI2JWMdwIqNRSyYMh80Q625vjTsNkJdauLJ84RottYZcJYdoDe
jEojtz3kKRoOL4kNYjkVCIuV5x7gt3BEnfw2+PzZk+I3MKs9VafDnNj/u0djJD1A
DDnkazIR+CeBUH+YZhXwmKKL4DLitph1/xk/mm72txZ8d3bkYqsHnVpirqZbjPQl
gwqkgGGz/I91VSgcsX4Maue8docLsZgBnVyeBoRLvMD6GBuXRJLLhW071x7OpzYF
/VAG9yklcs2sLGMTFE2Ct5Szsy6wvbvDygwCA6qUbvL1IFfSxKNkUoCeDe/309hr
X0aCYVG0BL8PtWASTAylp8GBLUii7A7OutLasT6tueQWFxbFiHtvrfWdx7+dRv34
IyU0P4oqwZ0Rs67+MCDVVuL3YQm4n6NtT0QYb8Lb04ixsvz/Qj4C/USOvJBo5NW7
JfB59YIJlkRrqICxJa76OR3Fp1On9QzXtkXx71YvF1YiThNbA95Gi+tVBShZ0Emf
y+DErRBAwavIOH+A1YkzC4HZbnMf9wNKjs7Y64FTH7vbZQ4J6wPjdKFVnlkdiH4V
SFFiG8oNixwQlOl0xBJF8+hvmSJJws6jSpUcNORNaYNngm3LBl5n8wowvgJkgS4T
lt4xi0bxanzfJrUG6UZiKATbLqZYwgsIl9r7OFQt746OH5fZtzKYTQazU+whGlT5
DbgM/H5+xlsCzZ296GvCOB2f/CDVuDYN7ZP5/1fBJF2RiATLFA9WUFMv9GeU+c/r
Vpp6YTOEMre54glUD1M6v5QvIVXRc8x3efy+3MiLuXtKXu3EXwNsB2fKYzbSmMfO
PLsYyubqXO5nppUGAPqvEQl1/jy70xLe4IZyAMJqlff+/8erj2HiPs7EeYWMVyfv
D+iuD+cj/t+3pJFZ3g6xkCmOq2uk0b0klK7Omcqdcq5Fidx7eAzmFkUhfyMNtlsC
HbNsLs2ixIrQZmDzLL9yiqXKLlJhte9wDDMeoRFKPVSyeHdvSELqooYVQOEz6XxU
LwzSR+26txorMFmbBID0zMkZoACUxLSZ78TBrwzVOAvXeE+OPYhtrZtb1sPFKAV3
frESreTR/NxTRqhURNAGu0+wykjQDIZdkF8QevIRAM+TFELEYl4J7fnrYLI5gV3f
zbU65A0RgKv3PvtzMElttgukDyFkksTn++FIagP7SB0thoJNNDxtLjTOkwV10Qy1
a4/8A7K/2d2jZWg7/O6yRvshIpdjVyji00ZisRbmZP749Ou1Sshb5g11V5ZESWaI
zMh0iPL2E34YpGA8KlxByc1m43KuVj0Ac6ZNm2bU176fkq+7Qo4Ib4DKHSIywazu
2ncrrrc9YTA7OArdhA7hDhAmEZHR+kdUiaXQMK5BWP1hNftxKjBPaSvinKKVdFBf
BRd2v2BsFFtvGcBkQe7sgor2qT9nfWgfnp20dTPxizd7mPcDLyBTcdq4FcOfc9WY
3SzAnLRTZjsWOXi0g3mgQh4iWsdNDeMJxqGI1kUinn0FI/bkoY+v8r8OC2ukgMPW
HwsaBH6VIr8jKGkauKquRUogvTxYeXBeMngt2yg2ykT/NjZNopAexA8nYSKcLtsG
YZ6sYf3dUyYYcxpSMGb350bH/cy/YAWYX9yIJbCGaoxwB99bBxikdEP+232Sv4JD
OkMJZX+JcD1ke2Og08mSszIYU7VhVhaUdcO4UeXYMlPc4D9AMZA6sqUyh+1jscWe
mQhCnKzbH8clGEBa01UvuJ02uHv2jgn/UT1QJ5gcFT6TBjVM8v5uKSV9FSiIkqmm
t/f3+zpkExfsnAyoMr2QrT53pva50HI3vl08xJJcfsa+kLfj2tSJkZzVK7YOJYiy
6tTEMQ7MEsNX4VoDjrSjKmDqp9UoboA4gQvgZEtPzpN1RpRar+xIlTGF2XNWAjj9
O7/XLbZEP34sNJg7vGwbsZ63ZnZFiTKpycFjyD0tiuPmK1DneKUyY9p+tuE2JMYz
4qHz0PcZPee0KErMjoI2IN5VnHqSs9M5o/hcfbmgOkygfV6WTjihl/AYyVGsK06q
DQMcMcwWWpxYYE0XWtvV91mQTwDqg2ocFElHjpnTmOEsO8qaxAJ5eCn86+b5EdwN
hQxsZpGqGJLBBxcSL834qBe74FOIies2hn7y8tXczeZOCsAWxar6pdX2ozQO/a8F
2GyGLJxkhWa7IFY3Agtto99aSr2K31AIoTQrjdfanNi1cS9uHM/Cw479zVObLNZS
gmGzDNVd3EKvqGSZrNDreB+ff4ORqXoNbISVtkAW31LNmG1voV7GeWJWAhPVLvrh
8flk1bqntebe8RTNbgAGpb7FlKa5vEn/2LdWFMYxJAuuKeUVl2BlB2uK7J5z8Vq/
Bs20hbYgSHcIosIs9tNqrhwRfKM0Z9sxbRGx/TMd8flFqXMw52Wc/9VXevzgrvHm
RMb8Yp34IaNwHjuqMiZvvMhsYxNokH48uV4HsmbpuxuZERHXGkzvqD6ZzYChVPfn
VnpArbEcz6zWRtnARZPzUuR+Wn8Pi1Zj9fTBb5Vm2jmRpcgXH8tqMQGyrKeXoHcL
ZffJ+KG66rlU4I+uv7+ZiLKqpMftp/e64B/zGYXVsn9hMOyPWfyCYoD8EuPndVoh
veQkGAWvXqjXy8gz0G82grmSfLlIXPewC2ke/vYnfCOXqPykcvtCZbGfJKf13Sjd
f1pN1H4atAh7Zl0GM4Qew1jREiNvBFLMcG37oYckiT7gDShUSw1Vh7a72PE+3hi7
8vUwZXyL1Z92sgTOMYorNIczJuBmcthIkPqJoatr0MCLQL69fEwW7T3JFmNFfD1a
AILApN9zzkYux0zxFRScvJtFMd8WvJJOubhn7wUNoh3XJWwN312TRO6RBMQ8HOxM
YVnb9rbew39A9OXEBpmbwjBoURmUraPFZ2GtV1j7mOISqCHgz6h2uPyRX34hPAqU
x78dcpFAm57Ld2SXVoXE5bba1wWZNDjfQ1E0AeJu9gsRG2qX0UvKCr/4le16JX6Q
GZzFqITos5rjkUi2vsqWL01ZykNHHkK4Fl3Qlh5Mx3C5CMwh6y1/zl74yqAoybdr
ogU0uqnZzI8m+2/UsF6D6FgOHHyj73wQLuJYO7H/kOeG/5lfI4fwfQ3f7xlLZOLM
Veom2iddkLWleCT4jzjCaxfyBeI4koQy5JwRcG+r+bYcKWCaEUFnSU9/j2Z9tzCj
2nic0ThwNXJr1aICHLgYinfvtzetyzDw2SZThlDwhiPKfTqliq1uMbR+02DHw3nA
EROiboS/uuIOh1tjPLrvT175K5Z7iI6GIc2hacuVcz/pAZOsbZNZxiYv59rRPGd5
r1AULktpZWKPAp4nZCCsdYuJ3qSwQx/2S2owHXBBoBB5wOHTwLGgSZK76wWCvg5S
OkGChm/osCSVLbIH68laVOLq51Cc5u8LQvaY+BCJ/hG7b4dzfFloisNnYHByXGBQ
Yn9/cYJMPqY0oiTiaghqUmq8WEZsjJ7GvWTWvszfgRsRcf2o6Qyfd0gF5eVCEgPE
z2DkkikTNBLZ693wadeLpKbN71BuOfpw9lbjffg7r70epufOxZfIibum98DOs9gH
afFNhjVBCWYLVtXLfq/iiP4Sb8va3OMCSviV5tgsi7ylV0rKnjLjp941NNzE2YBp
XkXOrX6uu40SbZiS4cCn/iXOo4w8kGAk05RFkZ3uRt6dQh44RnhsCSz233M8WgEu
bLW5mWfGE+ZGnw7zryhXe2f2HBxdNwUUSafU71ACpkg4RZkBd8Rl/B56fD4Ua/RZ
r+bOpb/Wg71WscGT+CzDDkQbHn2Z/M9UrWD4c0bUv87owMNMmhq6TGEbymiSXf4p
zANtF7fueATjWAWGSa48xl/5Mu+HUOKqQzcIWTWks5+6eJ20O0zq8ggbmT/V5qxs
dmoOyPMoo5NVe7hCYvx8YEHL0LVBztNqUfgLlMblWCyi5iGBtencU/Wrgka6ygdX
+7nxCoDQmc7tAyKUzRX82RB49UEIRzoPmNqSGVZ6AMA5tmabJ2SpNpDvypBUNS3J
S3Sq9ImtEDBmSr0BZtPW+tJjJVh9ewT//Cy837rac2Evnj/35bND6hKnkOojUv9K
zkzUmqIxtik+h+Zah0+BsFfIKq8i4RHcZ4kFM0zuby04rN5aeUv+Iu4g00/xd8Qq
pr3mQRS/aFzcE3NpaLaSbrsclXvKPWcURpgWzaJOHaffoDFdrE8lB6j0cagk3HWe
6f5lDdBJ2dDT1wpo3wraTj81QineN0X9LtNbVyli7nfLWR/qCzOMv8t1jJdwSSLt
rVF1xf0uQtQSlM9FtI5BWZehU0W1LI6OKme1jwwgn05ddRdB7ZYqpEM/k9xSRGNh
7XTZkUTE6L53OiRftF/GPmRqQm1U8OlE45JWfI7iD6OLo+IvnFdTuScgSk20WnhC
1xbKX3lUfUa8m1rOXjHe0FWcDHF9GwVU2mTodiXHxwY701fx9X9hpBG7awEjoYz/
RgwO0ODJzxVbOaH2yLoINzfruI3dUM5nRqACMY9suZ9IhQ3X4WPuvPDTcwiSLrWc
a1x14KqbL+Bw8xUqtmTY4ke8bQzjgVUebS2F2w4L/s8B6TVhXBqH1UjyVVgL2hoU
5OT/3swW09ol/YI7Vk1S8JkuCXubNuMUYXvO9JTZXTRLeSTa6ocHYrF/Rl7KxvZF
y3YsA7R56ys5ldQjz0elGZBw5TQFeApNPXy5Jcc5d8UhSQbnJq2mVqWinwSItdAi
MT8wT2X051J52WjEaBF/FBZdVKWkBCRgebNW07bxVaQZw1saK0arYsjENyrEVhKq
VVDNcCtdsIsR0r7WTk40UTg49bzYw86gqNRSL/fc8QmGYS8T1ZdmG0Mvt/DRA45P
VU9NGuwDMkQsfT9BMDXkRGKO2X6QwVJS9VdWD9D5ixDEeiPnTU8NwHe5VJF9+9mB
qjRPVwGmoM//yYosV9759jM0cx83iaOl4dBoLab3XIiA6IEn+HvfMWI3PrL0U3ZP
JSBniHXQFhZWtN2nplTbrzhlbEw0Mp4hPtvDIGke1vqOFjLgI1fZ6lYtYYqbVG4m
Pm2qhMu79IiQR2GL+kLdW/GMtvpcTfcDOX574EG0WOiQe/wHqILlkjDpMC93cIY3
ku5Ll0YeRMm8k75Xe3ey5ZHEZMpjAWyqkLeEWSXBYSPX9Sp9oJm4sW3xPiRZS2lK
Q7yk/A6tWKcqTvvoA/35UVad+e13AxJFdFNrnmod2J9CCQfiLSLkZmXcuuqIQAQj
YGf5sm3ZhummwanM1/8b833AWLpQpK+KdPCIGKzJJvZ0uzlZ2K4tfkfXf9o+wxmd
eYI5W9TufpATR8lgy4KfVYq7PLPrlwKyklyScsrkyNNqtHAWSZZONjDc2LRb/s/k
EkmE97a6ypN/twWDpEzk8f1UH8ZFswq3q5/0ioU+eYQRphfGy4272tRBtBr1YEdg
lv8YcXZZ1567QVQs78gxjBbrPWqhTDDQbQ6UFAsocH+HLIAYSQmj23IQk+rXqLUz
XSF2U1Qnerc7SHaeByNnc8Df9v09blPphtTBhG5k+YsXrVileowvAu3Ge86ZFGW1
9EJMtkvSyyPCA8rCmghBA2RxzOK3ytjSTN18n6td+On/ikrRxVbGSsF6UFIet/Hm
aHOWOXQkvdw79d9MapU+drRmNdoQfID/Jbk8P0e4FIEyfcUZcsWXr2nUBetjJ/Ih
hpgGK8zppuGI4s8f1piOBIYYBqgWsPO28L14sKynNH+vVdTHVTsX2lJOT+zjVgvY
v+kw9Du2vp8O50AVMt/57JZ8uUcwsIPuxM8KRhcbQPX2qMUSjC6KdTpNKg1Qn5mb
8hovPDXGdcj2jWwvhRAYZBtushzMaCYxORLsUuL5nlr4p41CB7/GiYcAQQDs21SQ
inMboYm1NJMwOTSRyhx6VBDlR5Y5s1OCjicmYcm9BJWNgdLIuBWdMxTuKEUR3/MH
O+r/xrDUxPMk81igaFBWx0muA3y9e24wuLXGpyjqXe3VQ8DDP29c3s6XK8aReJ50
YlZ1rVWaJ4ynKps+p3sTOaJhMpyLOGznEeBKz4AqCjc=
`protect END_PROTECTED
