`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y80GklzmbszjYGmFl/99wBWmyM3w5NMVhdiKK1asS8tX67TaXx55tE7KjRGf/wA8
1ZPvHLX3+KWLpav6GoEr7k4ARnAoni7JBl1uthcFHDGD/jq9+WE0zsQxOqBGI7fJ
/nZ0Vf9Ajd2Fp+3ypzcToSG3i7ofq3+2YgT+rL7r9ncQwI8I/K1Ck/rzPuIOIsP2
Z1PP7a0yAuXO5ChRi3s6tAo9deuPFC9w33IOqNtbdHX3GjEKfV9c4a3NLuh6U8fN
8rZ2FvIxJKDN1oFoH5SrBLA0aGA54OfTCL52WWvD9uWBuDbhTDUTvri3zL0sxbS2
meshW2aEfJVlMF5BC7I3CdQv1zV1JVyvcDM/cl5WD6U9ema9nWSgXcMrdEBU2pGO
rQZHkjPR42SUMkcU2rfyRw==
`protect END_PROTECTED
