`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aRd/v6dX4n2F8QCvZHLGkBwnN0d6Qv81gpXl0GLGzBW5uuipQNMCGU2JAo1vzdHI
G/eXI+2SKQ1Yz6EQqbkWuHN+8DJXvVnSW3/DAOPleJUiV9Sbrq+TnAvDL+7Lf3Ld
XVumMhEJUANf2mPdx7fUyIm8JVbmWq2fcOTx2ZpAbjrs9151zfznlXkp8It3Vo4R
o6gaHCfMcc6FYUoNsQWg5qlRBQGoAwkwCt1cqfrz+k7mTvXoZbroQh3hm3unYMD2
DSjX9NL9zC90SmwTharSrR0TYnGLI6nmtZTJYO4zuM2+pcjtI7km6jmen96cirD+
LmJaZqemCypsp2bLbUKXH1BWBjvLwb/uRFTwoAusU76u39XxYnSuobvKqbC2P7Tb
RygZodGkRPvaWc2ELryC++9bB6HNIdNE7PBCSpGEHrvYiTZ5b0QOi+zZPo4YbGoC
PVsGyHWKDeMeyu9SzLFeuxQTTlyifKB/3v+8TwzIPRB1aoLF9y467uuMR1LbIuBB
ibYacYNuboRmGFRh1XR+PqdFeOjRw0qWooKwp5LzuwFPPZIyLoC6QQdGB4BVy9c2
vdwFQLy628HOCZmeAg1n8zUKJgkuWQpMzOMiAVxze5YnHFgFd5D8xaw8f9BklhOh
L55GNNPqYLQOolmgjjGc3BOEDSXC2RSg9mF7m8kFKdre3hH/17wjr1+26HWglPqI
0cnA4TwDJsH3mRafEygbaZtoN7b9wo3vO0y3vg8g/ovSVQKmuG8KlAX67/+clArZ
cWG6W4+heNDZMfcukODFAYY7s6r5DxGsNJJR640M8hPkOPoL243qTop3obCHtEPm
qKS/t63pvb6bQ28Rxj1Rf/ewnqRyI2FtOuBYsmLJOH1HLKSFpD4E8MopjcyTiM0X
9VfQ7YlSuThMHCCQLaO/bA==
`protect END_PROTECTED
