`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hI3qOYGcMd0ETe9f20R4XplDRphuHyt23H3/Jcxwed1CRlV4dz5WtZG5f5C5IjbJ
P1pLtJ5hf+zj4XSk3IwbYYtsMSFXvbr0k5x8jpGKlKNv9MvpgnNH4oJDV6twYJST
MmRuybwkhGpS7sJ8o7pSX5+7SOI//Gvc9X0mDwyc1NmhZZ2a2fFXoyong9l2jqmv
ONygLzUpQAO3m5DvzpGYwaDVke1NnNzEwKF4IDLxUVS4EZdpn4Z6gk1qoaB8hPMh
XSb2G6GVFJ+mU3J87VH2GqMQbOd7LEPzbve+go6rPkwcCq6r3oT1SUQBu9Ww+oOT
t4/DZeiTtM+YZNj9vcHuSX9yW5ed4oXBz6LMY5V4Y+fgC9A7JhzskLXF4Fv74trf
fdJq6rJo115oeyZbJMOsCF4W5EV6RxR4jX3EihyNvQZ/4bDnzi7aGd3ldPy1Yqd7
/yUbVX+a8ngFbWxu7zax/MprL6qhU4hRkXDwf+xx+cOL4OzpjlhEuSnULzvdpCBp
wbdTZHJEtDb7lPLDVKKaN5Km70/Qv80zL1J/1RDeYxYcv9MO5/HGHlfTkJ4hr5CO
Qvy5xScDnQeUkWYF7TKqKgbOeMHO9kjgJ3q+e/JA3cE53k/HQ4r5EtNaLGnwz2rm
ZAv/70eUOU6QUv2hYknEeQxbAxCooHsAwKmEBUVwyM7jcGG7v9bj/N+5SAPshWlP
RDdc81aKYhkJr2i3ys65tU2k/eGkbE7G6rjOMAiwm0ekSvthk/I+CtKdCJwNZmNb
1qjagPWUJKqBnY2h9j2ERaH/NkXIs8Sycv6tU22BonyJGDxweQ6QR8t5GDWu5b4p
3ZxgGCvaAFX4HuCb5BDnX0CUEFd1Yn0cQ//NEOZeiht1EexrsW8nhKUSiuJ2TV9r
VHCeTHPXP9W3Z7DPmU37xCW98RSS4B152HCd5/9IVUxRnHj1xCqCanCZYT/R01aE
gDBDoI5ssn5cutGocmbNd6QfiK331gYEXYx83t2Uz4PEfjpP9C2K5OyKZo1o+XVB
pEOS3H/ovaA6ooRxBEVL67DdDLB/47eHrSKA6TzWHLMu+IyNA+bJp5iTyhUqZbeA
OzbCr4QM/3HP2lhVxDmoHG/V7rYoJYRedEbY9922cRx5Qy4Lup6/b6raKVr5FSht
PPV9hPX928zlRdIY1+jSC4Mp04H4ZkI1tAp48jmUCXCOJFPddWRN7TSySXSU1mQy
X45zNJ1USWV6kgQYMADe0X3wQX3Ofw0h/Y0oU5oyBwceku6caiXO9X0RwxR3E4lj
WBunCavePJbHrJ3ZxAxaTSIlvqVLhVEYcdh9m5fRw5rOG4I9YA2kIe8lM3QCvcTx
LpR0BdtRSYLhKqfE5w9ioWqIr9LHexCyMoZQJhv2v6qRn1tz9sVlVPe+KcxBk/lb
CQJVl7ukcg8cRGFTABUXBY/bCIqt5iBPGimbSNQE8VnQ8L5WSw/2UQkQXd8pgy+1
T9xdiD30bQsM04jEh6rEhM/PFXYlwW2CyxB3ZQSDG4XhltO4ateflxQcHOPzJ/xp
+SAtXft5vW5R3DSDRYAFRaRgZ8FrmYW+vaRK401umkZ1NYEVBGmIoLj0B+ivVe/T
jSZrMULNFkmdK0kW5G1xnoWVIUfHVRcvRkcV7FZS3azZbGiBrTYvFKd66dekebeG
ce8yKuMNc1BwjuN7nQagyyL/th5WvpSWnjuG/HaxLBz6Yq+XJKCS6p8wiwpK0JdA
a0EDvvwdLaT+mvy9R4u51TGvh5gwpAgUm56sydBapVuR3KEuohUxiCjGs1bf3Kdi
zwz0dHAd2WzxTl3UJXa41dgBZdU2iLBsGI2zYqDN5fRhtm1L+lstI0utIfdf/ynW
R8IdCM/t0nf/ixmX4L5TOlljYWnpYOVhjnlsCfw/dKIGhqZ6f0GdTBQcwqy6PtXm
8Qm2f4VcbHydFpRvVi2gABmY4M0Zc9FiYmVDT+7ryGwdKOb456BJBmfjbIHrdU8c
sXYuDfjtS3ZZ58RaK1g402PawYkYJu5PvTv59+qAHjRVY6mGUEz4sthuntW1eHMf
9/74L1HX+XVg40InxlVT/0XWX9LBoaUUM+1afHuHuuJOkxsCSN+jTJerIH0ZY7Sm
660QLUf6et7305ojn0sNebTidFVqx9liAl7/xugATDGp+ddVPSv+Y32Dh1Oh1Pc/
7EykvmFLAQccRVMUF7dOsraxE94GKEX1GAu+0IXpoHfcWUXRviGhnwzXxbq4qE1f
nh1ZUujEiEkhzfhMQdXRCcnZ4/M1/XEiDobprYpWIMgGlHnYLAoT8jtZeHwWaTh4
aXOS5AtgM6mGb+Y9c6HXMrBbmIUsDOTvq2/D/VuTLTJN4J8135385ZgNo6c+ieTb
buLj+G0rirHAAkCf/8gI68SjZshMqKKaA1ec31qAxA42VeCgVeXXZC9fkLyfeGWZ
VThbKfc/gtxNQBZ2xSuMGvB8KbiIzDwAB5LFqqb0VdVKfiZjYrduESrkNs5By1wP
bCHm3OU0t/tYK4WrDGoRhAE3HmmoYtE1KrsKKtSGq3aqguGp9r8m6Y1ziicKyHAK
DVD9VFfp0d5O6nP62YAW/sDxrfmmHxM/N6PKpHNublEWKsbOWelJftU9qskJMsCV
EjH3NPV6+kQpiZ9NMP7YRBoGXK3ahyr1eKcK6zyrqicMmaeZZv3yDO3V+ZOSLk75
BHw2hlypWujLCjXm9EfYRC7LVYevPU1MeOYvr0EVJj93U5W6dLJG1ZC70mVSgN+B
3pyWk+bgOeba0ONhVFXbwDimMnYwQvW+3AknPYpL5k/2xnIATWBNq0ZkoUGxet64
PkvkIS3jZdBo5V71ocJ5HmzHJRRE7bGj96113OJzUB8LA5CNkY8a4m0muFaO0q/n
pmYJlxjUYfyTZFcWA0ZF/TZ9O16Nbm1pRh/OsWMCqQjCKhFJSev7ZZpcmTpQLbT3
HuT7krYlt/PeKYKcJ/aFuI5VjYguZqLH1+nV36WHZDaXvXmwZidtAWhn352CMoAr
/GeUqqh4LgVotAnOlFv2jTkXAcsxi/fY0nt2emaYCrIYS9MFqhZJfr2lwplkvlC9
/Y3+UHe71ORKjkCO9626LjvMSlhXCSfp+sCcX2HRFkMy90LIB1nnmJh1xVZ+YPH+
iWc6Is+bw4r8LnAdVYcQaIGyfVI7OoqIBbExtrOBNhSAXAsZEU386rGJQDUCdBuV
14mQfhP4NrFFwnu2FslZIQS8VkuTgzqX+Di2IeLz5PATPcp6zFJ2+5hGs94OKT7w
fITdZIgTrDx1iE8mY/QsqOLF4lZadDMw9QqGP4twTjzlO+lanNi13OsVKWv6nRj2
w1omTJpHs0EATl2DchVW61r23yCh8pe12pcimUrh1XRn58mGUw2SCCZQhQ2z/QI2
76af7jOzN/1NuFlLXel1lcEhOBHiYWro8HI+z9Cnz6tCE7kYLoTeSWOMqaZNYj2z
Rbyzym2f3HqhosY3Mll+j+AfKTk72SYpkg2ekt3PVc3jxD/05aPkhaeO/fsIBvOq
U2fyUMv+lQL0YiKDWt96V/Ud9AHqxt6CI49qrtRXtJonUjE7fcYK76kPB0tq5aeb
xYvQ8HV4VLYv4C04aCs44RrWUGNF5UQMnlY+t1wFtpDkBz7Gv7HkEYWXGpKSPBbm
BhIzPO6W0pBimDJa9z72lIOuItKvu2GZpkVDjsZV0XaC+3xMMTeN7YU1ia/bcQyn
UMSweEBu+ph+fRV82zA755E8vZZSz0lCtPjQGC2/ove0+bcwxFGRkb2G6Afk3Rey
qyyDgumfYLsi4yuybbvZ9P/xo3oWd+fYsNPSKmSg8zxxVtNah/MLA0hR+d33AxTR
TmGuahHN+my2y8TE4jyLe8EfJCoPhQtICzUdOXIIGl3DYwuq6JV5Pb6dS+HqWPEj
BQCBnIYs7VPRa9LulN3UwRXhCvE+ShK5q5lQFmiUrZfMbwmIX29nycZ1K10hD/Yd
9UxVY7K11cyE1WvmiSeM7n1q6MjwGUSG+Tnp0dW+yBSSnHZf3M2L/rRpyYCDeRa6
ld3Ln/23DL0OrYmt+Dns+hlR8qIe9X27QPk1iLYoX74GrgNyGjiAPEO+S9u3/QFK
rbTNFJtpUt4dgMO+2aHvnxxJxDN3fn2YMDUv5viMHR4ZSjIzINimukzTmHzJE54V
USFgwe0SiIz6EDkSQ3HU9u93omFWekQlXthSrgiQDe3KZuwLsHNmkkFM1dVG5+bf
lSFB81i167IRu03IO3pOiIhOK+moLBWmPBs5VBAnplhFMVUZREl/HNCbnbsicqYS
Z+W4rUuGSLmhGEydkxMp54SQEeBvuqLPBM1odorzb3+Y/LzecFzbyLI2/agtWbsi
bGhXS7VndoT4uBOcfjYUH2YZbqTQz1mPapu3lmezhCHGsVBdQC62t0apOd9epKgN
hYnO3pCjed9F4lBfzUMrv4bQNt51S90+7MbMqL5fibeTJftMlnNoCZ0b1q+jHTQw
c0udv+pB2HN341RIhiUHzdU05YojmxHmi5DbE5JCndlC18UdYI/htGheFmDru1cf
2lTwjBBxqiUDTpkl5QnlGUswNlWuvWTXuzLqaJTbN39ci6x6AXuZdKeAuHY/WRKF
TE+YrMvqVqiMR77wSsj3iQ4dWz747R5CpE8TPb0XeZ9n6BCXGbWWLFkKwqJDGJzu
qGGzjNvtf8lTG09FCA/52AeG1tGxEfMlTW92jviLdVHq7A/0xi0dN9xNrMGRSDIt
1k7i5k4rtVcTWi3hMZnGw4pfolV1SZ4Yz+76mJEka5nkPSM0z/SbNtwKk5y1cyGd
EaRnDhCqM4PXMmzrJRxQNrmB4i22rEZsm8ijb8G45OdILDOMigj7Bw8xuy4HrjGn
PyBxT/NZUoqsp77TlnC3Jo+Ij/2dvc/1TbdEHTdxaHykhR7kbo5D8lJK6EBY3gi6
ISaTsWPVaI0rFwRUXlXhj1EsbcSk34Y/TQA8DwF6Tn6WcCv83jQUnsF3T13h32+W
L6waP/9GuKeE+bYyplFKW8fciVaRReFdYSBd2VCMerJLb2d8B7s2J/HjkznBpFIa
DUB4S3j7hBjj8QmhAxbzqzggeqKQkBOLtyFXgRIX8UEg7CLMf4wBmIzStAZQqvO3
WRF/JWzHxTrnq0bPHYYyxBoFwcRCVPrZPItKBPTYqxd4ke5RrVwAL3q2ps3OFTue
t7GiOAxyHZjIL5uEVIBqYNcD7K0dfBZnNKU6C0z85vgUgcB/6iNtThvGIqWUpBEP
6ZbCtdbMxMFlqLhMTkwI2YfmWNQ/nom8ZgzEnqnWf8OeqJnLSjm1rNFVQ0aufKGD
0VLUFYVROqBHD07OvteAeaUntRxiiHEEmHieJ0aIXoTqOSkauA0XbOeGm3KynV0J
//0aTKvscQV2K8VZL94pdJkYon514TljR57czO3fXAR9pJtzIud5yMkAWjc1lTf7
mIorVZjjtCnTRNlm2OO8nJIW+2Hr5nHzfO57ePFmIqG0zTb5eszke2zJP1T2NPVr
ZCUWr06VGRzQ057U5j0EFLcXJoyZEAf5DZcep0rsWcBnhexUKElh+TwGsNPQuNbS
RxxfMgF2lMi1Th7/dsraauy4M0GqO7j2+l5smqbYSo/IjsZ0M6Xieyo5C89OeOGT
s33m9nEGHOWqCUI+2CkdR026Mcv/Ltt8BcZAZw4QznEgfkmpNacnc3jd3Sp0Foac
miv+E6gSkP1R8Rd90mjnar9YH9wPvpcfzj3QvIr6FCg57zP5212QRl9MrG4B6NdU
zy6D8LPn0w4fJt3h3oZw5s4PZT5m/6d+d1WYWrWHHr+tjGGqTAFNI/TZhdYBQ6BN
Ej29IxrjHGZhYaTUZ81ng3Ux9Stp3bzWjjBlGgJ6hBvUjqMw4KosJUajKpHK6j7X
PxnAlocArUBZVzTPAmKDt9Rm8afdjyH/Hm//j1QkLkgrePUCzegvWlDgOwTcbZ1s
II30tfZj+gzA9XF0kUcoEVvYaErK4pg4+dCa/VHfb/KwKLs7bldbma4abazNyMUB
5q43wfGUajdOjoFEOP+KYj5yiW9aH2/8UVmU5hGilmJqyjcVii4vIE+Zayqbrbv8
ONXlgdRos3vu9yCSvZVrOhAjbBavUY6KSUOe6fkhwP1i5ZVf7SFHxMQHhXciYler
g5G1K58pfAXOu38wwNADaV3l4sENxEPLQbBbGxeJYj72CqnybUMQ61gamQKK6IZM
SXoNqpEyjZ+1wkb0jwUZsdhC09kTOlrEaEKNwMUKAMVQYuz4A7ncbjXO5e0nVzsM
2T5u6uVh/8bnzaqgNc/Gv8pEuUiGtxemkw4+pvN+fziB9ZxRwDx5OdDXIG5YrsWy
LZ81DzBCAJA1gi4oV7N5krRha9bdZolqge5hVRPMwYhmhK15jDrYyAQKuLxezbZS
Zkq8xmsk1b9qRfYXpkyiEuCjfvBn0fBYm6UY4fIhVO5fiqQ/0luhgAbokheXjb7j
/EvpQVhQ8+DsB0WRzqfJRPNHxMTY/tXxLdsnmEHaSQznJN6SNQ7a+v2n8gapSXLE
mha1pP8rQPS0yjujKzxOQD2nDiCveFgOebY9HWujSthWGnU3m2vOolkO1G5bZfQ/
/FItBSYjueRXJn2HtytoXeXrvMtPXw9M/Wo7SF1p0YqlI1mi/lDLTnJXVtbsVDuL
b80GeX5936hMJxDNtR3LNil/E0fs3m84FwuggiE146ADTvRV2zAUy/Cv08CYMjn1
0dBmtDAr2Vw+ZatYS2FbV/JNCKnkuh89nyFWzajHF5AJXOktN0AI+vWlHvcbdtvg
Gd591Gcu0rdA2TGRrD740ekPIgSQ8zPisvoBeceCn3JIxlYmXNPYnGMk3iCxzID7
tz6z0o9YV3zpzo7KUEpOQd9zCW6r9360H2/Ej5ZYt/TnsEg34iNFTp3eWGSSR2tK
KAPL2IADRfujei0LODFjfgnVUZxJ6YEYx5aNhfhk7eqRtr42/PSCCurdl33JurMY
O1nJb1miuqJDqX2IbhJ4/qAiQFZc58EOwfJVT3B+jx+eN5P681b3l6CTsrF4HupR
s3sZDFuv7Hu+Ziazzii30l129vywargdUuKMh1VvN/BlKTwtu7lwjVWK1LuOh9BL
C2N1CComD5pZwxjwbrbXfTzJ/bMunMr7L4OtoGXp/hpm0msNgkEo/OKuvBjXTV5p
rBhZ9S57LH8nAbXNmV1nsfgt4BONOxhnT0D229++pNFriHJ5tJ2q1UNq/HVeMKiG
5gHXwNUQ3xPA9AtJM9BzTPDD8REb87yEYAWwZxtNoqmKYy0/uWrbxfmTIL1digDs
1KZ7ph4hZ4EHzcuDWkfDdiW1gO8gJMu/cFzBpxSmWoO6q4aca8hsw+x1euy8l9hx
QG4SLcV4UdCio9jWBAS44KUe5yPE5wuXlfT9SsOAUEFZM8m6SLMSufFCZHIR1uXo
OZR+rd0qG8ocYiBQO0aou5ZF0pgvthqmMOOmNTMx4qZWf9C2HMuYuT/74CG/Oj3o
SFxIr3vPO66ON26DijeplTbobe6+ukbWX4GKUfXrQvj153JlfzpQDhHhx61eezlI
2sI9jjQxEFlbvVVYJG/ib7wmjBx92wbqZSY/02hjGZeakzMFc5U75dHG2jUVV3Zr
kavT7PVdHwmabgY4aX1KScRtIqmA1iNA2ao3/p5Gaf089naqWYeqHFEgBDKQKCSW
9Td7Hl2BwilYCm3/QLUTTOPs96ECp8lLHi4vEELA5tvsJUzDUx2/AbN0blyyaQKM
10+c13TuC1kzl6ZFD1fyJwTjozAxteKtivNb2rPyfspq6dMWN9lazHDwz6G7Bh3S
bdYVCydUL7+cx3J2rcGD5BFD1ePsQAkgkcEUSaabz50fh1YQ5AOA4oJdbrJCRdpw
uRxjFjVN5idTxaj1ABvj3Yvym1He4FWupzMY2QUDG7P9n5e4IcNCpZHFv+bejnpt
PfcBuDQgYKBdoTBYMZKSDPlOwllP5ScGw1wVkiZUdyW1U0N9NT30pduIc9rQprKc
BKNoXjE9/ZNXjsCRLvilLWbHWoRZme9nSLrtoOxR/sWzM+4nHNp+uIeeP1jW6a2i
X/FiCEMVPpAbrhyfYjBdHkZGBTQFg/S/qncvJgwSxntIn263aD4sZeTz728EZaZk
tIM6dcZSjWpJ8lhyu9e9cdHvx90afW6AlKST0mOwgOKkJXsz5u82GFfoLB2SBZ77
UpWtxIREKYcWQ8qmj4d7Cf29BrivayQknwZjOfex0ViWe2w+LCQgQ9Ai87vJ8ITZ
5m4bYZO5/7pmBkMcXTVAOOxuJq50g1n9PThZaHSClW/zaH6JhmAr58BQv/Is6pAe
R+zRp1uZIdIUP674rKQgIrr5TSMko2D+zlIXBdF2Kywvng1i3HFv7/c0rDvb73nx
wEhrYwpF9jlxEK0+Ar1XhttxxDKRwoa8NtyXH1+nRQPD807VeKFTHqv9v7xWbWtW
+e5FZxlJ97fSf36upN6vUpiQbSBljlvB4tlntVSV110cR1CE0ilCSHPb0nM4tD7F
V0p9yHKJb/+cImYl/uXb0hDdaLT2/HjC3q9FaP9PR1URVrD9FZhxH0TvHFpeTRfO
ijK7mXZ8KGdJK/9LjhhZYMHYnLlF3kYhTeXYohLw4s+mg3RDrQYg78F7dyaDWd1U
Fiiv0AmRkSrsRxaRWnIuLSmyM+f4b90f5ikiUWSWTyUPF52HalScE+dCShRJzJ42
KqjeDuusBYYhqj0+69YpoHIk7HRPxFJzwQuTVnF28rfmoDPaCubMCxxJVhHdr5IY
DUTr7ILivYYJhHU+o3TkrlAdsPJivwiOMOzs/d9R8b4SPWbNm/WGW6bOzOtAnVbx
M3K2LltMwMTfPw1BMsX6Dhfll+0+UKybLiB6FY7srggBZhYctrq4ic0C4gShDkuO
BKcX2NgD/AWGPKLFiY34c6+dDot9QZRX9z0ReZ/f6EUldshG9v50vnxg7gvu8Izp
4UqLiBbscVs5Cml5LkgEV3ji1/tDos2kr7EAniGSA9w2CTpQSs50mkBFNGhCsd1F
hlYbEaxyvQ0mx8jhEDZzzNyUU1RxNjqg1rsYVxiWAQIAOjPRnyIwag8XeVRN61/X
cdJ1R8xRhQ0Z/7ypT7HXZzobDy/a6sSvz6IzC6KrgS7eGfJlKaMbdVFPASv02qfJ
qjONv+rzriEJtW1KUkD1HAFHvPLuqwmJrKyy3kf7ftSmnyzrsivwmA+SLriOBhmY
HrZ084/HzzPCF+BF6gd40fttSf8ZQV+NZYK49MSABKaFHV9lrjAHAt2P+6bnzPIt
UWoHA+o5X00NFFzEliw0vnLNknniwaV+E7Yy03xqSi1l8JlFNX/ZRpA6jO7/w6I4
H3qJD1obye5dsTDy3hyru473kAkQdL61IsIxIInzJq/PSxYG2Ux4MWIYZlcqrSgX
mIAOxcReGgwVxCx+QdKZ56JhyO362Gf3sjw7dZDYvg3G0p90s9S8T+CqAeFOiA6C
9u5X7uBlsXtbbQZZJVbjlD8VpKONImRZuA5zinnUir4656ysSW9al7dw/iRanjb6
Xyz2ZvvaWoVCz0AsZjpuW4ztfS94c/juRlAjwXTdFmp8/IBt3wuRq11mpkKMGen9
4WD5bsiMWzhxc35Ykwht7t3A7hq+0eDg35MvMdxNKdGiy9B6ylI+hJb0IzPOsLu6
CVc8q5sanhwADr0pwm1cvfsc1cM7sDiKKYevICKjwM4HvvevmY4/YvwgD/dkedqb
4e6pBGmL8ZgPwU3dTagQoIisuVAAPBNo7uPhvM999AvRHzPo/mYG/sYq8EYgNr7R
uHZsWZ+ZFzpN9VK/4D5CeJG4kthifbK304ih8WletGDd7VYnJFgYRZmYl/HaRrbN
t5JcBNOPfTE4p2ik1R3e/qZG8VsLxsPI5VN9I8vZPS9XopZSLcWLeaXAm/Wdqh71
6Akwfn7sWRxzPkDj3U6q56jglnpeeBXrH5OeiHAqIUfHAbH41cmMnKECG/mwOBkK
sAVvjO8+CBdM1PX85RZCxSRSC3IGq/QC225Ud0zVcD6r9p9uWwYl7Z/9GJKf6TOB
pRVNHBKMgQ/2R/OEdJJFwTVDUuI1QCYrBlSzb5+UBvBOkgd0/WmpCCZM8BPU5xjP
FrWWA2kTcuMiQn9iaxgUq6P9ZlOuSZY8x0masNfHyYFBRzZCay3tX596zC+8V1aH
RS3pVe127cISQbQnf2cio18GRC3h/UdUU/TIW+YlpQSwcscChIoNlhOH/OIyaFy0
BOwAppupHNH9r1LuTlIXlKzXCeqCi4fS6GomzrO6C55x6rnhmn3GEy58DXQ2M2z+
KqcD7eXeXVkIxWMeMZtX+yjKBlfhjcF3xdSE8vEVH1Ox3pYaILitmCrx1Mfe7Pl9
u4aXoAXcJS+F7JaBZsY9XQdUcq3Lwtc45sqdvJMWfeq8sSjJGJmo5J806RKKCqNl
0/76eY6V8kzfpuDKtDPURdwFxKWlXTD40pgq+w1gcI1zemaYm5GAnGeOgvnKAttj
eK2sw0irtm8XlBWYmlP3CofJiFezMMQinoa3S2CjinT7eE8WPQDTCAxQihe+m5KN
wjwWqOsWNfu1nvlF3ETBUHH1Fi6RWdH1uUfReX5ZjBKECIp2pfi20nEujzalmR6l
g1G72OHIZCKZGZqGAks71sU5PJvUAjTMxpQ4RFDHWaf1oBtyyKwdhsZweISkfeCF
JpZz855SzybWK2Oh6AwtEBg43LAKLFy8B3fB82YPs2h0HMEIAwo7KnN1j/laYwPc
5tbyx/lXcN0n9Mo4GsZNWVkgGg0En2Cpu8Sxnp/5BuISw3dWonX8xNbqiw7srDja
CvfVpE7LNWvlKexy+KFy8ycp5E4TZYN1pjUHeQB0MUjnkPqy17BBun5R9YZ9X23p
WeQCKSlBZq7QY07XfkcmJvbuj0Ueeymb2EAsa9AiXTEIuCh0KZXvE6VAE8AeWoLk
fffx+BtqCesMGlBaQiAhVbUArbs72wWcznjmQ+mUwCn6XKoccM7kRkf+j3bEIj1G
2gs6iBOZTrkzbsDiMQhjlUPkxecftIaEPPaEtWLaDrrrOslGDfzSsRUS2W8JzBLP
S5/KXK2OMFXqT6AqND/TykgfO/z9aJDFMnI3kans1BfQtj+yQRhhwBB5CaT7P2m4
ofutot93AaG+/TPu91ub8t7X3IHS8COBGSAEt9ImLMhof312V1uE0bhrfDtI3s+6
NzOROYbvK3zLs1nvZDxVvvSnArCnixx8jXE8UxGgbKC12V/7Bue1No+QEaN7Y6BN
uHMY+kCVxKJDJMqN1NOvqcbz+cJRzSulJ1h/5ytsb0fX+ibi9P/37tuhhNt/DYm9
112K31osAsNuX/i1Hf4hzumsMozZeq9BmlXLqcYa1hZBqctK+3DbX8KUH1qnIIp5
i6Lkry/Yb2RAZuSwYy3Lu+T+4HZYZ2t1jMM3DAo+In7imftdYqN+JpB1bRIlnOsM
bxFVuUcpXu9m2WpZbSiQc9nuY/GSc1mM14ObchNHxhYopZub1vviLMcG5K5Jv3sD
e/7aamd1kBscujXzJOgpQKiod6HhIBoz1mI/TmW9bF6rmyWv8w7E0KLMVXxEcvpP
0tQlT9eU0+3DX/nolUi8f4N3kfdLFHBO8Cv5Uttl6pXffwr4BP6We5/KWB6N6qB/
LuA1HJ/lL2xpbW67D1+yhNBGLR/KbRsO80jFw5n37CDRDj8umH+azsy9CSQbmCpj
4UkEted97aro0SjslMvXqmV8rXhDDBw4fV7Lwxx7a/1lg7zQ+qzFy0uywK1pngOa
aUVTssXExI4TaZTJC2BNFLliWwgltS01zSH+mIVWL6NZyBlkpggJM2k5H+RPImtD
wIuIUIxMEV2wnkNc0RuAWrUwxHsYsHVtAWDwyH//5aSG0uZ+fjyHPinbTBtASQVa
KMbDXRDbVNdzD5xW9W1ZfD7vLHJFVZC54TCHkvhXLDhcfNUIcCMNq2JKEbGV64VG
DL/fxD4bPincayFg/VSLcJ6gIeG8rU0QGcc3TREgWzPYbKlKdXm2xS3510GUJjIi
k7pRy+nje9sjosEAfTWAfP/u8vjFhEW6PpgAuftYNZzWkzwgq2Dk31YGkze7RT2/
JQijG/L8CkRyeWHbgNfA+ZPnZrlox4BescDqYUFGZTiM3qDcUMKw7Rh58UMT1y8S
SD4Ggi3ONGxjRueB12DT5La5Lm0WhXg+FB74YeHFrVVaqYGFkLKDEjlGvyjBvJa8
UlDWBQZC+YqiQFtflhahOgMSA9GIR+mnB3PXdlxuOGs+GMvOe+ajxiDfgfD+0h6u
VbCr4R3dmqF72HfVi5rFLxPRxave3VRYWupxJNi9i6iXfNwzab9PmPXljXTK1V34
2LDwogPmwldBJ1lVKepoBOh0TphH86xD0CPXxynlQvr0Iftibx1zaSTmF0vCzpId
4fuOVrVZTYlpAoKrV+7M6c3QwX+0wGzTl/XjUlOxmp2lCpxVwniQ3Zc2kcjLLSux
oH32vaXdYQVFrJ1v1yP3+EdZkxc+IqvrruRBQOqKSBs/9Bm7Z7vwDOeokbjPb4gD
hDR4XWJuvVLnuTMH27SEIn/6g+3NsgqrgSyaykjdUMTolNHr5LXUWHg3WtMgwhhB
mWImrTca04CmsA5Az4DEi94NqIY+/8teYfgLb7cLgYUI2z6rjR4wOjSAz/6ZOE3I
LXvArrbhyl//48jA2wDaS7Zu3rxTIuMUtsSCmyXNiTCRYrt5lxqSibmooN6AKd4D
0Mj+j1FtGUdqIqYci9UZbquJvuG7JAhnvTOVVDiKpA5UP2vzDB4+Q7JEykdqrqIW
QgwOGcTZ2asYm/96MrjQdz+6xXlwB+ePZ3ioWrhwChlcEvzYNxqBLg9cFXknMp3w
29yDnyToew4MfU12iI6BDIsQBEomRV6Z9z/eSCa4Vk51lTw7wnWeVYCSntOAABcd
tCMAWBTT58bX4TPFncgLSBk9FK2csBJdiYyt+8bj38+qnhtt/wMDOTSCj9Mxd8UZ
Ign2H7bfBFE7uq+r92V294Ojh3/IbppjlqwbBGuPb8Gs4AQfWyPB4KEiuwIlP0FL
VT533N9wx0nuo2dhEvH1eB45QCYs/QXuaIEMfRzMkR37RMP9mfRNUlwsOdBjJcVp
E1QPH8bIjAeiiBESRFve3h8CT7MUdjKbkPE7wuy/CJKwrsE8FUYXuCPKvOSziDz2
7q3PJSor9mVAtBhVr1PpqwmSc/70KY5IAebUFADPOnjV2tSbVasBbtACfeR3KLyI
fc2S1F6miQy9puQKwKyuZCaCWpdIXEI3d/KC8aXuf4s=
`protect END_PROTECTED
