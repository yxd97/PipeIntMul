`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FCcomanN8YoCK85Ed0IR3zd3iEBEhAk6ij8Arb3y32zEBKonjL/x4xdqQE3WnFZ+
AB5MBOznd0/HUR9WGoczRJWj8HSSGs53G6tB9xRaZh9kri5HStBdjdbdFsP/755p
FbgMnBQolGVRHIbRqn6tzCVx5ASN0RhHeMabWyIV7O67UGVUufdK7X+SYjEHyL1U
oIcyNNYsogKTqGSS0nut7mJlhKufLep5Oqbjx+2E99AnF4spG3bpQLRGxVMwSbyd
GD/S9B+uRJeRFFMu8sEgphYueA8XNg/KlH+ZGSAZE8ueK5jAffu+3JG46mra+U+i
0D4IVayHo7lTfFL+Wp9JHJ5a1UQ0dQ9qY8zPKIxrRiQsHjDRI0LYh2dgIgDUjXmI
7+7VPPr7MQ62vuRMRWgyI1uojJw/Il3dD3bdIIIRk4V/obow8FcGUKM/wexHbtT+
i/XjNkwW93KnsZ7awAVIXb3nXLza31rxl+pc3/gErDsMifGz091yhTrOSfgunUQ2
UIatcdJIwFxcQRabLsCcBp3XrKn+ohEcGResLopvZQKPU4cU7p80tPbm/GhVpwhe
DFk+AKvdogW5IOSUPZGXuHN4k6CkmWoTUUB299aUco2ftArEueKn14K+Lfkt6o6r
VQPBZihH5P4VF6LFCdpVbeZlaBR0eWoWsxFvEjBeHdpMET2m7KknsjEsSyR5grjV
j+sXOhkT2ZrIf7/Ur4GBA1Es0H0oDEppRmGhICNkWkg=
`protect END_PROTECTED
