`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQxkAbIW+3QVaX1Olom3s462JoCpT22GDEHzv/crq6v2kn68TAOqWfuCNl6dYeJ/
MW3g0pIcH+aas4/6dh6KyJnaUxZgTm1uwL0s/+Q0nr0wNqq9oMrvtBMp/UEUPKCI
ZWcs0T0sABNsMjsB3G50pRNjWzejX+TGSAWGhWlo+qzxuVhZ4MEHh37Yaw3jzfbL
i+M2OTAM8ZBqfo+By+YB/t086RzbzV12FsP3vwTcvjS7ApPeSeYURmetElZLcECg
V90/oz26yDEGMC3o6wcvTC+o1FOcgpSxlglSCi9N4XEVB0aNm/fv8DWSuFs+gBi/
SSq09ejQai2CCGU6F23FQ2ed0ZID8cZc8Sx47RqBsa7g0ctaFpjrMgNcE7N82Ghw
d4WVMSudG24jeTiOTSzfeOqyKyttV6xt+kk1GJVbTdxU9yONmy0tSfJZDtr4/GnU
`protect END_PROTECTED
