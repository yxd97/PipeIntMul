`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hab9DNGAUB9UFCcyIOChm+sHs1eQOKYiXEw/lEpzq0ofwlWcuvKIBNb2W2mIByiG
Ec9aGxez2m2ChGOWguRNz5skZC19l5/oLXNiZLfPyvSZHHiw/U3MSXz6I0PcfQ7c
UqATSNHTwCocnzsSExVZW+vrCCvKAeT4K30Q+ZloSgI2AjLHXC9ATDMj0HuRUPRe
SA51jMnxBpVs11P5unC9f67ePG6BLoba9gOODeehfUmiEzOPfYdp62iDwI8GFMQb
5Hbloycx4fjBg8DsV6SXzrMMkVPjbYC+e2eBZQSvkreTZBmYwb+SDd+AF/RM7Wxy
VbLz/X/8tZf1aX2pZszPlSMyRZi2TPiwrxf3L3MDtYw0REE3MwNoX+EL5gMWw6Ye
kBwIGEGK6Zt/eyJIDaPSDwufaKpEM6N1LcQ9nIzcw1Fg4RDMa2aAse2TWvx4ec8T
`protect END_PROTECTED
