`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONkRyzpu/IuEmH8oSKv7rlSON8bVc9NiNqiCyTHCuTWPRaOhUJdRBDRRtR/pqBV4
cN3/1uE8lu+u/OgdDRetvohlnQZhLwQRXVgYP65yolRh0rti51XEM6YVqTw9X03c
1poasqVA8RyLkByjvasQvKj4OVnzh8EYTl8t6iUiBWuhIl8sM2MJIUTt0vGfNp6V
gpxQxs+jMJENORDxG/2C1qXUxe9CzSEndaGSFof5PdvKkHhlg8lGu9CtWxm5Wpf8
xlVvOzIvAYhSpo+XJScz/sq3IoPsyq+IeBK+aLkoPYhoWH19iMd/wKJf651VxHDq
aDlMIspjFsSyfiw2pvyJOb2Qo3OoU4rWEWUVe5lO/tsecXrmaM2iAL9AJP1oSgpQ
L7nmrxWgxwoNErJob6udyGsE9UIbet4cbHSsRnZUOBArgZMwqu/umaafnf4Q71gv
GL9BDvM+Ja/1v0hGhTkzqtWp4EEVI8F755LJgja/tiQVNJajgkR7Km4YjQ/d9Li3
oikdp2zlfaDxPdv6p+lwVezd9V7hUQSWc8JE+fRm34m8cLOLrhBaS0QJ9nEtKjBx
7AaqRRxsO1e9xu0lI9Xb7od5Tss/QnakQzv6SCE00A8OFdP8wZTxskFAjFdr3Dg9
FHyzbe9DfLYXx3DjedFgUUjPj+SgXEzC0i4ZebMmrQ8sDD2Mo9qV1xaYVAJDfybD
ZE27dk2xZdhUxDZINN2sA9b6fISpDRGSd75IBOQmlz1M9bhgrlDvi5eam/zSu6kO
OQqcKP+gcHU9m7bFyc55TUTCtVDnOvnCmwJbIZ0mfM9ULnywhluPFUz+WIIlLOSs
ZTko0qhjBPr82dr2BCc8XFEIk0TyR8w/RPTG1OySmvQDg5RaKjPJdqkNL2Xy1Fpl
VAiulMKQAacJI2cCnCGQ0fArp07vt00C5mVv/mR9Zp2q68rC3+adpMFGdj8UqpMm
wDM47q3ld/TrQu9BcHip+Fh8NSeTMWxa11Al3vxPJxUAFGoBbGVg+igPnH/yA3uj
dwJR+dyEmgVKCnpsW1usAcyWmtN2/jRSJtmjYdj7lh6vjEuc22gEEDGqLEbVHixv
GhfQaE669LB/J37IC4/JzaUF/7hN6RbvEuGVZeLEzlJflzJc8sp6LMxVd/kUdxXx
Z7p3nLy2BllfqJPZ34a2DXH8Rxcw8Tn0rpFTRZJvpcJf4iqr9ZlxmFbBg6yku6Hg
n/AnWbMwbBqRD99UtYuTXCHNpKbHEozpi7PkeoM8z+/csOmMk5gceYtCzO9eXdgS
TmzuKBNbGBfoyikuTg9JQYYyzSOSqz2BNTKmNMzkgHIFU3vg8ItEzLr07rAt+O04
2D6o7Wz0vAw38iMD9P9f8dFG1bvvNamWzmYTPTZL6yEuPIY/fpiuHyKeO9iUqQwL
pAT9iUsXbQxDYqshgK42DTOPJLTTMGMiLEOjiEHqE/75DwnA1OakRF57wWIB1GfB
eNEf5ZQ6nS1iBb8LCwQAHSlxAT+T6vUH99HTZb2BBv+vD+9j2s9D2PccVvUDD6Qn
u7JBaM+bH9ipJe/W4RFNT7EC/RTHSN443llw1/AHsGHXUslBV/+88dppipgcnrgs
vOsbybKKs0BKDbyA0hrQT4i5LI9lClnP6Vl1HsjTfJ2y60UjEEGSv+WhoCCjlk63
uVmhBqXJPHG2cnqWbZboPmjmv4IzUaGLaV6jzt3SR9GBACoimHNzKL/4XzXD+3bj
NUVrD/lTZsfMBfMOotmH93/czfs/zXs5Upq/6qRL43fYiBpQg9xS0Xlq4Hfy+HEq
so0LiPgPtGCTsQvHlfzoYq0nPZtHZaWYcXTNDkH3cVCYDSVboaQT9f3i0yShpUZM
4IqSzWp7h1qysOI+e64tyOzAN1ry11gVEfha0G12W+oidhPoZntKzgLO6vZUPslS
+jbh0C24D/9KCYUwePHsRRGPuG7CLp2YIWrl4BCz+eMN7cdb8HkSxVvwm5Cy/pra
a5bXZweunkuNuUtrc6Gr/y1/TJTYTBkINYePB9FxCbN/aZ2wJjPembgHiDoTyRjg
9XJMZJMxeA73EyWsYVg2uPl0S4iI8+ac5YojB2xPhsrXSEKxg4K4WIT0rqWyDFmd
en5pwBbRQ6j0A7IwmGN4Q19XX6p/99E0UlTrBeM3cEP/Tixjb+p9xgO+8EKojpY7
VZ/QxRvYJ7mpLDF3bx4nG7qkqk4+cbV84TIX69h31mtn5vYyEe9RI10/+J5OLcCS
WHmmUo/tDwTyFPAWFJvhg3Kf1NDXx7h+EF6gLdJg9fi3wsdivi4UJNu/UkLkfCK6
R5BUBk7PanKjl57QsrjRLhrA28QyQYj+VVNtO7WiX65ySIIHoWCwZduxuDL8F7m5
gDMrLyaLja2ZmQ74LWThFixpfCsLifKxOYDOk27lz1SDUHoej6TdOsm7lgKfo/BY
CFqPIpwMpxPunWOa5dXLmltt3a94FbKBY0HkuQuHgUi75KJ/TadIL0UCx5VO0d4K
IomuMNpe+oG2v0KLBlA8QUYKsyWDnq0UJH0v4PKQdrza1ykSlaDZaWX9rGIMEhyt
PYCga5bj+7IHCmpcsiYZtFDJeqhNizaCv6+NMUfCGoUL8od6ouEhx2GfKCPE+6vK
u+jl+vUS9DwcA1vnqZf6iisbXP6+d96YktWm9Q/UQFcCPg/KqqLywXjBXIUEyMEj
ui0McI8GCZbGpuIMIfvKg753QSKTrgqNKvUbyBisPXJwqX+mJn7w+mCgs+OkosmS
CVikdc7bjgM6rj9RnIiW6CeTw1dui9vUZ6eA/f7t+Ka87ghbTcxRY9RKlE4ua/Oe
gQsgUDpHEvSeUOdqdmYxrYigpmkA7Is5JLAQiOsViFm4RP0kVNfkmK3u9izfIQJN
ty5B+6EjFhnWKDplswujxlMurnH4Z0QRJgFdPdgrZFGC36+iqKJYCDersg5WhpWk
4DvXish8/JhJ4SgqYIPmQ8pu0lANEU4Hf1oPHzDK/Wj+K2sdPmvQJZMoSR+AUH7+
0N6vM2vgn9oaw2fpOpz4gB3NKnw0qB+ARturNs0JRcl8/4FWNmOSqhUPN+It2+wJ
VsJ0tTh50hxHd44VzH/DFtlzl1AuioTlYThSa9Sf3IgAxjp56kX//7syf828MjwY
QF5xzRnD+O3vLqdOliyjkqO7Xp1WWgGCartBrJZiIXV4ghKeE4sQIhKlug7eBZRx
4NeMTTOzbh9Rxa9Xg/+yqCRkA6ZPDPksdkziSekQ942BmE9QvxSUpBLmog8om7cx
4CCPbzWFlOcJBJ83ORI4kQP3XcRFBlZjzAbTYlFGGKQ3F9cr3iylzdDcRfWomT2Y
F5IfA6jH5DxYw75/x9A52IUblkDYhzz88zLFweyxGQlZUlr2qRM1G3ZIcVhkV2P4
wIndVu86owJPpE41Jbm9TsdazymhYXIQuoV37LneG8G0FZbYknr99gw3zS9+ehMW
rZrGmJkDqbU1BYbWIH+rsuLXqLpRcYbQNwfUj0YpZPwSlIXMb9/ZLdoDFDOdmZhW
7vDkulp/CgQptGzvsUKc6fK1fwRCErReCGyhdxAiwbr7n/4pWOiFsAio5UyAsLxH
Hh6B+1K+7q/RciXUNWLy2Wa+gP77s4q3SElNuvaCGsz23LINNp91hSQ+jjMos+HA
1EKN/hFLtyqsZJXu4V6OolKmusEaZJZBsdq1FZuTUoI22+6YtJzSuLOFy+aWxF01
1xUy/1Ur7NVD+JBDKXpTe1NzYAVFYgvOE8TEZdQ3yYKqcHoyFpwfIxSudLjCj+fD
0BePkuzi8D8095Iidf2HySY8eHxquLS4Q8hND/jI4L+ZmEfaAiBadD0U4b/+sJQa
e2gkye3F5vA5uLY8sfFqhYmSQo4TKInmi71Lnk/KreWDkvXa66SpQyStirYotvKu
943a0Q5QoHLL9+qoMi78ODlhQdIDRnTZcn6vGrF6dEYXmGA7oy/w0XoXjCIJSU2t
bC76fcH2R1EN7hQ13HmGYDU1vqlYRo4MTjFl6tDt4vFFpZMprtA2j2bGPF80I/0n
DhoWo2cm0H40/6s0nMl0zZFnbwxZDHdUJOzKl36e7dD/ldpldsnGcrXiKRZ59GP/
dllKGDKwJnDjwyqEwm87KCpBCjpCtBWLGiqB4i+/zz2nhLXZ6IPIAmfkoeseOCvO
l3XrEGHJqrQW/UQG2esA2OvrKi8VmAPdoBnRdRzCxJLi/M9doVAF+5Kg/Rczn8P+
ak/VTUZc1f9BSycptdCJ1p8fwdU5EjOnhoR1bZ1ZVbN4DX8bgq4tKZ/vhM+iwGid
sjsgUgbeeEr5s2hPBeQ01U/IlahYxnxCAU/bs+1NPJIfwnq1grOE87XED1OdZSIJ
jhsNpDKDr4xFZpS5/qUsJePehEkX357CGbn3+SvLGSrViRRV5YwpT4hl6VWpaZy3
5lOINAYiPojDK1q2GgNcSRK/NNztCBknZkTDfcsr6SD9Nlo4c7vgczmcb+DqjAOt
b+yfuQs+IIRghlud9ANMs2JbLFZuKj3Z+16FyxWYodeonB17JQMCKdZ0brZIIygR
OCPRJq0ePaReLJF0C9NWDx7Lzp+8tqDUQL+fBgOtga6G+mCb1nGLvDzVAIZqxM7n
JyYV52JNsWTjBw5ob/j4676JYxibA1hypDqoDMzvVvE1xwLLwnlZBVk8Td2RnUbm
BcJ0dleP93kic6Kr/NBnPxGrm1GUtEbLH2wqng+G9rYSFxzOLtjxKTnYhPd0QesN
HUj/79de/O0zTppckJGZ329Q8lXC/kEiO8gc0LZUaXXrfRTVlWEF8tQdDZeHll03
65+M/O0sliPl3gzRCER9XTDUjkKPxFWE8aVGTFWVYY8ahGskgMZap52Ypcxfg7qX
74uw/kH0JKbpwAS30wgdK8lrUbsuuSUSrLwH3Jr77FOupf68rVnxRxi8QFybRTex
2AS8NNb6NQChvXdBfobJkMC9nD0MTyR4H3x9cPtXznebLacuhY0RCmUTwsXqx7Du
TgkB1W6H5RpSIiWjL8G8H+ty1LYaKHPRdVZJ/actKoJHAfcY/JXSfMpoZi5xhvtM
J9uUT6XvCdv+PxkUw36wH/HR+IBvlq6hRn0YyEgGsPzXb641J/ot4SGZ+6Rc3xU3
mSlnRkw5SRclTTWvfU64ggVO2QYfZDc4azhaFw35+I4pM8hgDHDwxV2lJsncucbG
iGEcLegPdFKoGdvkWj0hnJ9CVJnSFHXBd0C8M867Ze6a60so6mdiYsUZhfAI0tWs
xKgL0leYOtR3lDyKIMfPNsCDwdthGnzhuYYFS5+G8rSJobHU3l/GUPdTUkee0Xuy
n0OikBWv5L4BFqj6aXMHt9MTAHjea/v1KyBf+CU+OzNEycd7KUGjIh+rL9snWy/r
xv7Dc5zYLxm9lw2h0ojSDis+/2wDKRMs1iOrEjdlFWksYUSI/vgsuJsBoxBy6HfD
s21ljn6p5uGd8Is2CXTT/49GEzERCqH26AqwnDe2YhXaNx0VrxG+/MDbciScQQD8
pdNe7I0PqvRd7dGX26WdQ6rImzmuf97ND9rFJ0j2bTxDshcDZ/ObgOT1ut/j9bLu
NtLPvlFLLmi4ULaXm8rpe2xP/Cf8QIt0D05eWg0w7B2synRVuA2jq4VyjO/o6qYH
INvMLn/ZH9gYC+/5bFn2jcJ8Fc2VDIEIYIQtnCKnsGeMaJ3RrRZ4KTxzGFG+xO1J
JhI7iUG4be4xWBvNoMhbhrQpJ7jZlobFm27PndPmhlVlyoWB0swR2Vfl7XYC3tY4
Xn6BKcG7ghlatVy7O3JkUi398IgMJTH8gZ/FYwiUrhfdRERWw71nCGGxYDrvs/tp
GIxnMc9KEIKym99/xCTB2/RMVZz2q843uu2tySF/obRjSH4mngtsNr1HzIk3Ibdy
HRVSJOpLmW9osjUgSv/kh0hhWyf5OWD6HYLvlBiD9HQSnJpYSYGGb0wyM+3vMfBn
lBy07gxgpyvaaCiZxHn2WCbm+HRknD7dVnhHScJ7stxKW2G86SEyoAue9KfxpVJh
NoWkI6ixvlaBWxmtPK9MFNjtd+zcIrbDHt0Mf7JkaQBN1nwbWHK86ycBTZyU3GgE
bAfXns1FVXjwFXisTTquEAq9zxM8DExYEo3s48+1eLzy0+qeKu7IALFX6jmQrW9g
ZJUP8ic4nafvxc0S50vR3waaw9r92yB7tn2CisM5zCQ5M2yOCv+cwmJFCSnv4Twv
lKybvWQ8oGRwpKUUZwNcVzHL9U/ytR1NTeMXWSW/YjVsa4bTPyuQ6wdb5ZtPgZ8D
TUxhmyNZBF40sRVbjXT8u1cQaT5Jdc4EIZAYXszPGTIwWMw6a0e4pw+BqaC6AeZt
4ul+k4CxA9BpA35PM4z7wPmR5gwmZipP5npgMQveUMAuz1KGkXAcoJoQuUXmD8uh
UCFrdWqOVSxAxdW0LZoV0DR8LKbvPenJR9wt1ey5aXjaphg8I7vqQJM7T66Ihxtl
V/PQZdt8U7gucUvb904PgYxHLIL8XOwsCNkulGh+wNm0raxN7OSTZwG9EJzsvuHy
fPr0uob+OZtCBCBkE3efwSnm9SNdi+/I6G0J7fwlsBIosu9gcq7WurwXZnHsM6ig
9zgnKuPC7z1fxhbqKzPrIQ3hLnH/wLbTQRqtp/KBWBfSn3TmfZYQE7Z9CTHpv/pY
z+ks66l6ZzQCwX3lfWlVZNaO5n+s5QPUVqBFboxdCBs1eSyy4bVbRyR3/f98A0Cf
WCfd4Wf6XyPWsrmbBzvRHXjAdqUlRxFiiP2i975rPxd/9DbhYaSfCCGnh9Wa7m7n
1zfl8txDsgQ0/hqDN5wVhELzQ5L8z/oicxkyRnpFcoznkaGyVWX5vChstLPcGn/t
4m43eAYl+2rOSx08Q+B1yun9UjzvHkthxaMvnWLbw3B5P3voPrP9xecWeGbd2f33
L/sbiQFDVnvb4nB1g0ixQs6jztEchL/GzETWw0LeJp8z3d9rdUvVku4ggT8+rAQS
NJ1OmxtcEXkI4KPhGaqycXDSohbhngdjsM5pkrKmyMezNGdKl9I0hY4pTOsNl9mE
6390296fUMdUNP2goOt0lK/Oj2ppsKz193NinZ0BhY0cZ9YzgFIcbvuJy4H+d82M
Hobz6B/CE+hnQmXmcAytQRQb3cw+ee+CYlX4mxMpJafQGzwiTnfQFMLMTeIkUnhg
Q2GSzgsTcuSs8RMpXGEfMqHd8hMmXRWoDGgtHXinMhcZVNqTpPiVUQlVXtb5hSjJ
9L89Ai8FNB/AQDCeyy6wectqLORLbQyXWAqyOk4mVRcehVsIGIA3/5+uDLokZEm9
DCaSG7b99UX/o4FZ8udjTw==
`protect END_PROTECTED
