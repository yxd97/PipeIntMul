`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ta6FPfdtRybhhrJeW/HaEgTu4Tj8s3x2jOKoFDtNGAJwdW1sy/I/DwxKJ3T1fGSH
ao4rGEupNUOcxCwGqfOagVDY9pbqAcaRpsLjNV1Ui4oaEdUCVHUL8ZWGzN+2pDMy
19mmjaMoJ7VyNmAY49sHq1ltOTesCnOFM3JryG0qHN48mfmfbJMFhrNQm937OGvR
tXi1vYuXvIw9q6rJA7hzBTHoaXKVRvZg0nA82bobFDiGgJf5Fnat49X/tln+8k49
ul4VUKTglmx7sqy/FzlObK5VA6TWRSdrrFBW2UzFfL8K8mA1Da9muZIvbilPEy26
JfHkaH3uhITbRGxf4S8xv8jGb1S4a/UCGW6hnHJdAqQrjfLfUvHsaeemtwtX4dYh
G1SSKtmkj1p/voPoCW9uj+uHjCzd3JXD2Dx4jlExuwhbIuTfjTsQYOQtLsvqZ/ra
bs6Ebwk0w4b23mVT+gWwwNTsiR7JeBE77jxiLcvF3UWEXQcXqRdUB5p46CGbhLuH
o1SpvoI/5YGLdxD6VkN79gjue820fP+KM6igbGjpetlg2PJXqKc4FyosxoTxJGYZ
YQyZQm0uo5srAMHKuzFVqhIYIiWE49Va2FQo/ze3mozcQJT24S++QpTL5xbom9UE
0GGVFMEtxtNB673353TPh1R094ZyZgGeSBZDF8qxdzhbQAR9ARJOHb3Di+0Phj4O
nlj2zfdohI1TTr1AG17Au+BYZgduro0sD8RHY7ciXghAA8P9cjZ/3/trGITd6SVY
FT9ayXoYhC5hGkN7BX+Do/JtDEDs/ri6nQhxfhWzS+Er2PrBnek4S6nSyBI2GlCE
hf+qkiNAhSFmWbKIrgIbq8kyPT/kDwoocMmCaNN++Eps3D+mo9VZMSzk81wQ58nJ
QYvymVFk2K3IfUg86ZJE43z3W4cuqUYyXR1dum3ZjTUlkFkiRJxhp0qUSi+Co+2A
iRaluTNGHSsdFptfjTZPKdf9q+UzQJsz8ALSts0MkOyORTKpMY0sxxql3O9sILUx
GWAQy/T3+BaNCmwCvTrWu0nl8o2GrpE2LTKG9DspedP4hrEUgAXH8a//RDAzgdms
52cFl2s9jvZAk7SwuXgCAStYIgflVC5fz89BtdIxiRHAP6buMBbhS5/HMPvIkVNI
QVXHI9y8LseneKdw1gCzm70RGOpfE4Z/+EXVvU0szKkHfYlS/VaMXJ0Ezo0Xt0k+
i0zpF6LFa+vA3vUnwOSdfcWUgjtH2+2j5fLFdkr9xqxSHjvfMxP4O01XfBsdTieq
sTgbxkEdlmEKc2zmS/uE6QAxbS+bGqzfHtQIeNdNPq1ZK+w267H6LkvXN5l2tRYF
sZRP8u56Zt9QG/PTW9/mrvA2/dIuNmBFKh+xqo+Lpv4uAiaEjTSaBQfULPTbgwMK
05pHr0cbP25Cu/WdkeJsVCd8vPMKS+elglawGY/YMrNik5u2q6vQl749beIuJp5G
u7cEcoiggN8P/eDDVGcJjOYnBUHfR4OsWAv8a0l9YKz1UNXmkAXWFas0TjGPT/47
FgQiC1Zwa/fOyRkNt5Wm5ONNQWC1zbr3o18kh/HgQrrUreQTzPbSqfmNQy7l8xGx
mfBAx8vN7gkCTnzqKco98JprJt9oZaD+1wXIjaLShCWp/LA9gI1Ku4feehue+cx8
M7eFzHCYS5iAlc2O4ZCoxANJ2GAawQ6rTtJoEkc4tVftVIh5JXZCYFI9hnxpqoJ6
`protect END_PROTECTED
