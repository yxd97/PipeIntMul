`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nP6nheKmpcxtDQktYTFIhM+TxnafWN0e3/oCy66/9t6xaMgOUMFA8nqphUs/llj8
/Lpb9zd6V9f7v0JZsOcIZxfiUL8jiXVkGjg9/b2UVSR2UXpFKH2edKqaUf1YniWn
pN3pkMt4ORvobJGl3OTephsiuGYgdij2WSTJRazDYmilm6vtV7oO6RImO+0Kh22T
UWvxN2pdSx5r9nAesbrO+zNK7GWXsir89SNtZb+sXU3BV4u6dyYEbLLMRxUAGR5w
`protect END_PROTECTED
