`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0+YK8+rUD+uEdMol3732KmLk1EnQa/qiS0MSWO0kO0CzUVtz3inDa0J++/sAUzE2
KLplAOMoAVB3C9eTkgrYcDLLGT7AGXGcjUjOVFKIqMjteH6LwHIrqz6PkJCvVOhl
y/5XDM+H/HppKm1aHtVl8CmGncV0qKqho4Ca6lwtGMHnG9XDiP3bU2/uKRqKwE5A
hWculaJvwWqi5xbyEE8VvGj/m7VwVrkKQDZnaiWPabPWWNML2ERh67imZP9mUuRS
moIxvgU25BAdCH4x0Gr1eR8yqNUSF4MDXF9MDk0haWk=
`protect END_PROTECTED
