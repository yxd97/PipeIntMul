`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8e3wxLb7IhIVrXWCEfeZ3bBZApQg9X0Qs0D7ZPDJf0N68VTSVi+hnelkw4P2GDHf
1hRKozvhD9BYfog9uytsZlLaDKOSRf2vC+mQqldKgZ/2bIgnLzvl0mWu0cinJRDp
hFHQjtrgUudGNj/OAJWRNROfRhKBPtkOGkUcklSUfUoVCiqTdq0BrLZWNdmxLOEg
7JtVR8a5U0mZEMQjfB0wiGL7VZpU5DO/kSQYr4L9cTvyQVL7DDpxhYwu6VToXfim
tyCg4rdxQOjbzVbKMdN+Rvkx1eHPNojbgv9UphsG9j9MAZMFr0IM5wyBcqxyY4pG
El2NoFY1zsRFIbUy0oyMCafJhkQgolrRTq653cu6dDlYrD+deiZnE8mbU4SxdMMz
ancpd0GsgwlpzDPoEOkxF8uDQIxAo8fF9Vp7vgBDn7DxFR1pWIB6jqSFCD4lzcTx
oijqJh4fbylIARp/qDzSflyMoW3bFl8nZYyl8oqtmE259OZ+GQyu7rtyQ/ZYK5WE
A/rgGVnC4Fm7Uztr3usEmUA5qrFl7NqdFyBuW+yJTbF0SMI+3/4D2vRaKZbZ0zGu
+PtQb4biuYkHYeIKkHLxQ5eJ6yeTGnd00D0QO5zvBjZKkY8N39SmLPw7vwreKG9J
LHzSdPLSqyy8SaUPYyAOF0CYYczM2LQZGt6DI0itDcKaO5gYLaMGMyMtrJ5pL+GE
4cKtrYVUQYC7kRjf6GUQSjWfkLQjauVgKYg6vwIQTHJemdCXampVcCnoTQesHZ9R
3tD5Q5e2r/oJy6u0fY/fd2SSDCCCZY3U81bfAxEIB+BoUL9sM4k6wRbzaX+xVMkC
O89c24EgQJsaY4IXT1CdORG0RJ0OHwu73b5YSVWsb/COqn6FUOg+jvWyv3DvYK/G
pxhfp1u75YhUXHqQsJNd995EvUXTuPok673VEIEkVnWdV4e93YQe1GHJW7xCU45R
IbmFrsbQU8Jmz/86p01nF3eamXm8rWqgAj8mmVBpX2rkhR0dSkSWn9Cv4OiNd2/B
Sqgp89cuDaI1VCENruRjom8U3/+zAecC1DLxjoiSi36n3kR1NxtXV4/u1q+Vj3/Y
4jsBFKlGFnKoZfIn/SuaaJ1ysS1QK/urlTBf3BOyLWFDt40Fx20TfW7hO6GEaEwW
ZUyaXiUVJUaDL41kod9DAFVhe/f6BG3JhxMWS6F/Zuscs/0Qro6rQ2BfvyUaXXOv
8dSCXwVeJeopjNAqmyaVhCbe0b/F3D2d58Kf34A4QPlFAm2fWsDIT+uX5QbjMnaR
bCu/E0cdktlj9tC9j9ptAjY/yi0/yfc2WvJL6T4dczPWMut0/Lc5sa8AxpnpBDw8
4Q/hyJVGaYYIVQvI8gaOKXlNHaxqmnu8CT4tzl0wRnTT1TyycoCn2M5UoIIUd875
vgS51y4UyrahX776mfpmafc+bz1vpkZIChRXNF8PGgV25qXgdjCo6V5jXQ2lokFJ
EyrWxTvT+ZBdz8ThdI9ieLMzpHrtWLwurU8aPBZ6El/LO16ebSttkC5oOG7g/sZL
W3PZ6meN0H4WbE81tfK9RmcR80wadRS+9O+SJfy+9LcpP4pJrxi5+2dnFhhDrarw
fMeDbPrsKcGmUD+/UyvBlz+Ye9p25uwbqTwJjAaFgsGphz26KKdjX+BpIeO8jLqO
HpjfI2YnIo/mUtK5bKLzOP3zKhpYQiH5vpkxXpDZKVg6TqKRibgBKETWHDjifz8X
C45w6g+SgbLi1ffUT1XQ5H2BbI8/J86cIkoNla4JYhSpAx7646PjT1udmbCQ6Uxs
aGkYUM+p6eERFC+9+uTVyVdAow2J6i4xJT1G4rCiuBswtiNiqYFrp77undvWtV0F
/wJaE3JgC5LJOyRIASgw1GvUIeuiqxHyVgW9QcSsXcFry4DAA9+4iPwCU5ngRNAz
/sKDWf+FvdWH79TcgO+bv+m7/gh/XIJ7TN2PIuxTKxsf8jOdYVRyEFwmsGZoETqn
tqRfI9wxvhkOWOIOU3f4WCTyzk6NBxZgf7mFChrDJOlOPGnKPKOOsjkocAhsT2eW
jMN2MchL+WLmWqhJYas4fywfIL6FK8LV/oadvhgLBNfaoKyJLfoOn9HDPMCij6+Z
ZuAqVIqP3RqXUa+AreaLMutY/qTr0JwDK2fv1qPadjKLW+ttRaT/K99W1BNlVJki
otoApfQgVcfy7K5rbVjTH1fZ6NWMjdAeyMecaGMsuNZfeTpWnD65yqLoPpfDqBIs
jg8GtLPtuQVKG3jYpSUBMyBhrSlwEc+H3yPHEKwl/3NsU7Rz5vlIHmVJ13VEBSKB
aoHqE7Js2TZgOUMYoE9Wy/wAZsQI+Vr2klDaNoDfg9nCQGPNPZ7xyc5s6TiWFPxa
1KlGjwfQn1NO+gM6tiaBlOJW7jp+AH2ELYss/V9nULyMpUgzWskgGhtO/T4Dtm8Z
KxT4Fnex6pskq5ox4r+nVTfnEFJPn1HlX2imGIz6/qJrwzTOFagpA95jDSQbkpOS
nys5zB9ytP/zu2u4NrVP6htV2VcYdEl5jbHqxteB3AJzN90wKPwAxTzBSPMlJlGh
0LA/3dvtpkpexnl35ryf23H966jH9ALviPFOmFddB3DKFF4rY2jz2F6Ps1AbxrrQ
prASFZo4wl8PHhaMisBtFlnTrCd86Sww/fq4agSLafvcxTJHrFZ4NWqTrUm2ifZf
wbLspk47Cu8I2yxhmQUWMX3yJS2FEGsNHa3Dy/ryrPjEpI6e98Px54YihXZJaYIn
9U5ajOLXcJbmpOK7uK9YXjzCrs7lQK2YuVjl/Frb7MYqSlr+C/iExW1+kUyeYNnz
4CvVlmvWjCt2508NFVEdSLlAPTdtUoy7OCMTCYZGGzFi8q9TMmqA5Bk+HZieepQ2
l+7lamHJ++Nxf34Xt9o2muZ0orsNTuKEPcaQasCCJucWbWDok7Bo38SaDlixwFoP
OUMzI2zDPl3MNCvFiw2ex7vlHGYJkk1UezDGLyL9/3EPHUg4iIWYAqQ1as5kNKnc
06xjYZWZbj9aeEnBavw7z+7ntTU645Qmqc0nu0d/mUNadU9K37c1jXdM/FvK/Mbi
wQz0+1WSKpYTZhA+cpNQjL2KNl8abtiUqjvb6gsPgQPWf0VGki8aH6uuYwmYBRPv
V9zsNcZpwNVeqZNTUJW8d9ZD+9gbnBD9miOizE5zyFHeG+pICYGFwNv/s7HKY3eu
LbBniXAMnCiAzug5MoMetQJnzCcDbPe6JcGlvxZ6MsC0I4NhVbnD3xUIBa3KSDeZ
FLs/TRFIfTCIWnaDaHPGHUIBJFeDHrF/Fx+pjZHGz7bcMB1Xcjve+XjelR/Z8Cnm
HiMq0gl8/hHL/jXZe+Zhn+kB8Uy8DLN/iNEtB/LHU5Hs4NPadervMLpod59YrjXm
7idoBW2AjxWUZ1smitIW0aZHpCe0W8J9+W7MRn9xw/cgUW5at/7NJku7zI3Z4qMY
z6gOPX1LpF+7RCAos4mAkLPQkm8SqcLE5OuIUVV8bFeVnW8Aw+JrEJZCF5n/0Tvt
+gSkHvTJ34LfCwWdVqg529nx+5aUolm2vA3biDGp8uo50UXiHfKe+yKD4WHVSyi6
RKX+qpIpuwT43MAOqK1kKbn98Ql5di3AW5qC/GrNDcF4FIQceoTcoemH7AjsVANf
8PJU0WO7KOabcJWK8f9BfXuPIzZ9eqtHREYGDsfZyQFs0dAxxPqKZ4tYihm6dQIs
bk7qNfEfB0KaQkY2WeSw/5UxDUFOZ/Z+EfA/Q3dOVJ443yf89FPaQOnNIpAIugg5
q98GmmlDzaZyDl6I1CK8kO5YoQEt5K8DyB/Do86NDg3EdDhLvb/YwjC81jwZx8yB
K/0ODk3I/+QUg80QlBS/BiudHt0rGQcgL+Yfsj36Y+lWfgA8Na+TsTb0QNCS8O7m
MkWBRehJwmjjBrngICcGzPshsiOmf3/8Gvz15eVsBQei1L0lwnz50CJ4nYiAS4vt
NDZHrV2kbIJmsNivSz9MWMUh74/QC1LprSec97MCpgciEGUFctua0Msei/TtQNVi
j2zPpMkNUkOc3GiOsH3Jd/xzwrtaXEpTWYiuiNKguqT5/EAi/efRNGhWjI5SuxmG
AWZCMnauDuQLfEScqqu+kpxrMAxP4TVcrEzoT2TQYgSaZJ2nOiGxhGY40oi55qmo
pJ+nscyXgPyg2caSsCd4lc4YItr7H/fZlWUPTppgBU0P91vrzWZxDpnWykNlmh8g
48C1Wf9UMnAuGXCiOGi15z5Rb0Ql0aIPUZDAJcro8XcD3ccQL3qynCNrUqoPpt0y
MxcP13oHM/Kc5PFCklzEPFk4rWjnrBDQthiH+F5gYz8DjAVWMREkz0srAEFwj78v
mDminm8heO12shO1hAWG5VQ8noa1j6rQO5XZPmKXTk7Npig518+UfNHjwcTWf+N8
4TCerCzyQ8Hx8lTvPEv52ytsXQJ4Eicm3DKgmb6U0FeyAGOWXjzrbR/omjMVZs+K
auXwyqhSQz4bS/5YD6jekVy3RJwUMw4tdpbf8/GVZ7gSV2GytOP9Krj9vQ/RvVIe
W6gQkA8Y/pl7nob/fTrgRCBjXspwfOhLKf8RDxtD/PdkW7VNk/oWu0tXk+4QHHRl
+Fdwb0LW7QUV3ZvORItzIn4o2ujd1DNJQemzrVecpyv7CJQrXcrD5kECsS1LBXqt
GwMRf9MMgrrczYBiv/ztAlSddOERjgNS69MQ3kf+KuEtV/Rh03on4wqCIzH2XJBy
FC/AnPuF98MB2EAG8WxCVEJacozhUSdW0MF92UbE3+eoaoUj7mvX2gE/tpeA3tTh
9OVglSN9YmPfMES94jk7UMfjBITBilUgyd5QQRpeA+fuJ8tkupJ9C7tPLBkVLx5s
fL9303g7G1B5dOmUeoGBbL2+AZsBDrCZCW2vxmmmtIS6MPGezxiCiJkYbSRwqFI5
TE9WjlOZ1hxFuvN158PawXLOvLJtp2A6Yh+yrDeEV+m81xgUzshBLnytzrotsV5F
z9KeiwCPfcYEGuroYf4OCjAJcsL3w2c8K9EPhqulXQLH6iyXfe2Wh5VspCIYPPlI
1jA4y4yhfaXsSmaGo3RP6d800Gb9GNOhJVCo2fDZQWkqX5hfFtrh3YlDwxw8Rym2
stE4GkTinqFkVy0S/fPfySqx96cv33qmgRtWVs5gXJaQiv+Kyf/8YQEJ3a4J633O
JI7mq55mL/JqKF07OW/SGYZ/s8cfn31W+hFFsh+mH+XONCsQNDvuh9MBVl/EBICF
BVds+/Pf8xW8wxyQ0wD4InJeKVnnU+LGEhxjMdBszK5P2aQ0rLA1BUfKjRE1kxJk
PQu0BzQLrsV2DpTQ9smU0hmD/3RTRg3eCZuY0H1OqDIUEc697ZVAhyBR4Iz09MVT
7hsABrFe3QiPf9vpcKX53u5OpUIxHvS/tk1fTg3VZ6+pRz3Yqn8cLpQlpeZ8ILEw
fnp8DWxJkSmXE3yuvOMRH9BpvMgtvup+I91bifdYnyUIM5Y5Z0ZahIgkXLSEVRW+
RWS3HVyNJXFtnqTRk05kE+EGnpkgNE5pMWWpJx30pqQ2UcQAKOY5Ec4jyeHanGzZ
LQcVh78FW5XgmLKzFo+rv5GMEkMml+bApFna9g2qAP8asxHODmjzABtPpsJBi0xW
J92q3vxPjVehOfjNHkR5nofupsmmkYU1+/1/Z2ALgSM=
`protect END_PROTECTED
