`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
208B+PxFox4OcU5c2CIumFMqEwGnPJqWRpadBEKUMiJjxy3aDU9e804IQPekcXI+
crtVyorLV2hOPpcBtUzD03ZtejrhzZkDy+rzwDNla0nxABrcmbC7atDdQs/qFixn
xRrHOg+OffF0VAIp5fkRvsQtJRnZSj70OFqf7tax601KqS+S3wUGqvazqI956E00
Zrt4VsLS0lyTvYQ2SAKEaLuBnQivd7UNCI8OI3CB6bLKn22PbTI/XJUepeKUhptc
iNZm+L0/N3QLUS600qdbINROKIRjOaH1+HCb+5OMWXxo886+NrL3i8KhDIZ7otRk
T4ekGQn6ibFuSo1+GW3UeKEriuxCLvTi9CyJnNKlUA4aaFapcSUEVt20bJL5IztY
Yf2UeBO3VzupV+DZ3Gb+wKCqAmTnfLSDFbvQeYTbEy+Gi0yVeDmu5EjRXHermQXK
v1XdUvz92U5y887LgkWllcmED/g3xRB1jzCZ1LVHmvWoSTFLCzup66Tm+JDAeuW/
oU0wGuu0nfnSH2d3bXWVfpCdRDNzTp8mYCh6vrgpzIp8U5X/v2yURxNinTMjSW28
sloexJrrx5PGMhBkhgkTloepdmsGPY8zpdtiTMU/0Xmm6X8cwNmlwMxOSWxfVtVc
PfJIJ8x30w9Bh+bL+BEY2pZ1zahfEa7NXe3UkhR508MZQsO80ZYN8so8a8OC3EqG
OVedHFua/xwsM7/GkFjd+uHrRLrxh/Mh5RDHDoqOexvGBv6ltLVFa9EGpGKXYcG5
vxEhZxp605KNO5IQoKlRxdSEV9bWnDjLJJDBCAdeUOyKibMbfK3XO8ZYf+RdodEp
6UO9XZFy6BbJMPdKtKyKgWEeB6dKRJzRIbefSxWG/K85AE5x2GiVIi/umIOM+mdr
LizHPhkk5YrVf2ksZ9LwIWp/WPFVNtnb9pD8CxhP6qUDz2xPolGG65iQNU3ZAbLg
n6bvkLrQMQx+j6gdKGS5NX1WP5wjIUhmZncWwJTc6GXTyBtgm/b73D4CSDy7iKQl
aLb4saQAB+lsz3XTFaXy+qAsd1an13G02ZufYjAFKR952R7oA4V9ieAMWy3U902r
SaSUrJbDMoZ1K7kdhQqIf5B8i+uifRyDfDklBCJPMON98wmruItCIJLO7wQhj/xu
U2dRoPqv5Nh05UsM4IBNfG9M8fLgj1r8zSNrm63rTKYWGamL4xmdM+34who5C/jm
tUTFJb01e17uRrGG8+Sq2FLyZDSPHnPKxQtHxraBoOO5sGR1msmblKwr/c8p3HPo
8pW/2/GJ0BqKf0VQVGFZK/kKXLvIq7wKm2aVg4hD1LpOIVirTw1uaQOKiPdoO6IR
1Pa0ftOxJ/6JAbcl36WZEve/7JTvq0kgKtIfbGeoJcyEC+2k1Vk6AJ9VMLEOLUoU
T+bU1gx7rPsVGagygOpVaQ86rIAIIajp+v0pVk8RNSQ0ME+LOBJPA78ULlVX21LL
SbvkHb21/3mK+psumhWfJNG+umRJrQ0mVV6k6pS2NXum9OcUmR4ztU1hHsFOl8gx
1foAmAYS94BbANW42b/Ja3VycC2HPT6JXaCVIBTSL94z88a9FVCJZUQtr/H8ijQg
S7g28jQzNwf17fMetrcsPpaJWVBOFWdPCuZG/0uUxDz3tm9xzoZD4xO42o5rIuMq
Pgw2EeZYjFddhKddpUFufn6HdjESrcmoKJyFzUZe0cQAhToRys11caz5YnS/HpKx
kZPUvhtRCSphAb0Npe4K7DwLrnViXS81X9nUSUbTC8hZlsMGTuY929TUDJ5ymzLB
pkWJ3jTxro1MXRGzKz/M0dExWDEDqDium+owhlFRHJx8HjxDYNPbI2etrzF54MIQ
hX3BCXEFpYLsRKzmtfbKKyxnFUjHE98p6QnOtLaufkNCnD/+mlwoKCpk+Wrotr6N
RyLKXZIn4aXwT4Qq8aqBtlIS7OrSt32eiYLO8B3ioAFC18gpLfkvomdmSmR6artp
HyvK0JfmWID46g0tlZ//H154rWAXWLrc0XdqhzqEAGrHu8v/KuHfJPjBD1r3it8Q
VDJ8zr4lZv0wtaiZ2tTZTujLnEyu6c3/WI2TrOeUYrE7oBHiQiVOjfgAnnf76egR
nOPZ4sp6gaRrFHk5ONc6DCvCevStGbG5y1Uei1o3YOg=
`protect END_PROTECTED
