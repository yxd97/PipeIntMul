`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LiwsPQ3UZbyOe93cvXADq15RC6yOqGzf3Ug8od/lORzQC1sDzwuB/QqpgvIY+DUV
rxfuulF8EkkQGJIR900eOtT9SAOTX6TpuGIMDyQ9HvoGNo2jBt1vfZCFAf9eXZnH
MGXe1bOzha722VhVnGY5yfxOQq/oWqPAI5atbYcBrdiHR7z+4gHcI+nkkK/9sLWM
qePqIE7oaocJh5MvEhZtMEWOE1+IQf5Nij/pvT//OhsaEDboU7Blm5y55a963QwA
zk3+4p/OflQCRjLenskSLcqHHe+vNDmEA8aQ4Gb9UhgMMTvuB8ZQundmV3KE4Rki
xzqq4LPMJE3vqAE2razW797Hez00QC2Gx2krl186ewRD3MADRBIvsD6ejg45EF8q
cp5KvrrALpy8hZjWLDue6J5lRhhHh+pboePhI4rXWDtFlIFzrSFKHrGdBHdzKwVa
4xNHsJAh645bgDIq2LeEXYSiUQzOma0+qN0i2yw6/eY3GGTfWEQqcgd63r12t9FR
jMo0n0Nwgbq+TKsZaMghQM7lGVslqsSx7IdcxpGNCK7rlEfHe/pwcE6cuClDcwFV
FZ1cdbcz4/EO27rpCT/gJI22KCnMBQAL8U+XAXoWcAQ=
`protect END_PROTECTED
