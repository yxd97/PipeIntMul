`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d5QbKh3JbskDCOcjHJ8TwEX4WOeb7aZ8tYvgITjUBP+C5W+sjCTVxd709ZPSV/93
hduqTB7jhhca2Ppj4RrDmVNPWPv3DOcWbOZoWpMH4ZwCIp5jU6kvZkH55cYMBYa9
PMgfNmOe7nqyHX9G9Mm7nsEw8RThS/pwbK7+eu9A+DlIJznPwnoz06vvhJH+sJZy
BFmyEWnYA+qU9Io3Z0gSXH1XQlwNap/US0gWBQwP+Fs+DYmEMm9/2Jy31EnWHTmu
p7SuEvQQn0t8ynkwfB55nAWOY58LTmItuXajK6mhksHRiaAnEFKCvF0vgYfmJpM4
zQ3jKVrvEjp6X4/8kkQZFtbuiNvxSthSGkzO+DE8zBb18kqjFwPkLKHn9jmNSIWL
6elQoiRXfO9QKf57YL6EYHrPIciNjyQ0Ekob9dtjg+Si3SAIXLBwA+jBg9KZjcF3
`protect END_PROTECTED
