`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7/xRiYUFH4ne4hJjakm1+Zfek/vFNtjtVoi4rs8tJr6bIcYuijrjs+khSUhmNEU
TXYGx1BDX6xseQO23n5jTG5jcADEoUzSBysBp3p3FprLIyaVgFupXvSm1ehp6491
2FMG7Qh4UFfMfc82k4ajVAI3MGnkMy4aMa3uqjZNPKYUPtGJfT6AMAOdxxExgIqS
IB2PKk1dkzZBrxax7iqQbJgg5HvjCaGP0prgI+g6qtwgFryRhQrQ7KDSWJLKXpLM
cK5+Eg5HCKYQ+mw+LY+zcMNaDD5jQlhjugW1Rf+46G3nJOpyW3g01cwwAB3B+Ga1
bCJq0WCjYtCEmeg4onxKEYV2V5qD7KtlxOiqt3Hs/xD08rVbVuNOQT3m/C0WbLrS
7SHdhfK/doDG7dmvHuzJ6jYX3q4JHXAcDJifcdfC1HN2uDRnjOUsfeSjuo2Bh7CN
`protect END_PROTECTED
