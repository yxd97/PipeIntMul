`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
igQcKOuEgzEBJQ/QRACQ0X27ztZ56/ljMEfnqvgDoUDIsoQylkc4h3DIys0oq8Ik
TxITfx8oO+hl5Di5bhOFQpsbnb2HH61vAQLJ2/jxZX0oUZdpjzjPbrNSn7YHFO9L
JDA465H/XtwnQGyggL9VwutsQhOv33NumSe0JtLsC5Jk4qkGqwjH04r2ymVE04NT
AblE9YZLtAGU+t7IxNKRhhOVCg7lufm5TJ1b+FhyJ5UKr6hb12Q2owreN++GkvZn
eWqaI8VYUdreXvxEMGfFQbSFw4tqR6fqQEf93YiVXFDK+pmw6XI2MN7ITXwirkpI
BVePpfFPsygPq94Dtx4FEVQcoZdm9mlfuwU+BIPHliodAk//IgfvwcOvzaLX3pY4
3L/y+CV3YpnYdtUghxREEns6PJUu0vfO23357c3EBiw=
`protect END_PROTECTED
