`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZK69fDAHVvaFTDqOu0NyQH2WFpAi+jztpzfm1VHxJ1aXsfiDV6frLB2tX5Ef5Y4
I1ow4K3b9ZYJsMjqb3Su/IVB4+C94HPfJ6hFmyT1PHl09SX3kJAT9KaW4njR49g/
5E43ydqk57w2JxSCMgJT6U1eH4mCQTk0NXXyOZciEv4YvmVBcOakHMW9O3X+7cP+
kX00WMLz5QgQ73+2+9gYKOV48LlMUr94qx+ZLY9GteHLcTir0iunR2vnECHEJmFB
6OgtQldNWTQSShUZ0zTx+U57LpsA2kC2o/H+KGgEgf5Q29ldNHHROJISrmc+rLwt
DMM2AlR6xy414haiE/gAwvxxpcNDVDDbka1LAoPNdjzd/3A6eQazoZsrUanMXB8F
dIENRPLx5oFOwHNcs6AsS8iI+swUB6o7Khr/YKifUSqwJEp5YPCKDrvl1Pa88k0X
OsFfQ9xSIr5zxNnksmFazHrKwVsBYouk/+9jpYnT24xdfc6m2b8mlhse10zI454P
g8Y9DQMb5PGZ//Ek8HBlWFSNZABo2d9omwUBz43kW8AEwuNjal8fRh/ynOupta5q
dgHwpbr0Op2VVPtCss5l2SAgCX8UJ0Yz1WDK12ObsQWVe2q98fcSnfhgeiiLnRzD
xJ+QzT0NwtradErHFm5patpYWWBqZNos/p8hLZjVUQ1eCmH2ZNr98WjveZgNREfB
`protect END_PROTECTED
