`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RajpS3eaNPuNIKj7k/7+d+3eBwcj90Q5n/mJD0LMJeKRodcw7SZAg+RZ7M2dmN0
ilKgkRL/Q+U28oWLZevmcL/bq6IK2vBfOWSdcIxwh6SaX1utkEgiXmqnf6/byNaQ
ifwvqO9ptGVvhUBGfdbpXLfhstp8HbZBZip32DMjXITbCgr/xdLn/5X3mYkLewXS
TyTRzyttY2YfiAx9WmIhB8u824SniekqX1X7mHHyqxfMpbE/xp0HaWyANXK4+p+V
svFNNy8Qvp9aU/iskLwYehGd+hv4pJVQL7NlCkX9N2E04x3BR1BuKZe+SgJYxRjB
xrugGblXqUBaWLoBn4tcBzBvr3HsvjKgZD0nf/4yIbmUpQsI2drxxfMaiRKAOFtH
gfWbxRguMzVO1Mdpeht9ji3z7+eQnITg6DPRSl4b11F4LMadNallcCOmDpr/Kjkl
9VrxCvZl5+o4ugOaHujynaodMFBGlJeQLmOu6bK+qtErQxlMNQy2w5nrAb56S1Hu
ltE07wK6kujtH6ZJs9JdvuhxLgfLLmFCNTQkBkNfNtTKbW5FGgRgJeGTDaiw2Ecy
Pj604n8ptoZVciOYe40PXvU6EOSYd1t7p0K+NGwfSY+NRArZaM81xSuWEbSPyf+Y
C/7dOGr6Mv0jqFLSRjn5k+530D7qeQxvFsP4eSxegAZAn5eMer2e5NaVEAp6Gi1Z
behMq+bGU0e42hv0qiZWT5wpc5wbORTAR/kDwTvoqJXmmu+3m13vJtxVvURdyQ8t
kPiZjcUf/bJw6MTuH4eIkgbLeLqKGp1H8n/koJICjAMxS36gMlUbJcSjlMbXEoG8
JZ1UG8+57Eku4pFgCfOuAQ==
`protect END_PROTECTED
