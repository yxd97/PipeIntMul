`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGSEFZfm9g57KQNV10eyAPqZS0qKGuJwHyJ6i7TpjjErYpfJ4UGCa28Azbrwt/Hy
fuaqZLBagWU7jHIwLQ16iN+Wyr7O4heSbJx4qW8KlJDnoqeOSJMDVbfgCl3qOV/E
vCHEX0Ku000qft5k8z0mYnbtdnei+laE9gymZDOP9f26us5HZgpaQRq+JeeqBSsV
wQnx7fWhGoMIhLwi4Hhs0TCRVwA18wREek/jMDWBipX5OuDAfUYhp8k62NwTH5Sx
ZxtcUjI6kAj96HfTMtbYujAdDsAKBMRuy5juSNZOf2pd5Jma8B7sdpL70PvwYmqV
XaP37T3+ji7/IxewPavelQQVZLAHlMc46JMxKnR6PvDYOn9JWMBiZLj7PTBjrPzR
tGD82iqsaXKhk394oCe6Z+jeAS4eiGmkIKt9/YCnmtwJNKxspmT0IPGgsfXg++Oe
uOselsE02NDDFtqP4DwYEo6rF1YE+wRYyOF+NZ82iJ8i1QIuBjUeFJH6bhmw6QxW
algUvyaGNQ3AAjqpcwoB9oJoE2L/6QAiQJ2yJjw+GVR0neS1bRgF1buKhhhSylkf
BvlvokS+aUOY+7AR1TyXNolB3cDw5SwCOYZx4IqqWIIz+Y0XRUtRlvp95QnY9LUu
GHVUk+heFLK8Cwtnt9xPyJ2bBr9hzJkusj4oUaJV+JRDQJ4aHCxpOrfdzBnPK5wl
Bv72FpHYLd01H7Ff/sTBZAr7qUegIN1h79XQHNW++1jugPLyeCKWwaQbYYgu/apj
qNSi7bEej+HK+lKLz0nWaY6Kpwg9b49pJ2cb62zZmuiBw6Tp/3HdqlbifBY145mP
JuWDG5f9+cJkpIArk37lkJlQVpj6IUTOLP8nrjgj0Q8zV8o3oo/3wyDOzjXOehc3
b6rLYcTGatFBeA444098Q0j+Bpz5Se20RCoopdWMjQIEgbns9ryb9evIqeDycdn7
FSNpTaOFCSt5Rd/T2toPcOnoFcGNJvHozRSFVOwpIWpxS5BUmSd4bwgdx2o4k+vb
3Rwlk0kkqWNwh5lN2l62rKem0rtqqmngWA1YX35r15buuu4KLqSJqzGpqN/5w1Qd
M2xHkgibDiUpCo9Xz5PGDqDNltLmr8VpNJIUS2F+egOQG36k4mIn1yPHUmSn13Vi
3jQiAO1hMkR2B8qwL9ycp5502idU2mjXKFJJg3TvInHJfVeGETtLaskOJDT3c6zk
V7llHiAOr67F7xLfR3hB2uWC5n5KqHn5IxhWPX9HBcPumIeKzYTcgEy6i84dpEBa
QZhMkH8oobykrMb8a8HMZfVw7y6mTwYvzIMvSWRXnckq//kABFEd6Sykhn8gJ6/c
zDalgnkh6k4foipiTbqUxobX/s9DSXXGCIqwnrRz8rFUpqwigb+s2sYMEoHpDEgc
tzcqkm2W2zOfiZmCtbBhZLN5PB6ZWm+NVneymVH9E4dKLXIl3qESna8Y0RDsCOEy
duJQ5wX3wYN4/dH6g31pemwoRQgVsMO/RSwl8YM7wW/AejHplM4eI83pVgqbPTgO
nWIpK1aOk4+xHUUP+WpEm2eqK/rZvMxCvg8EmBYu38Fesnp3HacLRggd3wptPQEE
mWKgQaGUVV78MU/rP2TqtpVdmxE8SC4ktnyvCbvUH9ct/pIZ0rjiyx+Ai9IEVppG
hagNRi6U8hOAKNIZ5LB7lEqLcHLcTpYNoQAJixriEHXJ+BdiTtRxL4xKpvswKY0f
cP1QgJqW0bUxPCjmac7vIZWyiJ1qttsdctVp8fPdbkJaY1j+JvY4irgtGr1OR6wX
FcTtbOgaDWMfQ+NjNyNcY7HpYBJYRX9YG+6n1elggLOxSJbKpAOADLJUMoYV68Bg
RfjnKdNEiVu1G5w9YUYSHCA17jW9mxCEEEgdO8Z70l5NhLTWAEU7BIhBZeeHpFFe
tPwVYIN4od5SdC3G9Q2I1tCQxWnG4pxeVD1jhq6KQ2cwbszY3MH6FYxyh9tZyXQ7
h0sIKUBMcQ7pAYC30hbP96BVk6icnZnJrwnp/4DIjJ4dVKzul7rMyqozQxMdahAQ
4Fnw1MRNuz/utVzoPMLc35gzTPJWDRHVUsCOTmoSFrp6HqrTieRuozzjSFXkrB81
CbIdv2BJ4Vgcgwj7FT0dPA2+LWYCOUq6dicvYd/vXtL7wsOiDjJrPHkNelnIRnhy
XJ7+gERsigyWHRd8tiQ9v6Hg8Ui+M2Rz6XwQ4i9puXq86ws6ZnmQllYBglzUjYXL
peXIHGYtSprpNxyk/N02zsZqtM0EsqBJp/wLL4Kdsd4wRhyS0xw2f38UoieuUm9u
SRsyU2o+TVDWQVf6ldBcRJuCCHMNQRHuWnEzSpXy/BqSfFeJZqFPbjyUBrbWo1tX
v1e8wH55H9AAB8lYe/nvxqueOt3vylHcfn4jRD56p7FoJCEtbKR3udzYoKctktpu
WJiRnyyZ+oiKErU23AiJOLbSJaDuE2l6YfVBb1BuwNYVkMa7ms3DzP2QSYcVGwqZ
I/8agbWuIcvzBx1Fq5EaWuRQXxp3kOsdh400MfatcCG15uaCLYv2V1SSA7JAXPRk
7gjkrRsry/AduC/BUekqEun4K88D/0KaqM/+DBP4pEhk+Q6FghuJdxNyBON0QAq8
oIA39puJCkod8+Ky5qfEDts4tAvSdVHdisTVgGeqCM+zz+boblqhtcL/Vgar5M12
Wb320PDjJet3QfGRP/mkvmiqm6eAk/xjdfOc4CX1qDXlcS/H2ibJzNnaKpDjtvHl
a0fR9JS8xET8itFMWLOhWJtk5mdqw2Pb2TrbkRhXNr+al1sbh+/mvtq2cwJvqPCp
HTrMVLMmOJq7ZUmacZrjrmd08oB3Zi4lLJp9TX+QXgeIzITNplOFDH2yvdzGAJFl
X8JDJDxJ76tgmN8GgivQgqRDF0Sjcf2vMQwJ1lPQko3128w/v937Jiy07YAFePJF
a828H5ZcbrMlQWP2v1qiAUtwab5M4HjAlZWIlNM1Fwu9WvRc49V8JcwizzaaAsiW
aUMIwOzUEnghteXR1mYnEE15XltipjoXGHrjpnRQYSebMAh5wBYvt6z8zVPTueAE
omtYNj4yt/UOKQs/hawq1vMbos17ZeGR5ARsXhz5vF3D2vHTjboUFrxxj51PVe/s
mHChf80MSuypoIFPJPAccNsfgB6h+Sm1JAfNg39e+Mpj023vZUtNdlHojWZ8EwtJ
hGpEPttq4bcbfI/WTVnwGgLh4p8UrXIOWlqGtr1X4UqLF4D9Fp+cl50+CQ47SCzF
LZk98CcwgKw8Nx/PsoD2EcQQee88ynAQZuGbbvVs+z5gOgm7PbSyX9IWM19aWGpz
oFEwLuGQpgf3CKrn7ITX7HtueyxZWjLDUm/b6MarWBVQlnoKtgQ8AzS4BiSDxb0t
JDrNp7tqNE8SPTm37FNekevugrrU7QEupkrL+xov2oAZKYJ6+q1u2X9XtOX6WSNy
1Q8+t8DvBkIcFvalaNkSbAMq2A99BCyj3GrvlZnKfer5AhNDI4cEQ5FsGGgXTm1I
UvR0VgicHqycLSxUSp8g+17Iv2t1Y/2io57IlsXA7tnsbA642erliU4RDy7eZXAF
VqF880wWNHDX97Dxbxvq4MY1DoxdJikUMrx7ymA15gq3ToqII6c14CvEoyY3/wiJ
dC+JExv7t4b7dZF3R6EbRCrUx60gZw/IMHq9nhZl9o4BckNzYxuD83XRUH4TA5sO
GbifqjTOo/Udkz3QVjkDeTd2CAm9HtoPrvms8vlZ5HtDHc605pbBewv5FbTg6zpP
TGKuq+WhtOxeZW0elMhjORg9k/oVj3iiH5+xQsZl/vkY9tkPLlwNPLQLvsVmkjFu
OpRcdLdHL7PQR9brU95diNVrk8zPs8+aafXdHNwXaAeiPj+WWn96V0pUTXrgRK+2
pflu69ypD0JC2aburvLrzzmGr7iiMo1DOl3ZOmldFdEFYwxPk/m+hUMvZLDG7z+U
46CNXF9KkJ+Hl+SGKVVnyofQ4oG7B8OkYskLM4tH3vTRVgSScUOWgaIXvGfFiiMd
x3fwWetvXhuzuCIWpM5jl7Ar4etZlahiTjupQr+upqfTWp02ptgYw274+EdwWsyI
Ojx9tXIM6AV99/6J3Z9NT27dzZ4x8h0piWQfrhHXWbVTaU4eyfcw94ZB981V1S+4
nIh31xFU5n3lXECod6rmU8sHa5PWrR/nRx5ipkDWi79eYnumprm7MC3knRsAILes
yp1XSvlN4t1RJ22bdVowT+W9XJDqxr91hnO5y4t2uDsUP94q3T9/nWr/Gy1+w2cy
TcAiDzYGLtEk1WOwi4duQnWIHCVLnYQW+C0it7PTiTEohbqiU/31lSFDBQREGsT2
tbO5B9hwnfkyCnyr87+Qxs/9ckqMIBiDXjQYHNRpcEFNQ/kb/COdZtk3vsSMc0sy
6hWUn45q8HKJ0vH1cXz8VBWVlKuD2LiPMQEM86OZGWcCTPQGq1kgXtzfNUt+68cL
13dHH2A2jDKgVAkYsyYdS290mlL1c7N91m20BGlEwjQmsl+sFAecJBoQVBwulk1o
M+vn2j0IweOFgS0BpBGKaX9jIoxXfK7QZqJIN2kEFLCkvQxZ5s+4iLWs7wznquyA
Eg6n1Uzg9Ltt4omI5rFQMkmdgSfpUz3j0Ux8i3lO7MYpMsS8+Q7YzGvgtdZaypV/
TH/dCLrAvwe55ltiCZ10nJmpfELfoyUcB6O58dqmHASfv45OCJFZuB+reIIH0ZPj
bmsDqzwPImUiX62Qcaf1JFGHl6JXicyylKxUK/kexPaFF7roxDPcmZtBswn8Y0KW
i6Ne6rFC09H0XJeC6k2U+qCLOwxz5Dq3232WdcfVHLR+H9PTsqUs92Gw0Lw+dbKc
jRBk6IRlG/9QEOfjvnL/yDczRHACbKypaXYx9HyikfF/STt78Z+N/cfOSsRfbbvm
mnZ4M+BZfihFWX7pSkvR0IJcBL9z556HOP4laYx+BAXhi1eJZYr/vCnxUB3YT2q2
FdqJBJCYv/cwOjU/KkuXcwxTtQE7ABSVshi81lSmA1iDsKRiTXLucSh/vgaHno4z
ikP2Z2xe82p8zyxqxPuBsJ6THJr4ei7QqR0QviRPe6dAusf93m9FnGZRRsBPWnvG
hC+5V40H9+Fnt/Qj8jYzW7dCapu5QZeTHAQQnqq3YnZzvJQjpp08joa4W0wyNouv
eOWO3tVNBfadjYJbE+1gnLobOWF1eJG6Vya+IBUbLEyORBwuuOdxz/3+vagHSh7N
y1kxYUgMtMBzKBUYWDdYYxN88mB0zKvmpmKZZyNX7CmLdDV9Wjvv5to6uoRZgtHJ
KpGbjbJUiqKm5HomP9tJVJw9B6x0d+4TARq97kN5vU/2A1BiHKBRXk9hxJ5be1Iq
8K3ucgS5tqtx3i6YCGMWS9wBBIQMCoqU5abOYXA8uBZMrlbzVL9aLunXh7HUUwPJ
eh/LszYuA9a5o8iDWibIS747sYEqkoYgRfiA4nMjZizuorGUlWXXpzIh2wbMpk4Y
uw4Gie+9FafolTdnU+wVadUvyjcNjky28z60d1l9SxgXaSLKQy778yzpd5ygpVzq
wJQNMKuT/5XQptzSFgYjuK8jWgoIHl/XkCuHVyV8R5IWKSc6QSIpg9ADThq2wDcC
H5G7nxxwU7INxJy950zRNnjVG1FMb2pTI1kOEbV0PsibVWgfjeHmcBV97Aii4MgC
OXF6mnMHz2p58IueTXdbT54ma9L4Y296BstNAWFUPDyLhxilVcc9e/pa0gYZGIHu
03xrId/KKIP7DOwyJe8gbrpqwmG0aF1mFpkOVMCXwEHH6raQpqV1GrozXhf8hFPr
VBhOE/k+rre0dQpxkADhK0ZfDDGmUDRjI0gl50+dB+nc8Mc5869VhICcNxbgYzZO
feBVIKju6oEzBS4TVUn2SE2YzhVg+OmUER/iRGffvWWYH5iCcosut0uKJcxHZueV
I+/QOWv+iBo78FJpdBsAgYoU2DTodPtYYDr2VrWI0jZWBooMhhoyxzpNBqkkLTzV
vzYgITqEui3g1YFw/qxty3tCstXe9AQgYgFKT4k+XDgSikv/RK3tnsffyISBGZ/i
E3+DB1v7vQOZwV6a5Q4PTeZzuQucEMU2Py0JsjuXzMj35oFQnKOHuJs2K7zABECW
fwCweglIP7Lty/ITvAlyofcNzUie9Qe4Zohnsnjy/hWhRQJaL+8xy9CgchDbcgQJ
+ca/r7wJ1OJfAovASHJ48RK0IdCvGbYvSePi94jkh5kZWa0N2sCM5atKArDcn20L
o2sveyBE/VyrMSx8JLGGkD+dSmF0P906R9iju7v1MNO6d8GplazkzoL6b4oJSltn
xc6VQXFc00ONeQ1TWOxYestwDsciqNLLYwPS4k0ZuhA2b6Dz5WWavgWPM5G9zzBw
z7baAEKfHMpM+qZv6uu6pb5WH64WDl2a8I7zqpEkKVFq6FRmABu9HIFq4Kc2r0Kn
Dcl/rPHbLde+B2zjAFERKkVGKlayzACl1vfdGwHeFy5XCIyp8zr3Y9sXSQGwDbtr
vG/EsH5e/stYmvyMQrzHnd3Q9qhNSJEBA6cCzAW1rOOZzPAQ1DoIobWu6AoYF/fU
/7ilHfLD5XOnKgVo126qk+x8DycWsp5VESvxA9DzyzmrQ9JwcIgxQ/lK2GzXZknc
yi2KFZYRg6Wl+5lPPDnYflbFoRCzQy5pbRYAhvblnnsZ2+0JbE/OjmFCoU93S4aL
SePNRQmV3mRwEmDRNTBTVeKhXk8Wd3rsjclvGVeVi9dxtfcKAGmcLlmz6WtkKVhQ
UKheu46g6/36OHglgc5Lg6t/OEeF7bcqUo9w+s1ZSK/HXqodkc0mgjxITQOm1feZ
bn+1tkA/f+j2poCDgb2eFvR2xRSLhfNsFN1DpKasFVlxFDZENWJkUk3deB3EVl3C
ARj8UYS3mItGJjMEU5Clyq2bcLSRGDbRbjFaMXuzugGlCl7VOCGhzSPHmxEX3RNm
HM1ZgYdhszGRRGsnlqcDr6N59tb+NHoUO0xsgLRqDmT1YW2cTIk24vJgU8YaIeH7
vPBlLSV0vIBXYE80gks6XdX5xpquyTYqQlkZ+zE7qY5f8GiLKVxYSR34azIfmhnb
xEIS8e8a6WHQzhbImDnPd4jUO9eEV4cfG8VTWeIbE+2aoyahPKMy4lgva87nL/MZ
Qju9UNscz+0/FUnFwLPdgGOle+xO5HeaaGQms9F+Wa2/fp9gz0WgzjhpGtdV8d+0
Dg+5Lmvcc0kG70zVWIPwieD9UqN8+bodovn7boHlOHcZQDmddBmpI5EmExYK2pgd
ldub3WsohRijnrzniG0eVuXoX13VVBUwa975i9WJcE/nlHdME6hkjS+LMdnhRP8a
VPlXKCbBYaIDnwGjHnR+So43601mXhrzrzhJn3WwsAwI9SSOIlAQWUZhvZ3Mif7f
/ZNaT4DUd0xJwJtjuVxUOpFR4V2nLjp/41BukLTukNQMi9sS11HHf88Vzzs1//y2
4SnDwNYkrHMpqzlAPp4cmECUT1bXrIUXepntKb91rY3nKqDkieLdLeTwcjIMScIl
WmhTRePFBTsJAzHh4fNxv7jZUMQdee1IFVX5OdKXQiGNE6QFSS8FXF7WUvhIO7qD
d9Gob+xTINwUqRtw8HsksynOu8dSw358gh3y1Lw/hSdkNIgY4SP/4Dt3nwhTa3VX
ORPwFDy5yeZYyvvNVSTHakTJXAl+3qxET7nqv7pTBe+89gytXv7hzSr/oN7qG3Vn
2Cc1rffpsCILcMkuLfz9YC0KJBL4XSFWT43TIZ+DAOz519//GwoeODhZ4F1lie2u
VJyXl7D1jNseyREk2uubs5PSerZa9mpm+400Qv2fGpuNIPeMNfNMz4pIakKUfmuu
Dh7EsvLrr61AXpUYkiKOhrXZzidhoW4qnasAPEKFipEUxhAiAk6l3jVBPOCvOwM2
Vg4EpST99hkhhIZ38QNNXfIU+BkWNgNbxRnnMoQx4Fz+EWIeA/Tc8j+f/bbVfdmK
llRZ0uAVbwAu9fOb2cTmvxKKVXPLZqJZIkxjlKzFkcGkU+GSiKBHfBSdw5ALgkvD
ZUsK0kT4WPC006Z6w8DlKa8EA0TVGPCRb5vmN9V+PmrUT2nI98LJ6ljxIJDmtBuM
PSoGqcutmZk+Et4kIXoJC7lOOQfanbQb+DksenBND7IH/F+UL0tmkzA/CJpQfE0H
8Y1Bzzh4xZ73b8f6BXW6DGOwmG8L3+wkynJ6D8RJthuJaDdY0keEo0fGAxNBez+H
7CM9794noFqcYITkzSMA3HkpehraLtJUV1WGANcbgMEvNipBvMuwwFz+KOXEjhjN
d/jBdZSyoT7aMji9Lp0gci4x+xQ+OA3K2aszhZqE3IF8fGT4FqLR/NVnUEMf+q2k
2fLpTp/29IVnC2CgCR69vvAN3JzqzcTwGiGoRWOSJCBzor74xtmgybfNGDSgYrQd
P7In35ki1dq1Um20jDbP3p6+929rTiY4fLeMDzr6j+nRosf7LKY6H36iaEJ7xaB1
K+dDjULpA/suaUcY6eq+imp4pz3f4V9or3DGp+B2h8ccA4UuTJK0G9CTepm8rdgC
6q1GKclzrqG5oQBOGiFhQWxmQIP3FrCobwhUt01pn8K892rEI6oOwJR0UiYxXpmV
2soRLov1WuIu9+2gLvkmafctDYuJEXt1UZsAW+WFd6qJrTRMVw0K/62zH2tMKWV2
TNYTAc3MrUel4O+IJ7DqHlBcUYBqgHRytRpJ121mmHrEZvKOjzF5NhrIq8JO53i5
Ox0phBH+zzMiotF7J4BdlZYvTVYLSJBgvZyCscNHkhhqRtph4YAn68VtFQS9UVWe
VwUGid9T4xcaNTrM4Jfs1nlmGVjEeT3bsuO14k+/eh1ZikB1cmvBPnlVBWl/SLv+
+IGg8fNG0nFOubH4MsJW23U6mDHiHQxGKNY8HJHE6JDCckuDvmPI4uD7IvYFmKj7
8OkLagto2oJ3Re3OyYhsV5c7RXcH9PFK60baQUbcNXWH0iT4+CdoC/0FBrfdKP6p
EXlj8h3CRUZQHdypBwp8Mu4Z91uJXOOhKA96V6HmuWJkEgWqSHppLPK4qgAkpuYp
eNvnaraSRdOnpL5zvFS/VPUNgYQ1eYVGCy852RoEn9HMMEX0JGJpE1KpirDLFG2D
pesOmDS8x8nAEUQ2lnsBiIdIrPqBYptkUZx72GVhVPN8S8KGRlBf/+FNjOxGbvUY
bimCGwIZhzrH/EFyxcxgqyIpxmgaEWwNtq7ubCETmkpJReapAOakcsEiQBI74jte
iZSyw5XIHpYscD7ZODTUaYLvdgi7g8aVwTIsWMrqKOVvb3TcVf5QLO+ixMdLL8vE
i+MRKNdMqeGqilBg0r2eDBTt2gujTJ+8Rfud3NiLmg2V6GrARXqbUS+0/l3/Kjru
Q3xEaouvE1R2WlNsJUKDYqouSIr6rY2xR+FVHwVD+T14I2sOYE8JspuyRSC1P3/A
QJ9XZklTzlzBEbZP33hOSA5MW45SlLeAvr8JxnDgNFD1+Y/Weh94ricoPex63+ew
076yEhQVwtL0YSel3hHwoOIv3Zb3cq5g2XOgAu9IrxN9GY6rQwM4Xw/BzGr6eA65
PzrrtDoyrETfzDdbfOTgm1l6eXrEBLnwsfrojFNB9FFBkLvbcoS7SSEXMmjZ1B+2
JCBFbZbWMV5ymJqi/hbu7IALVDrmXxBgDAPsYuq38moCbwEJi4PxaF01sU7D7ZK3
ukLychg+Nifqr+QZNP8+8OyfHBw1V1fqqQPO68X1OLdl67OF8PBqcY8rvTDZ7p67
cb8LY7K9ai+AGq2EsZqQ/4aWutC923SrK7DVQGPT4Zb/Lqesnaofv96ATFrGg5/n
J8YaJi1/ud2OCmtfNZaOBtaxcAAN2DoVEbVPql2ConFKN7FtCBseqlx3gZoi3TbJ
azNZk+CdBuuFnj0LUaHDKTQKJu8idcQpy2YIGsUDgeqpmRWFTeQtbz+VEPmV5rzL
fuThJ183Cd1eHfGeneGZQqN2guZc0LIGzJ+vvuew7lDpJM+SELtlSfBx2zBORzOd
NCalH7IjVd9FDGYS6WP8wFtBBv9+P0lTKKpyxCzTp9jPcGOv0fZFBACz5mtbPR2x
VG/PxmQ14ZWQUu73UT0X2eze9pRJXFGhj+DT/X1i/ma+qTEQa8rWBeDLjzu53YTU
QsJFQEbHbuslvRcFb6FlHE9O3Tgnj77jmvuRx7Zzd0nZF/KQG6B2cM2WAooE2WcR
pXWqv6wKUaAUEH0yk9a626zm7PnaM54r8ezL3mh6io5XwEQMKjBukgf7P0dPeX4W
x/uXIGOymlc1u+iIjXWOgCEPw5ymMvCcQQDSwu7YcVMwRpN8ugQFLrlooGtdFrKs
Ip0Wy/x9tJsNtQl3HxIv4MuGwUekU34q9ds7HSZkcJ3VJVe8ZJy15SBtAmTwWnRp
mOKmklizncA+umI275CHW0alaJd6128IGBKWlj0/VAOJFe/KxZdqdIiZOkEwjSM/
Foq3n4pAsUmwBmTf9CdAMxG99NBh+BNPOfCQOpdjC6CjZ18tFTlnXg7T29WP1VoJ
G2CKji/WlvSh9Ak16pWCYxTH5ZLX1FSmxf1gEBzJv+lDoWMJCvfCaZ7dhGUbwSNU
mTANdtY1MCSNh7ZbsiZX5OYa9tElEYPJVSpHBHav8CdMFBa1QpNrE5DjGZqf7eJq
yuAiSI4flYCa9ehZ+R+31orSCMtg0TBE9aR2w3KdBn7RpvesA+ub0WpW8s8gbLb5
0wDFgbHB+LJw/6EhIYgb2HnJ6GXE/I8mKBSpiRY0Uk7h8f1HBNkKZQ28UyM0T/nh
k7abzfkTec6lZLC/5o2GPFYe63WcySIs5mFT8T+e3XDnhnkt0DtacPnTYNlA5vX7
x1tg9nlqCeoyqwVD6uUp/3H+5hcz8iB6+TJFH6HX/7aXdju2l7WguhnMTHFxNPwI
GWIhCUYigLMBeL8kntI2puq3ExfmhbQ9YWS6+rCzOi7OKLuANCzfx8eYrJd9u5Cp
Z0QT5ngG5pLqZkQqlOP7Y/z7kMZz4IR0bdU8iHwOuQMq3uql7UH78WmXubWCjVC5
vBiyurCpF0Mm7VGU8RCjPYumEsf5Cab3AeuLMw6rgqV/XTd5pqGK/iFquSkEd2sK
JZPnbU4ECrsmu1NpdCxL1m0scyWEti606vrX80BWwGWV6ax4qvPyOR6zVN08Usbw
RR4MJWXmx/ceZoy69ilpjcjgkZa+vtAsaO2ClCpo4GVQKPkuEqo3wltfnljK66eW
OZ3nvgJqaypkBBXMPfr3kyiMFripcowbyL40S61Y+8e0h8aZwXzvZggdA42n1ToP
XSN5Qn/VgnAR+GC0nS3TNnVfXmIkc9IovpF2R83n28ItIR321/HhNLLsp4zR/vS7
LY5F0OpKQyUjskuidTyz08YJjg3TTQKhMQy3oMKl0sP+Yk5OyOERfT1yPQdOtcrR
Z7ef0XkN56ZS8JSUbj/FI+kgbcmuSEH6AcvKr6iBiP8QruOA8qEKaOfUL3LBUGX9
Nh6kLOz/b5y/OQw8fZRx2SUkFnnWvYKEv0T2hs4+9EzgUIooXq3HmrkIbyrI8lNi
380akZY9LB1eR/lnGSaK4r8h8MK3zo+lGuQLSjf1NW16QAUH6OqGgTO80x9NhA/X
pP6B8qGkAUhOGeMTh1G5HPPDG5jV2XRoCAIdVvkcB1/zeJYRHYmbx0aCWF2glL0S
VjZRmEOkk9WG9NWcH64UgZevr8izuolDjT3Rvwz2/eAxCYQzt1jkRW0zXGxhM/YN
m3lrLkeC3/aoHyzGvalhXxbkfHlVAZGJ3yBhLfvWCSpYLH6nSUUbONYM9ArXaTZX
419cUh0v+j3w4jABjQwaejoTBwY9gC76NbhVLsppu2D74BKd5OORWEuW+HyB38sr
fRmgTJPoXtrHfBLPQfyte+tHALqBK+i1SUowyfK5pgh0xUd9KghbbiBNUWeI542h
I01uBprBfzX1tM8qP6HijNsy1hlnUCZplDVN4tt00k8G591Gw2H/ywsvu0ueA36m
zzVL6oupA3Q7ixlAfgYDRmvMG2Y9zp/JK1kc7U/vODWQw9+8nUw40N9cI5A7lq2l
KeU9zBO5RxdY6l0fp1c/bRRr19ls4iOINIvKFCn/apBZ2aDQgGY3uyTZQyXY/hNW
ByhT1lqHgYd1Ntois+Fdn6BDGoaTrTWIzR6MhK0WGCRSVS01uPV1q5uFC2GPvan3
SOuW6aTpsWPoLxgOU48ZemxLncXrl3zqT/1/1kD9pDuXHkwOrKTVu5pOF4DTm2/l
boe1Uk/nUZBzh/VNESu9V+GBYpgmdFarLbOzrRi9ibs8cDfm/sNYXy4zE2ow9mO2
iKFNd9rtwXvkUq0ardNsXixuJ1Pmo+EYmFmq1vqdbeIRW3V/roLIqyOWZZCu/E73
JBx+7+C7kPH+8tWq5dAiqR/oQPQo7lBlC3oPNvmPzQOahgsy0x80X5fQrV6f5ZsJ
IAjxyR7OJVimxUmiZrQA2P2s+dyizVcR/2ndSFzAsGo0xE9QpfWrR5pAs1LRKjR8
eQdS0wBBCJL1WxK/VqUxGHPw0LbWNz4ktQH1TPAYOUhmXMKaKfqYYf2REh2UGUUR
YkfcFpkOvzJxLRJgY2sEPk47fs8joi2OSEDqWHc/B2DpEXiieCBaWGvaSCGEI0IU
L6qobUmIFqCimR1F0Bxxv1Gq1GTY+QXCKI0cGuSXpt+/MbFVR0D432AAHMeEUUo1
b0hjdT7zgLXP96VOKjkhzkHBa9jwRxTB7y9KPhWCPi1k2A1J8EdPJp02E0VoqxKB
USp2TuWAs7jNZ08pQcU7H1dYU4WBZ/XFKfYF0JA6XRYqpCgkE9H78InclSeDGJxq
0Bu16ZfkKndZVASbSK2QfP4ibaky1fEbjBxMdyMhUwPswiKRBzlc58OPlsq9boOq
r7TDcYSTeU7DGdd0Wkh+YByH5JnL6T3I+8MWM0fuTT/sFu3wfeXjP/NpBzmewzUj
4nPeP5h+NlAR+mK05zsmcl9orbSfb08tg8y8JIc2Ketd1bKUJEkGORzGKirbg3Du
CZ9jT+R7xeIq34n4bBK+Gt7hPMmo5znIzsp96dyzAxHJ0jx56v9AezxwAA9KZTou
pm112wbjnBi9hDz6HrcT3AZdX8aXmW7UqJ1n9lC9vj8a7bcgOJgDpXf8TqsnlaX7
dT/zytov6X9DSsUaepifW5cMDAewXjXl04DjzUGhR+1Ql5OqK30ydCfucqoInma9
Rzs4MehrZKyX1358XLLS2j45OfBKDFWBb0abzPUf8LV9KVwbaM7Zj/ZBLGSNss0M
Mco07CXwMDXUE19IIAOLDYyBFzXaGaTK4BbjLk0hCYVZWNQa1+W2ZHD8UQOVbWhc
uRRtBalcaI/Z3+Csq79Z72KrOo/doTtd9nkarCqN5djcDF9P7JQ/Tpw7LWtdfE1Q
Z03JJoGv7hEKG0c26D+LXAgZ+UQYLrlIiAsun8OkEo133Wp0a7khIx6dYARN9oOM
3vSOt8mZ+lajM3l53ygLUIKfNkmkkKRBXEVycOZQuNYgOHYVUORzfvzPn2SNxY3b
Tg5GnEsT1gwGentkSn2QtLq2OkOh5e0STL6btvseUR9sy/5f1Zy1kuM104Cllnrg
PHltWyEWD8lyLYdNP1SaziIghvkFDZf4lJwR6zL8kEaI5SQ9NlWDfpC4ttfMwbhw
9hKHGnU+S+3uUjvj3fhweJaorkh/v3i6bboaZxLbR1/1nOc/lcUXXamB9nlMHQB0
WghViYgb98YyziItytI1JU7FOYOXnbGvC4tfHTMt3L0qITj9o2FetzsM5kVKWadS
TboSt8P+PRgEsh/GmOx2woaHYOV5f9QrySnqdtQYHx+ZtXYUi9Jb1aAclSv6rub7
TIZMNl0ccVXvKSnhF/eMu82lA6DeLLubk2qnRiiqsbnwe/lmGqr5uhayiGP3Q8et
nM6YIB2V5+gq4VCfA7f+Ps0PoPt8yy6wN0H3tqnVVVJ2Q8IKLSzYZN7BYxen0Sry
lVpeqtLkCd8v0sX5g0a1kGVms2CnGqOt6Yi7aNRauD+ZNwP3q2emthnoxn5iOkmy
qJTPzIMjU5HHUGYxDe9/8vLJFNQQRUOKuh5w8tBZV8sW8M/EnV7mtPxmQGlj2dNx
v/UpMXtDq2w9JsvUFWDUY3VY8QNQhwFtUh8/k60l6FkN2PGLokTc5PguuvKLRhEX
HZSWi5of+nMgezSqH7HW6uRoXUWBp5m4akd6Dwj4Hsvx46KttRvpnF87ig56GL5c
7WzkIBM/I3ocjan1nfv+tR1adDIrdhjPd30v413zZqK5MpT6AEyWNWMU7g0zZljY
MJwQBifUCKEkqGAs6hbcYfN/kterna3I8snDiAaXVAAw/1XeqGd/t3c8xteD4ETF
HPDSz4mmxdxcOy4lopA79Nd2DEDNqnXCOHg3dIaqOD/UaSGr4RKzly0u4zataDBH
v6h29GXFJsz4RaLr8MePsDZdmz4Azl7KA0BTnM/7/EWH/7UrAL3YGzbEzY+QGsyV
U9/V4jsFovQLELg4y03Q5KlbyFQ4L2xDhr2gIHwG1HfBvr51QyKM8kB1jG7wSzL+
jKHVyj9VlDQImxVTqsxmoe2pFDi/g4ZXdOvhV/bHxYP8Q9oAHTyBPYEMaLHsOQjN
odOKHUk0lN7fhhYSK0cMUlHrnSBKdAMGVf2U90IX+QMZWxqGEF/iE9bPmwUkV72X
ucNL5bbIJstBluj3t3y4ddfXDcoNpdQikX+p06y+pEyNiGPMDMVxXn25Ji0B7ahI
WNwEeAd6X2HEQmLjVd6Acyr+EWmR+xjYPW5qwOTqqatWep4C5MbnOIt4U5/1WN0A
+3SYM8q9ULBcX+i3voVqqhCj9P/oMz+BrYi4s1nj7zp7Spxjx/oX0QJR72NEFwRc
eNWWjcAfAOpvdgb1wx9n64r/hMV+rkOAUGXCg8dOOLBbRcf5CgtgKsW+kZOiaLxB
LlFz1ywcL/+iJ8iogRV5RUEvmBElfL7oS18SDzNDugqE4FLVbAhYoC1FeKsQCJEU
4wD97MaDpIjuhDBEi76bTs+MjeH81U9PxTLiHC5FRzjGw2sNUmL4dvI2Jlaede+i
ioGKGjNdaq7zZ/RHhF3QtehNvWDTHQ3WGK8LHm0p1UxZFZZXN/awU2638fJ3gbBh
pw3Whdrj2OBdndOHxnpS8Zl7utLAk5OERrwFbCEsN3kFnoMOCSE4ldHU2PpbdqKS
Gz7uGEr04cGlzS1x11fT/Fs01Abr8L80xT7EDaVJmxuN+e+8NMfTZfbqs10poaYV
7iv0L+CMSpHZMmagAYfRzuFA1jmW6iG3E3G/JNpcYvPB3r+JwXD1nEmQHQ2hMRLL
T4T+eJNUQs3g+ORsBJyjYidlRufffZQ7yH5+QaFXMKADJrjPtipar/5lWibbqkfK
o01/9zApicpYvMOEbL1whufeTwx5B5pUgm74tfXOMVBnztw4hsFbQ1Vf6euYh1Jt
bgkNKPDnxthJKBdk9xO9i9iT1BvbMzDF0J1T3FxJQS8loE2eLZGXcMDEsfgX479E
meuF533PiRVzWq3B3NGNl970rE29xsZjH/lJU8iEaysPRAHfGMyKvUJDrpVDkU/1
U8mTtrosnLhgweZbvHYMXri8AWE48FyzLPoLnLzv1Flm2UPqyMpdfXZlrfxV17Fd
njj/WLt58KKlhTRYad6iuw0rxHUBqohhVaeEz0PMC1NhIU82GUH5/Wi8ylEkva2n
L7bWZqTqjmmdZNCIqq+hux8pSlg/n4NWe9lPvnnbkh6mBKERI8xyrHTeTBN8OQmD
OZq7l5znD6eEs0qGyNu8R0NitQhntxhC+aOvgMVZXgEXKUS5XY9gR7uNQFShndCr
uN8NNJkp0hEfzUlXA3BxC1ZICo3Ote/7k9nbzmFIZbBp1OzEIHiDwTH4ZWk/KyU9
e6v8Q73F4GdYRvKziDa2VZY6TFGDdsGfLMYGoJv2zY2IewbJ8Pce8JeoPrkKS9hM
4I2Xah2J5MW0fTJ0Ww9+/qZ8LLN528VtUZtm8TDUPdT2FZRX1HPHlsAlJqdNu/c3
Vdu/QJWJtcbUISdiWu0Op9/hDJbZV0GHm9AxJRZFNc2z0W5UGRGNC1iprZ2d1JIg
LeM0NPSGLCtN2VisqkJktNtx7UHGcdqkCEn4r1zql7AGqmjsRFr0jE5FWdP8WMD5
Xy+LPM/M0M17nR/H9RwT18ipiOKbmxhtmwmJpqy0i+mdJnLJk7y78QoU1ByQzyvp
3P0lCEjrPcaSVgAb0udxCv4HUECQSkyvHSwrzguv1CEW2wHg9m0XkqqOpZgsblyx
mFZJsGUv29YfN9X5VVt6is5pt7kuQLHj+61sVdQG5P6Smk3wugai+Lpo5pQrk+cq
tYVJTA1h9I5Rx1WeteAO+Vn/wjNIbtgGWZI2qDeRv3201eZ9tfG9MJWe1rY3S5Ji
UgQlDz19f5v4+bw+GVms3vDfGL10HYyNhaaTM2dBWSMmCyNIsXxRSu7g4QZsLYET
3nKWwA3YYHrD3O9XeM4VGv8LPj/7xBMwK/Gd0Fc8NKrgIlJq6iyBAPe9QH79XdXh
CLS0OGrMezeCAVx4k5Jn+e7EYoYHILZqQDvmBsBbQctA0kvRsdpKU/xOHuWquZ1u
XSudl1TFd3EEwXWT9K3cPwHJHzSJ5zlwHqH9Y2IwmjdhUBFBEpMPOafjZBAM8QgD
+QFpx+0lGotgS0mTDt7LymPPvUA4GWqkET+mR/LZPOJFQ+QbaxBUWPLGLNf/cjct
vTzFIaUMt38eLEAnxFDyOKLqm1u1r7xbdiXuhUHmLn/zjrModFYxhaA6fZjwGP81
/Yf9JwENMyKwpx7AfYTd6ct8mcM/VB0juNdqJaww3AvjEHc0TW9QK4WCPsTj5qwo
KIHTCwrkL1S/KyuCByMuqt6S13x74UtRdqmScq9DWfC33PE1X2mwZhy73+SsCuOO
BIQdvT+89piIbDTbJdceImyp/zDiibq79NWhTuZNS841AK5qRKopCBTq61Eano7i
eO441lzEuG5Y/7K19ZhSo13/YIouUCRTQuQzLYZPQf9ZnDd7/faY99Xf6NBrdBkp
vXsCU4Pk/6il2lXhUHptqdQKapWBzJxS2/Szuabfad4nLYkSmgY/88athzlJIaWr
pqZ6eOcPVzlce5tCtWXriu1gY3xM53ApPQqblPxtdVs0lWrzRQxC9IlXcToxw1XZ
7m96sx4rUpNCUTuU6uFIuc1n6XF13vSq1a/66HGA1nkj7q41FzFaq9MZY2tMc+iQ
uqCtuPsL+p2SjyEQjiIBDsQVHzpxuc5jYH29hFMvD5PZuENM52Luuw047zf/igaf
oI4/wH6pWJ9Ltjp1o8+6WE9FqkJYYD7cEDatPSfME6fDrv2LDGCTZEhjEEtxSIQk
9WiX2aO/hVel2X58FFdRwBmGasLMMESPvd2TgWJSCBTG0XyYRIhmx5FyOHDRiUpT
/O/XQm32+7RTbW/t/q4IgpO4JWs1+hRuNerooCqYJuHU1XevE8nf5t+EbrzNwxS0
nQAXIUTSALzllHHJxlOoCnvD7ZxNTv5NaO/b9k3YX9+UlbLOyzizxlZ1SKyaOB6q
wZoEeERjSHMlRwk5k1DX26xwbGjynmlsGAipy45JqYBjaf/v8Qr3Fa46ba5b8QXB
T6HESbP1MHwMygyCYHsKntWKEOfRaF8VFU/NZgtSVmq9IzdpCY2b1cJP5/p+nXs8
vJ3se4JsT1642w5hD1h/zS9qyl8pKDunmEfX1VdCCeneGtvvi29Z9Wf44IwCoZRY
7kkgknDXC9QM0pRWgkMpo4Gm2Hymq2QgzLSypVPJerGhmrMECvRPSfYViV7a+jcM
4uMj8qsdiVdBE+4ibShH79jAB2RNrAGsYNf0UkkgWiJ0c4dDqhAIuTVDytOyPIal
qJ4txFx/BqkIDqS/X+5IH2i8vUufoicQGnu8ZYiZfXWB4reJHD9p6j3pp4RwE4vA
ql70zlOGgYHglsuYlvYqIeVnKbFxyi1k2tKSblyBQhxPkU8q5z3uzkUzOvh4kEmM
6adrH1N1+/u8UV6LcM0lIoI42Zjb2NO7v/ykgeGMgfngjYNz9BzErqziCnn5Tbbj
CL8AsrYXahw6tlZOIZ8rlnG8xCDOUFgnFTEg6njI/rsH/+6vq9073I9VfAT4iZcw
enHQIfR2kD768o/xtDTuBIYDluRDVTKCFVm1EAK07A9q9iPkyssn2ZVGzH3vw99o
i6HWPtCBsCf+SdAwyW0j1eu8ronX/7evKqiaQI+ksD3cXhXjzH6pHgqys7NM95xa
RiiSSWLwxN0SjziStwCaV4TZISCIq2GYGT+qQ+C85U5snIhcLnrytWg2I5Yu9Yxw
gPoAJxbTMGrtfWAygpHpiuXgHhAdju3RFNcu4cHvY9OukPeFdtRWLLCnvQ042rnw
mw1IgulGNe6CJUCIH/J8ELtZgftqHk/MiDNEyS/SnNVUrSjb82ubvUxPx9NIOBRi
F+N68On15r0lt1i9uaDxVuOiQSPPV/i6XfDiV+/o4kMOGM0Yk9zzGCGTpX8ROs39
iAjhQY0T0M0K9IM+6P/FhDOH13qMNaQB6RsvovjOEFZCIYxTqrrebvJ35mHHLzwI
KfFBb7efTPRouRuem9i4uYsrkzRnofrN9p0WFYxEoYieT+kRPNagDnSjTxfQsFsd
H1rsjftqJboveqAQ2F87yf7nINmb5OKS3Qtyhe1phkklYu55K2Ymiq4DAJd6x5zj
wP+3DQdQwO/BNyUsDfg34P7yPPNaA3pTYwMDiCzytc6uyEiqV1TJE1wHoi8x6vkE
ExeMQk3iNVa4hj/bPhJV35/+m46RZ5ZHoLaB2BtHF/Iqx+anr3wlHmEmTxItd/IC
U8oRaqg7EJSsLf/NKYbWo9pMkjgoWzJrfOSpq7dAZuoMpm+rMhs9AuXtJAh1C53+
TfG0RYbla9zuK5Au+QzpwRogZTpdClYYFOcBYqkk540cyziqMYgWukWCjb4ZjiQi
Z5bH7xnYscEqEf1W6n3tIm/stPLA6P57CCXvoRREw94BQpM2+dS6gv+5WrD2Sv/f
6KDhkMrgsRiQFGQW9yhulLP4BPyp6QXKx2+J9j2LfqSvtZjMJluq1OVoNam48VGF
kMukGJcO+PlzLhx1JAXzCJmLolszAVp3/yEW4lSNJwNmxhri2qqfwNpINJJRQnlp
bA0U50u7hYmpz1JdbtLZAm1dw7fJPAFNRzR2TXGALizSvZdXOsEVJs0pYvjLkyq4
hHtxtt25P42nxZ7armjN8jHTdrScVs/H+JruK/iMDQcMQMb/4BCNOwteuLC2yqIN
YSqiOTiTnp7e4qaPqmLEt8gCsFbV882lqaDbWoOUWyDI3MC9wgCnRv1yTaZb8WS+
wx99tMzrYT4PXCec4fu9q9DCyCrh+owGPJZ4FAWIYkRy2+Q/zRsDo7i9zKToExSQ
dj/iSJeAt/Ecc0VHSxbQRnTtJBhU+4umJ4gyZIe3q1KUq0i5XT4smmohszv9aeKs
9XVNlYQ7ScWRvDkj29DDYvtqoKkOpluh5xtkErhXvKh755tM4DL/o05cp4a/+Jlz
WKc95Vn52PCwqA+Dmk+9KQQqDvPN/IVS/w7mytayf797cPAyrI085+tnHe6xkqlc
ofAgs4KieM0A0WBeetIQnOaFh7HMdVKkuLAsx8+w3gUX273ZYLdcJxNpeNku8Mc+
TFNEbssCfM08ca+74dOMlkMwVBzGkR9QJi4xD5jMDWHUVjpa8YeqgXFoJIDZMmK1
2uGWQC2kHAarMOW9PtPfnvbPI1t9uw0+ztKkndiLt7CsFNEkrMcYQddVZYN5Y8uY
oEOa+bogInI2LAdiJ2/W5VSt/Ci6Bij5yi5y0+D7Jle8q6S8asGOYjyvRXXKGNbW
ksD6eAMShubyBwy4LVK1d9Gz9D3yX/Z/IBsie9O/yQ9KmJRyzkJEgY6KyuQ0AoLw
BQ0TsUNDwq0lAtFrsIuj1TazAiaXtxToMrm5920BK8MmgREwr24xcZg8i2x4qRIA
dwbsazNL7UXGptfBzTk71I5XBBv4E1ozdu0HvqqAoXsjfYNI2eKmaby2t4ICvpRp
FU+HZvzVoLT0jQewutNe9hGUFrNnrKc7gJCEBEaMsh385Z4k/vzY1vtV7SL1WLai
PHHoRcw7GD7BHxMCjplctritZ5Tk5My+D7dZZZDfqGAUEeNP33pK13PbKJbBlGmL
ybnidV4e0zu5FwP8iwWBjff7SJR3Ree+4B82gc8s7OnPSIJE2rdDZh0CFfqUItrv
5NYRLWh3NhBZ/BxZ0og2zpGYKDlucvjryo7LsGIKoFDXPfX4tBL0DvvfIyopQ7Wi
wavlulIsAkEtC17s786ntm3lY0UFZxJR+8TpvEIbqOE3GUkz/lcNVwWZw4xGs0fh
fBhVIM4BqH38WlQwtWaNQbe5gJddoLlkbD1NtsOrNRWOJ5NtVGLNG8SPRBHtSw7a
hbOSEdrmKWyZpCu2VttpChs0UoeYkGHg8HJB8Ww1XX4dNDmfFGNzqxdCDTc/MCBR
B0NQIXMXWeF1inKm1xUjtJlIS/r2blYlH3oRBfokaLkjsqwUgcXTuaEieN09YFFr
AJgf+N10FoYJJzg2ri0+50HUA4CSSCIqZbEnSvmp3e56F5swJk4rlK1Wr8KAQwv8
8wNhrzA1T3hYIVwUgWWlMZfEpquCeS/apO9yiwwFJuTYZsdzmZWAFaEC9vx8KHsm
DW0vhHrz6XDRD90sQTBwPSpn29a1ZPmN9GyqLK7u20M/0ieABURLTMOfrZ9ADJyB
tHsYnBwHhBP0exLvWSSZoGKBLJH1eytgHRh49Jbc1sPxCFa91Ub4rT6+MPP9eu1K
883X1HHr67f4R0VXnbXrkyzzmpWDy32mac4YkzHvUOs844lxDipLOqnefemZ2/yw
01uIxAeJfdzHYAtQ5mE3bXAx3pp3+0oJtiSX/ZXUag87Y50UNaRoEhhdhBLAdNWT
MK7eKhDnzXDEW52nCvo8iBAOPPNZlsi/zLjWV6Oe5OUVkyk25FhqQtnbG0kew5Tm
t5b9FX5o5C9pDTDPK9d5F2uYnCWGIor4/1ekMg+4mSwWEnzSC9F0wVBUDSAtVJOF
SJD7vOlomTBBcrOuKsVHP1GwIIGs1uE7EL0jVnNuEXgKfkbBalebTHYTzfD+MRdc
CsXshvMHypt9l6t2Y42toH+SvhprxbplKVjAk3tp3k1XBMuG4rngloBlnJHSTnkB
cIgYIosb/6JPLW8JnwnP7bPrypkPrFMfYtRU3OFgZpwzj+r/j6ZbH7/yVvZJ1UNA
ZUv8mOZcOWGe1Rt7LlkPvS4X6cy8eiKP/3FtOoR9gOw0cxz6lhpouu+2FEIuDub9
4Ks9dy67UIj0FwPx4dJT31fWGZFBt9duHDJO85RGUoOAmNid3jJj5FfAJWlKCC7m
3I+sKA8xhNfYOPLzxD/HiDWKWDO2b3VRz4uOzGh1vDJmMxNdA7efAJDjEXLxjk22
0YuVV1a/H9dfTmFk/JY4sBWQzG8wcEDmM5yoMqzllr16YVXgZkl0UwZpqxjIqLFZ
eiB0sH7qujaeURcB2BurTbkszpzf4nl4w31QPrl8ztGl6zuRqeEjbWsv+9qU8s6s
OGrgUi+Oc3eZ5BsWJ+wFAlZ5uLmlJxO59h7floAKTDHEQTsP/KgmkUuXftni8Hx9
FlpE7BgVOcu1Berdnj33loWfKyKEmeawt2C80shZnvOvrs4H4Bz9VpgF9eloL7yb
PoaxgG6QLQZajbd1mTDGdtvXeLkgA+tCZZt1+TgRYd2gSLP+wfAa0XKko56hpVwc
lL4nfTw/L4GOG3fDAuQQp4I9kopCcZS37Y1Atdkn0W75zCJaZqOfGnVy9a+KmVH4
QaP2pzivI4MAUEcqEgQySs8ABNfy19QhlH7CaoKIJtVbNvJ0/r40wc0I4yf5/d+D
a2QwcpwQTyPz2RWwidop0hxDao/XTwgCfHW4p8CuSLjxJPJNyDUwdAEntcCIEaRs
G3mWMmrCzO5YnJUvuU8IrdijzhBYLsuInBwc9d6xNMPuKjeoDFGLEeBZnF+TmboS
Nsek/74cN19GbRaKqpkF6xYkc8O1d9rW5mmqQyLbA0iAakiElMa5MGxdmJwilWoy
bZfUGt4oTapxOq+YrxriSqRRZRfW2TrvmQw6wkr5P7K4f7w1H954+9hplgwtkNyX
c79xAdQt9uUwrn6dg82DUk09N+qbEsB9tqcrrAkA4zSAxTV6vta1CqSORPQAQRve
O2oamAgXnjJ5yAX4LYKzBjcjB62mx7j92mMhicytUS8AhtVfoXGV5M1Xt1vpKhHl
XD1w96F6wTpwzCLPFtmfHp+krmFKoZUwKwe41YBtI8ERxZZApu4FY3GZ3ihCr6VR
OwjF7YgN7yVCgDf2//z+2Q5DC63lrswO9nA9rej5ejxcNn2WrnEWq0beHAuPL64G
KjGBDQtLpEOfulyLtZBJWCn1wxciUhMFEuySNOQKbWm63XjUDtHLUFjzJhOzaVuR
7ePmdpCyqqqq+/y6Ilrr3KI/9/6eIfnm6X1UnRdYPmiQzbS6dAbR4H0vIjqbRRK6
H7acXMyUSa/HSwgWrpqGhFPbiN1uKYVGRkoTkmra1nBaBGM9nTRsWCxkNw5edi7g
rlCfDLot2FC+5CF3652fJ/TSyfZxp/PyUpNE6S3dWDmyYnYr/oKMre4AsYTxI42f
2d2zGzytc/Rsx+x5+FUBAQuFKC8Um2L14YlYl7YyblWOfMDEDGmroJ+d/b8mPz11
oYqhvQVDMdI56SHj+kDGkB4IZBUNaf981BmEqGEgjL9cfBcvBzFmZcGF1fB2q10u
UE2pFp6wbr110gmVMtdFO4+JmCXMycQDvF8LEBQLVIFZtAQtgKv+GDe234IwFgpg
JP3gISK287UCBQCtxhAz7eFb44HbkFhbpSq5xgureNgnceolpUyyRnXrIHADdLY0
mf0XvB25yP0NJmh/eUCfdmZ1dO+I0v7Gfv5l16450vZ36O6QHDm7WILTSF7Up67I
lcQPNBz9qvYj79SU7JRJv+FzSABquML/z6vvRhWkjBUqmY6wrIDMzevxaHvtrfAv
B/CBofdegqVR71xxO1cl3hmi+NUNBmJ5xtNSQU18uCDLw98dccSACz2Iy4q4Zf0h
fBcgGHtMpiN8Egn8zycCUqvUHihVESnHHA9bNJXIrlqWYgWipEgeWjAzpO1ILRbG
GCGGgNnkXo/8DM+074IY2NCNlHs4lAOCqdpGEQyDJruCZW6edJCbqu0pfELk2STS
8cdA2o/ltBNsHZwVcA8OWfszzGRBY2um+DF183/rXadmJXIe2GxnueWtRZImiWWC
sb7pzHq2b7jfHp5XWbpfa1E/h+i8AAL21S/vxJCcvHR3zAGSxG96Jgo6hWO6fQmS
ns8c393jAGwmLZed75XkMhpIK+5tVIt43jqsHJfdBSsXTM4bEXeSKgopBfdwY0N9
u0KS5PNcyrevcNv+Lm1pAlTotTIviunVdBmX6WPqT+Y6JNGexmeF3JqupG3konb2
Q4irpTBIfN4JKNGwh8V9H4hCSThmPdKoJT1A6OIhxzGXwKFnQlCxXqkO1yQckL5r
vvWu57g3NulkpcFyUtOSaYQD66CUjrYudKZ1Q98MHvAg7TPDO4/mWZ31LFHvUSTR
S/oO3Iv4kuxJ4ITTMffubClugfLMhm35VTAelqSANpdDAnbZJBZev2IAJP3ezr1u
Us30I4WZFiaN2QexVgyoV5dS+QW5Uz0Pyk1D7VAzrbBiFElw5oSNC5y+B7U3+laB
ZwTnot1eSq1ECZPBG7GRRnKiLEKORGP2m4pBLS7ri+sLT51fSse8J8PpzJEgHfGO
2H+5iy3A4RrJtW44Edl/6pSAY1D1Ua9akmh3+wK7iFW76zQFsFYQNO6tiv9DlASR
WtLhMTIcwmz8vU5togU6VA1ohvIxGwBOpmBE6Id2J4cDff7MJrcbTZ2PM897y6lT
kDMqR9JdgX+AzjDCpzai5jgNS2XnpMqaj2TeQVXHvgizBfe3ZhUZhatjNRvcrtBX
T/16jVlunm6xOPvEuKfkKXwTnU+I9kdZT4PueMM81Bz4GNgZ+HJvvg+aBUhMd6yW
rLe4ofjrGJm80DThNdMzFrYNb/J18srYFUX2sN3Ppz4sBpovCaxSWErhqjgQbyzi
glf+3zSdE8O0eRbFWD8EZomOjKT//jRQ+fI7iabcrM531YuB6PZHo7rj2i3lsvsg
LptY3THRIlB9bJqKkbG3ZwIvZN72AgiXfqvvNeDDE/A9R/1MX/DuAUt14+MyVRt5
f6ZH+q/SP7JNBf0Sdjn2UoCAElPC7+2UFS6DoKEwNazOizsd/HA+vTk8bJKoef9F
d3Sh2Adve3GINsIIPp9kfMfm2vrOWfzpeiUwY/39fozgFg9QuYwKRjBlKM6Zfm2L
GND8Np9WMr04u+7BlndNu3oLb6ktAmSjEw5Y3PIIZLKT8kiOB0MgNIhPp/hh4yhY
MLAx/wrvuWDa9ZH0Q/FLX3uJhZjffSGMTtFfDKrZu0ooopkFzQPMhpQsZ9co+DHF
PwHQ3q5X8aaTHtWlwyY07VLrk9mtazjmooqILXS3hUanviuk0vl5I/2TyF37M+mr
UfoNStrsL0O0wgpYkR4tZl6QF3L9fOFpmK4WNxmuNrbRB2wUh7DMNdmvGiQYPO7s
yV7N4077Bm6i8qOSEWrMDcIlLFX7GjffGdFyJLB71R40ZsfPh5YTMyLuDo6MTlX2
ioNOZiyKpQQ41/Bx7LPo8whje5FHdFg7W+2PYf5+ZxMir/7jIV92ICoNTjN/hNSp
2Nw3rv58N1xVGQu3RXw6pNqYGIHfhJ/jgVDcXFrOnz7jWbb5cpZ1WG1YaxD8OndS
c7TaXl6ccAqUmPXdl6r1t57+HqaMUab0ZR71BHrdfgTEjq3weKgc8y1mHcQV43N3
XpkujFX0NZVTfYwx+D7k5NxCfOcx+ctmjETMfNaJGwFf2ztGZswQIHPL0/ZWlIVS
Q0x1USz9blMGX0xqzv/cMyCMb9fwpMQyPqyhoexn0VGalt1FzTdX9xSJXfBWVZjn
HZreHIihBiTpobDyVrMDn697ljTt0OoHOBw0RpkgL0jR2vkl4s9hVhsy+QKlpaDf
1cqATecZOZR0hRiLwgBBKHWe3zymnrUOWOp3iUwtP9NoYGbtpkd//CEcwQ+s9svl
l1RI8q+vpNNz9NP7eCZftFzgUXIUlMohUfD9vPVcAiubg1Gd+GMwEi0nQcIZYBXT
IX/glgewiNMU+MeKvbSfPH8Dl4BnCFZpGszPJRXR7EXPdekr0AjUihg6RRARc3Z8
m5fYt9GwKpkeIUGXh/msk2Qr5qobU+R9bYJHHoBcnh3mezuP6dt1nj8zQkPG7qpu
zSWDR1AbL3HVOYkeCv70RtKdSdAOLrfuxxdp8eqPsfABvEPFON+AbxSfwdoq5xvN
xGVV+ZB02BEPZhiQPGTH1VCe8H5sxF5YhBLvuKYM9uS49MIVnfg91Ki/RxwO5YPt
sfGGt0ZSiDjY/msvunb6N5tAjOxtQEckpmVbsng58NCqpaXj6zT4eVJrBp1YLJBq
WDog89MmXjkkql/814w9EUC/1cjcXWFu7DFWm2/1yHTwSx0s7sKiR5tDz75OJhYX
M2yY0NSIY80jj83shm6lY7W/LJ4FTx1MQdJC0/xRUFw6y/ZvrOaKb3n/uxP6FmEo
5pO5ZbxHkNpBMyVz1yCpwk8PcBWRYpvKpmdq20EXF/SNhaDn8qto7mW0ZkZktX8O
LnMnDy6vtncES8y7BYPC4fk8hi31O40bf2jY+NN6+toEHSL7U+/JQ/LkJ4e1dIpp
TnhMJwZwHBpEp5sCPZ7Lx30KP4j5Z08Q3z+vXGDsixJkevVEUbWC/vfbnncLz/fv
X3z27A6z6dQ8w5wTgoIyK7kdlz7dB59z5knJVguuTJiKtqnjb618zsphES9mb4UT
J4LJ5y9eW6FwySrElLyYNI/1NtNy9Qevzq6/mBDWXSY/camscmZEbVPog+qeo61f
MX8/Dgzcr6ZFR95byUOnY581576RY554VOvN0qz5izqBnygkQgHKW2vXWCwTPhTz
ZmFy5BNZraHHiRcZ71DR3Zpd9641X74UT8TAqCkOxGkvs/SkyCGBqBnIcPrShKx+
pmOa1OlSj7ba8/zFV/wCtBVhDx2gIPKr6+texo42F6Yo7WZYIIDu2Hu8U3Nw67bK
psIvRUJevVJ88wf7Luh8hW3qdP4ISFkQDzECxj1xZ8Ll/If8cKPs327UMAjYBnPE
NN0fCj/RieUiC5Udwcad1Gb1JJsL6dkv0cptazATefw9VRP68k1iYEYp7QMtIP7z
eQi2qyWCUoS79mb2A81u84kBwwQqmqSQJWjpVxfFEOCmefZO3Q4mzYR5KlIg6DQz
ejpuJKVikslAg2+gp9tSrPptGaHpTti5Ij12Qsbw69nDsBdbpsCNrRoa0k0YHHDk
7SCpQEpxDIiPQGH14TlHqZJIoBnuOIG8/A/wRMROGD/azQYH8cdVChD+molcf4eV
WWVJsoHCcbj1q4RI/DcuP+6fnBgOFBAnOIHM3GIMZ7s5hPjtFkrVI2TksFnsS1jg
UJAAzTihxHYVRoZqWmCVKUXAYJd9477/JXnuJuRv1b0K/VS4ajFRyS/zfJ1hCWe1
ufzXNXB5EZjeVqx+LqRIWX65L+CSMJQrixsulg/sP/YTx1tkDnR+gMYSldxJc0bM
VszCKjHSs3uE50n3bcAaIpTkf1wA6dM1JbveTu0CwpFHy1k4dOyhM52s1/Npkszi
qzlJdmwZnDlMM+A64HcFimMx5M+mPYvmIOJ5ywUmeke8gaG9InhJiKm+kZgqtwCK
N5wcCKb3y3xJuCs4Q/PnaAJIhuZlLfCa7XIkA0kkVUk7AvzLemZuGV6dxqpXLuW2
5/s01o8Imy4WTmZCFfm3qISC44bUOBrwVqyApaOR8AlLroAgEsNYnseU9X456eVo
fxxzVM09WhehELiCX2CpsmGrl1v1In/W9mdLU108pcunoQCu88TjIUw2Fo1jjvb9
X+Ot6NwwmNWs/lXoNZidkisOyplI+/hBEiaEmtEeO5CQQs4NVTDPpMhnRUqNSkbt
JAZYuoTXdfKudQTk8XnudddmQ50cbKgIDmqwmd7lBjHPHjjf+NvIelzyEcZMfkBF
lMOa4jEeFRLxnUa7Bgu+pDVP4LFUaK0gtxyhBQHXRhRVbJgy/6PZTZorWskJys+T
aogIB6LmlxwwqXbaUqJQQlQQi1pnAJTUFqvav2UP8pmDIYBd6Dvi7XQ+zqC/xCrJ
dCKWBCGJiCJEuztQZR1HDWFEyLGmXyUsyZZZJGXUCVPGvcykyiuDNsbkO5nM7PIY
XgG9BzF1+6vR8rWF8klnSxq8MvnmzGshS5FWipcfoIlLb41is72QUIqBlSGaoa+n
SKUryIGmLnpekgOejWJ6lrDkj8h+lPjtdeidk2um0N/YdxsxwDF2Ka5eMRQC/yyL
9JCbbhW42dSSRu/nvHyrelo5IXH2vKLszDKZGWjWbR1Yuios0BSaXNz38sJyOUAc
z0qXb1QW4qXK9RnJedEQMs6szcAp0Aj3SYPU7gvifx/SNQvuBsDdj5yHLVYs1E8R
9Xau5ohvQwPUnoeN7ePvOOQLpjPJrFiBXEMDHffrLglxH5n2qaHk96nYHmDVUYI4
p/3e7fbN81WEE0mYOKndj9nr4puVI0Yez17gfbqVr/nPFrPSeVxP0n3oszRiPGGl
s6LKBIvu/JYb8xTvfe9q5J99tei6zSeWOoGq+5fSSjAFvU90nSJMURPyW0IPRqW5
Ie5hmynYeDTEG3sZTfBvscUqn/C20KyVHFsvLP55YUWdeapGTS3Kx7HTh+RSEoDy
WEkCQJQ4MBg4o1jIUroq4uBlzpss5WQDnO4y085YqdAbM5OkWWyZXYEfWiVIFCgn
9xigYMaX4VlrodJkb14htm2CM2mWSO/jzxa6M46G2x3bLajsAwA1mnV0gX8Sy5EF
3X1tnxgFLXMYU2/h/aHggRUhU3wmQjMubihXai3KaseO9Zby/7U82yeJtMbQvq3v
hCJ9Ttx0WmXlqd77X/LLNljktQ00enw96tou4bsBYAVP5J0JW/FcKZTlMhaiDybQ
T6cUZc15lMGVyHKhNhCa6WlFwNMGu7iUFCDbRumJATnBnNZSJjIqhUwb4k55Wm1G
c3biC+1yhlppaGxqd67WwpabIdfMNhNPEfKTApmC5G4etuR/mOjc7fHblq0dXwFd
TNkt4HO9qZtXFfNrku7LsY40Sh1zLI2xlJ7miOd+apGJIVAvULtLCSHA+XxVxz/J
rzCLp/JEiDAS1AVKbSYAULlweHq/hNh54rgQaAXiynIi9BKG4glY640Pvwkl84HZ
CpFniVOSd8XXHDV97TD5KFshxGvOvB/yg2Toz4JdSP/kzoYwu/2CQLaddXOOfBw1
k3SauDBQyEzSUeEgvh/mK0ZgU8Zb6PkxVSen6qWoe9/eAt0zXxzCLHYJwzC/HopB
34FzrN4QQcmFm7yWwxrZXXr8tXBB2k/w82l3mgVemr6Dig1OzFbTVqnHK5WrJQri
9++xV+RBqPx1wvdCcn7xQc5gyYURRISYo5tTzkeq89vgllOUwJDh4Sk0MKXeddUo
Oe7+jE42lkRwwmsscIIhRIQQKKFfE8GwbcK8JyCKXtv/wJT/SK6Om/Ec3Swo/ZeU
NUmDYswxrg4hyLhTz0h+6ddXjN0GXsebhoBsVU15hOao8TsTzd6y5eborjzU5PHt
WBbY1/xnUSbSELwmHrmMN+SYJKn5jL/13m/yR3BvM55qUFb8CI09+b867CoVcYNv
TU4ODabVk4o9ED159+oh24D7xHEo7sD8nPGQw1S1P2qCPKr8B8aQ7dQ8taJvoK74
/c5S9mO3H5SPYGGJvLNJcEcuEJ58Hf9AstwqsH4mP1WM8pbhhQGvhikykPyNHj8k
3j8e0S0Uu+gE4hmDX7FEshk7FgUfMy81kLgzuXcfubWXkbMcYrvFgL++U212Sayj
jdiCtO/aDC3+LBUA7e9c4XQ5sSBLJej5cpKzyGEqhZ5eF8EDDGS5qBAGR9iLyzUO
B/sK0bGb6KMdG9vUDZsXaN3/BP730oE2lizRY3AI5O+3Wyl7kZ5Z7UtNv07tIgBv
td/7oPYo8/bjOJ5q43wCi34EC7vteZN9YQVNni6du5ytqrjVMtEsPr/xxOfwzGZk
4QdN+vv9zMhNpOYtbnhiSN51AFwbZPL8OsHSHma7x0K0Ok6WakJX/y/wnqse9JdE
L3+dBHQmmap84+DRtFqluoVqqIP8PQoqb56kRvnChd7VR4zhn0W+y9ug0U4cn4gf
HO/3VJs5AbKvVF9iVW/C+LZl0pcJnSmQEDoqswrmOkzxpZmQFVeXhT/SxCfn8jjU
14xJhpQH8PkJN19TMnWw3vrj/Zv3TBPxsiZKkHYryc6naS6ecM2patt90vVEAqpg
3BA3/6HoNG4j7bYcie9NubDQRXv1LAEVxmZwZnQ8C04E9EhqcZVf+Vg8TEcNxM21
gUFEtdZoAMinDbvjY5q9z2kOIuphwBdkwWW1sxGxQ3N6KReg8Gcqx389FqumNBlo
uwoxI7mDqHE/si8lykWGoGJtfnF2CB6eO8LqsZAONk6mXelcLqSOk1gAvJsm4Y0H
Q6zHRVuxTbspZx39fbLDasK+8Wc83e2OhdrUB/+u730kLyJXO/his8lBkcNg+j9z
XNJsDA4LUH5rjBTxtxH9Y/HyXAQ2H+poKU7GgC84+5o+IPpU4bGjGSZzmKyEkDTb
WTumAQ52voawWlQNJ7kfI+NLxxLG6d8oj9EbC/yJ6MM3NmBG+w3/R2NWHuezhYuc
Iz9C+rzItWbu2YmAfViQVoF4oizFoh/dYAwAf0RuhrEEEK7LzmaUPrV3kLL38QyI
tiUsZi1KqNqo1wUuQQ3be7UsQLMH7RTaNOYAEuIet+jABB6kcP14qnG0Oe2g6i1S
IICW3+/tZ5mbjqKKzfol4lxGhQ21J5BQwO8FC0LbE9m3JvH/HKUV7mdN4wbWrkRL
1EcerJXCckEpRDyYRluHIP0oTubL9pVYNWoTI+JaDXi97cHJ1n00jIHxesMK/TT6
tI0HsQAWGligl7+7Ui51LFE6082rsbVKXdUmvQTPjqAneFnsuIHUxcBGTOeWcFUU
BTtJz9M9iGCN/8n7JPg6pK5CC6YeoVPyNs2+nIegi8XgR2pSDWbZpPi1Vm2w3AC4
f6xxgfo1Q+AcyIgUrbBkpX1UMVledv327NLNhrnYIXpNxBOquf3uZVNV8n6Ttgeg
pOObuv/+pG6Kw/ZKmJ5Bb7srDxutl4FpD40GVCQRhzXJd7AeWur+sxJtjyG5FytH
ZTzbyfKMdUd9k+MZFnQ4IU2N0dBN4d3uDDnfmyxOAIiSrs9ZfhSow3G92E+ri5NX
zQU3qahrP8w86nTI21jffKE2YAq1IzNN/lyNpPwB51jsrBaFgjtuI08B2XGJCsb0
rxt90DhZPxfgf6Ch3OlRG8XguE7TztIW6cUzlsLyYmv46j5zH0gq14q+CafPPPpS
8YY0hrygSksLAdp9BX5W/sy8CktK85gUEnTwxg7U8V1lREKWE2NcR7dfpVYvfiqO
wm+ayBFPmaXKmNNh7s+HPcKkcbU53/Z7zFuclJbkMPXUE1vp2huDVgnwC9NBuxSw
sPoSGxJv4qPgWOAW4qeeBEwFbnXVxn/KgsvpbgtmLWbNLrxApMrSFfPIEgkIZEKy
fsDqehIk5FvddCTV3t7qU1lN2Deuu+X6vQCdkmFL74jXM+DcpS92BlC42V6yu68y
2kUUP0y1ja46xw2YH2gMaJ0fBi5sBJdbVdzhZRM1ZXDugYjMVUC2ErbPSmnW2vDj
HCwWC29v0AaQ4/roLfWlMPwbXLcv885SL5oSwNBAPzs+BFavbaovD+iPsCygS0ug
r9UVA8Z7okK0W9Hy6towy6rqCP+bZA0qCWsph3TPtpNHR4/TqcNqhSlFemZGNUxk
lw0FIOg0L9htCoJSU3M+E8qrMKfoCWp6RTapPVMWiKAok/l/UoBUG+biuagtCn5V
FZD1fKVHCu98ufXf36HDgZAlt8Y1WUGccggb7IqxEja/s55gnNAgp24DdkLpt+7D
Q0FMJi66VIn4mpb6597ItJstCYkFIDJSoBkRJ1qpY8ejFEquVuOrg4jX416Vxgwu
tZNdEN/5+WCiK/FkEWB6FU0cIIYnLkplpoEkpTU+nIJ/YR8yH/JHBAE1LykvncFf
wDBzXgAu1KJIo8zZwzlYvkhXx2byjTXup2Bmp6FYgaQ3mdHi703j232Dh4L9Wb8Y
pTzgDu9jVk4xPa6rJHqvXn7tWiEZHGAnng/ofUDRzO97JkzWeMP4taaNYqNBE3nP
E3GQyDa4jsWyrBQaOr1IWtoyzaKUDZIR37Cd9K2s8r0JF983CIGZoleEOIQo/0vc
4spyWSv7YTnVue5XTlQFskBPPgDMxm7/QKRgEqBczTiouo2QgWld5b1jxqo7OUhL
t41kxTCNquQnBol/K+roDNfvIDBLCbOQ2qwGmrILpp3uXgTYYSMWPP9IgPjcHPdO
d/SWTCCp7E/wpi8eJT4isf7x+QrK2C78uwxL89jphFre82flZ0gHsFvZUFG6svcR
k4XkDtD+19xu7g2AnLZ0Jhph0CkEHXAM6m2rz1AwnF0SpmrTKYKj+6g1D7BG7NWA
jR2hQkDRqdi88b/CWQYct7Hh7bvT1/MKe3aft3EGCknMCAbyfCEAmmUFjYbq/lu6
ng4h+RH5Tux0eoA31I3LOf2P9P4sqDRFCVFUfjVBvZ4UJzchBeQ8DBiMgxSpd6G2
ptWRo8l+xxMjRslXvPw2UKmNqWRv1vW1sXFMmoIybGzkOo+Cbz/S5PIvmnzF2OWE
BPkCio8PDfSkPM/fi34c8/9H1g3du3rMCfpasLAxfoH0m+nnMv+vCqF3OPOalytG
pSECMjH6NCq2SR9R7SOlq7pynL5QyONsU8lNfW+ZjfR/MdjQPUxwH3a5js5tUHP9
KWMmE15wJAgZcJFRNvAO420W5rfGEFC8fBe5dScq77QMA1m9XNLRitL1DvdyVm67
g1mT2x4V4yXnQOCzW3LtetNVPmDiWpOw2LOvcPm/DgO7s4huNGJLKduV5R0OAULv
WfBBUsHEKIkqMJ3UTGg7gG3dAfP/f2ZoS21v6OaSekEO1zEX2NG1+UNysDqDzBA3
f6DizpB5EUohZbMsi/qUbftCVibcqMysjgtAvKjbk121cCa6+bxlx6r+K6guiLzY
EkGUantL77jIuvBJ/YoHWQrwWeYQz+62a4T2bz6k0FsM4Y0XXQ27DH3SjNyzDyql
ITJWvzKZ8YxPWSRzqwLoMsSitJdohsgd0xqmwbRuHzjPyg6Ydey5NAXhwxlbm/ai
CnVMPQKReUPbaoLZE4KObgFGTGEfWMGgGksUeEXon7UfYAl0nupVAptJP2skROlB
cFIwK8LPOExhRSVOI3Zqam6p5rqxbvSEX3WcQkISHbg0jeNswmw3YczzCutargZ/
qUzClLipJ4ULODK7PZpesIgfu0f01VweFw8+Gs4p4xsKCYhAaQhl5Ab6SdWZep+r
aHMJy0msAv2gupgl7k42OAHx/lEuKHDlUCyQzxJyfjMQ/0uyOmh8sLynrvr6XNb1
nRmbljsBQZBG6ic3mPsYg1XpIzoTuIvWwwMiuTdQPIloB/d8VJC9HtBe7DxXLgmp
8386DfrDjgISjF0ENpBpzK2ZHALqs5w2F11GcVYJc4MfL/FDhca4O+R8MH/yM8z4
czTAHcXbp864jrHOZOczGU9qF73fmI0ITPKQ3nAfMrFGlVsKP6QuCEeir3KjfFxf
i9XnDSWrjo5vdBK9upip723O6TY1qWAz2CbflBvBTM8bTzXk3vC7iG6SS2zSKymW
ZsXMvDOCEPdlW5sIajK077nvRzuqv/Vp+W/EbnVjDmR3bB8lD2lhfkQlj0JkrbgF
pML8z0k7yMDyX+hQ2vshl2DyCxM29Osnpu/1j1WRB4jNqrz+S1BLwt2B2qRNE6GE
DX5zlPsBNfoHHyMlFUB0ee1AZw7mZUtLreaL+FLmyV5E7C3d56gRx21nllT2iQ72
Kmn45kcib+vD5n2x6svyLhmyuGZsFcTbX6fy66V/x8E1cIfUxWYNhvgLoHlBTPvl
gkmidvZfQ3FGm3gX1P7V6256ASw1cbvaVgjHYhuc7rEkeyZk7P+EGx/Lr1sG9jgt
k84UWgMTx0I0ircbc/RR/kaCeD6mPNG9knq2oLQoBtmhvTlp9rGatRAgwpYo0msD
87AhKT5Tkxpy7o04SgemjxfBzHtxPONC9zE9Z4oZPrh8x0R+kmbDc64yQixxbGR5
6bZ5A/ZT0hoAho4mtXEFRtvqn/LS1fIzkezP/aZxWKccARybTuoWuiBz210U0D25
1TdTzZTSJu6/sGYXKC419GyWj4CwpBWnBUSyKfy1cLM5m0LzVaaiteSr+mgnyydT
bD1e+2BYPJumDpyRQDsmhkukyK9G497SmG5kAseu2R+Cl7CQDoXP9ut64c7nQLCR
ZdS6hHEdOzZvyxHSWDUCC9I3cxRm0IBLBXW+yOOyonLo/skXuPnIe9xXDpWQ8gfw
iQvJXb+7DttOUpCyZd0fdpKyZPpZ3TImN1SJKlV0NNL0O8K3DSwYkggWeSFi6cT5
JuTerrRbjftFS7Xa6lfMkkVlMzmNILE63ebLel2zEBbNBqaT4I/+EqxmMHl3bcPI
ZLSFm3OdWx0HLC8xfX9I9bxPth4otM8pJfmvtRCNy4bKAI3sBeyh+LVGVvw8j/mr
uPPMkYRQk1j1M9OhZsx1FmKaNbX1ZtdeEGLFSXVbBSUI1sXv7xQxiK5AIn7QmlcT
V1Bdmv4+EQXIfMRh+PqEmjDxxX1fX+Z698msH7GK/1xNWbWcEn51vd6MDPkRQbxN
Wjpe0iA8e0OZZNmTRzy0r37RhDJtq0CG6nnRjCZetiZsuDYQXGP+B/AlmjyMvKLA
k3CuraGNqm1JsWGo98VWBjGdcmVeS6X1h/hr+K+QcRfwoScj3VNvAnJ/c3pFKHez
63f0Oj/+BUEmV5lTybUtANkhir60Oh6+hF3By7s+iiAEIXl3550Z4eBnrCjIl4+U
lcgUNAC5//t3+NdnENI4tQwwEYpLZUiXySNod74o64R1Mad/0t8dlyakHZs3Tmgx
tQc+Tqu/mEQ/rwSi69Td/gyNhu6EPowc+lyzju8ldfRhu6lYsePrdhz8bNaphosH
ib9hhH9DZ9RwRJrwJ0oCNHu0CwGSGwpVMKtk5KHzvw9Gt+dvdoVPbnM0Ppb7bwxg
oQgfWLUUunSwyw00JJk8b+tgVNLotFCOyuUAQmycHK4ZAry8AXrB6lT9+Qy82/ev
+G0evdwdmBLiJBbdW+ZPml5sA3hdEC+59/44fOa37G/ftHUyYVB2BC5dp96roe3x
gr8mXfLAxFuzAQX0TJQJaAckWyJBQUo6VjtvGKv9Z1s9BwdcsbTBv/ltPPE0l9Lt
bs405DXJpDrae4XAjd8fEym6Kg+DFuoNPxGCCWWUJO5iXT9UdZugupMBAsorsQd+
LkIM9uMpWhBXQHvsXvTjLtw/o0w9zPYqYaNKhhhl7NXloBKnLtaU4DK5zaReoSNc
aZS1znh+s8iZiyCXghw2vvG//MVTKqTu1L6bKo+4CxmCgfitvoSgheCxqfxr2rPa
iv9moh6YXQBJF6SkJgaPDEBFt5xtEOMCDeDlu62XI261ArHOMNS2xYmOiUQX3jJW
eRtuRi2YoxVT0fgVqOucIeCLvhurnLytgDeevHobxZOzdQTcxx2Xz/xqpFi97nwt
YfNIcP3nyqPl8DjLBLnrZaAeEOjDaAPH/dIBzUo+aiHBB+FliiF9Xjgwylvq+VBv
s7hrNo9C4LQ9ryV6oDl/z5+HjQ9eKBci57NDSz3c+odzyWS4Mgwfo89zSVv9n+C5
hcKkES5XcK68muzeFQ/66SRbxrPXuy2ioHMtIWXHt51ItSrW7bJiHKAncEohA6tp
GnxwCOEJFhVPEbos/9MsLYw7JKtHQnNS/g3FQqedmJzKkMbac7pif2c5BrGXCHQO
CqK9cqaH8DFiUvdRzTMCvQYI0j3S6UhpwBkBTRf/8nd7CLfY+C+Sftadyys2x3J2
2rGxJLC+lZL2vtHQDsSFaZGITxrXTxkrQ1pIiyP0Nt7HRd4NZ6Ce6fMbNqdDt2rO
IBa8JTETMfD87kGtdwwz4ZcydEm3hGyKjyYnavHEEJMJGC3SPNVOYXsfxrR8y6Os
FR+qS6vcAj6xK8o4gK+mp/GcuYcHW8rPDUI54wRbKS0RttuVW7K1RRNdRQdGyytL
H9ej7yma0oGf8ehwkzhxHVBsiEe1QdivX5LNMZb24KmYx+XVvzGc0v0x7nsHYgM/
M4qgIG6cyNM4Qdf2hIP92qaXGhpN9yxJxI4wz4BPcLiXB4X+0O/MBeDuSJusvZd1
IOJZq8hcn+1ngRn07o/sBe/MY2EcOjVkSHxvZCce1OkvwkrdEJ8F4Gu0HtTMg855
Pr9X7exQKrOhJBr/m03yRpFTRroZ0r7pPF0Spet7+K0DVzPXP1swXDiDP7xlakNI
n6Qgn/CKnxpDJgtY/bozYroN/QKzIIptOdWDjTqLy6AdaoztdJKP2bJtGIDd2FPM
z6F24G0VFVy/Nhc1MWEXC9rPYjQyo1R9LajE6nZPeJe7wXLIF4bsRfl034e4MzYB
eI75RrsyfEvZozd/UxqF3BP7IxGWeORsA+tq5PuPDRfdpdbM6URe8TMc5GdNocUn
JN9n2hQiwbrL+g7/wD2hppywVkeRZq2lqNE4G5KOr+SNVC6aJkHB/KxszdR/NVEV
M5/L4y7vCgTKL5gjXt3sBe3FfZrk0E8js/iAfdF2zPANQ8CY8NiHb4Zue3XkeG+2
HwFTM3DFCgz0kb2llptXWvMVlU/oMfFt7Tnw8wGAaHViiR90Uonfa+1ERE7CEYCn
37LeT8z+O3bKnP2/MQ/g4tk/NJH60Sl/vbVi9g4gXPAxfayXLU730B7aCUyTF7/q
8TTZtC4g3u8nQOqYaaN8TGAc5RGuxul+Ay388y2oqMsIodUKxbYgmTS2kj8E7tMO
EPUXoFXOiuDobrYhpp4ERL4QkxLkNDf6RXGZZA6s35AevAvRYrCl+v2PO1nwiFMj
FoVwugP8yi4y/8HJX/beFQRqHsiMlnJ0PtZ/B6EgcHpBmtDHNnf4yVwpzVrCzKZy
/Hgeics6hNC7dX2EzMhy5KIUg0I5z0E3lOpghchJZQV8kwmjnarA4T5yhEa/35EM
qWvGYZcvMFGvcN631Q6WtIfvX2O1EioJF/XKPFHWNReiHb1UtTB4B8/AnI0vUZqS
z2wTsX4HsBI1Jo/shfwO/v6mimUcoSdIbAsOEsHXbD6Hq9X64YP5jgbxXODu3I3t
50TRMx7zuvgCvfl1/v+wN9esN8oIQnVD1Os9a8z4lxvMGwUR4is/mqflrwPnU1p2
fRHwTbjw4ktZDx6obKJ6kf/gy4v4cHV4VZOH6HE8FWlbmOpxNsWsvWqCWDP+36Qf
6RnluSMRGiUy6Ru9izkgZgiEaoS/sNQK0sJcCD5Oht1fPmnP0knn6szxqKKQAxxi
CTL06v8fJutJlJafP1vvV8rg56NXqzBrFEcdIzwv/Rqs9FvXO1s6wSzEQq7kFaRM
UAZWQsPmN8r4G/8j5e7bsVICXF7+csL7uB+wspSKHiHapdXfOvd7n0pfd9zPvB1y
78wAekiXztEHIVCNLGeAZHHWAavUTUxIOcMNmRBsXBqT0aE5vCE5WwIbnVmvM4Gl
XTDo3FIfYA2QNdt4L7H0y6Xf77Gxkjv+3Z+P3sYrs66dOqcQ1aTLMNuQdnHDr5+T
4zBTWYG4/43VPdlUZhys10uDRHylCbh3mr2+HZkrKqmYROG0WRk+wx2Nf40YIA6T
ksQU7GYOf2k1+ZGsiaIv+TobxfBryf9J4Sxv5vSVzB9iJ2hNW6rNnw6yWHxt+RMO
cRJdWgKoFXdKbiSOW4XMm3KEKbIVYd1pTjoSvooM3vw6PHRChMiR7PHs1oslXfho
gz3dU6uSSemjli5XaKdeta0ktyicYHTgrjExS8YcoeJd7J+dNE/xGQK8Qnya11YQ
Z9tGj3nA1NIxxeAR8QhS0TXFrIfi9PNPQGdFMObRHsN4k/zSAZBBLviDEIbipISG
ZwtgYiNcYbGdUXQtcSrkerBTUgxrhvfK2YHG0zTWZwTMPPCyMRkfYVgZFaXf/sFU
lTfSzGGUyLYRCae3hc7ABySoBNmPCB18yrNTmS1nLZpkEqS5V7oZfZIT/6KeODtc
bZ9MxCZ0bM1gpjRD1puS4wo3XVruki7XS2kubmKQECdcUyP6FPzPCbI+V/Bb6PvG
Nw/8b3k4asEIhCSPx8XJ8uR3bmQwOP9mGzIBaBTf7AbkXKs8HsF1uOggTDHEdd+y
K3i3hqHoKUHZcfDRI1ujY21aqvuBnEomP43+Xt10iFNVqctIxCVqjE2Oaa3PkFQd
F1Qu/iJFx4znOpWBiQWXzXlJVIk3MQhNOie68r3sPumq8GDRUk3qU4PuDadjufOo
eUgyiB4AplKNkX++W7rrg6fZvCGnFNEAXkNpRQmwLrFznBlxBkzL69twLgpwqKfx
FMIXriz3JycWaXyOsXG1tH/Gu0qfoR3vlr5XcoNM8oGSvQfUJGXITtTlpySpylvc
ZoKMA2ef45gMm4bQvppfH1kIOnbCdesu161Y0uK8W16SRCNYNfERV7q7kdJ3niRD
3vInJjVZYucQdmVuwQP7Ywidr184V6jmaduK8rlvgEs4D2oZgBNyzLeP3wHF5a3P
fVaGaGAPWX03LuUWHd3yxJMuTi2tiQe+WRPDOBXpewemtgG5oAGG2KeSOCwfoWXI
Q+c8XeVROOx2MC3wMNpS/0GItLKdm44AXlhZQkOenYsaEzAosMFzYFq3Kb3oHBNU
dGZIIcOaCbzYJM97HJb/FIzeHu0D5x14yMgGX6Y5fvvImexQLErXQ++lSf3tjcHv
fR4cbv5getwy2fRN4GsiDtyQfTKnzTXkwAzOyDoBmG7htzgxDVMPd97NKJNXqFlD
NfruLJ67zYf9HB47hIIQkRB31zuVXpvxNJxQAPOy9Z9nJ2RJVi0dP5H5lw7wxW/E
pz0B/EAC/yBQK6kSBU/bDgk93esOlVTi+MV08slhLgkF+ZLOJ5FwBBzA95gpQevh
kuHZZS9x7UJU2wR0RvJ+8GJUaqUS1Sd3eobTExw6ueRcUVKPVhHD5Frzhgb6H6ID
ED+9nLi1EOgTEMu7EISnBxfpPUfZrpLaQeA+Ve9uY0YrJLy2VGgtB11RSLfopNW1
X+6/ArvfkxBowN+hRt3MsiwuDa+dBr1yef6A7SqVhor8J80d1pF37oAvgVrwDjpP
wgD1JhvfSQhaZSWasVN/g8PvNiEEkiVZyfv63yp2bOdEvSds7J63AqajKO0dUK1u
1ytFIrqRrfhK51nrxbKBGfUBCVXysHxIFID2w8pXd1zKoh/sGy8KWUpdHmVDS/Fl
9dfiCXBM22gzkFII5NHfCHXucMfTuHOTnfqdm2aaFDMhmNLiJDWRmbkfBE3rbCtf
4D9DobW4N9lOKgZKrxN6p9nz0kAFzg/nIwiX1v4M+XeHQ39K0TrKPjAUwpFijk1C
xHQVlZc5tvp2GiEAc9A4dOtb9FZA0QoRDFa3R5Pro5guCe670VNdliMC8AEz+3bf
Wo2ANn0m1lWyjXEeYl3Iy4H0hG3QFH3ZWPBlHobGRij8FrGt1gGq2xPzZt0XkXYB
dbTTj6klxTIQTrnDvxVBL5qycocfF7GM25TBerW01YMwvHMc5lrNE6R7XBoVMBtq
MCcXzP7wjqPpHRDTl1Zhu2K6NorxdAXLwPZIVLmne9qNwJB9TgT6B9PbvyuwwVjB
NNFGSQ/WPTtbpFrEzNgN2xtn9JfnrglFjYnDHqDNH9UB7KnspBUnRtw5RUr9zZS8
5ZYWmI04ee8NoroOkjeMe8GsvCqY2axLAd7acDOBDtgGxfCuVkzzFdzmXrUfoeW9
nyiS3NfIBrut4LIKP4REvq/wYZgRwC18hHI6YOPueZjZt/aEO6/QJGpJmDUTiLGc
rTAoIKL9/FNfjwuSf03USwAetmdbCONdyc1njhCgHqe65QjpYe8YCKTWk0VBOOBt
epf+sCkhG+xn6IugNvV7qDq6TOq6aQDYN5HUZWh3UDNacUFCokXSoTjyagBPY7o9
fqRbD2E34QARBGeFUEYwpoeP3JZgitWw4rEscua6RyBe7eSiqsgGMe4N/Dc5FzrK
TnW7RvCO3Us6EcoG4LI4eUJWcUDxYr93Zi24OupKtAlQEbToRewuBirDkTa7xnFk
NRJLS3m+F1pxgp14cQZw6PBjWQVsqv3gYaVdoVjHM6qt1ScUyYDi0l/7Dtvf1daH
Qc01IRMkP4R0UNYUmdeiWvDS9D+rNFRVlAdvtN8C7GlemEW62sZlzXnWETTtw6rZ
Wfwo5R8Uh4tcnsKG6HVThxEFLvlhcdxwDzzQr6KDDvMFRBHeybcyDTpkvuzbq8Y2
yZuYZ3JMODdB3vw2DcTpdV+87dEUd1PXweiAGJn8pSIoFRYZG1hv4g38ZArFrRpV
tPVCv0KQyudxH9kQBfmW0whu+4j8cIicrdL0ofCBtiTYEEnjlg/MQkoUCJnXyIGu
1dhq7EeW8TAiXqgCsqfgHO5SCOyyjZoSSsOS6bNyb2Riuo/YlPO6kurMIWILde87
Xg324UTZi7p1jmibeSReg/1DlOtktujORGpachQlK2yI2TCSf3de7yjvJhzqx8Zs
/uJETha8e+DRuK+KLRr9sA0EtHmyvYN3G1KbnJJMvTl3Qi+zGTI8Ji5s3yqfryDN
bEgNzkt5sUr4cP899h3KPsisAxSrGTRQQXgA5GsMgHIRglwPy4434DR17fnD7CmN
0RwNKwsOr7Ofc1+B2AWQX6rxKO27Qt4xPJRe+6kSq1E04+YdjWoKpyWN5UMWQRUF
QRghleLIjSEUB3t3K+nbV9nlcjdjTs3Xu6Fn90uUaVN1mhdUF8OWDFH4Dj8dGkBB
H0DrPDPtpnFmPRJhE0aakL9mlTIEd9nILaJuWi+hYu/I8pklp6upI7+WqXla81uU
vUBMx12V64kRC7oO4+dqFBbCAsmJ0+Tx3pPS+NNWvbSUZ77hKmiSuP/ym5NytbuJ
VcedsGmZUQZCKGfDHTxw2X9yhk7iIwgJnF9PElBiFClDRBi9oDUQrbXjO7JCT2R6
CnFphz0odfr6Dvb8FaiaXNZDOnPfPbrNpN4++PwTdK2f11aMuzrAQl44A2TPuH8R
67eB+KRZVHnuFQQDgXM9rTI0uMQQmI+i7iIi2fFlOBW0T1/1fC17wcjhgDDV0cMH
9ChyxkOCRbBTBVbtYy53b1uuunyV1b0sTNQtTZ78g9KEoJL3MYCQ7QyTfyzQEKOr
IIKLWS9vS0C8IaMUrqjFFs5f49GQ0xsLjTmLpRWfKNLUpHFkyTqCajiB3yaN8oAT
HBbYjEffGKsIJiQxE7HTK9Lolx9vtgS/sHz47ucSTXcmiLQQ8WFnf9tvCsHTYeme
kNUAGfAIluYHNtoCpkjWK2xtIjinJRH5IiPi12wG3XFpYvprCLc40rRodcdMMAcz
rop6xVqH9ZR+2NNIg4b0YB2vX0otQdLftXCBxOpvvmxu9CUo+bW9eO+rnYRxsRoH
rv5leVcNTj6SGDUYQgIg3cVcolpga2DTwnIxhEF+S+SIOYQ+TkjdgfjAZBh12z9b
QvpTLjH0W01pKGb/lamlKsOPTkuEyKzOpzof+1r72yl7E3KPnHNd6usmQgkgCIPZ
Ud3xw4Q76/sD8BuM7+qd3T8M3gP8rfNrfLo2TBa69CQsZ5MOlHySsyTNW/ioBsR3
1HCKr4APUTphs5iSe/YZhxMyR5r4WSuggU2W1JBdsWaWxbZqhdUE8n3SLI3Iy/6f
lVKzJfM0sPVQfUH+j13lGc8YGpp+vQ8sKBEc6Axk58ZNM/a/W5ITAHQL0VOgUjEr
gIZ8YA5dvgO3gbOCGsL31MujqmE9sG8N3zoE9unl8lkRbo0BnavjzShNCbG3icXM
qyP/m3cIrqjJr5sFjMdfIB/Bm5khNDeJZnJhfpkrXHs4TlT+1oL9SmzlPrpBmRrN
sE7QyVbjFEpM2BXBGfiBxujRvV8yFNsw0qT1WqdfAMYSCj+aasV/2TCzx7oftKe8
fk+eFET1nvVv8SIAlEWDUnKj79ri78t8za+R5RC0P/8qFn3H1U0A1ti0xjUiAeqz
lJx3+nWTFD8pA7acP7ffV6VWLv2f1getMJSSytoCxNQ2vdIHNFPWEgp7IcKGYMa/
hr+tbFLp/3M2x3pEV0CsRA6Su6DipscXtcBz6B1y+EcjTMa7RH/S14ytThb09ak/
igUhfAjhZJ8CHX++VPQM18CLAmT+v00ZydXCz6jHFUTnpffffuSNNtyqf6YKt5/y
gRXxi8RWt84iGc4L66sHuORopY0gQhSDpZ6jF/Vm/5rxuT2AeXrdXNSLTZwrKNCE
M3+m+8RYaH5mbHhVgdMvt16yjLfc+iPGz3ZPHA3jQSLbW5GmtdJlhhtsI7keV0HF
YIKJd7scy7bU/+T6BgDfF3o5M6ZvRj4I6LIZF0Sa7lsd3kcJrcfh15ZsB03+l3Ga
olUtOPo9FRO8bxGnAjJzXJM/0ItBXkcfb69kFRpt6JTqPXeytulbNges6EhcUk/e
6v5SgI4PUx9azTk0L89tIujgXYOMO+N+O95O8fHgDindJDoVrz67iZdloqsdKRJY
FB9C6zrGRU38nKF/+pwLDEgmq4k5jlIJ8RkK/EEo+v6JwhlTljZ68l638ADaIQZx
NCPgJYuqLNmOKJAGWnFjN1QqY33G3lgTClKKs5/s9gOvqOaMEqdEAaX2EjL0VOa0
i1pcM2bvZhqpEQriC1FGl1NYLhy7YSohddS9pa3KxjlOcnQI5PSauu3Q2M/zqh0m
AROhvsa8HK1sdA+D3VUIdIvMhQQynJZxoBm2nGKOldPZyFXGabOjCct/mA8LW6Jh
8AqqP7d4SWozHwjtGBflBkLovoUNtaas8QHhAp8Y7lXUjAInTdNZ+JKpUJfKwUJo
YoW2QmeXSM64MiSzq0hEpnFBK9aVvPy9i3EeSM87VtKbA4oG7MAT8ngYZsNdU12b
e6zfCKI/qL7xnZxAgttLTG4uDxyh1U01MuNhx9oI2c/SBm75aAVfjkTos3PljZ/4
a4NInrThVvpf9a3c1wziTB4tRZkK2d4fbEXq3VXX6VBoLRbqAvCvYlQZC8n+RVGh
1gr9ggsYrKjLpPYVZ3eZik44Ugm0nVvAmFOULbCK3BenvyWeTYjtvH8PdJI6GsUa
VY9D4lq02EhHd7qnSSzeZHd+e5GKG5L/zphlQh0vw/1Yy3Ptv2ID5i843kH/JXx9
0B+PndlPW5i0y2k8KUDK3yzbcctWga0gBMLydOZDw0vU1rcltS61v6fJSA+SMzYc
cIK1gC92QW2UiwsBeWg6ergc2VmidDfZEsGsjsxcQj6Oyhw9ChiprAkXBhw70PxX
wYWSwZ1QYCyINjSzMD4mtIis8Nv3+DdomQwOqYPyIV27pwOmHXECovKf2SuG8v0k
D1HYEW5pDR0hmLDIaApQXigAfmSQDIhR/cmzHiimiUxL+tsPSmM4CMYB2uk6+4K4
IJnQiHJFvTVUQuYq9EUwuKpmYpmga0LN6j/6aEB+a15rEhE8geGFfGuTVPvG64pc
vRrNc1bAcyeM38JNpR3BE+U9OqZX7wZeKHe+njK3O1POZJfx9dedZgYVoVnpDUrT
GHznZ+bE5ZljdTokMtAJkIsSct/ZHEbjzf2o1JDXDKUjw8lotUE+XQmm174sk14H
crkWdgi6rKrElRu4Hm6HDUtPCs1cUUij33ZNo0fXbT37SSkOgVzx4XytBTwaonmj
sGXz4cnIoFjkzNNGt0srln3/jX2xUcxM0peFsmAceiU7TKIWUaoq6XlxwFzR7lCq
X5Yhi4lrESuFzu8D6WTjhTVLdh7sHndJ5MDA6NgrPJQ6VzVYgumQTYTjYBWESUW8
x6JWQCZCK7fTxRhwSyoS8NlRKH9ZKm9J1qYr/EWaED9HBEa5NbGj663xbkZvOAky
InqfTQD1J1NrvYsPzjCddaDOUALYH2/qAsX8tRL5lnJtfJWDFIvZPwepg/rz2QSG
YvyTEaEhbNEnqEXzNYzpZJDfPXom0b3txqv43lBDlT3lj+icEC7V3Q6EZUq1j1e7
V41ZJD4GlTDkUQGx7Ys0l5QfssqqihD5UTgtVabiaKsbxMMmTV0qSX3C2Yr74Mhr
JoNonTAypaKjUIXy58TLzEbc5oS/gz1smK4NgPi3mSD00SkyMvYXUIysY93V6wtA
4QOC1UkkW6wHFZqpSHpLrscUrFlT2eXCUT2ImtzpKDI07T93UWAFHsHEKNskcl41
OGlwAdUWab3pah5W+mRGmNiTBKdsRWABz8flCh/b8IBDxgw9ZMk0eg5Bha3dofQF
3/V4fnVPPs99ErCGXjjL6OJkto/bp/fJuFFVvJzDm36M92WbWr48y8fSwR/HfyFE
wHS+JpO5Y2f3AUR/B735veWl7BS6L0Iai/++GBH83NUN2hLwbH8mlGhEmCJzUUuM
hF9Wr0qVppKD16Dv4cYWM7luqPAJrJ+AI0IPfLnMwvXZK9yNpHlgNYe3C+HTsz/Y
qvd2K31jTpKGf6Ton2GfZAEEXhI9I4N0A297yF6RgvLfKcUfIYiEokEksSRKNBeb
u62Zv+JGN6dFbzDbTFKvOBmiAvi/JrznHqo/siD2pF84jIKIQ2aksV0IUoANbedE
8CVl6lzQ7TqLGQ/yP6pXxDIzrxE5ivMqtly4/HAm5/ms5nmlqzcggn7Jv64K8I2H
Kggwo/DHzYJX9j1oYa4yfzggF9t42gcb2N4/G9CV5AepS1s44tpLMqtDDH6E6pVI
xG1m9wzMhY9+IaWN397Ri3kTPBj3xP6iIPSYn4BOJrs+pUoaq73zHa1wP22dxTrP
nj+462T9qmLOK3JmUzTikYgA0/Nu6TWxsACDyBY0MDmKF3f5fg8jFP2x2k75nfk4
O3sWxCc6eSgvPSz1tFoachiVLD6OxoTkwad76W3ERcVVoPjM7qQ0P75IdeT4UK8X
Mu2BwxAOb4SfRgJ0OBoBINWt1XxlcJSlHDboLGfl46c9nM5/KCDXuKLFYnEEfFH3
Kkh4QUz8Pqo6dYZZGNDAg9KxHxKy7IGgd8MEPSDFNOPDHl/Xoo+2QJe40T2SNGS6
eG7UeQl+1JsLVviuE+hbO+h8HvjCpu1ozku2LQkaQ7oqI94mZ/43xFuhMkHywTM3
HKMpsDChLTfvVx3FDtaVj0GqedVDp66KXOm8bnn5EAMTPl/pqWCbMIQADMzNnarb
1KBQR6+PQve+/JRVNE6zRQdHxa39O1McYbkAf8YsTygKCUIvIN4G1nhb6ToAXD0z
tDYD1rc3i0L+6YIBsVGGy8dhmb89g+rU3CynjJckwofBTuwI56QWFAZiWoBYC7XG
M02LqzMf0QW4I0zFhBl5O1L5c5RCkMdNWNDdvp6mPDFANr8sETVaD4HxWOh1io34
NLjZjP7YKUFQqPx4rOBoDSub7Q3Av5KBAPkgDeqYy2DRNnC9O0sJWBmDb8u2jas+
5tlMHVCTcbdkuEatj2yXxPRbGswrbhf2dHN9ALs4LwxaxfJucBwCI1sYvaK4prlQ
ZWXncK78Gr8W2aeeAA4a2mP/YN3TAwYXCh89T/Wj524rGM4neNOIA4zQslEJ+hE1
vawI1I0nzrLp11vfKehwa8nno8KUlveWZziN/lrWGBqp7QeYT8AFzZ+2ot+cuIa6
uTjb1uRbeDR62q/LP1fyar7uE1cSRY5j7NTyjnZqcUEj1YUVM8UBo4wARB73zEvY
nHPY3XeKOlCt3/Ud0ye1XrpcrmhisIcGmO6g9A88Qm1Gvhnmg6p6Qzv/yAD+Tb0s
asNUE2PXLAie4kQbdFHZAVO3rf571mefnxal6sRTdRXANuYIRCjwxThJvFMfY9EU
jwOAOCHBsdcAcUOf4xyhqEdA/ByshtDGf+Ve6dhP2XwE2c4WK+88BFwiZCbHAu6A
SJWVaap9PoyqrtE1KpUe8Ol7qKtWeGSrt0D9kGVECng7xaeSTHxbhsvj64FDeH7m
HgraWfcCCY5TlPynchLpysgpnkhuhtBRCoroTHJ4xFrg3jx6Q7bLqSZeSZfV/vJi
3WQAcNd06QQQlLkFAMRNunzpKE5hZnTkyUW00gFHCecK2bSL+jnTWcKcTt5UL0/t
kb7g/S/2KcZxzGdhkNelwdg+WTQ+OGNXOfxn0l5uQlsHKyhFsfKZc8waiKjcr1Gs
fzFLCC0Vj0QxdmK9w5B1mVqWqpPBedB4j01lU2vDvvH1S6eHZ6IyOi0vhaaU8gmM
OzYr6brIXZJ5dXEdCYhmRhhb5dxlwX3O/avTLHmdMTgXFBpojN9+ONeK8SJnI93D
EjhXW9ypIETJKrDumVxDkJE1SU3hQos5ckAyrd+CXHBiAwrtiL4lm6ineCSfkgOB
+pKTMZse0iTJ/2oo1UMMlwc3dl+Xj7QNl1cA6o2nh4/JEXPdWk36fTw9BwoNzcmJ
NCA3CBHFPiOsmKTne3J9iOB255fEirokbcIDdHUZcpKn46rNqbVgTHWe1GLV1z4d
D5OSsXMaL+C9YThmgJgiURS5gNWpa0I8sWIJgjtKZkNVUV+gXQ/LKK95Y+X2StKs
143TkCUqDpRhUqgfLUlzzsHpZjrn8lzcF5pO6wXiGcKdJFjbibNV/P5yRc8MTSJ/
myFEg7LlSyiJaKefQ+3+TRsESLY5wmkKx1l5LSVIbCrQ7UEDqkExhJ+HA8lDE5F+
mNYMGevu00IiJTdEhuVdLr54FltjPAAIkHNrFT8U3ufELKl551O9PaNhYjnT3epn
ZtI9D0EJNWKx1AkJIHzSyOTj53oXeDZfrKFxWdLZEGbwARfObRdb1/rUEpAEailR
LKDkYkH7H8PefwNlLXuYY+hqAmRW0n9hU9P511OLqBxSqRlcyH2nkDIBqflf8cxI
6HiIXw3lyOMA6gOJOkqAy0ze5ULfVw8z24g6pxyQoqzegZO5wk+nGRXFwhyLEAu7
3b0G18QM4m7WmsVtI+VYo+71sg0rkycbs5HTr6vurFLVksB/rKj/t7E1wZ65FTIW
p0wVRJ1Bs5MLDcwhI1+fxzS0ZDA/XXO9C6ZC+lurhaPMWWRc2v+qx6OKGsFtoU7v
xTDs5/SZYXDj9Q9ev+UHBOyVh+Jev3cQa8/ujn1EiTubvll3YPAQhQGnSfeUVCpZ
laZZ85CamMobCdQHtE75vLXhgimUSyAPtUsItYTJUsA5l/0FHUaMuI0jfRtXD9CT
JTl72W5XSW6XWnzQbSF3lKtjZIhOz+I1XBYGLyQOffZNPu3fyMpN41dD/XCNyV84
iCqiqM2hT9qPaXY5I2LX5Wo/I0627y0TuVhwM9/UhC07yYCja8OFXeBm6FZa5EH5
8krbFB6Z5ird9AugT9N7Sk7Mor/lOscfzKqBj2SJ2R0H8QkrifR4JBRJk0BVsN42
NBMbpneHkQugdpcZo1G9K/AbF++mrftisUrig6OxG5XJb+zz0m18t4a9TB+MJBS1
RkoNZnGre+XfOUWiUK10ANadAG0j7syeGoNeSvXKknIhu/ihnxvY4n1jZquMoUsZ
4UfWJIOGIJ+WA5o4tm9RHWRAjMBXQFnDdMRnyM2poGYCKJfLxt0B4WFKJ1C69BA8
0vcaBx3lwKut24VJzFf2QEx5Qo8gG9XEVsSIe37xO9N2Oa0Agh54hVHVmDhaK1KS
kKxAKwtrVSuuQ4BdvKh1+lH9yZtidY0EHBcw8WScDT2Ptpb38pZuTaxAZKEvfM/+
81YCt0pCj1x+V35v5HomEMidCexanHDeS5bvdzKATxnL/manCG8Wj/82oKVa/wa9
tzo8tmwuJDzr4RrTBGnSH2ehwo194lwfa1UEYpiHYlraF5qPDQ+Q8q12/QWIaFhC
MaQQTXTN9ggWBbMswVmmxCMgIjUrdZD6Bm1GnuZRF+eUT6rpcRieG5TchCKmHGDd
2RbhD48ak+qQMHA95bkIbsRQhf340u6oBpN8nvnEQm28wjWgtKv6AIJ+pkpKpb26
h7oxGD4djLaj+xi2ksNJdqIAeNw5HuK+IABENRbKAuVkj1G31sVagKt3q7XPEVWi
VCph7I00HdTp1OlLgM8o+3hHCuOfrGVADH7826iz9mNtUguH6a+rVnexUJwgQplb
eQ3S0ZRGdjDPXgeJerTsSWus3fyD+lD55YMdyVoL5vNKMAN85tBEMCxUkf+fCIwI
jIL0iA2E/dmnFQBPZuP8nIQY7/KiiJYY8hSiK1xA2nYkLmhsmGIFg9HqDJYJx70l
lgabMPTx422kYk96zbZL8nCDQLPREC4kBw5K0TeZl+UYvmiT3+yd6NMxFcohcEz6
gXHM0X0dX+6lr0y78gouyQPXFxYWn8sGADq6dkvqgcQmXKwqPN+DxVFXMX00sx4W
qJftsK9qEyY0EzR9YDCGA4+gg65Htznm8VdmCeayUybRNsudnIuFVZr11Jf0BMJj
a5gJR3hSbHF4hW9PUmQ8O/kki29UN6V3H5qtfpj6LdP88dNE/2AXYqheDfcSpykQ
VryQh1XoiUwE89hTdO0KcpTouQ+bAWqF2lZrSkX4t3UtxSDYLukikZ++Nfw2PQW1
AFGHBnpg70NOrje5UoL7Ihjn+1TUX46BNuQ0Jv4ALNK/QMJfCZ/eaLROSR917Y9E
0X2MWCg6+37COod8qeVscx/edM3AKTzCQyRZRiD6YPaHQJ+kq0UOCntBOKdRscBm
5h9+LKoSLq/JvaHm9Af+8MaHRhu1cpNNxuu+eb13utcFJ5PKksuCfnadtLf2ztTP
JkYje2g/q96A+k/xujygPNIt3hnntkXaDsO8y0merNJ01THNQ56dfTap/QYvEHlc
oWglmlv0a6Gjj0uWS1UBBzhlx22NXwCQmgIs2WdbkfxCuqR1MrSEFQ23HSx/VJ/t
GR62jCw9AmN63DP+KpX6relRDT/un1+R4bxMLO2g+DGhMk7kyuJQWxVNYALFbHX8
MLrev1ibVCcKVGi2ewPLBcSigUZu9ZxdVtIUE3768XwtJxK+T6GJJnVzfU1zlIMR
`protect END_PROTECTED
