`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qa2WvCzJogwWw/MraplFVrvCp9ZbEODbujilQxW/+XIZPT1EWxGCNd6IY4Tu1NzF
ZIerfsEqKu2NGs9wTPiqJJL9ZgUD8MoPVtg908Sq0Up0e/b5mbCc13lQcok1HxSt
UG8iDVY5ie07yueeM/b2az1gMAv/Ud4wsrFP4RdrERqkSNYsCiArrboE2KLDFqf4
h5srk2TEy7LMcKaGkCck/K5ODZhadRi8ywbp5KKKi8R5bsqYGQEiEZ9c2JPvKfno
bjxBdcjgQ9Uh21JlP7/BKRp1EO4mS4KZU18me89K3TG8ZT5p34b1+Cq5P/zAPeW9
Z8eWZ/uQTM6do7ZFBVuWyFSkoq5l9aIvk3Wy3S6anctv9tfVQraojSh0gMuXo9a0
yHAVeqsVpF7kr4YSxFyyROs/F05Yzfa9NA+wRDw7D64d6gUIEjFks5wMsYPKGCaR
oRglx1w05h67mY7AnJhSQDlBXPhtIpCkPq3Sgn/mMsKeGb8yMPei5pBCj1V4qZ1s
SN3FZu2ikc0x/k8QY5MsTvw0kn6JrIu0tl8qG0elvJiz7xrvgQqW+gv6kpitNrkq
gfcesr94bq7NtNcVQ1gTUa8Dd4FmXmSVgcdQ7BKPjr3TNrN6XGjq4+kyT5MZ0j8P
YLbvReqjcpKir/rtaYoWjl/cUBw1kJxp2m7hQBNtAOzCRMnrHv3AQYdhMzHxnflh
VhQEPpWOxFTCKRfOYhxo/L4j0Ub8Ae9AGeVA46AZuyKMh+JWJQ7Pz1+qFI7V8pN2
wbI/3fhs7RuN62BYd5MIsVYnldOhXe9wnpQdm1N9JaNAOlUK6A0Q8oFq/nu0HlWJ
vJXp7ehaD9SPYFL+3Rn0olPlYTCfuitCAkZo8gcQrAKSgw1Z//ehU1rBBpndfzEf
jM1R70yFNzR2EB1rsKp0IH/bxsvODe81Pc1JRzcc+CNd+GMGbd0Yf8nY/gTgBCtW
yEOgv5MjWp2p4dsZQF3QpVtQvXMb3OCq8bNwXGhIb/bFGo2eCgP3UgwZkNX0NV/D
diLzrcTL64oYk96bwurshM8bRxY4fds5bv53qtUAHMOyKRIB9mXFzZTnxxF3obdh
uC+lLocnxtMliOoxxQKsY7TgUiwa2CyPbd8qEWPncjjzKlIrQ66CDAj3h4W/UuSp
OHHylpitRilnQhIvawupM7VaIfmAyKeZyj5oWoL/ZNjltFZKIYfUahmddZ+Zw7ZT
5YVAw/BvxO7al/KbLUufomQZ98zecyOvTdUSnImeic+Nx2CGqoGBnQzPzWO8eQTB
qMZTP8XJzEZPB+iDDj0VJ0T1zaCl9+0KoaCXIH8igS00vYg9nLoMjSwwX+csLgS6
ST2sUXjGb8++mDCg1lv8QJNM42KnkjK0ufD+y0/ryk0GajmkDfMvhPdJz7YDyrGw
t1tipY4oy722l5A3eO7/M/l4E/k2pdIXR/COSq9hQwF2GNdciQLlgst0INoERiEj
zFgukI7xm3Zp7IVYvS9h0H8FDJypicIh7spot/ayNlJbCvdFyO8+p4FB0WLD0VK2
xXkCIyECQ8DxMFVln31RoZ+HxPE7p+HXtBvJCUW/W9YPMkSsVB+r5GItn5wyoxEz
uq1gr9TXRoVJ7trv7NHGMGqAnZqt97XbBaO4ug1vSB0X3bJ/MuZdTmFlrPA5RbgY
hTg8jBxG1H51xCu21LV1SM4Q0/4zq07SIXLBATnvt0Y5SjOChDxq6YU3evWV9TCD
qJj2saAqOuXNTwszksVBLPPh30MoCZLZug5mxC0DXuCctBF2yxmHEwVl/aQTM/OA
Nxz+PRHqIwMTA4z257V6wLXc5nLFXAP3klspe6Er9P586NUZrIpPYW4iEuB4aSR1
IpEn+raRIyFLNG9Fpd2mIN0ruspFbqZpH+ZTzSiTmla2QwjdYaSNSm/udVSZgpYa
1MsDk7Iw/vXr76EMq/Doi3VpbQQlHLDBmi3zRc8XShapCzThWd/2DM7/tz6ylD/Q
BhG/+7J3/p6/JAtea1hlRW82OvBOHuxBzr1ROBcou6AU26e9eKPMCw2kAmKmOYmt
3YLfLEOSHj2Wwaxp+FmWTOtcXheeQqYqhcSue4igY/Y26kxmHecqMTf2zTSxlnsO
zYLAhQ0yp/2NesiE/xBlUGmqtOsZhYS/1+3QLANqw1Eg3UoLgK9CofGARjUMTsRp
fYAzsxXhemNyv9Kta1GF1+OKqda0LF+YzYrBfcYqgg0=
`protect END_PROTECTED
