`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GAh0PIf2/pmxVIACTFGsJqW9Jp6ewLT3AzcNhFmL/TJ+nDEVSQLHcBPr7kTqSM4J
tJCb+3CCY4/73DSy6SwOm5GGuHaGmDLLQfp8gPSwlt3dZCddWjo9h93zW5T6lZpe
KZRMI3yElIgASGvuH3gv87GS14O+rBUCica+V8ObB7DirkrhQy1uI3uYgMXhyGlq
i0sDGqfsBqKQEzl9UmfT2lqWR2fXOYCFNmyHuKe7zjKxIDcWmdyFkrB0RU3KTc72
1G9Jig5pQTucPuSE07URD30Pzo2A3RDJFMv6e3J8INjVGNZcSFIUAri9ird1xpF8
Q1O9HBK8KUKkkabd8+m9hiFV6rsQIhq8t2ArpvLN9+2NFXihfIrE0QyOhvuIJRYD
NpGawtZyUflu1vYLdqbbOCOk0o1p535y8nyKnGFcI5g227CO+TFLVpmBY58eF2iM
kM/JAVJd0DWjmhpdTVVIgUyMcDNYVJXHyKQ7v6+swLilJldxLw/X/f7FdPbTrf9o
P1X9fxrL5onn9w90G1o+Y7g6+8/uiLCLw5o9avoCmM1viQs0M9ImOyRwrsxHnlc9
DqEpK+QPa1KzR1qGPYEJJyD8kapqv+XWvq5z09yR/3Mx1LPX1c7tMzT2L16Zwx87
uolOMmSLwYjvlGo5/TFAzg==
`protect END_PROTECTED
