`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HtPCn8hSZw8FiU4PdVKsPr/drIoIjzDcI1vwPfvGPvC+GBynBgpmElgh0Z97cL70
4ODjRCLdx+xrWQ488zqa72j1CkzTrfTocgeexQRTp+A/WS6IFBFR1Kx/hBSe85b9
/ncEkkyp7LS0EzJJEyke5yJlQTMF9xWgqFeW5b5KOvUnCfXAB7HewlhDogG2VjWK
PEoqaEDO0Y/gbgP17TFVr0yDaIdXuRc70rueBkbes26qz/TVzQR32sHis1/ANJOE
1ebTP0PxuWI2mqyPpYUehuacyam1AemSu9a6fKGObuOsfYjsXGyoY7G9npGk32Cf
VC0Y6+UBJoGNO/kJcy+unX8XizIxNLwjzL07cqKiot57emgGaITmbOhDrTa8RMqu
yhGsehdI4LMDMdHHHD09VzrqWIfk12oeHx2AV2jt/FcDNvl2yZB5rLZI5rWlLRQe
Jm+aSwC/wsUYQb+zW7kUwLaL9hmy33f7kyy4ypbO8YgcP892ehNd5BaJ/gEENS4N
MzpBYqskJeGZzs7ZDQBwHF3U+oLtmlwhjM/ykxDp2IUfTCf2GwXZIMOYY+SlJIsH
PA3IQ5cOwt31Vt69hGfgD/uD+c8neJjkv3jV/1OTVY8l1h56AuBbZlU2s12dOWuw
6NNP4TfqN89pfcPAqP2oEB+0tXRquoXIiixdxxFKfzoqE4mdXY7bL6weHua3vAdf
L2kQ/qHm5wkUMcr33jbMbYjaLPbI+AotQLbX+3wIM+hSHYZFjREJy4oP+aMPJvM7
Z+I5fxkQf/yDb6g30GFTZt0nh+zTMcavl2B9bknSRDeMn8ejnqUr8FMSkK/Hnfc9
m3yDO9cDfx8UmzDQUivd/sqm7hk70lVoujZLK4XLcqsw3JlVmeA+y10YL9Q1Bxct
EElpzvtPXtB6W99Yubx4nqkdWv4MZcHbAolkLkAHzvypikVupPPMbfA16kaN48pb
`protect END_PROTECTED
