`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fJ/65mqnz6yfzacu7bAe2E2+iNUS2MRCYT8fo3CFSwsV16cYQJf3fE8dSlZM4ryH
3Yjuhu7JDffwOtmwCqpY85ie9lRLCnMkL0aTeDyarCa29Bbnp5PbHGdozlRd2SvA
FsNdv5zl8eMfMyWmfdkYgk2KPnyidK7j6nts+2rM2M+yfoz4j9Em0rZ97YnyHa/X
kcB3p+d4kxfMMspxWNzy/mWh4civIstMq6SiFrBFj7tIQDFL7DlGuWeHrv1BXV2u
wSfl6NBUKc0XxwTD5kSLVBRHAgcBlvNHC7SRzUld2gwxTQ4dXoZOhCsJ94Css4SV
sOyf4DqNeIktg87EV9B8l85R+cmXt1mSIjifHNmoGC7IroG9woEe3HEXROjf9Dr3
KX3x7fzl4bmpD3Xg0HrmCMwD1i/N3DCiXGx7otYq3lvovpTWx2MSc7Xw4UqOApNM
5UpHCigpaMu0gaB6UWDJqo2jIhPSx9nTyeaVZePl8OGSc5DLdr8hWH3wjYnyQk6N
4GPqKMI0rFn2TaHCAm1g5Dc9Kbdt42dhhhum73GFD7WH9Gx4Ig+kvZm89LcnKUP6
pxhHEAXvxbsp5wG+ZDLa9w==
`protect END_PROTECTED
