`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGHMCiHMHwFk/J/8N3lSeFj5tlSMyAKZn7t6IweRybvrTdZgQ3ItWGPF5oy8r3wQ
OdGtb2LwL8OfYqwnD/8ACNkS0PHgY0ghzbwl4Sx13ASFLWv+Q5lpCIozU1VmDW11
FcaqFaei86g5SmomzmNRfTD6LYuW5/HjRFOf2t9Tbjn2+7Pu1JOOv49EKS/e4N/3
HOa+EUh8SRDpT2Z1xI3+SYSiKtkSol7YEzSDIdi8rTHAbdlXHgYjM+qBjrCR1HjH
R/fHdZSEwHgRPXpp6iNAd3VbFdgLMiGM9UBu9nZeZgIx4FjK9R70/TJY7jOY3Ar1
NtDgHRwp8k8nbcjYDVkKCDdRYqWIqE6wFkAC1qKkP6zErQvGi/JkjYb+Z6mTDVGV
YQeZ/lAjcQ/TYp1JhP/cyCNs9fTcL124iG9l+Ov5jjgmMd1lapgapI98RFcpnbiR
J98NCxFJp1/6YXMFzwyT0ggqBYJ6BKrYRmc68jWIYZDN/dzx2wcUKNwdn9FAlPwM
qJYjN2iQ6wEFkNJEeSVw3SslE2lqQBP0Rn1zcgBmjxLv/5dQhOq6xCv/w2RdCKi6
kC4Y9ibowtJ1eIj3q7Jonl6u7gG07Mahq873DfOfqBSVHXZm0yc24YXnZdUkg18u
Ixu21AvnduT3+cWAyTVCiGwuxhrHz6jPH7h8XNIdUf+yKXFAm/fZLkEcHQkC3C7L
U5oagWtx2EqgnUvJi+BRIwzHvcZ+Grk45KYax0Ct7NQ=
`protect END_PROTECTED
