`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wu2F+Q4GDZH5qGtKx1pfiv/9w14wuYVPSLdTxNarUTOa6K5tQ+2EQkP5VgPE2KXq
jbRL+es1aSAE5YHZlrK1A+UtPBk4ASNzsch91STwlEKFdgAwyrTItJVBqA8Kn6Zy
qyAX2cHc46LEa6ahYB/CcP/+NA1yTjtjRDFwjresLgz7fJoQSG7G1wEammuLxrWl
oNFKzF1gS0QFFAoYFQx9P98fxJPrM8tziNjOoRW366ysBCOBnqNGOnXdT31EFfbl
`protect END_PROTECTED
