`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0lVYXB3dO9pb0lsKuF8tyMccq4xj0eVf9wCAcCbQTOdMRfsGQLFljjvJplg1d82
Q2YOEBAaZ8nOB8McNuI1LTDS8J28VJGJvVV9M8xOFLboA1ROgb+S/DfInFCIX5y2
O4KR+vogzfwRuUZLRApCH2gClsdh5gilSjKti6K8kiJEf0i9rP6kNUiYeDVOVODo
W+RAxWtQYt9TzVgKYAMwJUA7eMgPc161tfrySZ7YJSU9I4oxIbsDh5WHazR9J2e7
3tv3vUjulUtDkSaZvsuSxW+ZgzML/MLSmX1y/cRCbmZlf9SI6/yr/rSbKtRlgh7P
x7SMLLwVDWGxOQmwu2T3UKwsIJC4h6g7LrpPOedkrscJnm+D0XUwVFUkNrXjU3df
wqfiBYgN1lWhdXDTTzCj9Q0x44+txh0GMLAbO43TntL28x3S3KCkDWlm+eDVEr0u
3KM5yHxuC6qkBif6mot9TfoIm5UZbRnHCdamRZ3IClFs1BpaJxYlWkEkD0GTuGlt
`protect END_PROTECTED
