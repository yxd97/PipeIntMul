`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XivHGkYZE07wQeT3/MjMdZseSZo4shOxvR9oU7+HSU7+X1UAWBerxW7OhgDGszpe
OK9D89ZymTeThH1T77u4+M3h/Kf/E0AWfLDMoU77i28IDqdx/lDM52i7Gf1IGHA3
4pr1ilDysHWN7Nhyng8hyqPJyNbsJ7ryr8W5zrsjDa9MtacKRvq11jhvYOWZ4UWn
CFI8BcTnfPqBABADeEFh6J6+Xtnt+Tid+M6wc9W3oeah/BhJWxOoENv5ccDtB4YD
/m5DPfO9O176EY8WEu7x+E5Z3N+kOSlOcaukobPaZsKfPC+amolhv1K1oBc5TBfG
HDSIpCQ31We9qoIgIi8V8VBMQt4AnppCi51LiXDmN+Jusg3VnERtWCAB6M3S6vqb
lMZiIbIS67KnXlA04THk1U0+5H2h6aLYBYAh3ZqveVr+79/uIKWhytCTDISEcFX5
TfkbvXn+ztWM6pQMy2cf4CpwAq0gFAPm18lb3/Aqmx2D1aRT4fNZ/qhjyVNhl0pw
`protect END_PROTECTED
