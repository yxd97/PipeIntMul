`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MBRi5/PDJNCf5KybYyB/ogky12JrOQz4jKaKMgn0Fq6pv69UVqZi9uZobU3zUmrf
msqo2vZRRkcJw0nwsq11nsiQzM1vhoJvY4B5x7G4J3WmcRsrnBhTginsVjNQumpL
kLSGaLT3REAwq3HPgXC+BQrFIeqt0RnhxrlSSKdtAWLl085TkaP3fvD0SdMZRh5s
bDgVi5hPBhvtUm7+ucp/nB4RYKWzF2qqpVxWIEOa1iMjGbj5RZ2hU06wj5N0zGes
FLSC21ZiI+wCgUDDUpdFW7yQnfErj420VDrlxXJwEV3URPbO1hwQl/6KfEIA+k7K
vpaJfud2CHWMX/xXo7egQxJ4hjNKUN4tsxEPFl8r3ocrmVx2BhaHqNmOzY+/bTOn
+QpuBBgg7lUylyP+5ldzupVtfqDKd5ug9o5a9fEHylo2bg36egLeqQPRhJXp8N4N
xf7ndzc6cj06B69SxCRJl6B2qgoXZ2bxusizeV1RhiI=
`protect END_PROTECTED
