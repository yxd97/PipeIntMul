`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xgl36Kcq7Aara23hl1bowqSk2cBAq/B2EROCqxPu/HyuO2vqIBMtubQ1bxrhu9PX
0siZoofMAL4SUuYwdqagi/43EyQmsXWoFkb+guyw9Xh+JyKUEtNoYhUnSN3qbpn9
SVdoXToyHSiy8YcurIU9HHLTU3Ix4VGq3mKLV3idGv8k2EsUgPQYUvJ+EcAV7/yn
MkhO/TQzZpWNtLPyYuVkR1C/qrP2k/4+U/JEcTE2bCqdLmyH8NzoChqQs+KxPR+y
EhKL+IiHfeTuswmNn0VQqC0f15mZ2E1hLQLfaJwPCUZAaUrBrINdXbQ6QUlPqs58
87XD3jaL1SJyN2ZOyH+cd/E+il4gETl9x9MCAylCZUAEYojcg+wAjAR7HgzXt0Fo
1yxkRbwAT+zJ1s+WN1PmlA4Sl0llaRjb3szMHGjJVcBOo+TXJTPIisEcPVn9FQnP
57kcbswWpNLT/irE7ZoDu3hekj3a9fd/UOdeG6LZjSjQt/XHMm1Lmi+0aCW2jFS7
R5WH1ewFFXr4tYJDEZx78gvRVmY4I0u4/NnrZMPvQx3umUnco3iUaRzttEiHbF5v
1f+BTSmUIv4u9EseQT6+ltP0+gs8HZtXGhH8JNlRj6MmWIM69wkuNImsar6qC/2g
H8G/GRZWZDAf9sUMQwu2pAnH+Xt5T2Cmqau2mE8Bm6eww432QGsKXs9Jd3M+/S06
XcMLp1Hooi8bQvAnQE+UfYm9MkX9sQTi9VcZA6phomdMokr2vkaFccvcoLHNtQvi
0f6mzziBzbrPfDupcR3P8YwDL2RsY67b0hGC7nVCVEyY5NWkI6/PvHq08ddcnaUX
IiOEfQb7+z/28xnIlMfvmsb09tCw4WZUismSwdu5fGU50GOjAWFjdMJ+KqLeU7Cj
V4ofWNx5tf3hSrJn4ix0gZqu2hTmzOdugY9StOH3mMi1NqSCT1nTvlFtJtIRpZDA
XtDQpFwBQwGYFiF0tWpLP/4P40eEuo7qiHsKb+bSZ7KvrifVfwz8vSHVorSjoYDu
WbH8xTDkXx6JzEB1ju4WhQ==
`protect END_PROTECTED
