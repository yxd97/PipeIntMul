`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oNTKwjzH8qlRmAtvTGrSlA+UmcntjQbW57aaeFlzuRHNfDFN31QjxSYtsHEJUJrg
hHVQalG29rMP99Bolq4bjyWzZKpChcXOMn6gULoU9xQOvEooeEd3FCSC+5EmMjyj
GoD915XaZNaBVNlMhAYzVmffjyUkP99MZLvNseveIA9nVqwGYi2ncpapoIi1KjXT
kJxU7J/6J+8LyFES4Xg2bb2WcPWCxVtdIllsBr6I6nwQAuFJUZUrYuTyL5ZVR5Zx
/72JspvbY04II19mF53K4aAscUeem2/HhiXfDszaxQIxuvt74jNLnyoUdDq44GEc
r9Z417Ii4RT6YLnFnGRTXp/pmc9sFyIfA3MlaEHG2OhZppAW6YIXcP7emfe1NnGv
HOxQp0aBNmwPbiVMh9ymAlcWUurGRYWglMypD66CU2vRQU9GzrfZHmI7bO44UmiM
CNd/sJMuxeCjtyF2HzbRtYebwMMeeXOzjt7AC8aJEAe/41xfzIo/mr34RKAb3+NL
P1eax3XiVgGJVcuDRHlX8ZyRI5FaVWecCaBEnbWwe9XDUXAAqRpouAxhr+csRKZE
Bj7PgZNhl6rf83WisszZa4966bMSUfmOW+17rMHic2vdC+Jlw2RNzLiDMtGvvnB7
nOI3vKDBgTvHspFRPo7cxMyXzFb3/3QrXmIn75xEJjb8SSlvUzTb2eC6lkeZatf/
73nZ2+IYdRGCOhsLUwoJipNfAwpVTIKg4vTFT7z+nzG17N+r/6ty/oriNfLv8wI8
/C0YFcWbvIBwwQyjo7XhcjHIuQ/JuNuV94EFlR4HN/ehLq5cNIbQXjRajpbCr3uF
LAoXWZrbbS+I7+BQk7IEr7GFP7SUb2qH0IfVk9+e76iBfqFXfnJwrkbBLvblcU4+
8432ICzMixVsE1hhQzI3WD22iuGb9R4iDvlI/oIuEpQf6OfBZB7JBWbxESSiCjRP
P6ug2cvEmcVLoYdUUQXmlnRXRLoOwdal7ImzYByvXtUIZL2c2AXBgFk/GDQhzbQS
IJeScnxDkwWSi9wp5m1I4bXd8XJAKWClU5wvNq+RMI2wRdydfT62VPdRhd+EikRK
8jyk1qPGnzluJX/clyOAXj+ZWUiUadvMnGJp+ilL414=
`protect END_PROTECTED
