`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucaGcTX13LOmWdD/DcJSjNer+uNaC5iH5MYwvkpOAOKDkI1auJtVosx7zXltsTob
sHkJaALyiJ/Rf08YLOMzNX44MdfGdCkBe7OFajsia3Zb27oas6La7Ev+EZ2Gufpx
bTVdoTewjfAB8JxdbmYFf7CXBfqwRbAcOUt4YVvIfPCmUMdF76v8WG22qqNTdLbg
xhs32rmwlVZzS49N9QBgmKmnmvY4c1+Fja1MaRpLfBQVCyAYBQ6sooQZXEPRpuxK
cMdi5j2CX94uuCHRXZ+tz925VMy+iVkoOKdxBAfvcWepS8EBUwNrv7OJ09PVmhfd
uMGuJPWTW+OXPk0jaCdZRNhuwygbCSX8enIAf+5XB/CQcKLjzp+6GJJpwZYdBSh9
2rqfcJ0nzxkOfdM8Qq60XA==
`protect END_PROTECTED
