`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DX+ZVOmL7bhlD+eJ0NUSrt5sSQxVs06YrycNp/v+TK+kUxN2y06eNcIFNI6eQ/O
aG7fc8TEu+yYISAxO/uVpOZV5fv86uwrGdyRomne/BAf7ENI5XOToCp5PGZVNDa3
K7LUMShV2fv6py4ibXiR8I10rBTiFjgpSGvHlJCK/hwNsKiNT/+KTJ/CZyhZ2W4b
7q85xcLw/GAGFrLBoEwgENXdPmbgmMr39a2ns3sQk0Zj8silQm338ZmknHxknWL6
Jk2R15YZ9+J9Q6CNeMN50MqzTm2IKJ/p7ebQVFLyQdP3EGNZyNz9CNqN14YXR5GI
ZuDym7StBSddHxGNFhX5HNUt5F/QZOBbqEf8oXe2eX4/RD3aPREMRv06nhl787hg
MXUt3lveK/zyXRXvsj0hpk1nbAkZXSzV3G52hqixqO9hAEV+dGIAhoOQpH4sQh3z
SWKEGOPsqHn1roDvLZVjjd3bHV35id4pOn7yeMcpbX9ZdVJ7lojYb1Z1Ahz5z/88
QwmJxOBAI7hNfY/AEsncxdYwJ4wOZbpYXtKYuNXGJ5Nog8FRKPkgG2BuId+879xb
v3Di0+uFaos7n9xC1GtAC2ncb1Q6jAIrCP/yRNP4JoGf+QAXYqLt2GrIBWf0wvv7
0gb1XLP24TLSKlEyOlydN9C9IV5G7qO9UzUlywevvtu6Myo1S36zY8S5vgc0E4go
/mlKu++DG/z++XJX2g6/+i0lqHLCMaXP8eVNHntVkE/h9dgAn0x3Jvqex8OK5Vrb
dKMyqgfJTuhAz95untvOMbStm8DiZDuplxFoFYshiHMXDW5JpDiHlB9UZwHm6huZ
TiI6JkqrtaHP9Ho0dCuMLKOcTOv+XmGQpC75/acfheaGSIsVkea69ItpB0JH82yG
kn9yKBoCiENCH+z5T3rLNZxEBV5n3vEJ6pfoJ9uvF0GQaJ7wIP7yC0V9bwa/iRvl
XI6IUBDULigPV3crsGUQyUffOotSVvB8pBuQnZ3MwtbrA0fuATeSPPQJzUHdDGHz
BV6JF4LHC/IUCx0p/fbopm0Sr0ToCOC3IzS/psqgtcp65JdRaKw0cB6EJUQJY1/s
2oRnKmiIg0odIBHvj/B2TqzwlAbTjnJYIFgkK88wRp52B+d13gcbJTsHiZoVQ9B+
OPl3MTRQuzoW4+Ku6qZvLHHhi2sl05EUR5zy5xyJ0Vgd7KaXIUEcHBrIb0TDFYXf
bCm00YU0IsoDVxrLvlei6U85OS5SENh8B/AkxseA8HCkiBjMCYZrhbndsToFZgmW
iLm7t74LcWA2Bd2cw+lw+vj5WQ+/gIix16YtN4+NYqMNrcvKIc4qiycfkcCYD5ff
CW9Fg1gh1p1s2V1lj+hT3dvPmWLn17iEWt7a1mOnoxWlsprfPgEyvaPPUgojdEmD
+qyqOo0eYDEx2Q7hZiVhluQYbKtVi4zwx6Wet/iLrSQ8yBYvDDFxGacoDkxNimTV
9DvZ4/np1qfs78DOsFs5k6GcSelytpCzPw5XBOjl0hF00YMZS8N9f4kbXaW0N4YB
c5tzhN9aiIUbVc+naGsVQRLrI6ka5CF8/VoOXeCF0odNd19EBLLwpo9ZPI6y2P4h
NPfQks4n0XObhuZJi9G/G1ZzYCsMepdFpBMZ5qi6BBuqh9q0QunhKvV4PxxHScxt
Z+1YBaIgQ1ruEAezBw5z9fXYnxGJT1HfE7i8Ib12PRMenjC1/aQBtOq8Y3wr+vSc
C2veelzgAgK81qHFPN2TSpKaAWFkPrJ6qt8L+W1vMCo4teidfycpbE1YB5OKzUdo
lwZ2SNUOCM/oobDAnzS1NoMy/r1vlk4pIkZlG1zLJYobSzEeIPu0rO9Q+GGNbHZt
VenND0MO5QjbkQsPRApOprT4TxmFhWI7dQDFQU9IB6jX26iB5xJhMU5drYFxguBY
2jlYYNcuKLkU2ZUHViqdEo9rtrmjE+37ZGoouwQMu3RgQuPzJKQ0QGFIx8/OyPXa
vs+xTbii8ERhC3AtTKfHA0yJd6GOJGaTST1jK3VqHeHP3vJ36I7LPGwB+bRSVsii
ihDMmfTc+CT+qX60/PDDjXzIjdzY/8LVg+12NHzX861zxWmGrkqhoBt5iYvptuQn
y/o0VeWfEy7yFC+Hizi0a11fi2gEAuHfOooPgn/2wtrjXatcHrz5eYI0v4KiM3xp
cE8a7qO4lAd4sKugdhCfulrB3smjTZcNvagE2CJM/fd5n93SWEF63lUXIaiZbU5l
HZPNfTeNj3MPGgEPr70rFbGLtXh2hb3Rti8rThIKaT/nRquvOG+edbQk8/PUzzG8
sT3JFHxdxMuIfBBJWC2ePCOjt7aJcTLRt/nMQkvrbU+f3oZVabgGos+UIuaykpYf
Vf5lbVjKfcSgY6DoHKprQkcUguuFiPQZug/0DYrQuB/hGPcQjavTISFXHiNX5qlB
nOAohVJnKWY++T9jSdQdK6HmqPPYpikMMChGcKUIjNxLCJCJoZcNNDlriIG7jBs6
yYxozIUVzGX30NBhr/aoVIcBvgLO042EHHb2M7/lXAGuMnx9vbVktreG4aegUMvq
kRaq0TWf+oH8WzPEU/TVcf3w39eqUY53MA0cDv2LJ6D2jinVUqXMAMcvm3WaqYyN
QsYjaTcFYBKYIitLJsltAMiCcntuCQDACS8t7i1QgPXYgoB0bJlrDriMmojKfbDz
yP2HMsxyCtxosf2RZwoeuZ1PzjqQ/2B/vXm40/PFevn3eip6UMtx9w2bdceH3pMV
NW9NgcbjvGnMzakMMqf+Ld60KSWS5CuLXMhCWEP24MrCEjFVPW37ybn4FD3KXtv7
c7vhtq2MmDJFse1Z8Bv7arSBlt51UpAe2VAxM7G72xRLWQMLDD8VrozM+HoS61TI
qnCf1pBOW+1BzsDxUOTffeM4xKpCcrUGjxCnlze/rhIHfhg30TaXYZLbLl8UIaZW
dwZRNPmbOHSsd3SMLfMXEYgAK5uAxuGX9otq913XLD5kRsnhje59FXwuid4v3MhJ
4P7Wr8mccLE//AFwdr9XYb7H/GtnWEKSVPjHSMyixN+1zYidNN6J0+EXRKMjC1W9
Rv/KvemZnSpBTPDt+hLBKwqPYPtTzcSVxSViLCAUpxPKcALer6BSgBubmrF7rm0w
pQE28XmC8GhUbDy1V+1fSy7yc0YNNAOnRcvrUnmYoLJwkfPnIMDzTM2PaCoRLlln
`protect END_PROTECTED
