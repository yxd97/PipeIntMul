`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oIfoLjTVt57bzePEnMXDd9CSzc/TH50jPr0qGQ6NdWr8nhT1xP83WDJOjc0IGFRr
E2tlY+flXn8XvADJcaDqAxay3MbpUwN2ZCmOZjKj2vrCtrOwHAcO42rMPmHblEDz
S5vo5NITLQktfa87cps+INep7jZlxIwtDJmShovK/M0pL0ltP/RowVG1tMoOkwON
LWcDaOSVKGiNb4xmNm2ZHMLU6rhFm6zBU5N/DOHoCGFVdzvVw5wE/qQubmWdq0rU
oWxnPgdONlhf0QAAmEyLUuYG7X80EFganiBWwtFONe4DD2coG/aED9E8Ldz7immp
5t6cIrh6Ft4EfoS1PRreW04RYL+8PG6ORF1ceqJarFwHJJaDIRzxmWq54wUIU0A3
pQYIobla+6yltkmZrJGx2O54Vqq+bt0ChS1Di3E/es7xRL340wkayubOTCm5ssFD
/UkkqGRcvS73lNyQ2bnJzZPZ2Umq6mmXf0oucvVaKAGvvSU25RN9rQvxM+pjzsaK
DeZo8i2urpP8mlSaWScTzRI4iMC3UN7jzMhP/4o23aSzQsMZE4+ffBihyJkdtfUG
vh9IEiXDWzb0omkFoiB9k05WpBu0yM3tb4p8gUmG3vZ06MVV09mFyXkF+gFspbHG
gQVVEUUopficpTV8xYTA2xEFbAtSVQpoTRWOABz9nXia/OX4/aqkOCalI+5knwSH
XrsHszc9qNcKtiWVIVL8UCnKbGO0gNjNMUWdTwJZTFE/8TBQ85iAZq4z0nVqPr3x
sxUtjEfCLm4yuy7rxs7RtspOzfKtJkjBS3jfL59aPuwZhpkIQmnE1j2jbLhBWayt
Gp5Id0lMScftUpeZzCHwuMdhkg6CLE3atFbldbWfg6Yi+wD0en9FvqkplMT7rmL9
b6PYIF9a51CqI3egR8HU0HqK9Hk0NIuWMDY2Ucclusv//QqCcakFJ1szqQTe0mmK
rkTU/BfQKTd+iIT/Cf0dUS8hIXH19b2UPKp+iS0AUxziSoJ61dzVNCC71EcMYIvf
Na8VyqEwnoRvW9Fim2tt3UtGFK38hYHSjV85y5N5YY37ArAXTlxFEMRiOndWj8U9
7Y6aJzfwbcG0Osg388si90AOMlB/IfKM8y08z7990vCpY6cbGc89NTxxlDIkwZR8
CBaZWlSCLLs9X4VhYLY6ZFASYHN3TYmaAQtDqiHmgXPBXFwIik8+/wXOxbqBuCZG
h0HrMl4OZLp8OA+sk/amWbM46JiVHqamhb2pbQ07itFzaUB9pwhgxC0Z1m8GyAW4
GZV13xmazaCBaqAdl+h9dTNiBdl1t5FwUSgU4IRupwMu0zbookz7PWvCCcOLq5Dh
4cwiN++D5DuTBuU7FgaRsFTnBXkeMs1uj8KfTmfgclUquZ+WyosCFs8PeWMoOseU
e07xwrG72/ET8ZXCbDgCJP35LGgY5HejgBDVkENFrEW6AflwsXuJp0R5D7Kunu/s
wJk/ktAvuUwrwgLSEUxWOFf0TpXmDCWA+6jAgYDz8K6qPnzdp50pfaecpfK5tt1y
cwO+Kb7G2GI0uVzajWeZU60Kwc9oDOZxmsEyvZOPBdAHKJBxs7kBRH4Wpo+Ed9Sv
nUQnT7tMmcLiMGZiLM2kJvMW6zlZHH/RTCKyUFq1VvZxrqWWpLUreI8sR/2rlTNd
JkENlFB4y3K5AMXK+dew3QB5X6SXGpVmD0NiecXr+pCx1fwsdZv/2kyHZwiGCHQ8
x4GqC67/pWnXMyfVepykZnv1A9FY8aGE2zoJCGAs3r0zSBxJ9ziaTxuRzIueAdm7
M6QeiTBtqQov/mAaJm5UL4Fqa92CVo6A0fEPH4ziw4KTT+htaxM3o+yxAZWg55Z7
UrDv7i+uxfxj/aUKV9tmDT1ddzYkeWQ5XNtQoKGo3BDT6c1VRJ6KMk4av7NLWHVJ
didbCNoDTi13iznhrNWAf8kcgzd1Qhf1U/zouBekwV3NxEDRfNOEeEwalVYQYxZq
k1CXcVxcm8UIWmz9+VO6dtaGbjmR0MrnV0F1NVWlxInDiR0SCBMkaopiZM3+OX34
d2f4U7W5c1nJXwyNjVRZNSkxSVckl8W9PthGEp3yCX6uDc6Tv2Ie0/MjTDBHOFz/
z7EaQ37W1qIbmv76kWW5jk2q3+HL+auznYrklZdhlyCBurpAd47N5aL2mG22yDvg
/t5KW0sY0pflVySgVrRpMLOlt+Dsfa5dNRm/2PyNOttvCIcL4MeRmdAX854l0cMB
C2Rt41s2wmqPfJXRyqQEGN8FwFLP6H2XejU+QAkkdWy3dVO++es8RzNgKYixJ8pY
aqcMgxDftX6JkYCxNM4EO0DZuvBzwizP8LoNQVdUJ7DeHC5kXt6coI6qNDDPDeek
T2mio5cvNkZI3qRSBUJcJgxJeGD1E0Ej1xA2B0mbs2A1zo9iJx801MrFlfKM+K7E
E2BfupO454X3uxk5uiZ8Lu9wfkBsMyRknqhCf4NewKw/K/0zL+f99/AX+1iLxAk/
+cc4fB3WzFHrzlydKDf7EHG5UftJ3tO6IdjRHqDMg2IFhupRCijhhVbVffYfntGh
u94SLcTqvdZrQl+EcMQasRPXzXGTnkDtyS2NNZ3czAlZmAe2JSCxbGXX7p8sHueo
kf/KSdF5pAw4kW5VA3mo3MS6AAHw57C6PyxF/BDx5TP/7S4H9v21qLT0Mvjr8tpE
F+uJUJTuCEgGIFAxqzn079xoBpkmyd2Kv6oRKVUYcEl2R0lEt38G10aw33YF01aj
2GW6JVyN8qU443Pqe/qEjRLR2u6dsB8UIhswt6Wc0BNG7rQlYIJwefr52YMzJ0Ey
6kmodnghX0SAnWr4QWKAu+GZu2aBY/mlgqD0quiTXb1p583X37PUso6KZDjq8uMT
0YQZrEIIj8zAUddXAU0fcgK+kEmeYHKWj5WdeIRaWcgW0zuAjQf7r1cu4HqLM5pz
2fifp6MCtTQerhY3zcbXO7I5QMRlPldxfKkbs5CWMk5t34TzfQoB+bYi4+TYb7+M
ovKUrLydEn8fTRf3xeyQNiI4AFmubiygmJwU6h2557JjTdZlInGFbMJ7YgGQHaK4
4VIV0WiOA0Gg5FPYBsJkg/7iv35jfh8FuRMgj8M6J4Ncvdht3nxFdz13jyVq7FA+
BX6FaHQ13cE4c266NMI1TJe6qkr7ZZ5pF0j/KmMtT6UYCewhp2VIUr12nQcAmiig
djnmZSsp91CLNI8IY2BTeKt7K+MLkiBGEVhFSt2ewjiVw7KJ2fRv1EweDXt/B8P5
YeUK8trLi+YY09mFOyzcz14j135P7cMzFucANLL5yrTmjISLdChG/oDJ8AFJtKpD
EHpdjdsJn7/XmtxR9sgp6knl8U6b7vV6SAn1rhSz6joabAxIt+mmXS247IIzw1Nx
5UoSm93jHpayyqOX8DRZxOQu1usnLYQmuWsgT9Fnqh7OrVS5v28wZguTC0cbpQZN
isdtqit5QsntCyHZii5zARREZimmWCF50/Keg2HgFFAwfWwbY9DZ5M3nTKV8QqGE
pZ50y6xo9FTgPXcXB5N6pS5SKj/p3lzqGxP0eaRV5pw/1H9kb7OPw5yhKwDkvgUh
Jy9lEpdm1NMVDVZLS3FRRf9N7qu3rXcm+WowbpF3fOOUfNVX4tvlAanB8yId5KjJ
JOIXQDE9vkpl3s4vaqqGwzC5cm1gTKsZfCH1Pw9M9aQowAKsT4hjvSfxQBdFrv5c
tzljtnS1E5cWCwj/Oe0fOcPR5FgiOlfPQbaUycfEJeDbXi4dNg0us3iO0GFZZwzP
iYzBOJM2enzm0+ggMMEG7teAIkf5Jn3JzHhgQG6/xbS0QI1bcCQXZTjVCa3bwddu
uDrTrm6qcvfCIGFA3PzLo8LkXZ8b2HDbMscaqfr17nhnTSepHNyPK4ryQkRddxCY
wkM6cM8FnyIyJuTawt9PfJHtPiFfhVwUtXnauB2pc1kuAWfboeKHufhX4O3YkBR4
yzS3SuRFsl7whP4kBEyOok2LHvxLSSMRQuS0HNG4UhU2yJ0zDmlwXs3mNkAbX8NL
Wy284JN6xjVElPmre5X6cISxQJ9qOv5gayhEN9geO2X3eV2o/G3CryDF3HFG9MfP
C2OOxrLKAInQ5/YQpinGzAA0EUazZn8++UIS/lHTvTBuWlQoNosKxrbe5YE7DaVF
Qj7BNlF+sDLI1x4furYwQ2cHhac3BrXdAtMAA6Ao5mb+W907s8jC0lBBWRZ6VGVs
K+KOyDn3qSH+DdmaUua0ZbTt/lQ6ZSaJmB9KZfh6qn32/f1KY0DIPIrwtQ9WV0CR
AJYzzpV9mZy8YzUSI8PZI654JzPWdtp9Zx81pM4+3rLjMpgmkABRp6dh4P2YvOzO
/Y9qauwzJI8fe8IRAqlm1YNAyZVga6zi5PMoukehauyGcVVGcfPD2KnJZSFu0x+v
SC/dLvvD8rstx66N7Ai6XNjLMeRqVeVOYvtKKyBn6kIWR1R+AkB+G9P2wdDIrHIp
eqFTTCysjNc9t8TbiBYh5NGHMZ68GIs+W/4++Hdw1Fx+P320CrbOud7J9vejQsV1
V4MruJG3tuKhrjwGmwGbQnd53VydoWtZQHeeelaSm8j9wUUalaM2LPCFHbQ3ekl5
0eTtrMgsi1AT1za+fDLDL+knXEnimomAGI/XWg8BkUaw64QAs7eOzFABDVkJEvCH
FS/yzr3G48YhTzQIiUDggqIxhuYPLRYkQBt16l3gmyUp5ua2fZ4/pYvl4/wL452i
u2rWgphZuuna1d3HK2tGNgU0V704HbYVS9iW9HT5d8/M2YTdt/1LR+Vcf8xyZU+2
Ck09Gmcy2LQwIhf62ewyHGfsWpfsBFw4LVncjQ3LOBCcBFecCTeUR0xoS08lh9ht
2ix3O66bOSUlJgWKxc+uI+RwZ1C3MKtcQxg5RhZ1lGBuTLKifjJLm43QXQxEabmy
CugC1TVCM038kjSXahR7O4gUsnK4W9+PJ7ormkoJiLQMLSwRPXSU7OUpdyG5Xj6r
s/QrdeAb2L2xHiQWMbckC08M3xl4/XiPCLj2dd3bjOoK16EWivh6rXEmNQfHPOJW
77hg2tSW3MoN3QMEUJGsvUBjTMpoTxGvIEoc1OuVZYxAuIO4nAv7W0q83nJBWW1H
b7wW45BjxtLI4OzcZ18WVeGs2jqNp3uKrV1OAxwCNZuI7OrFOm8eb0i3MrhoT1D9
+A0eXTHCHAsG+4XCTI4dvRupYZ96fs88rCZ2SY2/9zd59Kf7mGC6fkwMaQE7Qx4y
kZVaTpJNkElFlIRopRHbGERT0gsayhIsyDBr5Se+8v7Lek5YtJp1Ewzve+ZvMqWQ
1TXKjyJGNfsoJiSSZEJ186pu0YgDA0q/JQncTr/Wva/L8bKJwo3KJiMiaYWX+06c
xRlkQIT1ribkX6Dikp3cuV1nmThktKUd1bpjrnr2sTeTk+Nf3l/WbHK0VUn+T0QS
JEGGlepuFlW2PQXH6vCWtBzeF6D3nwG/BdRoXdpXA5eKVE/i1CgfzcWqzpLIJCTL
gH2XlI61pCVgblyoKrQvwuzw5xU4VUj0zFzEOSLMtTVPro7I3c1Q/2jywlC+112X
defyK01q7NYdZrnunbjNl652Xo6mR6k23IgdydzNJ0ULsb6RLYlzPdnXL4cfiRlB
+x4Np2RotOw+0m9U6FOZ80qDSaVRQX8glYcUDMjwvUex/YFHCZhmEa9Ke4YuKV7L
4qfP01o+gW2esjZdBz142o2t5gEDQHskxRkiHfnc3KkxFctBbexcHGupy7kos6lX
s+z5W7k59H1GfQOq4VbynR/znpEdBbyXNLyheeqYdUjZWopr1AI/TGMYdA6BHuA/
BV6i1JyNrHKkqYG2ngOXuaGf+B2Ek25zKJVNxlAJXoNmZXwtlLjZ8J1syJhAVAkg
YqwR2s2IjOasSPMsPel8TDtSFz9BecvEQjfJJfYu0Z4+oopD/sR22hHYJs+iimgK
rUNSI4HJ7kDScgFr0xz+CFC21meqn8FJ1R4mj+3a+4Ee28QEsd5IYbVo9O6uT6Vg
m+jEUwCluQFBd4SD4j8mV7z0mIOXixu38AQ3073rCcEfeDUfKv/F6PqQ99imcHNK
yaV13NjsoFgJQlARL+eq6znE/+9KMe7zk4mJlRWM62ihjMGW3QoGwd3ctoUieyyu
tZpWPwfusDxYOPqeMSOqNM4gYjrVisVdn5eCAdi6so5Zq0040Ny1aGlaxV94eB2L
HZrqBd4JCEfnP/FWNpDZGnzvVmBWvm8bsTRfcoZiFAu8CDSPaGxyq+NLGqDSGsvb
7Z5Bcz/LUWO8wIHw35NQXkCXih84XU3/I605BSr/OprryEuGNC8xRAbjhxVYNOMw
mA5btPF4/afUYQH2VKNDFDQ3q0ZSWtRITtf2JMkJB8d5A9pSeD4el3oONnwxp5py
G8z8e8d6ysW5MucyieX4Qp7jBk5yKtVMNR8H4bhfrrCM4c/28HWQUhrUJsQukGVI
0BVIvEyZ0vB3B53El6iJIxVaJqypaRygspqJ+aveA/kby0qZo1WEgJDCSVlEaki1
b9rbI9g4oYR/WRWZqW//wBnkMyEn2Msdm+LNeej5yqfuWKNeIBHopAKjlt4JwuA5
p8sD+y4dfesKcn7blNNkN66JGok62WX21IbJhLeC6NCn2i6jFV7mKnIthqucWDwr
Hj/mow75R7wmW9FeCUyniR8fC2TzSLERIjLnrrpJ2ri7uHda07oh715+vhfL6b50
w6PiUcdLTYAhiPMzFdZVd7BJ0zsZD7nUXc3JND8pt0nAW3iGSJ0WvW5wAkXg5OjW
EcIezRh3Pi7m5/b1HyhLsGIpepigUjwdsxBehUeBXFDNcmOh7gAU10TcEpvr6PdU
azbLMjciShgO91AphTw9Llw5fWGy1CWTBOFLf1kXPCSrWENj+F+hlpp+DeVxyFzf
d/frLt4EDPomNbHqbUG24BTIiFol8WQS01cf/A49koQqIfEhXGvb/vjDUJYkHwsh
T6afDM0UyZ6UsbtNDCGHaB5n0vSMf1NcPZTAuHx1qScgT3CAnrzEv6qOHCsqC/mu
UIbsXfIIQOXvfmEELUveJSt/j+FYj/XIQ8+oVPGSHf2mPh+o00gpYqs+nj4HE+w0
Ql7xvNj2tpa03WgTPv8Aa8xVB34FYDsNoczWXEFjPkjXPKuQmA7qxDGwELcUyXET
GHGQlvPCkFGqaDs/VNQl+pP38LiWnoo5nkVXyhT59BfS5EOcRnl1X/oFd5Gqo358
u7gy+my7e3cbroXfpxuWfyqu/dIAAVmW15Awh4dYBQ00lidF9/k0BG0Q/Ccvr3Pr
FFiXwjmGUw59dc7ZLT/qb5+7LO7cH3Nwam68Idk/LBHDOZtdeS1ohIaTCQPrG5It
VCrOq1/bEuJPrHeEjF6M0BqMVSJkM4oAuNYkIZNjkBHCRa20Rz48c8EOVfUWbzmA
45qbxK7cYkf0JcRMs6HYmaPKcR/ESiQ7cdQq5qGfxJljDN4BwmF4kdFwjs9btxzs
yVx7MKA9U95dDmQeNBJ+U3oCrGZiYX4av/KL3WRg8uNTIrI25oEUGeS59XEpEe8B
WQRkUbIY22nFXugzJmxqOwQ2vlj1u+3TtHSos4iszSuvOy+qsU6VM+vsZFoKzK1t
xDHejSrf7ApcaouYNAm0eRXvGi2j7/sjC7Vbd0WyShHi3JpQp3eUJkFQ5tNRqsGX
fWa347/k4Z61TbNr2Rp25wKJzoux7u4bDIQxMUh/TUg40/ThymNBWub1pBnGuD20
X9tCaOEbpjojZ4WVHediAOX0fcZHxTgGQFwsdLQZt+LdXIpXH/iiKAeFSOlC8cTl
0sehy9xsLrzvc9L9qGlJh9lZdNzRse+R6jBI92Gh6oiS34ieiqggmwvlBJuUyn2p
5oaJTNriXfl57q6ECfOlsPFod3liaUEFd4zBMhsZzn+1hdwZ3ZfqOWuQvjuEAIjP
YtAirYbyfy876jEZcHBFHjwtDaEtXaasu7EsLfyu0b+fpbYcNVQ+9ZB5fx3JRb44
e6ws8Ocstye//2p294aXwRos174YFhrP2Vkfue6UFyiGXANguJTzslJOeKllIeWI
kbVZJM6p2u86WrBsYTr/Uuy7cCROfjauybfNMRx3YXmnpWmjmpI5F1N+YBj9zEAf
0JYRZcVFYXcqK5hZ4k927Z97BOzQGow2j/6cdGYY8KThTvwW3QB0LlmyOv19hP+x
fOw2EZmq5Xb6TBpcXUnzroCkY7N+F7FEONi4IRSlkTvrdhlCuMe0QJsn51kcnoz2
MeiXeOC5ID76t8Np1Zd7fOYTB6SoCprfAxqkl5jF26eLB3udlYP3VVUlMDU1lhlA
B6QTPl/RdbiMk6Ky1+iaH115g0jqFSQ0DVfo3Fkq5nnwnUVz2FfcIfH1Agl+afVs
ZCiECNGJafljL5pcp62u2Hv1nc+vTwEvLzM1Y6FQqhHkKBLxRwp9j5DmfBxtYTwa
Tw2rkGSbiVY8tsZYjU+dpWdE1Ok0jJmjekZaTZZRzw3JOQY24ags5LLTlWiAQDf/
eGtsHlvt3U9ELLsFIDMHmdi5vG4YPCDZcQu/OPphcMlAsABgcJWx70CJyJIXxMTq
Ke8hhokBExFANIdNGDOOg4SssWtYgmtZo+ieJD9mh7AP4kfnX0i4fxs8QFacTfoz
LIF5oci37ricXT+xG/kMl3m91+3lbi7xZZngrVO4fuuApEfNHk5UGULaCH0/9lV6
N6W7YgnquVzHuvMy24gNURuqTL4VvxYmnG59cCjPL9UNkOtvWRVzUqa6x2OaiR7b
1uG4uzBROcNXLT30nC0fmK+Me92iqMABFFK34eMiGGCtCx/v7nKasmgepIlbC5/R
g8Yo6xZNSjsfqMfpzmyhPTPRna4YJvbBvUwdL3JurUdWi9MM5GkNnTgG7vVd8PDL
Dxgwm8YnItzJ5Os2C9yLBUW/upzAXwZw1XbkWbZyddv1j8/pDuDcLf+J4bHBsON+
Yk3flerq47kHJGqamtSbopTqypZeUuVzN6POUD3lpP/vcg8SoZoXNbJZfwOcHtV3
O5Lig5kGl8IhT2LhoONeA9zL9h/sfmD1p0tlTbIsHwYgJ7jmzX+z1M0HQFWluq2Z
KdmxhzWJUULEtJUB9qL5eFmSL15f1RUa4YTKYioSfk3WJbwAmXLnK3LN/iym5cnK
zpDv4VmJYOICEstzCQD0T5vsmwytKE5LYTdvEoJqI+ql4fMq803yTh30jLoJyFwH
KPkX3eLJfn08kRgxOqEuA5kl9VZ5u+YPlO6mW0Jy5KDBmehzv6uGx9uBP5rvvjts
YdzhZSOAkGosISFc0H9oQdmNkTQNA6mdJQVjiO19CrATlyiSvEsemK4q+LBVI3xd
/Skn7pu4atQVHtJnRiHEIyLR1kE63rsu1hh3RMR6te1eQ0WmKNqf7EZi4uNinFAs
fM0M0z8FotvFq6hEsIiUil2R+9DHcZvmkLZqYMs7FfB8Y2nFbOdN/YMEeA/atdLF
5j1DOwQAMIIzla9QieCVG3TRUytWBl+MImX8zMUZ0++MPDDkVuFU672DtO3dCfVm
PKZ0L33GNKdwJ4NadKov8qnQYUr6SFFclZWBULwgOrZAhJEqVNgLuGvpu8ktGFDN
NuO8aHiC/K95uf6A4hNK95BN2rwX36bVAfjvSmZD66OrRwSWe2s4vQCR+X8KETN3
y8lr7OatBHTMKgt89bmsPI5nmBX39YFyTSHa2IUiFQGLZZ7j1ux79uhqKeMc1LM1
0p44YeXiFTvvq/FsmV0g04WDv4nxtYHoZXSkADhTPsjcAXYuchMzTpCPPRUhF5Wb
25oFsKtP+DSsioB1wI6zRRttTLJNcxd6qCzpJN4mUu59JvYw2Qmzl3ZsJaBdinyL
HCTwe7u6m9gbqcOk1ye06wezGffyPxUjwAAhNSAHDWq4zpdl1RShXAfGMU2OzLCS
XIjiKu2pEXbpwu68g1Y1Dw5QqZVmXV5z/OjnmZnnU8PZeNbJXYn8Q34QuwuQp1ZC
3qidljHm45L6SjbaIqieotguSEpmZPodHQp63IjmBalgxOE0fiiLCty5IcpPpgP7
L98gP1kgVpLdUzv4RxryakLgSD9JqUUfr5Il2v+12NfxoRa3XiJfTNOChVDVqvsf
oN55EFo5CjrO8S/Xh7+8kUoNNDpfozfAcYBQZbMbmqtOYGUFrznYj3DcmMS6atpj
xg9OeeA81jHbpIr9t6o8kw4Z/6yUStp+bIgt8r1q216gSFhFIeAZ5vv/fN6V6wfi
qm0ikq8JBQtJpU2ul8KKCso/KMdG64eOnqgsVayU4JfY7qQlIt5rUpPGts5oJzd+
G/ciuoaiLOCNrQ05Vx617TE/nIE6/1J348jZXX0YCXbEKGwIDHbjWWx+jtxAm7S+
xGsFtOFgx+7DoxZJ7w+moDo7RnpQPwDC/CMIHa7QDUruWJek3k+/P32fdsGI9lJa
43PGB+bL/RMs8DyjjDmRvP9I2U3QtsJq2+X3dTbMSQN5MLxwTzkLGgEfVSxonoIv
pgIGczgX9x+OMty3zOC4YNiIJrR9ZaOL0YjiCeWYeJzeQLIdrO5PWW4xi68s/AXF
MhaX9artpwSawaM6r47VbkUxCwGaW6wwdS3htGfoYkbWzrCkU1+uJ0/o6XuW5H9G
JVbErx5867swIlXhEo10Cjfwx2IB+rfKkMD5k/fOrjdw9bYjqHkZnSkam1lvSNc9
Vf3JDEoTui1ktAq3ysPMtSbzxh5ouSEG4sJ37eQQjzyqA/uM6X+hhGvylOkVWu94
gdANQqxk/5avArWFyIp1/v9/IYe4tj07M06n8orB1yHca3y556hddtngnh9XiOem
owCMJt4giz8ooXJAS7YpnzV5xu/fi26k8L5UrolNPTW428gT4fhQ5PB4UUmNgS62
bnlvGP75GRYNvFwGfvbsmurVxVo6ooJ3s8VzeQZVfFWUxYkEi/AebFSwKMJcKQEL
FnDDrPmwogOm818NJuTc7EDES7uu9dQgJU1WwvglWXXcJ+jrDfwfPLkKUTHKmQW9
8wnyr2xRb1wwjmnc4t9IONbhkqdCINHDl76w/18jA2T/U9yPeWWEvWXP7T1XT8ix
4Fr3K6STRUurZd0j4YIR7cC3MRcGx4rfxoM97RjJ34oplcizJ81EGLi0lKoskN15
kqCnOOKbfBPb+BD94qjkMAF2/2xv51bn7lrfCqqwiFXSGRDuc1LFB+VZZUv86isq
BeVEZFo7nsaKOyazFtfrP0wjGBhaELaUX2cjFWTprju5LKRteRl5zpEdiYF7/R1Y
W460mcpf+94MQNgeXHVaDiKbdSTQgouxSxerwO7KOacMnCdmpneLk2h2BDRG6DZH
BEC1VtJzEOu5ulRdSej2IE8mywUa4280FDneJJFjnXEae0+C1ZAQHumfCeeXbrqL
VBi3DNNVTL8ASSSdbWFsyJy/Jxxukd4Zj2KBOk96EtOlekojHAGP7HXKsc0ReOcX
gjEVMQqF+2Ts+N0JVqbxvGIpjv2GzVKWF3hF75O9sSxgW4CzVdWjeGPkkoHM73W1
vwzcmfe66P9lSr9+BVrUkQ6qoaNhQ/cEGaNLzFOJdNoxtze3vc/2vRCLkMU1gsPP
Yi4SrXPchySogegfVyXPneC2B4IcgRIpsS4oWdoSrQJom7hucSP4MZKa120+hrBA
lLMBICJJRGfCaQsbXf1M1xP2YZ2/G66rMrkYT9EUKI4vRPJM60rJkBDLqPd0OILl
bjgZ+AVgSbAsrG4yqQcjwo2zJr7sgZ+sdZ+X/Lbro8PaiAOjTSiXzVauHvMi5Z3S
aBk8S0WajXMRBCGIj0fSz280W/A8Fy7zlDv8RjPU991USTuJJ2bXWcjsGTb4Yls1
M5T4pTWHMuqjhdEvd0V74gloRfBUNbDI+jwnpHvvFdmOEQfi/iqU5+jY1ofCO4Pu
3Es3bHqAbZdO8VepIw5Uh407FjYvkIFoINAFMXoELiZWAgorihRt3fXvQGBHtpwo
157mu/THTUueu04UWXdAEDVXmTW6RSkphnFiSQuNiRB1dVE3ALYOvwnE6bxs+93b
6fdBG4c3DOSSn/sSpHxhlKrhgkaYO3ISZ8xfMd6VvkFrfJ0OR5fz7k1hUmrox8xb
V+W97N3FyOUqymjstsPQq8dfEA5QyFXxcRT3TkI9iCMrBc3IuOz4DefSG2ueQFmx
XKEZ0bsE+1Tkzdn4RexMTng/PNrFfAdpBXDx2xuCALHs1/tOhEweTu6vb9WTl8MN
oCX4df1JAyzoaSYmfRL1Suhq43bEmkkM96gz6vS83Rpr8nYxepBhW8OWJfyvkfm3
TDPXEngZvwT6SzP7drdCWt/rGeGHAFG5LExChgbFElnZzEa1TYUYs6N5QCaNB014
M6FWY5T5NcMoQ2xN62tKzi+awhXWRXf9/Fd7ilmUbydqUSEU4bAfTt5pg/MVWPLW
Wqhc+52ZhjzuteiUsLM98ByMM2TwQCte8ZdDw+Tm8b/Ku+3vF2grb3KmPOZZYQEr
ddo/vCu0gd/BkpoSlPF8qoBwLNlwo4r9UPy2XFBwIPmzgZda6Mb1xJHuIEqctJk+
BtEdjspRXvJfBwcrB3vEBWAQRIPa9i+xheuu7SwwaRvATPvBufNKqzzyk0FMLQqR
e4zGPiZ+3QeX8ix2aE/0tGhEkBdIGZckxQTMwH/bq8m+DeAGqXJ4+RLW097z3pVa
1+8cUdt9/ZaZN6fheplPjwxFjr/wJxcgPaBLe4gzNyCOSbV0AFEKa1o56i4WdGkM
qhvYtep3GHZK9ZVm16jSbkZAMAhen+fUumM3XE//pYuIT/Qvy5vAFOH+z9V87b3X
Ej9MOcQPhCVEEG+wKofDEGk9nZ1Kh5L4Jh/XRxyNB1JhRXaKEAzqK11DpQEYryV7
iIWNQNvf7G7Iu0647uhGovj8TekK8lHkyXL3XUiZgZLdxa2545WwK4WD3JO9TJAT
KrP6cqLqVgq0IVHw9IG2TwcG59m46qYm+VZYas2OQXyaJ4LrpQ7fNZFv5dQXL4kN
kXds4J9eZUscP12r2mEFkuZUmEHBFdm0l/JqXR7eDbnHu52BE65CE3olAYIH2yEO
0XtQeUvv3NbjoJWNX/7neT8BSPdIBAEsjO5nH4LepMlNa6LXe135UsFtVJGbZ5Gj
+vgomAYOpn0QP+Xz0Zo4KvvQ2y/WuQgzI4o+BI3AFYwBi92bvgYhQKnkDgBXSrun
4+iZ/Sj6ZqiVzCUc8KC9zCL5OWWDgCcJUizHkUNhFZwqmLI09zUGCRdLTCRW7eFF
POC/NiC3rD2VIHa7xxGTH/uq21W2Rg2AxClmfhao8zFAZT6MaVXFGIu37zG9rMqd
QEGHNjHtGhJ4FsgYspxT6o6i01m0DLIAD6kfBVpLAXywbG8z6WPFLCgT6S/saG9J
VQyqr2/Ajz3bigXaYhTXzFq7IuawtamyG0J5Oq4OJMCJiRDv0MD+OKlMNuK0U73W
dtF75kl3DLMWUo2NrxMDW5RbihawT3jFARrXnsYwGvSU1PelvdUh05e8JTeENqdL
prWfQ/LHwQrmCs1v+dH2ukNo2gEMPNFvoTEgL6iDqNI9czc17YK5mt1IS5BCHKCS
5MkB8jkuyv5uMbqqqQdEjtHsV1d4t/axDVn5LOlVm8dE5R44raobTaINunDW9DhZ
mHap1J6xkC+fqF6L6RFWgdN8/KtFgkYtuj9HmPXLWwYPXBVfrPSARkhLABjFFa4L
sE2/yyDjMzzaU/S/43UWQKUc+s3DT4eEe6gNZw4kh39J6C6sZJ3bK9ial0DaWzbS
3xdYdG2ImavRj+8bQyH9Yu6owcDP9q06SfdoaYcL5m02O5JcnKU8XMofbsrFwlZ2
bsCModIreweAxSx33yaKFxouWVMsWRnYSIwEj2KeeegESEkpdxESS0r1ZoNUQA/q
eyFqVFSXc39wY1jBvbv6fpgP5MsrOpXZa0xi0IZVNbRWN3+dKiFgft0IVK5ZY1yT
h4EvgQmj+TJ/Epd7q8oYJuNKvZ41u4qz606SB5OAcdJ6GaByHxftbmGqmSY41mZa
vd5ElX0gbW0O3jxy4wmj3kLMEZbUa1IwX1ill5SuAVQsduj4/8vd3n50gj8fV5OW
aaQ6nviv/CWCoB9C325qAIXUCtlTYnPFC6X1LsGV0QSmOA3NbeBCGYRX9aydxJSS
0JuW3C7eND3vIC974YWRkho/HvJOIYEC1Bh16WlUml24Ej7DZ05NvSHEq2OR/tp4
zHTcoS+WaI+5Y6rKeUF8SFqEt0QlCS955koemCTvHNet87EiEwyzeUJS2PbdC+90
crmJxKwyuK2Y/B5gwLOI5wwyvo2Yh6myIaMgWqIH7vGnnxwX6J0NvnUrKMjuOVsJ
IsDBSYVPH3WWHhHjjcPhpLzNv05F25AAArXlv5kDBY0DT7uBnU6XtYf0KgD51uXX
0M+/4edI0L9LvCRIHvwGf4feuff+AQb8wtMPTmmM39VwKF1T1WFhjFJ8Orm6itBu
fRLsnyHVyWi2yDJkUMhVzG3SEz3NIDHQkOa19YC+44WVqsreT7bhlXuOaHzK7yi4
dSi6lAh7r1iHZA2/VocxkARJhRcvHKMb/ryHLf8DTmTr0Fi2A3eilxCJd22TYPWH
r3c5o/xQ7PEr/JGf8qRpHdCstHXVX/w/qSDOaSn/5DAG8QJ5sQAu9SLzjkod4eW3
77rXcJTQJmJdB8cEEguu9y6uB1tC06lumul16MMUYEfWddBKWE49idW2jCQRoSpG
G+VX3o2s0jDtjyxeuhhernIEknDFgoXazkyHMRsL3okZimTP7Fvzzvlh6oZWeKdt
Dk54VqupTzZRHaWwjC45P68VLy6/pwaWD7sMBVkwZV4aE2PhNtXekp1rC20D/CNz
nttwhqaE0v/6nkIKAgslx3iTonVGSuHCT7CVu9ArgIXPIUZtro9juZGiBLf2dHM2
5uaq5ZM9530JZxDko7w0g5sCWJM62H3okTyVTp+bDd9x3p8zQ9t8dj9P+BkPxpZy
aZhILAL4ibkEz24L52zaWUOwTAJae8kxaL5PfNu9gBm+7XY0Enusb996fP+UKjC4
9QwftCIxMf4GmzNBNnPn2Rw4XU7XASJjuUqusWpq5o+HWcAyPBVvAy23ZV5bWAVS
QaDli8OcD/JVEJC2A8OBsihbYtYqgqsFlh8qtEAK1WK3e2YXxykgEs5NAFZueQo8
7IkvTHSgq67WbjaBna8qbtpiTiGu/t07h1T+buu0Z0rZvjwp8gfyqTjlKw4Ia2kX
CpGAjtzlJsUW9ywQ1g8iG5dQSxaBdl5BMTjDNWEfpAfILfU5PzBhYrDcDXHicZIh
ARX5eBPjNrhjl96S/PKLFNtltIMKoegQiHL8h6ZFeOuHrV0/PcUnfeCIy4ZUN77w
BiXjikMtaxOY8mG6X7dae9oe3gxpA2yneXmgOcmCT5ZA4C8cTMV/SQQJ6zPYsmcR
wJMxTYTX6yv1jkMdMsKjuQEg7bV+Q8olp3O7ABWkLWqCNkjMdAO0gE/ygXAPRk7G
QPqPpkdJvgb63pXx9GmRbbteha9l96SgL6p7n8OrN5reXWiCEtVtQk0qILNqmksy
c+j8mPV7Fz747b9XL+iPDhgOca+0wzs2mELwZQVfvuP/IAlHYx7lP8XQwTN1xs5h
j4pit9CZQ1LmvJykAXQsUyqkogSWIDjy4DMYmg1DuUSeHgvQUZr4L50Fws9sCh2W
P4s2WFxKRCM42h9/ym7c/9jYf5dqhHMbXMRSJjVInS5L+j1nTv69IVTk83nU6Bsl
kJYRQ4oF5gnp+o54UEhsOGhOxJAr98idljDnK5bOebdoe6SufqUfKIbtMjv1Br+a
WXFn6bDi2YW/KSStvzKutzFT87gPRBco36bolDMpQKNiYn0xwEMXF3tWzGKP0Hl7
QA1HrIcWnnXeACuHwMFL+fAvBUJcfrrVdsJSasYIWahnd3XrmIJXwyhn273rGsAN
znM04xrlivmY62XjXQZQLO2Dkx9SOkBShuIT1LwRnPbcJKau1/kf3/HjC+rz9sFy
WSeKl9RqVsjLvPWRdLjPF1FYQDBOmEYqncuUVIA5fE06kFfNynv9f6y4o7Il9tv4
WgBoJR2nqG5+mtf5aU1+M94EEqd9Az0VCXFCxYI3Wd4tUYv/pDE5FZ5DW74hOgHA
f90PaDFysdhT81BN7lbEJLun5y3f9njJZtD179EQLvl74lWETdpsWP0vcxWz5iHq
I4nhjR21ongWrJS0fL704tCI3x+D3aEncCgxNJwBWiNsYFcyBY0zDne33SacBSSy
sehBx653VvnNz2TARok+wXLlJioWH1nqIHromkJScWAEJMXghIkvN50ELrnd7Yxs
UyyuqfhOn4i5AT08+HM7JFzT05a0fHU/dX1o2moTW9HeNikl+DSxW9hJGUSoR9ds
soLDx84XKzModImwPRCvEMwP/UP/ad/sljyEe2x/F3Q36SrPGLSoTZEMYh1uI3wL
oQmb9EFaX8VnIgZMmyihvC3dovXAabkMJUAC0I14SJlpwumy3bevoFJWzhmgzOkL
cTEFBLJEaewirq6y4HhGGPZhvQhBWgNBG+CmMkZ3trG8QhZT+sY2YEzmv1/lpzlI
dol30PuhuyKpwgDP3Ujee/gZ7Q317T46nRxY6TRdNcXMFUwWe3mXGrF4Dzqarv/o
ZzZS7+0bsM2t0d+ML6POLTPv0Z3JIcqL4h1XLRhRJSH0P3HaGsxjf7gpXWhASXpG
00MTOhJdnFOFUrlcyIHJI8Pkw7OQXv9tWs7YfBcihXPja65tE7BFL4fuyidB+6Xs
n8b4fo2QfE9wGg4XxPrK1I/XcEJHTvkvGjVLR7MzSSwDUqB+84QEFpqQZFTid1eo
cJWOzbj+gqK0JJzQeOnPPVkuK2jfi1urhydl90sTgrRQd2JUhpI0cFfnF+IvoAtv
DM7ad5H8iXML0cwA9CS2YzGoDFNZIXDyqnv9z7+NKhiqKB0r5cDbrkO866alT3Dt
jPF+DWIDeVXAzKDqH7lzA2S9od05ndqzt1ISiq4HMniwvbY7x7ogziwuN/U++FbQ
Ozjg1EwyCJn9Oluv8jx9wBod1JVlgj14MoEDVTVnXWmOKcJeep0Ry0oNBoglMmW7
NfDivdZ9zR3lL1iVDPyYJg4SQpNMU0NoASVpf3MU05PcBO/iCRtnX1bnA4EIjwJC
I1iTXqdqMRn/8HlEudq/Oh8ZbdBCZzeuI8T1tg1l2+LBA6oug04APjfUkpxQRzOx
vuwjFgaYZdcx1Ou4vpMT4fOuZLeb98dyrzPXrMBFWpIDlRzoIJ5RLZCADs94m3Nh
8Osr/9GCETple2LWEQ7pMyyVkKRii5eFE+2/lsL+ZKqRaVKNa1klU5iPdV/xZfa1
OoE66xWezgpPf0638TSHjKgoXpOri1Zy3+bvpF7Qh8N5IrJIzR7DPS1tTK0yaxwn
i6F3tmpnBQ8sKD1sS8QZAa/R8hwGhP+pjiWe6n66rk454ay9OSkC37eYnPt0Mt6a
coTFaRvAR9jCqxQBbZybGjgywnyWoAuYMdbIlXsTJi7KqJrFMF5nlFYeol8Jdx+d
FTKgtdGrdBaJHwJpgIANlUJwQd7GguJEkAPsn65vphmVNoZDgGcRCZ/Wpwj9SBm8
vuS1u+qfmEuP/wiyAbKAl0cd9uScbnEViyYmmknQ+ctx5XgEaNwUq1rrwzTCXZuK
0CfiA4yRZ4KhqHC9ssc8vjTzCRaAyWMdbyvr+m6Yz6OaNWhjdhy03GkQcIYgmqfS
v0X6B6GTgxaf2nFqzojCatJzDr/jgTqBWyCK0TlyB9TLFS0EuO/YZRdjtJqxcTSe
Mxx5CeWRkHBgZpM3VANCiUZ+PxG+2X18un2ibq6iySJybUhf+YOUhGZqnrNFdfJI
NktA1TrYxjwRiUE4dbKvkspTqDyp05/TQF96nMd1YGYJtY3Vtqrd3G1rmJusTopQ
N4YT8jKk7iXvR9Rqa7MXOJvUCo3BgUq+Mkl/LzUsG9KgOaZUh6YkV0NgWTB7gWt4
hcuibZtlGKwWrAJF+sgVAWjLXffP0dZTCEDp6i/nYf7PEVuZXdt1VFLFXD80aWXH
y1eic48oqP5XA14blRGopc/aAxGMjD7Xcf84Qo0GsjK6IWkaEbRDf9GG/83M6OKA
qTc8EjTBpvXn+yNkuYeTFUfpquqEiMaOMrGG6xpvJsYlWoHbLTWwdUDAHot/TN2m
N91WG0kjp6ZEbdTpwwou1Rh8KTfQv7bp9kObjYpKvKFcFj/ZXrwevCyNsmSYVoya
jpL1nuphwexnPj486jAGK0YkY61H1Vsozz7K+EfKjuWXfjsYoQYHlzMvGZwl/9iS
xDD/nqeTp96BllbtahPqOT0ABeSl62dxRO2ljAsQ3dZBm5Oy2t9wMmacyEqmSdhh
5Er1SJi2p41j/4Atr9xpA+Qx0A0C7APy3asG3x/gAeKU3Mzti2iPTQg45UlXxSyw
iegTilwAFZNem0aIQYPV9tj0Mhbdy/MLXI9S/RD8MT+OO/V+ZbvsuZSPH6Zc6czN
c1Zutqbrb8atTo9RBSIpxn3hmRvjH7wBf8mMWp9fu98IfRQ73S3pRgZVcTaLwOK6
WQ81l4uE9yxy0ytUGlw39UO7dP47rz3XjJrcnH2f6rIlMNlCY110LGXWBOvS3ZtW
Qrw5qU3+PgZAlbQd9qh25Dp29qAF1jz1SlmuW1BHHbvPUHro26VrlE+cc2z32b0u
Ot5qSCUbeTujGyKvNGDOmIsPHRhBsFsz91z5IVAUsnMDsHSYAe9h7gsGO2ong6I0
SlS5JXPJVPzIabkL3bOcmn9+v8XnH+gbPKHdST/TMnpS3qv9MHISx/dm/YRzggvF
MUL40vCYQxp4y8h4gM6B0pAOYJ5QOml5/6te0X4Tavjt3GhQX4EexBdQn7IIGp4Q
7djDgMiFM1wzSvbchRMteBlJ+vItbJCbMxK+xF0R6PfoOj3H/rTAfPvw8851Ps1L
KBxay5Rlgn5KyJcx7I4G9XE5hiFQbPfv5o++bvv4cqkYi+/vZzNyHjWj7lg8WQnX
hVYW5NAeGvptzRlBuJjMRHJrFW0PeHRqQEr+2cCJBM5hp38MiW+XLEPtaUR3a40F
ISaVLoBtlGP+85goFoKLdbGi7sLB75uP/Fv1Q1fqteqppnV/q8sicJCE1ODGnJZo
0uaLe8VyNpEWCE+Z31iCLf1eaUf+GVI6uUdPjtJraHOnzChVYjimImSd5fUYIdZM
MO9giy1OuwwoC5oN/hzv6Ioo8A35+XjqWYES66BKwJ9kN5WcqgV0/9lfWl+VYTHa
if/SWZxMHDCK/GB50clAVF04ql/W6LtUVLOuxdBnWa+0cgG8gw0VAzM3J7jAW02E
2y5JEcoJOK//Q9PaCv56p8GqQD7y/X62NxyueivY/AhMfEFEjn4oQzdABpGgDq3F
TkyWrgejmxZd8ynCQZBUL8sS1FZ28KGuz9U26pHW2xqFQkpgzI0Eap5Cu7jfVOph
e1VRJxY9Zkq9QiNxdELQJL1QvlLldUKeJJkI7M27lBs939X+mlnsc8XT850ImnZM
E82qPSqizLoquB/d5XU7LqiY9yeE2Mqa6KQQ31YooH77UTF10bFXW3Y45E43x2Uk
/SY0HpA4NTtoxCcCCv5fJw98c5Ys4HyK2hDGKteFD7V01f5CM7w6nw6a8/T5bgXo
KE3q6PnPkCdC5XLSBCSzyJLNkzS3tinGRNKH2yV//3l1yVSRve0OwPA2KbMK8m9t
6JrZd86CgOKO7SDjZdNrNwbdet/50jyUYd5YWxyD1iXLO5gDxhRMQ2Y+6cEDKUCj
5z9nqVl9T8bsbpIj6Mo9UNsAwAsz62RQ56ibnefYQnrE6nTL0gGXvgNGAlvu6aZU
uWoj3JUPs5333huoLsMaeN5TZpkRoD/tYb8dWzmZBaR0urHx6KYtO0lZcWW+VgNf
ABC6QtGds2/YZpvesfi3KglYUrA3SUrf7H6j1WzAVMQ0GyTy1znlF0Li8g+I4OLc
7cf3CZA0cIgGksU1nySw9eLsV1ZmqvfKkH+zzBhh2BO9urZr5Pv2KS0olazqZsBI
qytQFH6Lxn+YNHHj1FS0oR4KLMcVQJFG+COTwIyuf/7cNwTFhI3UvZn6a+mKxoo9
Y7wRWNmL40u/WHi7AazdTiZqfjIWGa/+g58ywSJeM/nOj9i/0sEMHJe3Eki4Qv4/
izk4k+womaIQcLUHRqMuFBIqf1uota/fBazaK1/DMtX8/lXS6GhEvX3zUEi9G/Lp
78iqz1WHevv/aEtvEkkUMrw0OSZzm59aCKvQpxWEPLgISRoFz1bplL9X5oG5WJmW
f+6TeAi9eqFiLECtIFGfV6g1XmZgT8ztYMlkW+ZsN/sSE2O5QVofo1OqQjilsGtJ
DHczoVplsny0smCxllwkMBATyTeu4drDY04V7IiKT8vREfZKdjFxebcKglB7Bnvs
E6KCQWq6nBu7Cyk6GoAF3ABfsYJzGoolPZpHsxm0NlmSAwx4vY6cr6WwRaFuUmDi
NK5SV4Nz/jrXuaCAmnRYId5Ngc7F6xjmjROmTDUh7CKectKK+NUHImh6SsXWTTio
VQDKVicW5RzYc0seiujKpbwQst9aZ/CfV9tgrIoZxVxUBlb3GDZbhvTJ59qCSh7V
czwtzJK2yQkz/+aBslvr6cPeb392kvn5wLDlRxe/7y4VPCYijX0aiynW2STC+sLb
Cs7GmZjdP766d3AVc/5OvakfO4qIUmNTN0yWo1UAQcVJ5jR3JK6Zmy1Y+A1AfZVn
UFjREp2gC8t7dWkYk+dyNNp6euUAfsPrUW7dWaUlCrRTx0h074WrhTJskziiUnrZ
aHZBUoeXl98cwpf5nGbOCQLv6QWvXE3RC8MeHJjKvuujSnswxnh00dbxQZScUcQU
Fa52FuR6xxrKWzrD/JmhtdpeiO8seoH+NQyQxI4wlUbFRH88B2CesfhH5HfmjtZG
kB+a8mysiHtZT78VTXedQUwHuBu5Ehp871cYUDSQNYJ3sELHdHVKGeI1d2uuPoru
ERXf4WHhZ+iq/Q2l9YyGlATFDv8CF9gxy8CLSVQ5UdujXnc7tepMrOPMLwhonC03
MfYL+vb3/5296ZqxeEUJpjJ4Tdp6moX3nqdRIWFZFXhyc6uIAk8owWhnXfgYW5QS
9VBI4aoVEb6766V6VuJAMrs5ZszjOHQnWPvYmfUZL4bnh3bwFrRRPWXBORWBSSBI
TihXVDAbX1r3lewKuinJCvWqA0vsrRw5nbFRIQjrLTvwOrBBm2x9/OKte6YcxbeG
DWimJLJh3OzzU2L4zjuFcRKH2nyxWjYccYIbfbxlEXDw8/xGWRR3VVB992C9ijHE
iHVii1doRHszJIBkVwrJYOCAhCYXeqHulG55d1MD5yQCRL70JeUsIg6GnU36k/f9
ik3lmHNGCDNvQ4d63HEFwuuU3M9DDVicRzXF28iIu2GufFmvK62yxcbpqkiX9W/K
Yh2EFRIRsKE6YfNlyJ6KsBCHouto4OR6KTCGb4lD7iN706J5i4nq5E4q0L43D/oy
UllXSl2a4OfCUNaTmnIqO0bvR3TNnYzVqJxslUf1MTXdtiMevR1Lo+W1uTxPkdRw
TRkhdz62iMYS5b0dDrDpaceEFCjKsiPmgcxeqOr30qR79UdtnsWvcsDgCOZUvFwX
H5kyJWaafdi9Zyl0J/bAq2L0U7Ag5SdQUlwemijPmOuAtsGwbBKhN5dyabDRvLcT
YYmksF/Wn1IZVrC2053SBZmzAzcJb4855J6Hi5sVzuAU4AUu58Ym46vsAQM2+kLS
eKmytZBUxWpdLiRf5KnnOOVcshue3LuqIN8yELrzF0BarSvZUtNU0b5BExE16Kfq
xcuTngKikHzjT9d4ctiWqIVpvZtkCkFp1VWx7wRinMAs9v4EPg0Z1UV556xvPjFY
RuPNHML/VbKaXKonOcEFqqcHcpTH4t2EmQXLRUfyAEX1vKGteBtD71FzDCZIaan/
n7MVpPbNS+wuTdHRNUzndj++YqLUrFjk5DGgyRI2rP9JB0LGeQFbesNPOmkkZGRm
v+SGwDsgbnWdYWaHGWebPYFmUmGmTJHnrWBaxyXAUIV6G7XuQWOGJTS1hoHYTBE7
+iPPaeZ42IB29Qb/RNPFyRpmML5CVrcB/+KRCp1T1c107dMByyg7caiMCpLpf1JU
ziVIPeLW6uWga+3KGOVZ8lygeM2cTKEYGEOLuGyWab++d1bAqlo6lcgUDuBVj8nc
7XvD4HKTkt56EsX9jcvwYcm/L8WcnFZXm98U189y9RQtncAVPq0GOV+x1pZMl1KO
+vPQ3nalZaBSEIszxh+EvlVUgdBkF6PyH0O8WVq1RL30ZHlB/JQ2fkSjakeFHR4Y
Ln0r2wRdceYZb91jDPBUnuCnAr+D7P9fK0igaDH+oJNLrEoC1onTUzhX8VPe2zlY
7wuc2CBrKqQqDwctfwjQrncK+Y63pcz38fa6AF+VY6GX/mstEAuQ9zd9p8LQvCSO
8yqL878OmiI8lE9RGLmvOK9lsanf7hKVLkJ1a5x9qbx2vMPiZCVHApn3XAUj448S
Dxcp+qoC+wEJ6yTdcK8fpMQA3cH553ua7WwTHG745r1dcpt8uLmM6mdWbiIyOIar
yaI5trXgx7Uo4RAjJcPbiZiCJqG0/XUHMdmtM5/RY9gTJ6Q/Gg2l5lMZZiYL7ffe
QM8u7C///oaYij44tf/wkvbsgA9hvrJpOwqGVCwGZoDzNBZ0j2eQTKLA4y+O8Kbm
oSBH7r9r7EVbNXF4DVVnL6ndnX524hbcEci6K85VoW0MXFGYWoDAR4r554rOxNon
ZZQKjv3IdCqHypY3Rf7LUI7nf4UnIoqBU84xLROqDfKbIu+Z/uw6ZGfIlUncKL1l
DuBCmCu4SlZo1vNIu8I67sck7Xp8MTQxFHGPaZMNmKBL4CihahybDm3S4hbKXhrt
yav56ZclFsH4/oATFoF304HXXeDgXWQCWHlu7samBqp0p3xnYoFLBhmMzHu8WYff
Ohz14ireKCTpSPMkJtt84kktdCbtdJHNPpscoTBtWLBhI+J+YATwwJQPB1sttuPJ
IT1j+ZpIc+Fue4KKNqSpbaYAoU5lotzO5irQCKPkM+prUEqFFAyPyCQjNG0n48b5
ZSGV6LTvGiVqR2eViQEcdHBimH7dg+5hbT4BsPD+zyg7d8cq615fP8O4foZri07z
Dn/d7qxH8hGhyHZNCD7wj9HHPgThnAtrDHMs7525mUfclHFj60Q5IcyoXTLboMzl
2iNseIqBfIWIKMzs+6BthcP2UHgjAnnOKJYVCfW1mG5soQ4Fh4oOSuVa/Ugct2WT
1YQXtfoJBSqnvVQItBm2GSWW7iwUck4Twd5xmohQdExjLFUaXcRa0bRHd1loIrk3
c5b4kOvwu9cILBjk0T1nL1PW16qzOPWdoDFhQpSTpRHaBWU0uLCu6TZ5oPcPMTv1
exN/fPHsW1hLK6JKHwNcBj+dOEShDt0eZvdmEkwC95lQNAGHTS26p2rZT/lPJiem
PFOi70Sy/XH/iNrYi4cpfiLzMKV9mM5y5YVADlyuwLp5yobMAV0JCUM0wLPeL7Qi
iMB2RWqE+4CJ2kQaxddOB40Zxj3mtfucXIhsVQpQKwarghJnaKoOEKFARE6gvhBV
/dVBqkdvkPSd/z4xhwWq4fMSv/OHNwPhHJNQ2LjzzJOb9AxigCd+ysF/47bQiC0a
IsB1gpXl9n/ADGu3TFe/ec2UM5zELuvfzXVi3+DPBSkV2mh5QxLe6dQ5i4WvPsGC
V/TnU05UCAwns6c6xhTHJQgc6kBTM2dcG3Dg9/CnIYMGdfRqxrNmvyUpkWIcMvt9
EFdJk4SX8yfABioh42OefGxrzbWXSb9S4I8KHunSj9/WJyR64ZrSj9dAoUJOX98U
sBHIvXJwnJy2G6QhgGNe0VZaSKYXiPguv7jvg/dcuq0YFRHCtqtiq25Nb33Bmywq
XwHbEfNBzO7tEYYOFo7d/BXWqvYYryWDgPCn4RJDSBzyaxREsJ/dse00/skIq4PM
j7R7q7AFTHLTZnRt4accboykTI6xrbg8dlS+RXw0IjobpfH8lkygF5ZmbsjkVeqI
WREKAj35FGwSoVzAadPFRIomyYTzhAULNJtugUV0yIHltVeuwGYueuyUt7vO3SHP
6FbKP0JG9zd59aTPrVvcj/VYqNdRQnpnoVQqYv/5AVVLmfgoj3ViIZsZ9MU8/Qy5
oNKpnSjJxQypv5ZoeOpcW8AUJxq9H3AW9nJ8TS+09tUzQI4c8Ch7uK+8QOp/dNAv
J1AM/cIYhucmOoqYLqLw6nBt7LlxmWVKMMaLBjYe4tZgaRbM34yjaaAtEy9c73zx
8RJnunTZidIc9f7TxJKOgDw+AOBnLFhY9z6qeJYsuozb/GQz2Ur5GXPgnaac1Juc
jJnNYQ8+l+BC/afDG5bEPQPpasx8BB0cfzEjwYrrSW4cT/ZEOjJIs4Tuu84AHVTt
HruYjznw8674rQf8ZTNnvUmJuwUjY5XU2JdDt+69InCx+DLO5ItHIxW/5V90Um02
5hNFeLRHNKYN3FxIEJL6IKPmEiT3V2VcFDfyN3ceZUSuyV/s2bLaBYptTrpGsyuC
T8j2UKRj4501CK961aG8PhdBdAF3t+2/Ct/uuA1ARrb8Ad+ffbCUEIQqJ6A9Pzue
aax9OHQIp189srMN1m6+CZIUOcX22xXT+sQ6Z+HHnAdJsowOeLwd9qj4LJ6Hyo8G
oM/6JYHtBJPunQCC9riCnme32GgA7det02ulym9R40726LmI5XHb6Jb/TMEW56wL
cHBR4LJbRae96NO0ioDCur3jO0yG/mXXvITX5rggkFOM/PEDl65iIVkPbRvPYBrW
dQHs2fzQI5Sp+Gw2J0fkvptC43tztnfs/MJpFf28RcWjxUWg5SeaU3WMf/nEYZ/f
kLj3gV8KEsUiIWCgsD4Rj4hqP6QY7vK55W9rfUQGxYu5RTJbTnFsUbkUxovyuVWo
H5SCSwoOOgglj3QbCO5vHoFvujgsQCuLmh6g0cc4AGK0UgKOefOs6zjjQClWbbxi
B0wUj70boxUQyCyZFkkupQ6U0F1HwXx8x++S28h6gNYZFaZK/sJbr3KB/aUJBlK/
bxjHOxqsdbRV4t3WrqNYnYs5EivRP+XqS/Cfl9FX2l3JXDmG9KGkf4MxHYOjHcG6
e1LxaIZvb1N+lmjS8KC3bHNvT5cAwtJczun9odNW5NMEhMIgXwYmNF1T2mTcXLyK
vO7nkmxRGocWSboPU/y1vMJ7YFugsncw8LztfvAahXqJ/1BfNItlfdvmOWACBwqK
f0oQluGOuO7I+4O8d6AJJpNXrDBcoK4qJxFDuo5uTjghVcU1NwcYcqdVpTNtsbVP
KYumCffqs6dVFqIEaruWDlYlCFKA4PzPNLicShixuAurGA8GsPyWToHA0N3/U1XB
WjIVgsksrwDnNDCgUwI7XLt85QMn7niczOYRLTufNpLztY1lA45d9UUGjhypsSA1
C8y4UdSl9N/W7lmnoDWBr+PhU+rBXIuNAeX9jC3EM03vGX08nid0JZCfFOjBTWkW
mVWwodwQiBgdS2fMMWr62cpCDJ9OzbrsEtHOitwuRPpb71wKhtM0Yx310ZsfCz0M
PhY/5qUCytKFs/Cs9fNpe/inOzOTCnW9RzLrGkmxPcOF4a15N9gnNDgX0Mz3w35+
ed5CRZe1+su1MJFNJ3miq4SBdHQFC+5NlUc8oudPU+WHno/OSUOFSNRFa7GbE1MT
jCNmqOPMCLUUh/5gD4MtEeZVN8ittf2D3T/kicvzbScc4UyY+yyNutaqJ87tswnv
OeZeKL3lxjqMlPYx3XrtBoYDtT05dwX6tNPcm7XjIP+XZj3mVR1uRm4L+2x8diYl
zt9R4filzLKmGrzGzvBuLHMNzC45qbD1MihhALsIcQTIh/lwSTBHpE2mNEePo6fI
SSy7Hf5/oBNZcLqtK+ZiIWX8Sqht8VTE72a8sNjV2d/nh4PAbkpIXI8MW2su5Q5s
edjx+GNJs7Oib7emtkwB2QPnkh5T/xHurJfvPUVF2xFdLFrCdUlj3aTpQiP+yOvZ
eZkMrQyh5GNiz1clT/UQg+JZ0dEvV/lrpaEM8P5rke1WPEV9gXVY+e17cLDW+KJ2
Cq9iVL1oWNo//ystxA81XEa2MWXeocgLSr1AI1R51icI3cmWMZZN85dln4Zd1Ual
kWy+sDEVyXiZCLwhAfe48QjaR+xPxw2lZuocnLGEowVwNb0ZCaxUXj6MyrFTMEy/
i7soxevJkDk4BCzIy6HqFChQPpkifoEbtLoufSPrfnAnKwmqNhblrn8jG8S4BV3i
yueK9QTCxqcmZY3pSIBEL9qhWUodcH14WNEzT+jTXg6kKe2kshgE4Ra890Mt1IpR
wPeXMFYsTU2xSOhBrxAgr3zhaCuJvgUMOddi40DZIENXt4DGlt8fjOd0qD7avN4R
eg6wibLpgy8fxiFxYw2tViSDJu23ZxPx0bhFOAn4ZI1lhYSn/9kNi1r1A6+7CL2b
5EI6y4HVpR2CyhFsa3tA//XVLc3qGdwzwiMJueLa1Z95aNL/ImMwC3KJBmRGWQnm
VyjQgjfBOrUCEJrMEuZ3X0IY17S6Uge3rpjOx6yNOaCvY9aK5GKpwBJvudryRDOc
J76loM+Ze0Ywev1bzL+zt1yyKfWlgDBHSBJlM0g2PyIWEAWbR0i+m38j/vVJoFX4
k21YlHLG3wIknMMq7vPaEHjeJRGW1NaeJKAEAOAQqrCBETiAyhosTkA67wVtT5OM
S6r6OjkX/YRYKwrckwi7EW6SwcYBnjC+Kkv1G01OhLdo6GDTJbF8F1xQSNjAE4UW
VoZpkmgDvWMra4UW6Grgu22s+juv8mVs1NDR0RfVhV7DmwbIcw/kMVJ336krTF+w
Sok/9F8ZkRBBpciPAIiKRQGJFQAloBOb2vZwLv02d3+cmHeosePOBSLpcDHUt6v+
0TZhxrBe6qk0JOHbK0TMBS/clHPTDGTQ4nXuBqKwhC2h/Yka7cmgGzmccX90lRgN
kzX8KNiYlkIstJlnP2v46h+x+a0sEo8OQpTtBe3653XVGsnF4rTVqhCnOndrdbuN
pUZv35ag7/fd3p9qRWwHD6Z0Xtc3dY2wx3ynrrlRDAscWFfladTJVMhpaMUrNLDq
Fl93K5eNElX75FHtmqTxTnFojoa2w87QHk3Vl6YFk/P3V2X1qnryRndF+/l1UzH3
BMmfZ6ZispbFfc1PJVRO8Lo4VWSzh97GRpGw0wR3+bek3Z4fn7IGiduNQaHGAsEr
kc1SdecdhHtwA0FLOiizAHhLm2Le21ounmpQTZegITvfsiHZfhwXjOdFLvtPOrJM
CSYX0vH9o4b08Ehz+ZRgCquir+zWZyoYxol5FzSCx1CJhvZNWIE869fB34/oGwcL
6oNQN2TIK4PZtgzW5re6clMusY0UXLevtFtKyTHkMKTDLsibQ7c2bjPiDgh+0wed
UPPewtmekfXPNoAaZTDU+6AHuflzZrKLgqs4VGTMcOICkto2etVH+fum+5UlEQy0
tEDF52+I19Z+Me08vegyBiaYW4lz9PuIX0AnMBJ2BU5jwygSmiANCWgr4LD0uKEy
u1Qymf8DVptNQ93g+9kLBURIRSjFddnl0Y1129uiGd+ZVotOAp59hElbvklY45+D
tOXLC0msWQppL+e1CM/VFZKqIUTwWk15Lc8LN2jgOjCP7ixpF6Kto+pxU0u7T94K
8vbYG+l9GL86cnKFTN/pjIQ2j+fT4u6mDppt08i3BlVOSMC2LcjOuikTDk86m1iT
pq6E+fckpcKwAg4StnVpNs2hOfXCeOdWA9w2ebLsNKqH4y3PUGwd2EJN+In67hkq
Teh0wgzRgODTMFhk8R73ITCYKFzyrcIv8aVGXcQkjdv3C0YmDKWcXMoUyPc7Od+e
zvnr/Y9XmrbMSgglO2UFtU5DdzN9MNOm4ZoZaWzbuapJfq5QnMhhmDJUphC+Y5k1
IpQss1HSUZOParIs0GRbkPbnTSvVBISFaEdBHrY2tLuZiEFjBWQESeuGMSfVJU9M
KpI99yhcEidiIb9ol8VOQvGmdaPJnZzYDC+F9GPiTrNLyQBVqsraAhCnj86eGcG5
btfrnaclw2Gq70LTHgntsRhyzg4Y+RsYlaK4dKrCRRbJXKv2w6vCMNdcxfjIK5fV
CdeI/uucAPMEu2RxPHhu57+rI9o0Htxwe8uXZCuoTt2/YiKbiaUpFv89tAXN/s6H
wkFNToKkT32a3haN2ZhXIAOK1wiVHBAlhTXMOpaXXza9obd5CmqepMGYJA7jC00D
kh1k3SQrHCcAUul8x1wfpyGJnOgEZAXix2HvWD+ho3qyCVZZU6KH7L+JPYc52/UQ
VFKI9VzuKeev3vW82p+uMSqO57xEUd/km0tqft2zuU6vZWrwUVIoWJX7CEdBINo3
pN50nEaDTkO/Bi0HhiAHkaPJAQxFIqJwIYwp84/GLGkcXD6VTDfIBhAtoOnBx5kO
lBHs+YgT+pb5ADSBQCBoD/KujPZ8qmkv7I6h15KtSPqsjuyT16KLvd1kT8jVxZBA
W+NCCYWgpJDTt6o5Is8Bpz45iJNxR8E7gq6E5ai7nCUuxmfxk2PzrdPgrNuOUaHb
4wvgA5vJmfVDJm8J+48v5FA+D8EFW3r5Q5OXCu3pKBXN2wxW2OePtrCMpCIVyhKG
FMVpLHXpkiHh+cQPvchQiBPsPB44OOePKG9dJu4nDfGhP/AfaiQpgfHy9UXo4Dm3
QBa5/9Wp1GQuPu5j9mmoGKRpvNuyxGXbNc1BLAFaTLT6WPPwKKPNGbWJbhel5REX
SXaFgp+5J6B39cFf52yp+ckRfeZ3FO03xK4kcB6Ippvyr/4Ed1iJGy8nlrUuGwCU
BSQnS9VS/An5RnE7FZSWoW/xs74kNWAnBIUjIxBkZ7g3LSnYWWCW/sJEhIkBv/Ik
KOtUUocvBZdzM38tvFyjLr2GLCn3XN8uoms2+g3r/o3vqXUBKiRkIg3mwCbvq6bc
0jUiKL7ibhw+atcECZMb1jZsPdgffptz3liNlTc0BrVBAOLuaQLDWAzB5xp/uU6i
K+cGzvTWIIgkd9iPZam122+pMF82G7qQjIUeDqBE7Lau/O2b9btdpsl1yzOFpL1t
4S8qvtwjgEh/UF3pfUsCOth+JIXLP23yc/aP/wxHAm1WQsIuFEDPwyw/Q60l82dK
Qfkmey8yFYTRZtD8AbDwO3DXpuTy8htfQbHuMYqya6yJRV+a2nDd8ytMsh3T64yE
9sZwL8O1y1njjfneHj8dJSGSBgZAbhTUWjFGjeMwKsFTthnJiZ6uZ0H4g1kqU7af
7tA/WwXmsIwGHLZD+fejyHnN+iz3mIudBVuZHrDjl+dcv4d826ydhptXAhabOa5D
1IA0EHsHE5toOq5+R8EffA+8415e08i+kB/QEAouUE+ORMWZw4t+5k6ZgTbOUAxL
Djl58QxiDTB/m21KlSmfvV3bz2hykqvCqprFfYHoUES5U1cse1QAftZYf/0e/9me
ltXWTIwEGQLwD6voWrie1TNBzTLBykHj9g8Kzt+nSop3NERcm3hLN7wqxiQl1mfa
nrCkRJsc/9LnLNNpH6E5YdAWMpVxELTbE8VSwpQLmc44d4uRAvX0Scmc2tUFYt64
cgLt/VBL8ICSdqDxay9mSOz/Tto4dSuiUQR1mV2VvELBGESxUti2+VKk4JE3RfDK
ObGN3XfCIevlxqtmLNiXJEEVDhxKbTS/SgBtFxPBWhb0y1GSN+Pw+LqTjuFi6Tmy
JNhC/65F/yfkWgyIb1lOl2SAzxQuBVx5zn3+TPTITCyVb1jqOCKKe+AnAeZcmqgG
YnVhacMrTrUooZRSMN9w8qAks0BE2SGcjA7eKbdLJGd2aiWccvf4YPW9fKZE/9+N
e405aPF4SEH3iSSu+WjbZGOP79ebKg53U0VEvvgEsfajzig6JEierM2Au1hkNx+H
CDM3oKAm2l/qrx5PjtvL/UaqSXWa6lffwg8U/b/RIkFvEphQ3dnI8Obe1SAXIwix
FTbacvb+JzUw8gDIjwsnLuw+iceUZ3JJMCBKccSFSRrX+52gH55gIgGMFEAJgNv/
UWrgNMz0ggKPWhnCva2xApwTwOeEW15cXSLrUa00KvhEyIlWQD7F63hkxkCr1Vm8
8Fz+4RmGH+hjW/oKBnvt59LGLTBUxj8ELHi0a50nE+L7FKLhN9LqGSlMx7upaI0J
67BjnW9miEjjfWMscRYUq3haJZDyQaLNOm+BL+PaVV3rY6xzO1nkd8lLxvBth8Yt
3yZGDAPsAv59zyETH8d41+pnWM7RH95Emz67iLxcCCCaupqvduyHq6zCBF6PnGnf
/o64P/a/xOUxtt4pTy9Eis/BCwrYabKboIzCvEeq3JJir9SFMX6iFqUsgRMfZLkR
izA1PQWU7ucd0wHfzPJCi8PYjngJ+QYpG5m2yVo3v4HE2rYk0cyYvGbsRaCiZXu6
m5G+WjbrJ2Alkvw30s1jWjPuhe8rivRkXbi0kOsrIuCBKfavEaMBo7RM7eNiL6Ux
qoaCF/fe4hLNiNmrQT0yxuuX38X4f2CmwXkQDSFQPFH4f8pPl2vbmFayTdazry3y
7v2cxf98SuDVYvXKagARYkCR/qGhQH9LGA1FzxJyHWcEWZQSz87mDL/F0GXqdOm+
woVpK7pg63CLGQlcL5aH0hAsOF7LKdHZrpOkgFURkK/OKb/uh/dTz02sYK5/APle
2YyP71XvNssfbLLpBTL7WdGRlUcWWM26EL9mbPn3G1mMvPSxn/WBzfiX3rPrAj/e
+dVhuhD0KVZWOp37YMiOV7aUiEsM18Jn+Chr7M35Vp95YSP0/cKcYK7UkMWsvOYz
II4jiDtV2QMvdgNc8y6bnWbr2flmyPnicdy+37r4Eu5J5hjWSJKoVU6wyY4nBMVc
ov/JbaCT2vZ47s2wJh/+Q/ATZEKF/RMUSKPx8NSIyWsPYmIYuHnHUgMR/OoFyK1i
aI5TQg+pJ5PXpU4W/HRSrqydcBLBa5I7IOY0rlLbe0Zdlpt5wt0ZoEhzAG4lxbW0
dLS0gH7REFTb0Rutp4o1SqYu2YvEtgsSLAsViFhpW5NGBWsYqCwmb3E7b88sDKSh
DY3JQRxVTTXU0FNEHO5WW7Cc66y2ad6qEsqvKvQVA5s54el7PAremG+g2jOZG5ex
Vv7Q3SW/ftumIy1G2qAfMyX7grGXhppq2ic5v/Mvbkg9Y9h2c1Z1+8jL2X7MokjI
54ZSt1zGwWu4gcoBSvWH//d48+cStxUT/tirTdM2izw4w3RI5zhGPGPwqL9rpUcg
IttVxbavxWFPE77hYW5MYkRcO/uwKrDO76ROpLUjzPNFCxAKf4VcBxz/EC981rh3
WvRMQR/rM+yw3HTd9k9DbdwDqnHFB0CVBZLiacVVcX09jMgYnuF70k19y0nQ47PX
xw62PW42ZOHaDgLs2LLVTlqwahpTgJUxz35k0BgqStNWNYh0vxc1ybIvEnbvXNvo
qbpqSrtbxN5IPGW5C4bG0gzTFIg6I405UndZuIddEMK/4ohTKR0BglKvehNH41RG
IPGHkJprm0V0OvUAgWB7BXD/NmGY/rIK3uStPKh+mxzz8Q1NDjUwqsk6HMgrja/X
zfxOaHpqeT55eMlwdq8qz6QNPOqMVxm6YqsILSmh3W6TinQaUomwH600kGBkr9U8
R7wfBjSv9jgYOzKSwMF5jgVMjnvzQ6cKT+F/sHxsNLL1N/epHEJjOHvEfW6yvZcP
cOvB3F/tX6NXDifeLXMO9ZVQiyo2rjNhJ0MBVwxRmuxvA6WnnotU0tnt4ISIZkGD
zP+me5JgTxYHXzjH4rdN2bz9qB6l/ZZMrJOXIja7Vnsh3J8KcsMHUXAoLvqhOhaR
l3ZeMWWE9yOlkPj6b0khGjvmG3GbIwK6IExKiSp9GHNR2cFTkbDv0N8gVzZHa5kY
PJzrp65XAxwxqlf1dALR5cO5D/m3Tu9UrQ7xsYq3ysU6Mc1GNbaQ8hJePUFv+KVJ
hqqfsBmFabCIveUX11sST7Iole99inUQTfla2DqXaYM8h2DkDsLVaOH/v2BzNTcJ
bbuyaQEeeruTLLXKCKnMEEWl+6kneuAJYAR9scuGbUjZFSgT+H9YrWXtNC/b60ue
0p0vBmy/ddtxYEIvYkgmCsPZDJIxraZ24sLye3CiT1ho5QOsU0RJ5p5EyVbgaozk
NwjsueAdqQYvRMEWBcpSMs9ExJVdvb+m/UHhcCnpXzONo8+VqGUgjqAkMvv8lTF/
9dJF3aFG1RmYW+FR8aOPeV09mrrPYyKyVaSIdJGi46iYSrv+yAmFAIUiQ1aAd1gM
vd6nqNlGF0NH+Fz6wY2XEw9Von/O6QH5K65QaIc4n9mMDqCvK5ihqkg0FocGVFNa
dZwfF5frRdus6YaigH2vSli3f1xaenvwxVCj1LfOAZJI9bhXqCocoaugBqKRhWS5
9n5bLyxfm9zEiKJQz7fHXYrFJBiB5Q915DSKJuAhNehtHPZ5KfrEkmiNESAYgggd
SZbrfBTwWdWLYKPDb85sgA6hYDH2Sm5cnOZ2TwUKnQMjccGL/tkfEFaEmEhfDDez
NbMqa0RfPJDGNFwvucwhy263Mt9Cuu82AGlCqw3KyXlu5Aeh43Axb+t+AUlCSxnB
uWE0xEQTbVuhyQkfnFPuoDboKmccZ3rTYdAZhm0Uw9exAOkyyWTrG1oRjQv5uBNI
4W3DTZ5YlK0tJPNCPvi1bY8g1X3gwLYs83vmJfkRCKWqj3fNFGbO6Mv0jiLIknAm
zjBEoKT5QDAd1fQLyD2cti9S0xr4xGCXAGjBLcKqrZW5+TOL1c8hE7SdlMR6eI5c
UAB86e2ByafdceKrrz1/GS4jXmK5gsGOn4VU7gfmdY431yHKbfcw8wqetQ1q2N2X
VGzBsQVsRSj1tvXqgpSNM8M0a3e2f8ZhGdhX84b2CPvjY9V+vmUT/VK4e16eZM3+
YvkU8TOVoWAk0f8V1AtEaUlHPTW24b/5+SUIreOV9X9qqsRfEOVegGHaYBEESQGZ
c12RkRnAIr1xFyHFULg6+/6WGzdW8DCdZitdjxDpOyZLF+5rTJ59+GRmvYt3ubE+
wGJBKakwn500qpTHpIjjmIzzHifVt71ByrslOECYUGqhxy8q1MaKoa7XYZT69ekJ
JFFeF3Jy3dfUeYyzqAXpZ9d6LQCNIdX19Ss2eCI7fGu7b51KZORlILUthEIrwBJk
8C3xjzBhAhmEPiMVevlf62oT1rASfv8tsbno9jPkV2UwrvuAdjRCoUN6u+f5RD5K
Zl8m6wZGXv7aUThJsugJNk3ksmg9LQTyG9Q7mQWaIYiTVtF/x8c2yZF2/x+8hM+f
bnI1joHaavkiTeEdJ32ENg83KYEt7zDJh6xwvZfw3hOhAMVRZg0/NDTPYc0o1VVf
2aU+P5ECl2IrmCs0r1ehw1JgXFxfpNjMtY0BYy3os4aZYJJGRq7pfohTj/h26mNP
/UotU4JjmFZG4X8CA5BhcwoJKqnITeW6Wjg18TQgvt44y+ekKK54KhyCAlxxCYLW
ARs6Ezd046WEaJZ5RfgvCl3NHsboPDH/d7ze0LELzrEea5GfieingPQzHO3xHCS7
6HYpFCaTUoDWXoMedylzBC/tYb05r+0UQTTa8UxcwoBJW6GSqRLsc1YbUBCnMJu4
hmK45Z3KL7rKfq0zMRfzou3SfPGqgrK6u6VXH9Z679pGIDZOivbIyIbug1gN4fd2
YFxxqbYTC+Srl0sfwiJgdKB2VaybOnemaNaEPJIKo4zUwTprDvPGufgDqPUF5jYA
c8dJt1xe6XjC7IdXkwbvOtxHOryp/6R/AYmEaLsJpw9RCFsr3tEYar57MroqA5cW
7wqi09t98OLkhz/lvBUjPq7yzJy83UPnp2eErIA3cgkUogvErNiAjXwWrZepJx0N
94xNxDG8DGNC6TWrxNeQSCfjiCd/laW1n4ED8z0I3U+2muynCqXTbE0DUBxYg8tU
uH3dGyGHr9ivUZYbusNDTOTggr6zMPzZQOP7hs2M5Mdobb5oo7TrE30o2RN/caBr
rn9f6CVqFmLX3yYeltBYIjQ5bt4yc6NyeHPzE3pRPOKGvINvwqPZIUNpG0CJeUHC
FHFTld6rqjNymht0hLIPBnrVSvjj0cHM4pTigvRsrRNqAUsWXQ+43eunhWk5mKFL
M8dY1wsJ46bGFSmHC0lvqsoXxWxBzA0A5+WJ6lF6N5KdzlAH3nmtcyE+i13GsyzL
zdzzGt2Sr3XhFp+GL1QuUXuDcue0PnALm3/Mmic4f69/raeuv6UjiEdxIY5FdIcV
E5oVH+IlcR84p6y9xZrx5rKET7VJSge8YU8LkQYUAMOvn8ov/hju5cWNSRhM6R7q
4rF3B0Poh3NQl2UmQZhG5HgMOebdDYZX01VlfHXPHcjuyBSgdRnFdG1a37LqUeUq
Va4jz8fjcthTi1WwWluRWmif0I7JxYhuL8UJFBJD3HTg8tLfxJjbbRh+h4VnsAt5
HhcS/C7DGOUogTkZ5EJ7Nqq7lixjc9YcMcifBOJ+rXKi3NfAb1/erdE2XW5fbxQk
JpedrKBoCYL1WfaGGC8hWnV2eAfhruc8l/PVWDR4Yy0yXzmUI6bhrrsoGb0Wb26K
uae1mTdrPQpOm9mZKrfTkJTx4R0VeCMFemQKJRLG1vCCeUSrbVccSLmeVAAn4uEh
FE6n6Z3B43vVunP6E3l2bcjv4IRFH07WVLRxZG+sjwUFtJEkFE/7LMcbnyziShx7
182rV9gahPRSmPzQiIztRDD+K7LTp/TUD/3q6GJbih0bnJO4TBA+HjFzVy27x9Gy
KwGsffvTP6AYeNuHJSwF85WCi+ilWtnh7AWgav24doKYwIvR+Q1H/LYsYp+h+1qJ
3XWm4gwy2JJx7CI+TJd3mwAZ3xlccs8inalWBKAYEM5RIDTZ67qFkzZ1Ata9dw6b
e4fJn4ig2Up3LwZeowjYJhNh9iTBNfZ75ycgnaSdECH2nyeCa3gfX8qxdi4s5nT+
N79TT8Tf/1vLmPLp0FEDU6j4DYxhWy9qv6tUI9aq8pGopYnJVZYpPTWSTkfL1zrB
qBkTHrxbf0i+8HxZplqbnRh07KRL126vBnqJSS16r7Js4hX7k9MdY38CppGEi8m+
KY5GC4uX1OQa7vVEo3R1qf61tsYqvcwTdtI9stHLNvtCrhIXRNeUFwMxfeN8GRBg
tHmLmI35KUgu4AahtqJdguZhwMv1q9snaavMOSFE/KFtltWz80n1RzFEM7Dolmz7
RcSvBZdZhtTpaBRm3FEV3mnAie7+50wfKStfEW3tWTYvTL9ubG+rYxhZZdlDIH81
nCQWe4KrvuDo1DFpur5wI7nmh2W4xIglQUFs2zamGjsc0BtEe585x8GJW7OqEgRk
AIIM3tjUFsEXFUVyzv8OQLjQ1h9X8dApPF87rnQ0VxAvU+1j/IPeY4lfaxUio388
PHA3cU2KBcxYtxGDUz7UI9cSAuxD7c6T5ssGqcD1A4jdnKzTvVgFwF26EvXvTuWy
t4JnWBjVn+oa1J1jCb4i8mvp0M1oU+ksViCOQ3gpIWA29M4xNw0Y0zHcl99qAoEi
Dp3pxpPtdIZ1Jc8aPh4Vc0oiKlqt2wPLrVYBxp+du5hy9OlvQsfbQZNaB0UeClXY
gcTpb8ewVPpHPA6HKsXAXJO8Gz1J4eyiiIZR7plEbT9NDdLUCLpcHN1urFAsS8o1
B1Ky6Vrv1PT7G0tfOgb3nob5NkOR19/aGFFTUztU+8vDYEEMaE+oBbPBtZqF2FHX
tZJ7wS+oo4VKeFaYOMjJWjK0MIIXoU3M6uFpXpQOLp/3qw9Y2u6KyUXvGO8Ye8Hm
4ll+er2cB+KX8QT4IY/IDKwpQPUmZEjkQ4K9/1CZU+jmb7mnQmkzeyVnFXGCrWxw
maqbJTuvrhydVKNBj/gjrxd3Q6oJYp2omCVHs7+7KTk3XTYUF8D3Y09J/tkTerV2
U1OUeaxlf2pllOLuOEBAoDmDxf11F3bbuCNR5SYXJqPg1MpF/FCVrWABT0Z8gN21
CFJkxnz7T8FpLNW96k5fyJxWHl5zXFwh3l4cILrK1eppiP7dib5CNmff9IpBUCUv
rZg0PJsjquIut/PSI08QiEyevQXOaOS0R21Nf1Un8Q9bBFlZjAaaiGI45TvHu7xr
0xsWkN342sdNQBKE4hR3uoQNNQTxsGdnjjIOW0Hx1ji2DcO90VaR8vUrxzX9PGqN
s+ms0c3N9t2I3WQbFBRoFrTR7cvhv/xij5kXKLu3+wiD/HLGNHfSbTG0wqefQ/aq
CVu7wPEVv9JEV8sjRiBnypLH2NoNkob2nEI33wM371KSSgOZBcoUNe5a/6PCR4JX
ULHS3Ig2acwDM2rN3Y0fdn0wMdsvtZ4uNEE6o/HrcP1IZpoWB68EpqJmwNSuwDQ7
HUCG3MiDFPwNCrZ3RFlVWpiWcloSgd7gQmpULPDCo4+Ir9saJXW5HBLqqokHGWDe
cg0r2Wmq5nhFewmQw1OtVfPr18bRZZ9IlQFw1xq4RdZb8JemA0XnAGqBEvpruCPI
egk5NXgE+MAz0Z+WqBRGy7P3YDMhqZz/irvnz5Ujfc1Dq6c7FjhvIUrcfop2Eawx
lFVXRbsJr5NuYcSKSs+vU/DAAy+0k//cxJOO+DxKtl4PIHHaq8XullvzXej0gB4S
h1rkmYoAZQh4FqcbWORabFxKHJQ+6PBaw9PKYmNV9eqiMVKvIEAjP0mKWsOnmbVT
tAmBfz14ce+TDRjhDOq/DFyW9SgTor1g7w4Tb9VrVCTJ9Fo88/LgK3MkGGvUVgQ/
iz5FM7Hzwyle+3+yfWwvUKfaWtP4WjQL89ZOuiMtLzLKuGWJ7zVrQPi5jSM+CE0S
NrwZfr7TE4wM2txyx9UAExO0B/bEkdAuybthXMO7lb5tLyBoszLW2Mp6+7vDQhOo
AZpKm6wX4V10nDnwGVI1CiD2SbD+YR4TPYMlkwj6W3LXont68rSbvYvgA93wJpXV
KCLfiyih2Ikj3qkeWlwZVAukLpvz15JC51y/goZa9kboBRiqzZNEE5O2KbEo0EKf
DoqWTX9iN6Wdv1M6QMYbGKD3gPya8DWF3lRDigdxby9t2h6UQ1FQgxUeAb8KOl1q
P3Sko606jhpGUQxUKYbwTtjvNa/ZjNuZ5ed3IHTWzrRlBS6v0Nnd5ymA/TO7XaQA
fTaKDevV5IL8y9Zov9yTgUBAuCCqdoLQ1WMbThBf13DLdFytohfm7LGC/xfMwrNi
FhF/c2FqOafbeHy8rEdTnLxceW2SWoxr3CMRQX+iezhPExWZGgyaEAg74Inp9/3M
3bblNCkdg55Yo08nsqk015xY/3D8m6s8ssBM4gv6JOMppkqSt2Jvm/CqTX2mvHzA
ufteSz+5PkYuTRlebFGqND+JV2Y1ZpmHYdiueaCxRiSYAROX+8r4J33+PlOTAOf+
SqeURcGAKin+S6nsn9Io4Fz5Y9v8AcpFrCq08LjZzV1Kba+z+c2AKDL3UP6LP7J6
q78hl5emHvzy431Wbe/pCbaj7C7DypBJGMRDYxEuQehZoPt6390CzJRW8Fac8QOR
BUlCr7fH6APraEW1Pp+u+vT95o8fQnNLTc3OOTYs54N8OmpIll+9pnx83vnI69WZ
DGrajS7gJqCaQtj3qW2NPhpUnlhbQSIzq3EMGgbqdnjtRtuHlPyQl3nlZIulYFGm
OOz52lXCQeM8k45L+uBcWZmYIExEc06AF0XNs9Uclys3/w8yCaVnM3z0NvSHnlp9
rEs3kI3s31j1I9VI8f4TxkWoozggAHnXQCl1mVgxeJZzF0kZ84uH0IRVCr20qvk4
3ks1hZHlfMRn3ulJdyn2NGm16/fMfBsj9Mx8Ve123adQlF7+i7zPoTeSICtGLNi5
y1xQI8ARpicsck0755Ksf3Rdt2TJhP4uEahbgkI8tG+QLzPFIoeOKMfeCnOF/dLQ
cz5aCyJK4jMAM6eLdvbhOxMe4tSi4GkmGxIVWEzyxbU6l4hKikvb+c21u87zv47Z
GXUHXuLCy1QKouFQhuYDdAZrDgVkZ/IX+XW3Khx1bWIKYD/FEHIK6QVQj7NnkUG/
0hS/VrFrHiVhgx+bU0kPiH/T5xCfZYCpyPDkgwyBFxEu1S9EBwcytw/SDPJowpVW
WwUHO6CrKsHSXPS5Wzz8cc84NdeWmRbh3Zt1+cmufTC9bLsrzBPlHn/ASUqmceOD
s4kpBv+U9nVL4yQDlcLhT8/SaumpnL30vvoxRXuHSF/52T2nFMq7SuVFtuFFVZOT
Qt4zRt0aDWW+v0/bAsJmZYXkNZPlMhqmvRx1XByDZReJJRGDWLBRrQU3jfytgS1I
9gHcBKJStKgJW1rQWfPdytrQg+xnUiwuSgitd7ccDb8PokpvcqFMctS+zKHlrU4V
mQvreDTUnbKUSFpsBnBESxi2IxepW4oxxnK31IwUXRO/bfP5mNdbshAna2mAU5Mj
kKX1WowfVPZOUsZFFMIsW7ga/IE3XWElGQFvbywny5dPSOpPsW4HXrfoTvC1SzX9
XAvPoG/R1XGVILpJ3kIpS4acELHqm+p4OBAnLOMoPe0MXOkUQNsW5eWW2NvnaUF8
aXUjrDxPHmlUi2Z9KhjqofCHuP2od4ZIHZRe/ZcCIu1r5k30XHXpv9I6XW1ANc2i
fOt0bNLQxpYugGG0RdMOqBArJFSyg4MEPbagKZuX25to1Z+uBr8ScVs7awvstEHD
FBmtTF99fbgFC/a9UKPvR82qNeLyn4bd3A9AhZAXOfr7HFqoJxhkHADTdY4Wjr2V
/Enr3iXqdIsEescPawsrEa20fDmne08GYqQbc83Jo43tW3g2Z+kqJQIj2qVu3zjy
/A3Fzud26Qp7LVMbJ3FHPQp1rluLWTzbzgpnVDrXBASM8BcctzaJwoxxQBZM8aJ/
icEgzPrSYDzM8c8Koau23I7OpH5nvFAKJKY+YLILRuoyF6cEYQwhZ4+s/pHbp4+Z
nzS0aX8h6nFTeZj85eoThNfG6MKiD1U8/Kl9dc0bGXIEYLt69tXqgKgDrJoKx3Gq
TmjKadOQ2fTIosMDcVgvz6kMqE1jabANkpqzrfrVSwhtDJzExF9+jq+TEKDhIgDL
8azdffBM675skjshW4GUD5+bwClfOtYqpRqbZ41O8aAWicu0GVr7GZYyTRDn6kwu
irtifn8cIj1PZj3kIf29Z473k6Y7UGbJ9CQpM8DIEdu6N3YVAvfwyNoVwe3sSrgY
iT/A+s4+svxjofdxnQSXpondj6q7iJXgR/Bkfga89r4hiwtwB5EVB3577LWkhpCl
9mxKruEJ5aLzn7d9ntlIErYdSsIYuwfmWcZCRIeD7Lw/WxVkS+fRZeU1xzY5s16z
pGJ32JujBnLn8eXkz6r9SmTxIsBHqFKlGWmsSVSs/Pez4HRYEnCskp/ThkssUNHi
TKREEzxMQxs7lrOO6Fs5VI2BqPkuGsCsBncSLYnIp+phH8Zytq4jFAqgN26/EWY6
Ae5jgdZQfWubNFz/Y9mZfaVp7iXduqUZ4yE+DYhrOdw9dPxmEQL8Q8meJjlenofl
gVuFyY8TQGTnnlTDUphK9Y3IXx8DyCRnb34glLjE49bi9Bdm8W8XrmWuWGUF4bfV
uU4iXScSTdUM8byAF06OO19VcecluRftEZn61ze9fvDCX9DBGqyZS59BZ2gz1FwJ
vnhSVO8p4uiNRhcIQim4h6l1GvZezr44LzSZVUtjocsG02KoaF8Y4Ct05NpG5C+U
tKaD5TJp52IExsjblhp2hZJP9gS8xlSlSUmIt8eyMp7V/S2yJHLybhLqbPuIapHr
wcJYw71w+sNM5TXU1IspfLdCTPMKqZQ775sVU0RCjhQYqDqFaUkJqkQRAY7qv33y
bfTpuSdtjUjNjtz82XF6Q5ont42Cn4R52oqSfv9Ov5HnlcTNSH5um5+CrxYPwv5Z
z+ZXvXY8Mmx9h6qMqCIJ0lrKTCkvwVukDMIRSI/pkv0vd8K5UxSEMM6aFnb+8Q7F
2l+FUqBHKoCinXmRRsmmfGzvPjTGxorw7lPPpzhN8x2lnEc9dxcFY38rvnRIV6bn
7k3Ci+PDwdSxRmFJhkvC5qDcV2hWA9OykFVRkv8fGLCDnOs4+vgBKzECbM/QJNvu
L2ovgmydQ8wdFm+IpN8kWA1tcyS8GchPDrYK3Hk0JCMPK5r4O4MfNrWykq7/1S0U
ikMrAjsmaM4t9QYKXbcewGJXwR6TmErBhVOEO9KfA/L+XvW9Y0rbY51+3oI6l1Z0
jTcQyPLYAfAd2XimDyaObL0q1/tObZKIs+4S7xQOUO5njAjYvxiTJU0QMnLWvVhy
G1Sy8PncsmWJlfcKqwnmyUKv8JC5ssQdJO4qHlmka3hg2dlXlGdo/b0Y4i3rgbIt
G0FPJgjctDXF0pK7n/hhxfHLRVjT7q0fURBQToicg1FRotE13FGjHEDzbw0Sabdf
0UrZ4SpOvSoV8rLVaB2gWDXXa2RDOSTyV/38fpCKM3zqW7c76qIauC1uAAcoR9pd
L6Dv/S52fPUWeKiWlu3laZdOatSnqA8hFw5y3vTrux6WyUhWdmdMFlqw/FFXV+j0
QSSvvbbiiOY4iIhkS67utASPj3pQCM8wDDeXLEmjEo/AHh2a8cSCgjpzIWGdaiC6
bcNOba44ofBdCttSe8wNgjSl6sioXYO6hNrPXGR7Y8XV3F3duMX5qleHcQB11wwP
WtSinde1Z2KKqaLtPPNPcXJaVJGYuGfxk7noGpGxaWaPGv/7M7eoE+70/qGs6pYO
WKSje9Fpnbsb+81Ww4Ft4Diq7tdcdosKlOL2zEYQkNytzCE+28iluG8nRvBhif5x
vzVF9cNBWicH9rSH9ZVzE4PvW4D8VIQAWkGvD3h5mGCitrjJvJ7MkbonokgemsgN
KXvSc3g0gnUwgYb3BaUjD6Jltgm7ZCGxOm8qu6xdNkrQzNgXn9/O7URaVynjDUfo
MFw7iQ1zmnXHcDJjA/2KFPQjVfueV8sMhEyW5Tv4qHrjGvDLPLg/xW8mFtNHD+sN
AOz2hdjztXvT/Z+z58A9jFd3aIzng91fIEA5LH5XNBJc5F6IaJtjlM9iZwRxMQac
Aa5ZMPdAuNh46FzOzBAF2GEx0LdKxKQF0OXuYLemhqMDOUWGhf0NNNvzwLFO6sGR
dkK1janh9uw5WLh7zbo03R/f5jIMuoNsVlsi1elF7ykMTdNFKIgPCM/F3AkglsJ2
/0CxrfN/UN2UAzp2ftNGOi2v9oPCtzncrh2+tjCRiofuI7JKLBzHiShkIVOEe5k3
AeE5S9uXEV7JyvQeVDzdeoRZYGYWivwfH+n0qvy5hZqmJSxqMyCyte5YCIGrFhp3
Szi6XfTvXzJ3lfvIhHR8DpJvDvA5Q38w2k84nDOUIj7Hzgqm1N+Vff+vZRvcvXZk
wmfYrNNsqBcnmwavtnodTKLnhBpUaITGT7VnH4EG7koT/xiLFKtUuGAUMT5KWxFF
bTOLD/cukOmC2k7cHPi/lOUSnY9C9wZ1FXecwWSvnTGI2n4SCo3VtV7AMzpD6MRv
eSs5qmJmE0XH7m7iLpiQqqiN5Dv4K0VUsV0IJnFvf77jsufvIUr/dK2JbNpCAY2p
B699w6aVYnIGe0bpAKHHYJc0NYS7Xs6+FJxgyiLML0/Tbs9K/RDREoapR92B7k14
oCCxJcCakFVJLNqHtG9IgymnJsP5wsACt/SaaZrwbuj0KLCGRT6XYSfTnyqypmDE
bYMWXZek3O7zw02bgeHAUyKBlMiqAp75JiDOtz3/sfmAK8HP1OrzoAG3jiKuuPZi
7kWR58ZFyXWmguIqlhzN795n9fIM2r5bErFs0RqU4axlhzTyf03/+s1GCpYgwNkO
hQU/ZC6j7nWXNGFGtMyVI/k/mIa3lf+HHwGa2B08Z7guVR8OVB5s+/XS3aBWA6Hr
fcwBdNOCWdYfY5TMNcMIQ+wktyvnvqkPHHEhqrrWMlNSw4/C/uvqSwBs1i6ZfLje
Gq98CFM4XDx8nsHi5TSIER5iYbhbw9Ak0ccJ1/C3MHtxwiE4/GIFtQBIDqmEeZcQ
hegqIPmD32r279iW3RtZH/lQYIiias7D2p2FdmcYKAsfcCjZgkv0N2Wah0LVSuLm
SKU/eLDVXyD18NByiAqS+Vknb2NApdyiz2YaZGPjas01L3DmE+Y/4iWxZg5QxGwc
D5JYaPepNN9Hsmg4Wtc5t13GCh7/bjqOj4qrajUoOhiFscrlWte4ufWvj5oxueTe
4nsp/XGhZX3KBlpM8I1KKowpHX+1Ug/XRHjV3KcX4AZoG2K15LAqZraNlH/iz2uq
7Yhe6qIM8q3bO5ghZaBGSR88lPxUjG2vxdbgoN3saPcUTW8p2gUIZCz8S9wJIEtQ
P/0jNBnQkKbd4IlikVJoSMmwkqAHPp6yxQK4xAiY80Oa28UZjmYtfUWDlhy+l8+V
51p8/TfHKKsJbr8VbBM/xT5Z90cyi+8mXQjtkwY5Tc93SFqin4i8Sk13ajfVapb1
aEKp7hMnutPqOWi+HDJs+QI/5T0f2ti6TOzWIzipYmKDLrizq5MfKwvPVRnpCo9n
iwRDhwMrApgDzNILQxAnFTiJP7bUrA9wFMKTZTrxReJtgd4fL05lhh9w7XteuqWk
63i5t4VTdh3O/0ni4fBSSMutvsEMJr/i8OOR5XNMCWo3CdO4mSKeYgEGMT5ZsS2R
tuZkANVa/Nox5ovU5poQaYKQ56pYCUFHH+m6qrDJ1UwmEpLj8qdzmvkgkjgjtQWk
109yl6aiD9URrjC5NMQ0L8IJcgBJL/EQO4cGzXH5z9jmZpX1kDgDkeR//NYJhmvp
IigCzm75TjnSN3/KTZDyp2G9THf+qMnoz3OkiAPVYc5Sceufvxu+uHHBw4fASeA3
nVRYYKoHz0UWOClW5Mc6jg==
`protect END_PROTECTED
