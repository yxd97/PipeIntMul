`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jbYW1/61Ox3D0DCeyHIYBT8jPAfwQ7L7fgvB3ZEjabjGS2Orae/s6TJrtBMoQtuH
O44aMkDPviheex0R9hNNxyYtAePk7zSx9NeTnKlsbGQMweisRRmzuCoWliGfqhwL
YYZGyayOzoZGrCMyCevy5Vr3MH/r5syGPxCgE0m+cn0ye8x1IJnYlMGkFSWZj/bn
rjQueeNxVJKlFbBqyTxZPhppsmLzmZ6dIWklZUs22Z45co6C28ZJ74w9DsrtrQG4
CFo5pzFUVaA6Zkj2q3qU9eaINUSRkC06NZc/c8PChCNaVul9dlCTBuuxC5/7FSZZ
xnvNiER0rrvUc0VQC7+wTS/zqBJSnWlKMii7KV0jmDzL7n3YQqLgVzYqQfW6HAws
j2TQfAuzm4r9N8OGHWCFh05PU1NfuwaY1wBMbESaiT8oH8RcfTzji6hB7yHU7p+r
t5Z/bWNqRlovUsqvcO3F5kUTRO63Qgm6WS7CkOwShcI4/BwhrRf0CTmKbHRvB5+i
1svvj7LJ5Ndw+qMSfFCqJ8OXK3tiExARyfvWhpBTOdWa8Cdyk5EnNPPijC7hOyO2
MeIl6r+WY/itS8Tz+TIq0XPajsasQzrhR3UgHg1ZdNR0izuZ9M+BlibgA0JTd2rL
dkk/QXc00gQ1UMAenWbO+A==
`protect END_PROTECTED
