`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQQSscp6s+R0QIcuEWMaToPoJJ8T/QwFKbG7uksTp+jW+f26ykt1RWckU8pGFDG9
lofWr3NSPbEcO2+LyqkR0+ARiiCpoT8Z1ES1F17fZsJofoMLhonVnYD5qUzMWnVr
tTrjaZsPeYtnrmPLdBXn6PYhVg4GzxBQGQ3TgaGHmLjGmmq7Xf4o6ix46tgAf28+
gZ230k+sJ93OmH0nGzjaAbg2IJQ7FkjG5IHqhiU0KMsD7IJW0rrHCZYEYO+L6N3Z
07vkyvAVLyjJBcMCtOMZyWvKs1kAjuJkKSWQ39kO9BLWe74wZhubNSOtPA8CEY7D
MgImcRrcgGubQZ0kRy9klRhZPRcisyhekETeqwBZr+97ytPqDVlaIzapM9me+ts0
m/d3Lf4IZ/3wGLpg3znCW5ksy2qCI3WBmw3fxKXa4gN/yWty6Cls73T46W/X7feW
7rkpaB2DPAPdsP8IdK8DQryeWMnEYM2bR0ROfAQrNjZS3ppOzWMSoYqbcaxZTV5f
p9bi6Nbw8KITKpQjIgwTSwT8s/SVLn8ER01IQzPacYl4xXtwVxSf5jQNfyZt5Qr1
HS6sIni8FYF004Ems0HmElfh3zGr+dpxlL6D5B5gvBM4No6TbIp3MrL8MbZfK2Ko
densgVZszAF5W91vQMF6Li4ufR4RDlCvb7ORftISGnSAE0Oox+p8d90g8PyrekMJ
yBP4NekpDLiFm8EKKlvVpjAMeqV+n15C0omAcfwih64UhXFzdoDa+NkZCvEE8sEx
JDN0kRNgGJGJXEA+h/3pLX5O9g9Qw37KueQ03QXgZl/m19lkFBqRPIzEQy+7YSm3
vUOaFlq10MLnFJzcx/Kk1ncWkJiDQrmgb/H64VdHdVFMvkl89NbKDcIiosKsqheS
kI6iIvSEDAnCmqNQKXMHTh3exx+VFh2lB29eG3dc4dpspFQUpuI7qLWtESB16Tay
yENMbpMiRh2qU+xp9SqNk2CJmFpLPTOeaWM9r0MytDJMlmwjE57wS617xN2iWY8i
VhEfRo8fVJYNpOzfUn4v+t9TFWv6Bem0fj5YvuSeikdiJtdNRTGcCkrpCvx4wPYB
2SREpO8PaS2gpx/ubsLb7T/PmEML54bQej4VSouea1eaihuLZg5eAcFUky1uTC30
YJ3CZYiiBPsG9JfYfDMlcHc52SOfUoKlxNbIW4tMbIsPsB6MernMpGmWyRecQQZt
hhpEPYwN4hXQCQy08mKhwhHjNiXe7TZXJQj5z/TKu2CCeQ8vOwZ+lDlIiobRLxAg
XRsmYiNMWWnp14+39JjVxP5VyTMJtIzsbmWrc9boc7C6YcrmVJmajiVqMf08tBGo
9uT5+eg6c7ZQ9LyhMj7WxHrdmKvhhlID9DB79IdthJMzXyx+izPSU04wL5LQOcH8
T7BOULd5V4DHxXib/Yr9ZazFcrN4YvLDc8pSl7ByJJAeMjYv/FNOEu2Vcg6Njliz
GzRK1iWjowUpMmDx8NgaZ3jsS+fbAbVItFc/pxpeW4WA0JypTGdI9uucf2u7briC
gxsbTrBRgTuoJ6dw8ve8rW+150t44vjxnsK9lIKADdXPq2nQALcf3kUYHmEZfOv8
AA62ytlwrSFJbBuZ69PuDr03dxIyBHJmvkM1WuhSpTgWjyPP7+XunDTuSFESERDJ
JQgRzVPF6DqKO0yy75Mv5kBYnjcvkrji+djOIcaUHjc3RQYFwKzuaz7lph/6Qyhl
viVfrjI2Xoq5QyvXZFsikldpV+Svmp3PVrL9rAN55PkImaf2ee+tMBTX6d3LGWyH
e0Ol2HoB/VnFCZWdBaMkjaxrimq1BMLuNbJw+bECOmV6OBvaksWqVkmAVTUsVlvd
Y9dHONq5TSblN/rdrYZVlKHtT85Zu3qWtc4y0laWarRTvXdrb9aWI34WaIBB5ZyS
S3emG16OkRt0NPSH8ER2SKhEdwIA94w9oMCBWUBXEjWa+kLm1gsiLd2DNcQfrgig
ae44o41pC+BfLkQU6fVOgGyTGqU5Y6ubPrg9NyZDcxXdFjsMzyos2FaVWbokn8Zc
Q96lsf4vwPxz0C9nKf6ughvcAQd6fZvVQCvFH0BerbhKbDVsd9d0ohG6Ju0dcCzv
adTdpmqYMas1lPV2vvO1gfDjx/CVDbehJ0u2RwdZRrUYwIKRUnu13Crz5gxneh5Z
aSRmjb85W6unP1spl1INGPGF54KSgHBciljKJqqFMgr9SDG51um1WbvaxVzOYRR9
zn0zc6w1p0op5oKAr9mDz/ETDSt6wnwlIzd/0uy5F4uRu2k7sLfrgWuoqTX/8C2U
R9rl9KO6KZNrKwFAS5CxErSBPzjyNWz5twkISQO25fw9AdJjhDlEuUL9I0u7E1by
`protect END_PROTECTED
