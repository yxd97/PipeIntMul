`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OXfYt2vcMHVtn7Z1aNmocsQ2v4sZjpmldB+/7A2/BEzElrs8yseLmIOw/EMW2ePt
4MxM1FBJUDyknsFYvQFOu+1sAnUt0x2a+8Ei9+rRiT+9jAczvxtvOlDB5ECoNZzz
srLbSWCpuj3jAoWggztoyMKIPNUGQzaOhqGQwFf82+nqnOknVOONZOfVGM3E91wq
4pgJ/EwAklJqLUfF5Hi8EyYDBu/rT+/XhHt0sUh2fV6KZlNMIEZgGa8Ok9kYnmob
WRz9i/qRotSWJgw+MlfNrclGU0p9R+29fb9V4xObM1j0cONkE4cHH5xfZFA8z23H
BV+Ryj4BQ3tfrvP2e++f/Lra5wvG/bZq69TAv7pDcveTXoWk0jqTwJXbjNre3+oe
6esPDd5k2T50npVOqDTrYqDHoDsdjRbQjo6GMiwVVW5c/doXI6ln4U8p/AZdrJp+
ANGPMFT5wITquFw9fvcQJg==
`protect END_PROTECTED
