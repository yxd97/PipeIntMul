`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5ZFEERNlUjdCgk2lRbyoIHqvjFVktFjN4E4eEsVdIYGQl3BCP67YNYx5P6gAbIA
sa11JXkL7tVDSKCPWH80YeXV0KjRbYCRs4WoM7DIzTnjzIJodDGViX0+OqsFHq4A
hI0EirEW2o43UbWiNNEkydseOxX2E8lt88JBJoYC52KBMYj0CLMVYiYVvpkpSIlm
+wN7hYZFZS4GmlpWXqMEiF6qqna21hMxswJS/sD2kR8KIr7xTEN47bEsQR6T1/F8
k0qiHps1n4vPw4heX4KXZmWyTfheemThuXY/An4Wmavgiy0qe/opEKDlGBAT6Hvm
3Z7iI4A+I+GSAk3ZJyMuOgEuLUBuLvj0LWtrDVHlf/y2Fzfa2u3Ejbrmj8MViGy6
4CbZCFwmCt3SrjXuvQLgOnBTxbA7izorMbTYOqH6nHQ=
`protect END_PROTECTED
