`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1d+KLdXW2R98dC87D+XMT3RnpEHKbaR7kvQTtGv+iExixzU0ioVZlhffi9MWV9rR
3iAcu0fIEQ/2u5HxVhYONnQVrBG/CMu/z4eFm+wjhAfN+HmsSkjfVeA0kxGLCV6e
J4IUzx0N1mTWA7D2AL0augEeQmh4iaQI0E9kUtTV2JhhjfeB5tuAIBjbKF66PY1B
U/S8Jz9iRY4iEHOIHiDMRyLTgurNm+zbiDZ1IpMDRKpZ05DgiND3lpd0IY2L1mKs
1hYW3r8gCcjbHSzSh9LP/JquwU7/xoAsenPLcHpm9G7+IapDHkM0xCcGqM56lxcB
xfMHnLAfcqebbz/bccDOajiaXO3XaeuUw/qLS3AEnA0eZIA76PZcegDncTDle7pZ
dB/f2RLOIkvhfGat2aFJsM9WJ1g+YC0/YuVX1AChhpHKVQ+eDMw6lOC5RcaXx5h8
PiiBIjScrCZmH+ltMsLyDmcELIA08NcY6/xJtXDuY54O9qV6nANC5EsIt20SLUqk
KP23l36zSjoShJ4A2SZb8UZ51ni/YiEObof9kNJUWAh4sGN/KKyl4ln+3xh2iHG/
yyVk4QJu3S+EXV0FFvAsR3TJTCLFcwtd7MVQe2nxXLmOi0kO7pIDBLAm9mA4qTNX
JFdUekfwD8BSHIetodsy91APDJpCjpviOtUJ4TY+bv26XogJxkxmPJfG9ZbfuTkL
GkIUQ8VlO3fFJ0uw4jw00sCeDLXxQ0sold17/Em0PXaJ8U6Ote6Xcg+4uYoHC2pl
HS+V00UMAittOTwUIq9prbhGYHw5gizRAomUNfQJuVHDdLwvi/UdEp+5Jw+a8i9E
SYFwFqNzBolmZxxh74TUrbKgpmAZw7nh/FNJOroqShSF1yVJix/vu2I8EmXjmaGP
/q+UbkiCWcTbd8E5mg1R/BDdhecUbz1JU1gR/Jsun7A=
`protect END_PROTECTED
