`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VRI9Fs4cN7KmS4vEJ5g8y2Yl0EqJigi8L1lUKPYPXJROWjLmsmR8M520+2A3PJof
EPOO/bvTSTo9NQ1kcSFFB6JmNPmHnU5hv1zycKsUOnOwueiKy9TjOel/DUWnGkIl
BKt2kmSgCWpN86un5RGw/MG/H49Wr6VqTXZpIRVV+DNm0MA4omM34OPh1J928hBU
RCDeJOmD0cgzVS5Ew/zgF3321TzZ+lxlgKehBmwzKbDrC23cSfRNg46yRo64Io/F
qkQp/h+Id5TdTKIpxteIMs1JH4eGRlFJ0T9Vq1qRoTZ4/rBDIT5VyGfyef6DQrke
DWmoJH2hE+zl504/Ar4b3+yro2Z8zBA4ulmir3VDGLzMPE8+oBFanqcgzG4PZ8hI
3Gk0ZSCt16HRL3P8MiMnSGCzbs2t5J0C7k3RsoUIrjlrkF3I7Y7VEHozuZoxNU8v
DqJBpSnTMbpaehR0BpVbaqddvIA1cecS3ao+XTgRvK/YOKDLVFkihxRXUzLc5d8R
5FIeAabN6hpM0GtyHYL5nCtfuTsC6XbF4vKWXk6njEHHea4EkRIiZlj+YpgkwLAr
uKorWXbWYmkCMzqZnS6U1rmh99HhYXAt2JQYa2DYTzYStgIz81LFWujs/1ICXUeU
DuYrRvs+MSM7EwkFzMV9Eh7mALCaf19pfMt/CGxxGLHgfjVVxpDi77xOT/TXtnnb
+kdozBh3oY6h+RYEmax+/gz8OkklYVJ7Zhr3rC+O0MItVolDwjnRixAQHNhaVBU3
eFlhA6cwUmyaeatFSYvP9Q==
`protect END_PROTECTED
