`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqoUaZ/e/hvIH/YG4b42wTBqEO8GiBUWH3vR3OAy4dq+zwNP6ONHbCP1a+xaKRPZ
Myl+sTtrUtPsQ3HDoD/BgozRyMZgeD7NQ1Jw5PdcydaxYk2OC0IsYYOQPZLrUi8t
9W3hzqlxlaQdnQ72PPgIvkEw+TEra+gV7mHT2bdleTIQZOIt4r4bWi2O8QwQoH0s
Hc/rTRCBVEuVbj0qzokPwLn9nfbwOs2iZCiJT/LH9rqy++yq5jG+SDktDNx2q9XP
B/Gnce5Q5bD+4hohZ2maHpR3tzjBurU8FfDF5c86HUmcgxGJC7VrZ0p29DEPjU1z
pQ67Rd4x2zku7dsiPHChZAAQ8mAKFwOuQ/4A8+VLBJrh3AkrJzLKqMFAzJz6ltWa
DTu6OpBhI1leBzKgXaBwD0UpqideApOPdxvm/GR76Go4Pt8+cR6Ls5FCqIDN8eRP
Cs5Loq8AJy3KDJUe17Q4H+5xiCL/e898l/HqpSkcsf9I4nQsYO0VUUKI1AMcmQ04
lWA7v4q355+zSCKIESWejqv/3KzW6FBygQNLZR7p+HU8BFT5qnbqHUiZyxtx8XYk
Lf89422R/eZcvKqFegNjE18GfInxe/JQkB7StmjSjozpCKe8zHc8N4cdN8EcVkp+
Hjrz4KroG6ZesNDMCpyrmps2llGgH8pPQLEIa5+BooJ/5wkkd7DBi8iNqdYhfAxP
o9GBjhT2IWavrsb8fOb0RWOvpIrHMCfvOO4A1YmS0pnE6MuHBUsDcZHK6CFqvejp
P150F9UQA/R7r/+8F+pHp5wR9578Kz2gDw6SLz/8YwsZ34oG0T+wHhMefpByx9Bz
s+8w0ZmvGBsyIv8mYcbLPa1vnjHIujDsPbPWiC5AmPOMRzeGr3ew9wIK2aqnEZ4D
wa8IPCj6j8y8Ra77gQVGWmog8Q8WZ1U1qRk27ulU+PCQZwB1DlUZa2RZTiw/Js7G
ExJKGgPL2WXWT2gntxQG2nOrhjHzciU/uWe6oW4jUK+6mtOQkadHc9EzSR9OY+gm
Jnz9gpE7+VxKUtaVu8m+a8yQtMc1yJj3RuEMUcaxWEaZfnqP07PvDw3ikNITNQoL
Pvl0sCJOmQQy0gHbzB9QX95POuinzWIRYrXQIid6b8XZX2LgioG2fDYwTTgR0vm0
H9jaeZ3JruwLd1Ug3zuxPRdIBR9wzwxbQo/WKUDSTIE=
`protect END_PROTECTED
