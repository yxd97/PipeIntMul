`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zWKVMu5Je+vNein7Ua4rE/ASMyRDupwTJmTzujVjsGbAZn01uPSL7FD7XUdnTmtz
084IKzVlQO+IZouz5G/gk+3wMKt3bfmX1SQTQAmeD1jvEAnYeh4ZlEFnhyCFcIKD
O5hutWgcbuKQXRxG9/GGjrGl9MtS9iYxmoxCdcIyI0tvDHUjAKnZpAVZQ2yndKhn
tPQ5hmSUIqsGp6GEwaBNjQBB8Uojy36m5+rYySazze54kZSOE7/U4lzFSBWTofn5
WFPAX5WP7MneOho88ipsz5I5wCzPKOoHxbNMPa6jrZ/8zVdtpPojCRblDMUdB6xG
9w06c32CBwV4pE26Lw8yIbXF7YbXTazAmN7GktiwSk1EA6eJWDu3axsbn20s/NmR
fusSmeq66XhGCXhNfZbnFA8LkoqVeIFDhKCLVPqGPCYj5xu54sxy6sFEqVPHyCTe
X6V0E88V2Pgp+oB9b9UFX5ntokeo4mEcIUwyT5ZXZaSy6+XLZ67Y58x/K1o1WYaN
KdzXadTUZ7SoeMRXyH4sdKQVsVya/0KddbB9zPBpO6zRDIo1dcjJupGaCmsZ3i5S
Qzq5bTsakBTA6i1a2o0hSL2XpFVrWORHSIsIxSmV/Oxw9qMRsZaA1uYslylGuD4b
iS6fsoUbBRV+RkmHpnylPb7rIfs6gPtG9wDgIkHvOczaNikjsIn8UMXC/8YFtHmL
Mp1VDBVE0116HLi6FOHSo5SaAojTLxNOiRGRAMp5Hp/nu8rGavzKTaHi7vRcTeWz
`protect END_PROTECTED
