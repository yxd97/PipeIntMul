`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gy2xBk+GJZ7yfHV8X3oqaTbgwRLLcas3rFV7LU8GZ82NL1BmX4AkRId76E1b5KM4
tmJKxTSCQkscP25y0sXlc7MaymlbX5LQ6uST5JWSbxFT47TOQvsKetK7riOS2PAE
v+gd+GrBDrEKDGdfn8jcwPt2uqeQxLAWhg84y1qJyRDG8uO5puYb6G39NfOAjcqW
Km8b53atjTvtmjf6zSJkBShcwGRFXNloEpGLEWhr0k24591+GGRgWF65xw+DSzvL
BHTiqlvAiwnQQ6rq2Dr87R70rATJXmvIXs7azx52fkH2V26/ZkD+zSEjsZvC6dic
230i3A3WJ/35dNnGNnPrXbFP+C1k80zBX3Y7Dmf9MYlfUDBf1FOVBZQ+6tg9vk8i
HyopI6oDi80vSp9bICewPEHPdvDnpvIgo76Z6ePrD0y+bnqtGgfcejK8E/j6ai/T
5X3nCSMT2BKZhlU9pq1G13bGLCllM+EIYDQ8LkayYDW7qdbw51NPif94+KP96EDB
pYBiLEd3yQVQhG7mFvc8Nw==
`protect END_PROTECTED
