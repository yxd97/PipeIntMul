`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/Q7jung363VnVAZwNb4foaho7ddzPfHNCqmItEdno7Ri0OxhJyS/UZGRQcenUbU
5JxY90w9giqJ/tAyOhuJwE+eVbTuv9N4aYkdq8n0hZ3PGN6zRyGpsWkvhu50l2K6
Pa3Q8lQX66txp3cWGp1gPZY3g+WkbsRmLJswogfiZsLwaZmrxHhupldhE1DQTOAr
qzfvZovxDVCf4ZM5vOpYkRNaP/8ugN8NoS2H8xn/D4gNwnGnlxoMXQXa7GLuKio5
8mfmwVV9rsdzBfIpV6lpgT/fcK2HDJJNrsn4xJXHfsJ4c14CfIqevNSZ3zZg6PAb
WmMPYAg1/KGauOjPpU8XWmLoOepBpijOitPKnD3IWTEJXXgpwMTWX06ytz89f+hA
6YfmO+JBBk0whFWozEvrP3IvEPFfL96inCkFsAFGMhp6fPemfDFN1ZJT7YSspgOg
W5gCuE7urxCiCmlHtx72d0XtUWRKqZuZHFADWTreqBbQSlyjniQufgXLDP8xN8L3
MundskFJIEJlAdSxfZqfDXRKtrIQKhUnA59zQbazKcjEm1Sf28tyYAYGdngXMMDc
BYLywwmgn9XS9jrq62Gx89vFrTW8B4pt1yvvgBiyoztbOGVSRJ2QazdsBwbd2E2a
1J2ynfP8/elseBTYIjU2XliqDzhzWYF+DLcdG5EuP9jcbED3juMXc6JQ8Hovop5M
7X3p5elFtCfYr7zEkN3S9HTkSjCdgsEishtVMKSFzWDQ6KkLT2I5GvTVN0Mqh2EM
Cezc/hJYCPFKvfTe/+F0rw8AvDIG013Kx1blJaCTegfbdFN1nlNJbQXb6fn3bB5b
3xL2gUlJUFmloQ+NAZLd6d7rW2kpOhqJuGnzerYrEleQj/r+TZQJGMFCZCWbjB9Q
H+aIJOQbiGcwG6vTWuUTxlueGrT6cxjCkHA/5cKmsdIJuGKo1aRbu1mP+BRUT+Wg
TKdAocl/Mz/2ztqWGdPtq2K83X4ja54t2+dZvw97sccAbUl8HvBMEfoy6vx7HLvN
vIriL2s8cq8br1rHXGn4PQEGONnOx7WgUBz56cbl7D2x0lA/7GP4NW//+FDq2Xrt
r6AQIPVwBAYNzuYBfsu+EXUNzQn5E7T10HQxe0l4Qs/rKW+oPQVZnntw7gN/hQTB
reGbTlyUGafUHY8SQyfqFQaRFUJKoRxgBX7Z+PfdHJKLo00JCZtavLrviY1sk/eP
kzwM8+mQOLahRocA/+/c8CE8s9vTo0Q2pi9Qu3CwjcWE6EnRLIzd4FBJPnPj5DH8
ib+4I6Kas+JVlovbc5Ty/ZENA8fqWsacPwJJFODsuWgUmVa7InqKrh6dAnSqnUxl
mgDPcs8Vo7iMeNp8gNmsqQx6r5r7219Nh1fZxGGBsQu3NqvCXIVxAmN0f0ygj7D2
cmOlj3p+5PQ9pmRB9Kt+HUq4j7fjeyU+47uX2JqZkmBmwxLtW2sgfnuKmQWViWeL
cyoliUp6p1UVX+Dy44CsIWqvoK4JDnIsbd9a4JHzbkXiCoLnaF8A7xsoRK2hHS0t
N506eE09/WwqtC0eCCwK7nJ2RqXl0IgFHc0VQGntMht1pgy9C73lBC8Tz2uYZpok
BwYWWQ7gJe50Gc/iymTc/y6HFSdsuTO5o6iEpWmRodQzU5ZnEkv6R2AwxEurD4dd
ff7ry1tOFwCnfI8baMIMktyTG960Mk7a/zpAYWnAYleCCeMxqZjaWNEOcB9SdFUQ
4hUQOv6E3KofiRw/1oLAXmZfpGhN1HE8VFZRmj7YNpBXoEUxbSO2g7XOnD9lhNAT
rD4+NAN63MBRcz7EJ8cHVhe8KiN5ydwh+wWHVKJgko/3QQJUJxVwCZm2XZPh7EXd
Wjsmex4Pn/508xGfI/eWgm2bOjXCMGCnR14qD/g4ysP+n+3JRMcl5xEsZ/PnYyRr
d3PidwjvVBmN1igbF5DLyJlH4M0P+XtVbnxah5h4Skqu1O+WFSL+AjxTbVDIwEyt
xuhV0Oo/a3TAsdYZRMi3xM9acg3mgcqjo7z9l0ai0bxq1T3CZQIzLPqy1j0RPpf3
S8TWxeSC/BxWx8FKAPmnjSEdx7Scrq00Ot0bvttivbtUemf+tN5bZZvkyB/ktI7Y
h0sD/gm6cIZj+Km4CDgu5x43npEwEEffEOd6BsRHFdMdQ7TMGfzL6QifIRTjQUfk
x8nVb72aagrSAgXEWos8TxNE15WceVHEgerrs5QrcFLS82+OH7S3d6CXB4xiCuNe
15EXkkqp5fN0xbw1VvjqaOfgPobBRTvSprgv2vJdSGcdFKHq4QIuq1Um6cr0mSnR
`protect END_PROTECTED
