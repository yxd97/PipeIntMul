`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
14fL3PlQM1sZDsiWLeDpcsEj8FW9FlTuk/TvC8efn64FjYSQyi86akFPZ2ZSepGp
NyX4KiMJp2RynrbZ0A1DDskm8ywB9Y1lFzoY2TNh2mtVfsAv1qasSMQ115PNxM5Z
vYz45PKzkASlIjiPiX/ojHUcaiCSBIphvFSGGUxvIJNCkTx04yobtS1KDXZ1pjqy
vEbk1DSbE+9UTBB86YMxRLOLC3ZGgKpWEh/+c/QKc7MKYIrFjgegHPu6teiejAlG
9Y+AYMXKjeWHowH1uHWQ5h8V+DR6e0cQYQU+xf+LmITTK0CRQ1railluIWonoSIP
Fcyi3tx7la+0Ivn2NuKt0Difo6F4mWblYeoJB+EeNZPRZ6fIwMn+YgqhJJn/K1FM
s/pw20yU/XYTvOOMxFmdxDIw1RO58A4evRsSocj3BLYhiWiE2v2Rk4IIUPLzCNXd
89moIZEWvIkB6Arf8dW0KRSq/xAtoU8MQrmuAIg7AAVfRibPmXz6OS7nLLMWhU1g
Hkxi2ZWWN+Xh/ApPlctICHdm7V2FyvL1PVLLMusf3WKe8NbIhFuG3xhwl28lrv5I
ljn1ZAenzoVoUtWaRpABiytoqAZHIJJyLB8tCjuaL7MtmAVSrkmJEcI5hYpydBMj
6Kvhpcst/pAIPEoxQOs/8Lj8L91/SlYtsl/RSkCdD996E2uwC/WBQ8VDlXukywIL
U0XnCatsaHIUxuU84fE6hs0WUxsSe8p1B/APyb5mSE5DtGvNVkgjLW6f9r9e4Gj9
g8oqQmiTosob3IBcxUtqgrVyQ0ctF+Nn9ZiF6gNsNs9lsQ0+qHC32DCup5Ir42Rz
u+nniMBDzCnrwFZjAD93MuYXvFgvCQzNH+t/uADukfIZ7fxIrg0gNMA8dYrLvPC+
E7aOr0320d9k2yX0FfwdT/ZvZFbkTT+9igHdUkvj2msqE+0ubu7uNtTq+oqC/Jm1
tKJO6snL1A8C+Cpke8rof3ox0z/UBhHL7hU2pnSMJ2ST6JstDOQ/qwxH8ftbNOOR
JRzsGjNdi+wMCxrACQ50J0QZ47DiQ3AulRCnJfwD0d7umoNiSz+sWMpDqppkRJOq
EcVFrD+ZLGHBnqWWuJ7yfEbLzpwmJ/SxJrlBw9PcOwNSjBz/K56Zj6NQNjcrk7RU
OSwbUwtS/7Av6gBOWwkvc/9VEYih7f0vpBUSA8MAFVAMYIaqhyui4/d7m0o2q/FL
JciQPXURcsXCfepvtaYqR+p0FO3WqVxoGDN4ypt6nr6C/wh+3qGKFLPXwweOqbeN
ZOPblNVzXcFh8fMm8rw85cvkypWbr68ifC6Gdb4sDA6Hw7GvxEYPAQvDYtFNqnDl
KhP4vrlDRg6uxy6EJna+1hpO0jTJ2Jej9On50HatjHha/zE8nGrysB96TUTXDown
KOVx+ys9NpyOpYNWrvAh59lP4WGGTpzhH3AtC221QSx+yXTonWac5arCtFFHGgNu
DjhD0CZtiGbWnyX1KEeRxRtLUdYAXM9AoNyBLWnmLV3CwDUqmQUWawyua2MrJ8ec
pn+qF3XuqT+utrtUs0r+iTOsz7JQOFLxTLnNl0gnKG6yApw9L4UsdqkxvD/Zfdor
428FwiBehveKJJ3WAR7yVYc65gRJNvtH4X80pdI3Ek2+mcrgYEnVZvCU+7JrPCXX
hmyxcQHrJ7GWoQl/fTM7Sf60FioRk79IIsnhzNv79Nb+P+JiqoRaS4cdz/Dk/910
yC0FNvBun84kq2LDGBYsC5ryxPuzDsS2yfGntAxnqUTv47Yrshsybtg5lnr34ozc
RAIh1pwN/BAJQsbT/5012K1PzJxUd/83+5+rAU30SLhWqqRbUnsH+L8byPQGm3gK
I2kMia2j0Akp3V4iGe1m8vOfEjyqxIqx7w+1ggd6lUcNm3xh4qc85xbAj0tYjFNt
KWqiX2UtmNx/oFKszTwMntK8RVWIUTPwjn2x6+StK7hBIsdH7CY+vB9W+hPsjg2/
d5tuQepM0W2G0ZPWd9jyY/83gBSwcJZAhUfl3s509XCawnaJnDBTk7WxZlE8shXx
hrr0PASaxGb+8D3cBQuSGXDaVX0Mx57IhU0wzH+Gu5p2M4+ccmndktoryGoXExdu
EePLXQ3fXyZZTcZuFxmhITd/iAUgW5KmMH6MFDZva92IYhn9i9C1mtMUtNpD8Wul
FqmopBbKkjF7mR+8wE/ux6tfMmkPfb+qYKu1AowOjBbToSHY/wa57eB6Yeq5+YPT
YuafC3aSmSVORMzJynYPSxXt6yAtJ0Zw0pA1KvvpvvfYCQctGgaKNGPh4z+yEx7D
NUimnQWePpULC3YxJVMmg7tm16sf5moVuDKJIT5K6T5jwP4V7SFR2u26wkRv6arS
PQebvdQoT//zT0QtWgXj3IUdobWmNFvA7CRCKb6r9JHy/cnqdgyfeoXJsk7LuFPY
QREolpM30IV2bIpEkqw0Fy8NF5mT6BIJAvM58uhiuYBlHVld//iYRy7m7c6exW3z
E7wRXfAGXOr+qE4AqkZsjWXUPwPbWIwCqEuIt8nH8nrYVbBjSQ9FSoZNl9zrTX/w
y6QbmYOd8MXe8U464k+AATZbWw+uurEHJi3Phvou5HQFhDHpVjpEjYYplFjZ6h6k
wrcz+TMdOM38qERzjJhqZE2Tgcq284iFc3YuuoLq5GYcdCsQbjiankhEjFGGjjV5
4Do6m6pNaSnSVZ2LBbUIc9moE9sljzZert4r4Bvr+PwaFA8ocbUjr0DgxE0/gE4X
V//Yrl260HNHhVKHQh288esS770/Fuy3Fj1sFEnAP5LV2akqOQWeedm6zKDbJmhf
MNASgZhfViV/4ok0oWTg/e1rRTsPWU6o3+LSYxeX4nyC9B0YgBvNSdCIa/vLDyt2
kHo5uzDr3CGGKd2L2Q0/DGjwr0HH2XSroJ8CGKXk/fSmOMrXrUR74R4OEnRR2EgI
gSC57FED1cYRV2NWHixxPxnL98e5d4deJYwQBpATuBK8gFkpvWZ1bXtlAsy1Pcwk
JElrsrSrkWMn/JUoe/c4owlWEY2GaYzM6YyNDE4C69Oh/0V51277tjIY0v4aabhz
5c8+tIEYKaFCAV2EQj+ABtr0K2esBAeygZLnPrjv2XnvajLqfb6dwakJ/+WA9k2C
G2hEt/BhIn3vYrBxD+OVQ1GvDAxAe6i87bpnQMhSEev1uod9mVl7+l2ZxYda/mGX
lbnypN07N0bigFs6qdzT2kBTxf6O1Xd5QFcakwwI+Guzk+WlTd0sowNqA8G9UEUZ
DL+tOQ5qaljEpNeO/nxjhW3EFm0REBB85EkcZBWE31tmD5v3KRsu0WiL1gSI9ImN
sBE5P0s3bbj7DB5q6WD4MbLKbtTXmKRTkDjpK46jr3ZrOO1qEC48nSuySz4Xh4js
rYIEfkzf+bgxQsEQ/R8eo2apd5byznDHjjfvR6iQ3hMD5XoMzxwfjOvkShxJyWkt
pQOtZQ6uK/nxxluc3dQw4kq74pZ1UGIQ+YbI0ecuSgyXDvfWCj7Ib5HpKMqokSh0
ohPB+g/Z1BjdkL0tpCklxwoj1ihhv9buzTr5v3YroN8P/WfMwDViKbI2X5TN+Nzb
5Mk3rjlVFg3RzREOk8uAOzxisbAX4GBGZsPlvO3lJMTzG45godDSmtLSUTcbF9xF
CjKDlyAAW7HXdYcLNLXRbfqO/wGtYIfPB1uxRJgHevOmM5gQ4c3H4o0LLDlhCVGr
AWKrxDyIs9Gx+sa/8mlvAXB1qKDwDuIGlaFmYBy+3zTBplukbcXTBOfwyMQOVZ9a
+Y8VhIjLCYAoc4K3EDdzHicIvZF5Gl32tKwt45Z4+bKQB5Cwn5FddY9UnqdgGbmH
JpNZwxe0Jwh08dHc31FLqiMfdYJeavX1EWdCl9Q04w/ZNL1SgGnRKvG45QZc9xZ7
cR2RFHiBeC8RQjXhplHIedU+G4ojFbJhUdQyzhneVVMFVsrHw6GR6Yn7FJp987xz
950wKDB19NhxGflciDf8qJas51oTqDvvr+DbYSZxOhcdVmv/uW2jLgTL9h0aQ3BW
+2Ao0MtL6NvW1VwKyTYb20/nhNsFSRYUUSm93UlTdvaFtuUHcNkiAQGMQHUXDvIM
Xzl+DlSPcPVMkfzTuX2Y39EFRLtB16QoYN3ZiKxddNiIZFwgveY6ImGo8Z43MK6E
jd/hVFboHs0frPYBNnt4/LL0Etz9ycBmohN/za42kQ/BypVBkq3V17aHvizkLdBl
P1ZqN7YKOJeH6GfOOcB48Fqr1anT0bEJVM05X+tHop3zr/h/ux5NmjAkwYKcxMvE
WuNtwMXeMRmPjqnJNVNoY/YAudQkuAZ3YEowTXBsQfk1J+NmEbFD3IGtLAAGQzfi
BF3ONgK+3ePIHxehF8OzxASI0rilsWNknMv/TFRpL82FsKwH6MLlMMCeX57VjdvO
Wqnu2NoGWkIVGNos7qUoWXnsK1jae7QsKysDc4Ee6V4JAB9Ew7ty0K7PsmqotO5h
OC3TRK5fhW3vQPUl9etZg3eLAIw71xcIBpvyjiLKpjage5I3OZ0+bFCOz1WZXk8O
avR5cxZkAGGLycs+vXToIiXXP7RVIjvbyM+sxSBWNeBORMKMJX7yi8blAfqzw4aO
MVfmfYPmANrmodzJ+3jVhdwsxms9/HAUrNukC0bJZ1LzLLFjWyMW+5Kv0FKTacbI
O48U4/7x+U1e8KxcLrdd8rbwgaI7dR8YLWAfcuY5ZG/vUhYNWUiUPTx1HDRFJsvg
KD9HpaiRne+GMV8sU2UItQ/8Y3SbE5YfmrZXjPCK4anPyGOrunsqqUG5Um1TZnYr
B03qDbVOj1JJtVneA6VLYMiFF23muA/lmkvFjqnylEFu3jKfq7VSD4mZdgAE3U6n
0GczXyFsLAGvXOK1WCiYWU72u5scMG+ZTiqyfIpVkzSVWHMlrnQ3BabrsC9iJiRo
O3zR7HtIf4CmKk7GyKqPDGTJa/Cg4el986EtHVm2NuVwbwKyb9Uvzpo4OXrPrmBA
U35fFQ/nCryiJfS/qLwtnn5jgTnJv0dg49ipf3/KcE1nxDxikJu76h/9NxTJxvr2
ibn9xsqfYIzdEc9FjOuIiFp8T6cwkrCwpPLF/jYoycfQlYHO8jyFXs8KoaX8Iocz
wHHPKomZHHBiepw0DdIqfxu3bg5qQPitZjxsdhHnLwaBXhiz/fQPa/rZaAxGwL0p
oyzULuWLQ3TRvOx4F/eNO3YdEsvlylIO+D2X79q2c1jokpAyWjutfc983hiZ+PCx
j81QFZ6vshPTO/Op3bY568qJOQggaFDIA6vPXmM0pBNUA5XJrqk2vqkI2GvHrRYm
RZ7FWJ7YWybV8sVgEOJ+oPocLoLIxS0R6aK5pUNg2k5Zr2zZzjsxV3aLU1MFE6T5
4Irxy5b/QpfOrNXwG5EBOhxjJDytrZn7QTZAmqAKxBwp3rgTh3Z+YLSn/EIlEEF7
HKu2CEMaK0GBPweNAu9COe7V1VULM1sclBYUBA8YxBkdcchhdKHNbwi82kk2414W
YwrWj5Vk60Eu2i+IGid3Qwlw27DQAmSnOYYioVH7pzi7hy17DBd2mf7lKVFz2vjf
JI3BhVb9dWhxugMjIj6TDk1DWJzYUfDdTsDJmTy1vPc5i3nINZyC0K/3/F0z/jTU
5yFUdmGxBQPPjz1zr6MUbZHzwKaC6NnU5swS3qiyfR/FdJqiJAL+eQGRgeFS/n4g
NPSSrLng7QO/Nt1SVZL7x0kxj6lKRl2Ttyf1ngQS4nj8YZQghsfN70oLeOsZE7Ni
yPBYFpJibX0+/xhyMZBUXMEhZ7Lq/LLW471+cWXY6wjRbH/8nobFs/YBnCBlkp6X
/4+biFFIJPIdci7CFPVhAdAqdNClb/9+wnxyh+SkJLQGkAg1nLyqxT1hSxlxDNTM
MNFeWI6NguBtH3HTSsdqIRfZkXgOpmrL6qbIbY0lxqo8cWCQg8Ed0kAjOFEgS4ZS
tyBq3aMR1fy3jaOhjAQaNrP2K/HKvwTZ6J4y2q9bsGVJyGo76HacV4LY2MKlHt5Z
9O/dL03U+zPIVg1T2501QlNvgIGkG5FPS9v4nJKdENv/g38shOd+GmYCZuA1i0pA
csF54V6I97Qn4q39C9eF5dR8enoz7uDI8eGupMuSo48SOVQnxm/UjO2BDuYMEu8+
xBM1HHTv6QcQqphMdDdotZ4Ya/qU5QzLjuAJL+HvcuVUnOBmrx5R5OBin/c0a1S6
aIGS5omdKnkCrjH4O0XbMSYcgKNr7Ar7yeXfp3gVB9WMxg6Auw4t2YSXjouYZfO4
y1PsSxBN2Cj6gSpSmxXypTR1qD+qwiC/pWiBPYMyCyZ+JkpM+Qu7LdpxJcl0WB5H
qMs0gQmuGjRE+Gl77Q6OGcHToUzzgKgyitY0QxYFapiyC+smbRcNYgErXJMSiTws
4w8q2sEJBKofWMofMxAXEPMev4wnddKD3l6weHM6eUnC3IQ5HZcJd42G06lbbktR
Xllk0JgOjNcnBdzwlQ9iKymmn3mzXTxsVhsqwE+r0OIGsda5eu5GkCxUf+WSDuVv
9xIAmnQ3ZtsYMwlIS5oaJMwTRZ1lMdK4QTEhZ6793Nsr0CA90Sq5ve3X9ymywttb
7qQXvxvwWdmsQkptpeXmm8mCIZCyJcfX2drbTdNTop9/E8NgCfogdJBVNk9cJ4mw
Xbb5v2rfC/k3PH4mfZXPGtb6gFlkSS4XbMBicIKG30z7xNENeGiijs+VqU43LeAB
MHyCfMA+jy38v0JrPvMgyYL+fA7dEc2Yt4Dg0T/fNl/H3VcKeTa3DrK7B90GNQhL
b5efzwrd6Vn2NY6K1ermH2IsKH+GOuW7i0thaDylBRIdQkvnVw2bClNOdE3ThzoE
n5TZeiK0RAVzOuI6GJnfnxDPY5Iq577KFGhioQ/4bh6yqF4QHdg7jgGTPOmAOtYn
wFSSKjdS7bSwOCJmnqYhcjeApDorsDIxrXvUTzve5Qt+rPzC5Qjf567Ofuc82bcV
8kw5fMC2BnuEadsTkxpdhWMo4bGNeEWtDVFoM66ip7/vGYbGAfeLQG7WoNnvJAcX
hkQL/vs6P45GdZYMYAEJnJBsBdoEVufI8N6F9uW8Pb7n9Hw80vhY0L4AAKvjl5Yq
hxoEpI1EFYAwAI7V0HbkVuRic6opurL38R941oTNbTrrqbMRSxFWXw7ooMlp38jB
pfLN3Vy7rYDgs/AYYwqlYDod3afIOV7OXrjyxKrCNahi3oqMcJIPI/f06McBtYqj
DvVLftRoQuny7B/BZi8Q21fMOvzACHZw59TVWdkgWYR1zHfqN9/ojiAwe3I8tVij
I8Sap8LYFrbzuF5FGSyqEWkF/nDQEkEM9m/2f2TdYZ0w84tA9YPAo15ppdIcSpZ3
iDuJxBNbJ9d+PPzYOy+HjnwK71tPHmYo8X1xjT7+Lzd0ZxE61RYLYZGDSMX0aNFe
OJq82gvIxtJcKKUb6a5om+EUA9/Q/cvqp2B9Kj04RMrfv1FWg6LYqh+aD54jWZEd
r+xZ1rLmuf7NpblW9vS4EkKYfgXZKwHmWP7G1CNqo9eJKpVqS2+HhNZrFefZmM+K
p4IFCzZ/LG0LkKhaXQniH9wOfqRh92YE5laXMMEkxZbE8jY/R2u8ILSBRr12r9Im
Ip2jvWrTnGrs0eMzdJ8G155fzOPpa7iD+qZYOybr5nPDcHslK7bcVOoCZrFIjPVK
QGLL6hHtez4Pc69yKbnbkX5xzTb4IIJVYAEliBMNsKRvMfu6IyzssfqN3/UOjrfq
0oL5OtB79cYubscEig0dQqsNyrQlEPdBsRFlKVongzjjbmYJZcmZW+fn6wxCzT1g
E76gCPz9M2v58L23RJ1z5eMC9nKZW7HUvbukRUb8GfN31KiuND5pZs7xhV+vxc+Y
kMcrgrMff+iANUm6uQLLNfpTUOLXiQShr4qiPk40ukzUfKo8jKNZKGa69p7tcBx+
ZPGRe+WRfn2zo2zsHMKjPAUKbquOrr686y8ckzcdh3aRLsHtlKALORZtEts+qd81
YmB4Njg0y8BX9dqmL0tVrXptAFbKxDnnmex8xwjaW69t1aoCCKs3QkPEPDIbvVGY
MMnLYjSvqOWRODfUm7pHeBnxW7fez2BelCNF5lUtIEL5gTRmIdquw8A+/CpsjAIE
ZxqMYYKVEWt6kcYRJ7bm4bgMSm8NmxG8J2ulnH0POr0PPWhpLx0hFMjCUgQXocKi
XgVAHsiVLxQsGYSshH4rtRvgZrzi2dmAa4jjw57V3yeYkdhZLIvAWJ7GC4UkFkyI
HwsLwbFPWw94hiYb4xJMnSmTV4N3ECAHVHR5J7em5O5pRZBaTklywwVaQN5txdzG
nd4ThSN17R5PJqs+YXKOKgxDmZ7nXF95XT8Z2exPi/1lEHUnWCYY3aR7ovf9QCot
hIDpaaMg3Xzssx1N80GVcT0sbOGWDYlJniDfcX3PmaqtgVok7NnvDOHvw/CTrKL+
kWM7PwBd3avP3dTYCSZrkf+uhEl/B33aR/7NCwUvPIYqE95dZj+BB07Jh9hmvx8V
XsVX9JiVqAFprXc+cWphl+tUrwV6G6S6tUox273Hp9YqfpUSrYfBDDzm+y5oHze3
CPouRcOt8DutISQ3MY0VHnkwHBdN5ngszihxZrAodI+FlSE/p8yvlmhDMpg7kXqA
YdygNeliuUyK/KBFtE+IGAIOFnUCCt1pIyA37Wzjm61Rhgnobir3laca6SK0yNUe
WS7uEIoO/boFP9pHnHzhOl2LtxIKygFk7xlW8JQGZqf7saRAUpYnlgwqfsuK27bF
foPTQ4m6TSw+Kq8xT2DT4Ul8eAteU3tPgBslvzGPmwWYRNQpw+HeG/VyUc8o/njw
7UL337H6Rbv54c+TxriqjEq/4mR1MYDGbiV+/wfagviBSfsrTEm+XEcI9vdmUSA3
gvOoiwpT+8usGgJF6eUWL9NbJquiaaAj++rsATuC8dR+8P7yzavTkfFVzf2Qc36e
dL0/D+Q4uXWuWUW/RaOpCGpaz/rkJfbQkxIq5Ji/R7dSaEVWo7tzNN7D4RjMKMM4
ogsjsFRTzF3xKgd/M08eo9zRmDye/1HqP9e/roSF0g40KQHZPwt938Rwadca+PbL
pRt/gaN/a/hltyZ4scT3UFFDYH0phHzLAv/FoC3mmM0ccrPNqcT0cB8dkD1xMFgO
94I4NOflSVPZJxTeWthslLGPM28oSAXHpyNGnMZCUnYWnsyZzmeFLOSLUTgv9MvB
wvUqmPa+4w9BmQLpsYDs2MRRk5ZcqiK2qGqZE6zxyYpYfzovmmhkfid4MhzvwM5n
3RXfCfL7G0NwzdLFslASi9q+dkP8+8lR53vZSo4leTNEwwjhD7EpmpE4uerrsgux
hyB+0biD1ZZ43zldnY69U6GMSBouA1yliFoevEYbMnAlM+ZItY6uEuFXjsK8nt8B
ni4RTl9ODxaVTFUigA50uBWahloMXBVQ1b1FjBzXixVRfFmtmsAsBJ/LlawHmjaA
SByRKrB5Jkx7felVxPqNT+oTWO9z3wwJJrFcuEULKesMKBV7vVDfIp9gP93GNJg7
ALQimC9y11pyebrr+XPBNFc36OdB6YwD+/X495lv6wb4TeMHjzqauSQ3UQMkV4Cd
fdwu8YDG/Mn//mnkcUk53O8YNLmsOcbyzCruxDLGCjM/hP85wfvzUxWofkAH5L6j
l+rDH2Cte5sj/MbxKOnEey7cPuqpANPnT4HX+gZ9eccdA73n8tKK5e/fovDR+k3E
oF5u5urzPazMYYT767QWDz7VqbV2VzUaQ8LbdZEqYE+g3iaXSDutcOblP0clq838
3vskYJ2GfOXEuBSftNFn8IBQ112v2wtWSlaYMaxNAjnDzA0gYsWvYU0wTukRel7m
X/PZEvKEgEtcBoauxsR2ou0g0vdoocDITie754jwfxe8YoKKZtVcP1/IUiI//FtY
BQttaQqB0wSq8lH5H+V4Dy1Vf1YLWZD1pDTJtKMNeyJN8QDuG/tINgBipdrGUxl2
XSUIqvYEnbx37GyBj+6vjG6SujU8r8BhtS12y4X1UePTnRS/a3hzXa5WwHpCb0zo
k4IdvS1M/IBQ2WvHpR9cqe30RU9an02GigXjZE9RkARprsDQd02m2ONCbFbkTS3j
uoX873pBz+fHFcMf9ur/VptGps4DQhYpiLG0F5r/krY4PW0DkHn2RJyg78Wr0BBP
ibBjbzgtq9i55Hrm24ow8Ubr6V2ijY1FskGmRa01ho7N+3GJMPYV0vAuwxVzKb6s
4AMtBDHlFRg7T08dOFCPYZ8J+Di6soQywCZNhxe3bTe0UqjrEIIuchG3p45qV70m
KuDuwDtgZhSmvTxnHvO5Z90KOl2ymBIuMPCL13IEEbjDAv03bL3JbWsRvXSMAHPJ
kqasNTdRTMPCGK1Dj3Ye4HpDgt0K7Qr43DhBEaPVxouBq0UO4xzGyxva4NMWQabn
p2prxMVnCXV0A5SmIEl52mCKYjw65mvTjFpW7p3EJ7P+dzZTofDbzmGqlwawsCmu
4YjuR5hnB6wG4AUJ9hIMSzgYwE5nbPWbrfc+8Hq5eSByudHhEde3tabIPdM2B7wz
jXs8PoIVF5lk/i54yJe0Phme6+DdcjP2aUF2CYPqJED/wyRMlEgf2jRHBlAQQd94
dwtDnma01jSn9+C0KrJGBNAmjKLNIvYZeIbIejp3T1H4IxouRrIYoLlRTKB3vqUB
xoI/b1rX1lMicQ0u5ebXWi8WK4UwWPtHJYMzAkA4841v76ecSgVm6+agfkO8i/2m
zxN0S4sv7gbkerseZY2ewpq636j5KROHN8jPlaU5v6/F48qhxZfm0KyjXzV402ED
zt4AeuG5HzmLXZPc5gsOgLG15AIn0giJzQRdDbEDZSiHE8TBmig5pfXCjWLk1OpL
FJkRarjDHu/jXHnJpqdkWe6sYaVzocd2F/59Lz7HWdYkEtGbjqQpk+yS9iCof0ts
le2k4UIz6MBhsfbwNuL6g0g14ybK8/00TPq9M3tmFwJqgmqeh3ePjoQ56fmLJyQV
Uo+AGd4rhO8dSQZKrkS9QLXmRfbxGyGp6PbkmpKO4pfuBcmn5Fgx/zyNxpb+kMap
XK6yliC6QfcBvVIuLCgnwVoZUvkMK5AVrM5z2yjAA3s2nmaw6zRe9n/BuIVdp/4u
Bkvq/C7DiQ+vavLqIgB0Dy4/thYkKhANIUw8/bdqf3w+PZnNynx1F4MGr0Kok/ZU
2/2/dkDDNRNVHKtjtFgjolQBGOveZWT7XpTUXiqBdZ/By3hYqAz622wXtdMtCrqc
eM2W27RkLv4+sN2zbE8KO3Atumv7NgCUD/4X6megws2KOJeLPJsngnjzZszhtggB
ORyoaBXSLIwn+ucpSWekZK1cuvpua+HsGWlRYoIkYJjZASDfV8uUHmf/pSvycLWa
9Ir1QQkEJ+MYFCF1pei3J0pfmYi9Jhgagayw3NQT8Kjl+EK9NTuCoefKiYMPKCXc
D5yC8UCNNM253sXchPEa8SpB3Vp1NFaQMkVdeNB5c2ewF9dd9TcDShPKxnKV+CP6
k+UbgbrVyQZ4yAVUaaeW2OkG25wA/AvT89HnwJy60WY9a/32RsgmWyg5xju2kJd5
GzX4p5GlvxaC+KP65bg58oV0ZITVVjyV5XaaC+JyUX5QOtOocdCWWm0m40Hg+0NH
XDc4Z6dUNi/6AMEQO8I6lflw26o2CNmWrUcY/2rfKbxK9v1Hs0SHGQSdI02cZO16
9BHhzknMF+V5P9W4ooXDEtWH1RkosV0Ottafv7I7Q3zZrphL6/UQACbvV2yYC1JX
oEp8yi1DbuhalC2Q/yJFFP07Q5h0Jwrpwa5R0MN8mVCC2nbj1GfpYSnrd4NHxL/G
pLoCJKnSomnVZykVkJ+Cd60aVNhhaTK5vtM9Nbjd8b1HbjTjHflkSlWYCDaPYZvP
T+lqw32GEqxcVYjm1VPC57DJrSmYjjkpvpQk5rVxjlnRtYLRStapAsHF7qS8+M4S
dISPQ1DExBvc+o0NcQF1hLXbFecI/J/xfxAhHH3B6COyQ8qMUg2g5VEDNXAh1yHQ
YSgOurT3gOdtlpQ/vh284PwV9sqp6Sn7y0UgnnOTnRDRFSvwuPzUVD7VT+XfQy5l
j9AKb2jB++uJOCYwtlXC8Ac1ZJfJrTCc2wdbF17drFki9QyodR1SgJW5QQbgzQnw
xWXPiIsQrP6voJJsjMgzGiW1eFF3gGsIbh9SjZrqA9mM8T8CxrjINIl119hTTrl2
2udOkcvweg2DXRszv2HMqp9qhdMDwo63M+NbiCZ9LAJLnSjC0PZf6J6tWLwy8pMx
iEVoq/WPAgmPcU43T7wjjAxgGzPuCI1NfLp5BVwSomslwVRO/aY3D8BNjs5XrZHn
vWgb/d3MufdmvbuJ6DFB7FZcqAHfGYzS2ji6IGQOsDIvtKmDWjOhT2hnQNYyEC41
VX3Pqwr+V6VwHbytO6Y2i8i38YRCytLE5iHL64gLAMCk5UioEqjs7IF93SB/nGMB
xi7xNotH9SRwOnhoPs3y/b+EIvWfHLoDKeqPLMOjBTNYkXySQ0KOFCsocTG/79j+
ZenqJBYmjrDJ/lxGH6vdsUU2ikDfzK1NLFVRHq3nrAELoTKVfFdi622vbHUaBZd+
xAA+olRMn0heRdjTF4pPsA5HhYYGb5ZFbePhkScS7+j249McTVq5nkV61CFoWvHk
FDg98y6HjK/HNC1e9DCN76wZi8rMYZ867tndDZMdOU/IRdIJzenUecshpgOt0zuV
YmJRAr1FQzIHesrq1V+67OYKMvj3cIygxVQzfj5mipWP07X4SP5rl4MgHc62Y3sY
xuiGUCDb+yodrZRYXxa2hYfGS8fqNctqyrhxVWnrMFA=
`protect END_PROTECTED
