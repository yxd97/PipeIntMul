`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4XSTFAhtw14/8DrFWnqFdP9qGiwBMpAEe2ONk6whkoky3m0bZNFDRyzxb8SOk7Q4
QVgSQ5loaE+0/peHdDfqR1wKfVHFc8YjnOxf5tLzhwjWRHS99NAcCUCbbe5Fqxdf
GcSF+BxjzWFbM33tvCwcMm/A20RbVudG5u19qlq96o6x1woOxP32i4eGJ5joAsY5
emlzztceCuIHp/hc1kf9HcgPgi/cD1m4wBSaAVx0jUAeMfkGkYm3bIn1OA20WvAV
gi9eXyfJMiOkjcP5PwXdCPVQ1RE/n806TGqNIYHAlof04IrULfPDLNI7VRV4E8Tq
xv6WWm8TDLODdNWsY0rp4/2gZCczu9G7KkRXunKVSKdrACODogvvs5AN7Vx6/stK
NxfaBJDaIxLF0dqhomsuZmfhw/FDBOOh/cXgx9Zn14FRRbkdYENL2OUX4OPzMm1U
4CnZMVJfDMiLvXJcGQr9Y6UMuBRK6bWnatKskmgc8T10QlOUl165icnAZL2oITdA
Q7ZszALof4f2OdgpTSU87nRWA+qLohapQRiFd74kyhSO57uhvWYJYeehBGPK0EWk
ErFxxUbmbAQxrQ+SUTnkEEVA1eB+g9Hf3eugqzqmv19WqAyMokZ+f+JFAulYxoBl
0AWyD52w3V0uJ3lHJMjZe6oiAII+s6huz/9kkP81MNNKJH2m4rebbP2SObJzOOJf
WanDQAnbzPNb8IcKgU4Bd6HNHyJglYFgSIHodI7HvEtFADzNnfzeTk86SlPVdcSK
RA/gTDdql2gWm/B6gh5oZx+ORSGVj8gIbGgxbADBNbEu+ONBT7lS6AAmdwKT8Wx+
aGgL/AvzfBM+aiFhFJIxsNmHZg/9I9zWWMLudPLEGw0=
`protect END_PROTECTED
