`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jrSOVfRvKb2N4k1VK3pcrjHM+BKuo4MQpz/bG2saz4Sta6xdsA7OvswEuU+MJvfp
ObTEF7Ik1xdC+wWGN38QFnkCtmNPIrJ7FubbmrFhJ+G10IMTfddJdZMcMcM4SUHo
XEZ/LP+mYcTksb3DL0HamwP5drao2l5e92BJPv2JAhysB/UocUE3IvsjXIFWxjOR
kyVBM+dVCf+QLYZjZ1dwypSmIowFUejmIrzhTABCbShx8DwqxflKMX3HCKtU4NLg
7XmdI2ApalDg5U16UqnI7cKpTqrjDjzXdW7Qwz+1ZuXKrrEjeeMqbfwGLCqvfvFG
u4Q7esZIx1Vl+kzL8pN3s0BUf5wG0ciJ+5R4Jlf/hHlrsseTAEP+N7ipBjgpYBWF
QnN50FLLWVvekXjF2WJ15q8xrVMlTEC5Inv6qEpKJfZ0ESfqwzK5Jktuf5thtkNy
vbmrKyfqV6vaw+EZWCYngeyE6/BS0/CqVDN9NQzpCp3g978e0RYgSX/Qb0Lkzme8
Qgs5zEby/S1IeK178/pR5ToaThk/XUwGpvHNGFqaJ43s6RuLnG5ZHwSTZyZRX+HO
qGA+333H2uQOp2VK6YnRzRoAyhZyL/38SmJVdQnpxrBu7A0Nw08JHU+1dJYdgPkE
kkPUWi8ZgO2OFq7OSp8ztx5lkfXkzZpZPJt8bzHEy1JJpMpj7jgFdeKzrk5/Ayle
sr8i+DC40FkwTbzp8K0a4sLkdHMQLzjTBSVF3mHoXvWDYORXv4zawD8LSY6dM+A7
cWYFwH5ULNYXPU5xTuBrxasrAjXKjFVESl8U+XAZ5sPn8/bAl2ZeqeHj6QjTdWni
4rgjGF8Pmr2sXRJxdygcMkB6/HUH/rFOifCgyw/3gDTfmMRS8G/Mbr+zLB+vGc07
6aE8MHBV89luMwICC5sbaZLB0JOKJ3Ek3IwOTuQxHYtCGkmXwL0kmlnm86lUPutQ
GCbnO/b1MnUfizWMHgnV8hpBtf13kvssZCxEfjnXPktzCvcFCox8zlOX9cAXIPdD
Ec4Cn+QnTnFcRkwsixNS5KxEbaQGIrGe3X6IXbVa809USBsDD5Ohev0xm94rAPMo
w1mMz9uws+MgAVXqT74xh8SWQXZD+7g4H+3HqIjlt+x0A6VIfoBlAnJku4zlLrZe
9HFuwJzF9YzsaH2ycLNL/MxG+jpXGKqOCE9mbKawaakr62cNV0cHLcNBemlBd/+e
tDT/XZiqO4w6PRjp5GJIlOylP4/dKS/z63abCNTsEQuibMaxQRnkMUo51Vx7M5tE
aXJ898JL46GasD4TEH6ZDQjavyOVZy+lcjonOQ+9RjXwI63C5yGzfQZB/HCUNaYV
0w58BwiMqrWSWY8dvPT2R7Ts99L/cKq1HqE1a3e59XGPyNbPU//weXQOhYURNDep
zTA3wSZ7jy9QIcLy30E1magU5K2Q/bWKo1MI8ng8jecYDhLJXbTg2ZcWO1y0x8Hf
KpLTRgZRbJ2TKs1SBsCWdTusC/g9F2P+8n8FBdsCqjO5iH6B9sDo9OCTHR/7GtyN
hffWv6HJmrpKt/3DmcEpgHSEnvQfr9T25gD8L7QZ5NEJlKhvg37w0mBMfQE8YvnG
9B1bNOofoAtbf82rZMBI730YeWQB9mMI6vQNj5yFd5MyLDy5/2n/XGKkAf0Re+Sd
he5l0uM7+ZlMHhepGOX1P1VVHbnmpuOrJpAZ9+HXDVN048cdl3Qcxivyx4160Qld
ixc0pSWtYUlsIVuX2MRRrHhoxUFUCTB+SBgMzKKZ1UhExLdRSEYpfsoZbJ1jiY/D
Gj0FV54l3x99Q9ybIaKhYCJivUZe9W9tc9nZpAThodkxYq44EbqympaTQ29aidBd
cIMZbWD7Hi/2S+qyuVMjtBvVK+NSZ6gAnlIzeMeLYs+QOqeZGLMCLxF5VMXw4Oq2
9EixynMSCEFpx6iFYXIbppGjVmcOkHJq+xaskGDO65RpFt+3bEA1RsINm1yz7Rbp
UI9BHDBSARUMEQkNuxKA6iH4a/ZulC+0jdkxXWL0HrPJsAsOhRwIQUl7ywRsHzFl
28PCDMSKJrhR6PKecsBe7p64BGP5X7yBMn12P4rB/9IhkOLWN7PuxzzTc+OXMYSS
MmYxXq2GXxgHk7QrsqUL4XSr/Fcx4G88A8WDsKEQOfHMRYX76oVyvrjOq58miVPG
Gx/5zocuEWKsgMJ1AeJ53nFlP9NlMKVhlSc+CO2wvS9bkvHlwgId2lvc7EGMkXf6
LlcGcAUnEEyd63gpgdsjHTSV3kF1+FT/CkY+iAkAmRATSGxl1bNvRZsmDRvsd8Pq
xsUA8q1HFm4yMMlIF8e+KAi2xHFw91ShsZ9mJbX7djTchldkqQjsUeGhNx0xIhxk
sIM8BHV1is0K4FU5RJD7Oee5dTGaY6uzRI2BC7zEB7bNTs+ayUkL7SO3kvYtrObI
aq7eEOL02wH4AZt2cRn//u1uGJBfjensPZu5/QW43iKBJiSNaBz0xcqWg6CwBVG3
Z1vy2wwo2+lk931HP0D41kbkPEM7Im/DQksveUk2paL5SNvaKjKQNig1J6fjR9Df
cCO7JRKQix5UYZY+WzfOuQFp6AP7kApGpELw9b/mNNrOie7CIAK5uUn8N7fc/bBU
krtGKC1AJ4M6dySapMzlYg98PrQKmBvO5IHolGaEmmU+zqAXrQ7p8BgI/8nROccV
ISIO13zkcg7O51BwYC48+lzZ6lCRUmr+wBzRxI2BGhXzoqv184Cy8tgfNJSeppF7
2QKtTwCjxpUcU9x8WMw3ULBXPmK2KKn1ZuH4Ccqb+0Z+bUjCS16YJeWE18gH/1D3
D7Zp3tR8wOQLiCsVsGt6k9DxuW/TmxLnAH5VSsOtbeJnzTbcpQVOvasvcPdL4hsj
n+NCNP3dVsn5VcwtCYe3+t5I5Wm0XL575k8h1zzNanP9f9GosYheESkNDa5/x/1i
gNKsh43Uq4liSG+9rXFCG2clQvnlAdSOQ72rW+PLLIvOA3q0MFCm766XcjF97k4U
rHdoBJk1sGlqQfd4h3Ug3KaB8ywRF4w2bKfCwvopcXYIynD7qcVCO0BVUhei75v2
AejGsXpuJjuxJdCrrVYrI+V0Dnakdc93Rjva/3EewoUeIy8c9apdxNZbI70Eh5PQ
POr8bHqh1EnHDEdyHfp/V79uW9wiOzA7nvrvgiXHTeLeojvNjBf2kQzNyqJXWpYi
ATDhkNjWCXcGSFMZbsEM8tlCL9qoRuzl4b6nngIYHhxJ7tbH9381XMawlk32orbH
Swg8foL3aU3i77NblboelDtiwEATx5wwH/IhQJFhK+G2o6u4gXIwzxctWNY9SxLk
08RK6mqdIomK+gBkBqa/R54gtiEh6ACcsMV8NFWWlmvA4RKA0Rmb9TLndCOwj9QR
0iE8zLTvjlofStEHiKzNOJYPhlmdkcQDh8XuO+nLHL2WZBx6bZd8iJUgqTcah0+N
ppOPRWOisviAKZyM788+EX3WRu26wll4vHVMZY2XOfyQIlfTgE0RKjnEX6MD+oU0
tGZvNXbbFJWbTp/j39ciznvYk85mwmlw9JbDfBznlvK4IFXVgn8cNfQO1EZQLtSm
brqD4pv1mtiDGk6gXmAEnnJ08XMjqVZegE9o+wtBro0WZH/T6tk6TrclgFXA45f0
Oca3rqf6iupyv5k7NOpssdACXdrFo/Dv6ldo8B07B6veWX93rnrDnIToCpOuzfTF
YuVQ/4u3ZJFTCSGmCt8si/6nL/nNx//vCRsy3H0uz+efozZV9M2MgTqOECX4Lxqg
991jva99pUksUACCqllYfZC5/LMoIvdanL12r0aCyaJbZmweL9IwGhxsG+H61bwj
L4dr9HfWHl3lUyArLtarklGo+ZszoG/m2eKbwNgRqsukGBBVqcFsNHz1BkDZ0vxG
d75NjlWoHECFXiAFOaKAACOWeMLeQp2loXAapeSbkatLnusMeGnA4ExmAUUXYOKs
PZnrOXSeVOil1o0RaeaRKvxiQ/BByzluQNnWFH78ug0XAEj+CtcAmXAL5hIrO2Jv
5FcRbf/fmfH+Wy9DHXQwZqhhI66WhC14/YaiAD2kw0bEX8nJJi91apmpQ/SR24Wj
mur0Ktds9yXdEXFuKHOCzS31XLiOFsNYbGbP+DQFssxYDAHHtrSktuAp6rKzGUEE
mgeYvMVrda/7U1VcPCXqVMs+zh0hcL9mTIDevMd4HZvAX2FP+UNaBWsE1GrZISjj
1TOvC5n528rrIeHoYiSGU7HHB1Fm0tdOxxeVwjUQDVbOVXMFzmZJYMpcFy6DIO/A
rSPCTeZbOZvRw8FjQOYxdOAqLVxVxsB/0nWru3rSL5rxKPPQaMNGnFf2cfHDJYvs
eDGhSYVqUUKv9dwkiw9CiSdAgD1m7Umlvzfq+SwUDh9P/DHltcMCHdip/kOkXrZk
3EWaeLU8YOcuv9IFALixYAr/C40rxUWHUwQ3UlloxGWZKeNFgZ6XpDYwx/MwNzkO
Z296BrzHyGS6VafBuky/ByyaOVph30sks1sWom+KRmKJ+7Qa/CCrg8IrC+04y6of
u9lGlBddUBLyV6H0cZ1qsVBfC7+BrYhkrWiHwf34Fmtv/jxBp0P4vb4/hXXXMG4D
cOFRkZTCTuRwHIG00YIZLy7ubSktHT/MpAgqE55EHXHg6a/w/k2JYVM7ZSf1CNKA
lMgStdhtwzrbAitHxoxiBH4G3tgduGmNyURa2dAiQ5ygVeOq+IAe5alJ6CVQ2RA+
DLfzILVXMQK6NUrF+5kpz7vR6Y1DAW9OZqf4WYOGgtQrKMr4PAT4F/VII6OXnbUd
MZlBaM4xlu/bav05E+m+vZfiNbyJjV1HH5Hinb9RLL1G6lcR/drGUHEK/jx17rP+
Vse7SSxSW8zq8bQmtZfSBwEWXvlUiw4IgdfAeH5zAuP2vmYBNsJ/D6CgHf+IySxb
Ajl+k4rL18ULqoGqIAdlXuGxZg8qoojJ3T2/a6lRhg7XMjAnAiFQi8imCplAaRuT
PbwfrugPGvi3DXwGrKL9ckxaQZwdPuwP+0IJ2YY0jZ3ZRys4aHCoWbSULpUWMed5
JbjLXwYFnxRAebHiiIoQAmxnqchhLx1CYJteCFzklsysHaCfPlMaGHr3DM4+yfZA
Wr6K54HWCqwL9FBQfPj48dDuS4riMTFehRdzFAIOKnM39G/hwhKvQ9r116W1c8zB
aK3gUpb+dQ8kaXn3cwZDA0IEMkjXSgx3nxZkS1s6e+mz1TUYcJhA0U2CSReeaB2K
MUW51U8ezh9SOyjf3F7ucyObd1hBEKc+yC7U5+o/hUJ7Ak/3ueoYkabqVWoJH5ki
lB8Po29MMHwTSx2iYWqiBdt31eqqOQlz1NaCxx4OLSUpgQxSbF1ND3M2g6/TRtZE
psjL6A+/zNG1XJbhAOgDwvoTek9tW88iVHAYKWX1C38qudjf2X1lpO/O3xJW4tb5
jittDWfVHFjv+QUGJPSi8wdGh0ezPJypWO9THNasqdDIaRmOejCp8QWDMkuf361E
853rOaOWkl2j1A3RdGZ55GDqJbiMdQJnXMVmS3ciwB76vWg5bTzIufZMVq1MK8rh
IzXXs1fQM+W9Kp9pqOeQ/ygNGqRck94sRyDKcfUD19xQkpBkmCuoZENEkTXduNgR
d+j0YYNHJG8oVL61PfW9Seo3b9XKCw8yu/wA0ThWRAUb/VQi7LRTj3IHSfA//jBN
862YMVDXIOIfDiIvyPKqgEOs68D3MYFfh+bFyp8lK01eW0exwj9RORYF7QjDsjfn
vL+p9dJmbM0LxNXcwKK2adU03+s7LUbtYOCU1uWp7uC/BT5ezk2u7brwMqIjz9O1
3L49mLNAxedPNszR3LxCHW3oau9XYVjwDFXbvmUj2LGO/Zp/PZAW0qgsylK37xgN
A3HWnpT3OQaW8JZ01up24yguTzPd+DIGQGp0ksXfx+69AwRcJfFXdh1CsBvtNAR9
u82p63nFBNA9LfmHfqZdDDgwrvvQIgYBgeoVw2UtoZSd6J/Aek5f3cFLD65iuQYA
qIoRmeUg8yndr4OTsSIUoezeckY5a6z2QrQTbu8efPaM1mRI716OG49f5wVWVi6e
Z+Te3qeTPPT4KHY7GuReS5xgXz0JKwJB9uPTnnGqGbsLO0xSwoO9x80uOKRIHdZL
FXXXhiRQOWUKO7ZbZcWefDZDkPC1Yw+9R6nVyj2jc558H2Tal+xgYORuMof9Uhyy
oeceB1qHMDwRjhZTXyA+TcjwYvLDlCgALbT4MlMLXFpsmnAzWnrNd4DNuTKlDMD9
3XoixmZhopG0ML1uEHm6EmY2yrRWBGYVLaH0lRsjr43GNgbH3NKdya6iVdi8O45P
MdwCWv+M1B4nGbCAIr1IXzlsC9acy1ibztAnwSRqd+27gnErpMLRMHr7lHDrLYY7
FrhHMUsJPIoS9mr6fhabLhDih3QR7ZdBLCYsRvTdJIVmdVEzn55h59PuXarnANwP
9Doqwmwc77pjmi9V8PTryiuUvEPQExmeAgzFyXGeQQuKGTxh2DPuLag0FevkhjeF
TOtV00zzWWf5JuaGHLVSuHkEfS+/f6wdzHNYEHvbNbDPhaA9n03hjBFWNLNpxHji
lYp5x+i3ZpT0cMvf7egyd6vGz30i/Sc0NumA+GMF3TL/O+2kLys5UZPMCj4614pr
pJYSs1jc9EZwlflCnHSjlwsVPEWLjKTx1SEg0R9FbFXpGFtamZvn290HFjLH4Cc1
ANwCiXXS6H2cbIITaKyKi61PoMqkDwcpaCq+QPMTYLaluYdIOWKExqQSPbLNEJ0K
0AzpNRr+hwAR2XNzNdq2wupcvVzUEXTw6ol/X5SHbhM3UaIlGvsFn+JdccXhVjy9
0ousVPZ5of6UiDp1rhNfjFhL4+Sl1zliW2YHOh1MxvvGsdhWIdREWp4oe9oKcPVE
LD5wa9Ut1OqM/+kE9Df5motg3mpU+W4EPK/rvuiZP77NTkOF6EM5UhFphqcqEUed
fO5oOLRjTbqkPFLhF12+nPZd2ig3OnHg+CfNAahS0pPCawuKx5lDXncJcVCuwC69
`protect END_PROTECTED
