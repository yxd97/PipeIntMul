`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+C/CF2gRL5vc69uQEdtT8SLwzSjUDVseagWqHx07fhcqG2kmk0IrR6Txzp07a/3
dELjEHg+y7M9fbKKuK77QINXpttOej8Lj/DUZGV+oQHy5KNv1+SQAvyPF2yWbmb/
lih8A1Jz0on+KS0eJCryZblikDA9p2OKPHhyHkyNYs2WR0KpcZMO9ET0/AAwdAem
8tyx0vbNBOEHgdvFUqhwpjRSFv+ru1LAXxbRuV4AfywRgyVQklJepjWUsciBeiWT
PJIUVXjTM8z9EyeudpgWzwSZXcc5MB9Ge0/SoeTmgOPfvsNwx9UiJhxHwolkXNfb
sYtJO5g2l+lhpr2x49yAqj5W7Xkg1iC3XjlIhQQTmbKyi3ihz52OoGxISC1r99Oy
SGzPT7uB73EkSxG/JV1zPlZeIyyc2KUVR+1CdQCTPSW59s0uP5Imp7S3R+LjHnaH
`protect END_PROTECTED
