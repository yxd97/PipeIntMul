`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+rgYJ3LbZlV4FzdzRtHsGd+Ybo5m0t3iT/j4BSq3jxXcqW8TibHRYT/OqsAXKrV
vI8bseAhLYV2luAqUCaWMFuLsMaQihp9uTchzwao/87YfDiEgxkl9O9JYVTpjd8G
cuDI+TMYczKORZWxujN4oUeEe2QJND6br+4+ubhRUOgveVn3hoB2ggvOrp4B91sJ
9ORpnHFD4obhorF7Q6lKhjFoors9cpBIkgsj5r7R20rG/8dBUF+Fnl79uh61z7nM
jkjEX/M24EsoT/HFbmwIW4CPoYh+LGrusIW1KwYlQh2srRJROPOEWKtMzXfs/xRJ
rFVp1rXFdR+CF1ycXftXq4yKN+mNse9dLdWJFYHS0XuTKA+MlH6ItBgmA0V0qZ6V
GB/z4MXXDLHiKHSeYkYI94ADT3VcuM3wvsksMPhxH89X7OUbHVYLM4pu38CUmLBI
KWswNgnQB2SoNfLBGk+RzxQMyMV5UnyrwmQAJG+1kp6dqrFqvmD9jESPL3w7y+dK
q319/rPd8rO+BID+sEb5zGjJBRAZB8/oKcun81cYYTmVU/FTuZlDcCzVmDSCGfqg
c4gQYSOw+r7LzDZ0bL03uw==
`protect END_PROTECTED
