`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uL4bLB7wICJc1UteJrRPdhIXRupp5pyy4F54lfn93xFd6GP1BKIQIoFbEDHNQt2
4geDYtU1vuBAsv2L1wNJ2VG/K8qBuAq+cxQB/XvLxM5lsqliXNDzTERm5dqxpwVc
7qA3KxXgEbGJnGlURyCNLwa7O4B9DkU2fSZQjn6fLIODTfCBWvEwvFoD3pJpIjgp
HslsULm0EvscNOZM/36LDqyvMILXOdrHHi25Tasr7wBVLdgKz2Q/JqqCAp02W+rp
pNMU2GNozy4ImLBvi21iXuEAc090XE+wWr//Vld52zaIqoFGSjFQIzSq/C8iop00
CpcxuHjKwL2vx+2UuQTVEA==
`protect END_PROTECTED
