`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
08G75joL4IHdkBREdptEKDwWFpebQeZMLswNUi8ujE2Y4mNog7ciGbaBSthSjUGI
MwHPNSAE9T0O1p5lUVdN9euJDfES50FqV4s4DjQVxtNCZ435Henq7j5sBrNBTl8A
/VsxBpFthxQcOI1WQbPBWCaxfbUwaCPZul19POFtDhAUJ1G+2pqxL+JGIdfnkq0x
uHGtg9weQbbNCfAD/JDX9vTYgKbEY4O8Z2Dlh++H7OmQNLNxLLddW/g/3T8MxayL
CWQuuEK+qX0JuAJzlukbAT+8xqOZB70LgLPzD9DIj3Fbv4vD6gXuiHRWrklEZeS3
dP/gMyDpLJD1CZwiPZ2AB+1cm6d9j7Lbgfy/0zHh8r/0kZW9SRWYA8burkP6EnwN
YHP+v37SqFzmAuOOuegI+zrM2ryq1Q2AH4U6bN1CFpRtJaNAb/61BvNvzQpy9Shg
iy19onU2y1XvSLwwHgOtusa8lg2NNBM1WAAIYhgbRC5JnZ3kEk2rds0ZRv0BmyIy
`protect END_PROTECTED
