`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+ARwqccjEBTHjsTLNuQN78+2BFXL4AKRwlMOTE1hwSjvd9UHUoXnDVn7+XL1zDu
E8XqHcIQWgBFWTlxW8K1VowiPtD6YdbMUdM5+8/MRHWo9K0sV9mEi/KjNn+c7z0i
iO+vFs3QebBS6nbI8THAw9z8BrSdoFtqPcAGr0+a29+c5jkYA+gA1HtKBAoaK46L
XaSZKa7RdhEVfgTsG/T81jedAw9cxMy/j+oV6hJ4FktW3SiPMtGPR7VV1pnR7Xjg
4qstAkpQFerg0U4DJNIU9SbRbkaT9jw0RtyJySL1uOty8kvajvDD5GNQPfFTib7A
1hnGUAz2C6fDcKwUonAGcVx6+7TszVE5z8XUDRsuxfFUU+/8+Xdl0gl9536bPCsw
qrCH2iEqiGmkAXPbAGcw9VhX1NDjuSsC0vXuVrnhpUyB0m3Khd7rPztf2dGG11lZ
vxHTIOEcLKBg1NSvRls7sZlKPeThhHCHWpcRncvZ/8bmAMn4xT2Vomsw4v5f94hZ
s41a4ftDG59jJzkNQckGU912f5Qzhadr1ga46FwJ958zh2FXQaemxgDCIWL6zI7h
0NvXUUUZBwwPXMEmPFibxbUbnnu7JwoeWUZ8xarlhAZn7zgqWe3iuA7YX1mrwRiq
iCngX37h1jImQY1jb7F1FqJDGKJqrBOLhnz+X2b+vOptgGQhBJ+GMLMwrumLEuBs
YuxkTAWm9T4xkJIj9lVgrcbWz5uvM8ZbvRlyPW/V2ZIwM08/ouqQ25EQWcWSvSws
n1qa+C4g0YGofOEYI2RkajO9pZLQK2BAf10gunpg5Nx0TKewh2lbcRaxHaWSVIWW
O8l9rHr8tRBT723XfRnCjiEOPszhxed2V0XmENT78CYNG1D0KrVwY074XYV8Tb3/
xlg7zNCvJ+K7I2yuIMptiJp3q+CVUIQNcFN905PsGFNfPDc4eYaRe4aZeDJ1Trof
jeeAir1MvL3UbtdJaZeGg6pYuBlz/nuwSbI5CCDCWLkHgQLjNP4Iz3PhApf+5tHU
E8GUmCMMaB9kuoRCCoX3gfboF4vUHXM/O1JjUA42hRCRJx5VfWT+YIni4Ap9knCN
tOMM8VfemkiVndBkoF6TgvMW5qE/ihyMYLV3Ly0AD9zwSQAjdCOmw2oz4VA0wCsi
ddFAf30X9rVobLa2ro1OxzBJTsJlumIQthPihyONvsES7o/s9qSlP1C3slf1wW4r
vD5xPLoth5TAWs1+8d1VNgucIh0GgSysydtflRPxYnRx4BQZql+NHCbq3sVgmQQ0
8ZbvE+drZhPtYKyNROPXKiqlt6Tz/mcXQwXYt5WqUOml+y/UvydcAx0Q3pI381CG
og4Q0aiBx6PR2qP095HFD/sJ+VXGSvANWvuJR8cIBND64YiEifHrMm4ivhgcu6MF
wNTk2P4pLqmciRolIRbUo2/pt6dU2OeRmfCWfZjhkhZkItMEdIqmmEIkomU7jOU/
vdGl8KtgnVv3rn45MAvLfxs9fYnsU6T66ch+veUoZn19tsPoxU/O5uwHFXVMqDsO
zCBzC7ptz+0dNjIwUGElTWmRDYha5JMClsvhzo+q+kI2n9VvpGD6UWJX9FlKqzKO
T8uZliNgiWPXv0qciEaQnUuWcth8fnufO+rgX+P1GvqxXHRLrt+f0lexmAniRQ0J
1AVcXnafq7qKfwzPTvPtjZyr7Z8JBSROODu+Nwylr6LQRltRc3rq4eJ0Qw9dylR9
TfMJaeJDuYYh3Cv8JREEXSdMnHqLPuMJLgU9Rt4l/XbcGBcwildt1DgrOG63nUMg
YiZ8wbMa8btLLq835s3Www7I7GDJdJYHVFCbEcSgYg4YaeOZkXqgtGvAje0afY3C
2SKmDzxIcT9zHhXekPLKXxtP1p+j1oiMU1m0QjzS/a9cQrqG9nXsW79btibqGQWx
t8ODLQIGbENZnJxD9lX1p33ptfNGfs6aqDImSNWvXqp153ifNtqqZj0ayVWIdd41
z5zxFvZc3feagtQmOHN20hkN0Wh2pkC7mWjyZ6XOduJRl18xas3kr6yhFYyF++HF
9pca20cLR5YHR+H8OH8Hm7tcofOLxI9aK1EjaR5l7QRD5iWbzFSpw3uB156wu1nv
jdGLCSyG5vaoLnn6OMut6WzmsNYWDSlU0VMlY6a6PVV4OovnDMXA6bbqFZFTqskG
apcXz7mL7FFij3yHUk7/GcLVm+/rxMK1nYcEggGnmUP+0xO2VHbEWB58WIpC+x1g
zLrhd8hJkDS5cGj7VMF91w==
`protect END_PROTECTED
