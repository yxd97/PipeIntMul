`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s8hdNKSIMTEjrXzGb7nbkXxQ2owO6lwVD9up6nSz3yzvZ8PF6cT6f6LVKdkRkZy/
2XrDpPYIfx2iAJHBzBOY8JivWKSBbW39Jf3vz4U8gaDQeX81Qp4XIaKptKw5P7x0
tzH5UM/Pe/TCfB4HsM3nhj87HqU+N6vdCqobNOBnWjboaZC54m+X81zXRMpirdgt
E5yE78wDLhxtqwAH53nNimf6QsS6VYmRh98hg8oS+wYViuFxbLuPkx8RzzoFI/hY
iYnZ+9wU8K6a7um/RkvZ5N8HR0mGdu0j6RZMSHYOAJjypFIGJt1hUC5xtu5DpjIt
eYyMXHkF04QUHAkIy+geBFa4HPYzX7ub4hXuV2OFeX61JGITeXZuMyIQuvGQDCUd
JU6npK6/ax0mpTgky56jnrb2552ZanH0p2qpysjLMoA=
`protect END_PROTECTED
