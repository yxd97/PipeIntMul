`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16Jtx+o9qU0QQYRAeY8NN9SKoXKUWnphUMvl+QWQ1Pqjuq6REUmQ0oy8QojuR7g5
f5iV78XBxxG2pnkSiUpDKv3Eho2xblGoHADqlsJZ6tyYDyMiRSCQ8Q6OVHy7u+vN
G3kl2++qJynlr7VBN92bJVG8RNVPa5U/tRAmtKMWBGgw6wzkgL3UPcO03FYoMk81
KjflVs4ywyHZniNGD5dnmlYLIyW7/YIIiml5g7ny54Xbw7vXoHHYre4rikj/HhXL
9HcauqLz8FGwa5uYSEyh+A==
`protect END_PROTECTED
