`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdNno3ZxYax5Rvd66L8IHeSmnupWeAOgSFbmsLA+VOL3rB+UdUg4U0TWEsEwpK6l
lf6aadVKNqeDTcNf17M7hWmmkztQ5gKnpFR8nHIaO7S406ZJEiTKdSamY4NtYLO4
pn6dT/uvPimybEeXlBP/6pcWhHq0EDtcOUJMwWRCDEbHM4dabyicHQFTHzcAYqxB
ErzWgKeLnlP1VSeUu5AKjsXtV/mcnPOZggCvq0WAetmjtSU3p3wYA9Ec0OKObsar
4Acv6OyHf2W0zdWIySmMdD1Ce4UwbW8Wjsq5rU9M/2YAqNyIr46ow8PxIuWBLSzr
zrae1H4332Sk4usScQ/yYAfk+nbls6/3HQz35f+bSb6xcsBtTqWAZzEody+EJ8PR
OjwYqcSz8US3twCk5riQbQ==
`protect END_PROTECTED
