`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lVHzSBvrdPy/cbrUkjG52qgG12Y9PtpsCR9GUrqUggtBbzFgTucMzmfqPRsUw83K
km0/URBL9DcqGqNqkIeCFuJb3ia2V2/+ApYr54SC+LhxxIkUMg383Df0HEPxZVSY
5AA0ZI+7bkxAsooQdWAo3549j9t2qMrgqSCdtaGx8EejFZRXGNhHetzRkKCRosiI
GkltWMEJthgby0fZyyb2w5EzYJSJ2RrolA78qeReCU5RnKEooPzhv2ofGYV0uze0
I6URAPG8x0OTIQ21kQJpEinVzyf2DB53X90IQbFiZP02+vdwbemqVb7QJZlvzmry
uJtiJ7Xj/MC2Ge+BtdEU2G5oxSwyHeAAyTVdUlhPNGMq/ycTl0NaRX9btj5u9ExP
foUnOH/i9LUHr2mfLp4JSoRA+//lH2F7zWk4CqkAMD+4aNcXbtRBy0j4cD1gap+m
6sb2J/qjfn2hAhvOixdjaIZp0xeXwAhiG7+qKzLKyHlKb9wKmVDLlrjkcno9+lx/
7rlsQ5+H0OBNxCD+y5J6PIUk6M/Nc8kyDzAnLjCD1X1jBirsEcjUkwO5KBJkQvVC
`protect END_PROTECTED
