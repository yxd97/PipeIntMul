`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mk0JSG0Y3m+eG+U14QR5g8Ev0L/JArHXnEu7d+sJYSyOi0/ha3QK6uccSFKqQDjm
uiES/kKfJAnz6b1rTgpFXbYoHgbabR076x+NVM5V98/i4qustBqVxdYLOGG/wQco
DDJnmDFvF3lEFGPQOLmVW1AowAhf+CpSSdRIM8ytFHf6zIG3c3PpzS3z5KLdHYqH
HqfIAqnjNcFeddbkBi5l6B5t1cNKiFHxvLv3yOCR2h2TMIpfp9xafLArZJfvQiT4
QIgGVcGGB0I4XalBzgMK/YFHwCjvWtCCh+qEGYwvYPbJwzvWB87M+BZywv4WuSf2
npkp0NxOeDwPGHSeHPhd2FDEVcpYUUprPCyDgC/WAdeqNsOjHTxGSK+KlJ6cJef/
Sjy0701vWUQ07KttBMe82IYgS02WigXDCwrmDNtbfDOs/99byX+JcAfiCrENNOZg
DYJ0VT4ksGq5ezXPBU0n3AL5lXadAyYSzhhzuzJ2oPF5N/Wk21kSQL2o0mmb6oe3
IA5/OoOUnIzgHcDCZp5elIpI2OkK97AwsS8kTvG2hTzJPYQKm5O49PzQ7D9ThIum
vJ4Rt7w7tIKC8wf91jZuOCGLKlnFb57H3q4JhByMTPvizFuJQRSuD5TSlCn7ODL7
3kSsnLG/x8l6TjEkN38WpA==
`protect END_PROTECTED
