`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+ByCNNxyUW+xkRHzBvS1cUAKd7ODUdCMSQ3407ojNGtXOUtJYwis+puXwkfLevg
a8eGJNwj4hgYgzsNsaRBsUDXOtLK8yq0d2+jCM1hWyuRy8XmIb3fT2/A1uSIwL7m
oYlr6tAJ2W4H/4pT5iXOtkhoNzooFOth6XQQ8vbg+XHqWWCASiQEdUJPIC1mxBMh
9ilMstcsfYQOdlrXk8bZy6s05iH1YNNdMfcwC3H6qI8VFKcRYZLQ9FPEEbhZzZ+I
/jH55Znv+6DYcY/T+QhJbiDQM6Xc+5BhqTKZpDKD6ImkCPxwV5URwDh1tYQQlHg/
bjyGtukjw0xVJqh4d/69zw==
`protect END_PROTECTED
