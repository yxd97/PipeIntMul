`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKvuh4p2OcJ+sb7yq97SQpRs5Du6yUwSvDGtiS9tsRab+VbOIjLIQQy6uM4QxVSk
EfP1OFG2lbA6pc/5mrR8HFWfe0b+eY9lVFoRZwKqwA5y0ntaQlSu5Tc0AFGBBakc
ytKczdKgRFU4+kyL+wyGD+0hK1S8o3oVHLSjshjfoyJedm4PCw7Jo1NEHy11i14S
dqh5IhHFGxSEcNhkvIz5QZUSSxE6NZW6IsgRW6Wb5pPoPjpQ1FoK+XNe0OrHFp9f
dnmIwoJRID3ZK1se9G0vP1ejkgwsxIfgqY+qezD60O6gH8SfGmrF+wS9rYVa4ga7
kljnbHC6FzrBxZKWQ8PZrh+7I0L8ahMGn6cxlm77kdZU8I30UERoMqge4mhNr/hC
OHKjvpYJeP1V1vf8SXqRtJuVcP40kM5TgprnR7zViEUp9diUlAOrQ2Hi7TtYFIOZ
xB8r8WT5bwCwq8FmUOzalNSx0jLkNGc8zBV4TzbfvNHEBv3SsDtdAj5r/8O0l2b5
cxTF+Cny6LCWASl2pYDqDzJMJKvbQ5Qj9TZ8dbxXIQNUdLk1LZLMHD8ocfha4a1O
AXbTppPfx+0Ze7AN9djVR3mMlu5Gi8ccTwMxIiwfkxFhrQjQHUQTHuqzhgewfEzU
c+QCbWOxaR9Wj8RGQGt/TWqG5VNPrZthVFqwKUelyxM+9aoZ7EC+bzHcnVk4Dmt6
p7HAklxA7XcY2pUqDdJuHpzLg702i1/1iB9tZhlrbazwnBfotj010vVZ4KsyWGBX
iFdlw4Rme5MksGNo+MRu6sL6oPqgaUwKmx1KG5/YMAg0whJV0SN+b/iIZpOXc3iG
fIn6BlQYgX6SVreoIE560Q==
`protect END_PROTECTED
