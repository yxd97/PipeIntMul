`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W5DGUsnHP3jZ2Ne7tzhGJuZBg2KDrfEWE8zXs9ZypNabBthoANMhiUBY9ghrb5fK
P1TrOEtY2YVkELGF5dH+aU7joTLBpislkhofX5e/25B5bMD8oUqptSmxk8ePE819
PUFyj2vhU9c6iMUC4+8vKQE5P6d2eHYyS4HYaJgMHGktcE2oHSVIENp7js/aRsAb
OqZS6tTUxEx+BW3fMj+9Enw+76eddSQVxBlt9eaPgKHhKMzxjh8l/EqdA+0H8Bkx
axEWyvEukBofWwexdZor8F4nK65WGGEhnMnOYd6rwUL7h1jgUxFUYu/Xwl7Sz220
JaSPW8aPLv0nTrO/rmkjiPHy8d36sUPdZztuV6ySxnYq/TH/TumC/SrQV8gVB6rd
Mpxxtb/5yODExvlefrkTXwzRdT6yxgI69jCea366+XhEiTPxRNzDKye/ysrBJ0hg
cwt2/CK+T3OzM7qyEPdM2FHWThfVANkQ1Z0JX/EK4Gc+ezcppJyS3wQ7PanH5gCx
EtiCm733Qtzxftgi5smFFLOZhAZyzD9EoIQHL0rnP4deSTpG2D65KiHlMGs7USLZ
MOXxMaiozarJUUn9DysV8uN9iOV2oWCPY5S7Eg7cascxMEKQeN+/waZwVgoZweMg
DnYgkQe/MoRSCGKBTMw6b476wKGc0zhw1Shx+yZWmKqg6UGEMoX3QnPIgP0iomx6
`protect END_PROTECTED
