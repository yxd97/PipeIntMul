`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FN8lJe28TehMhWrPMmIuuDEp73LN/K5V9XuncQ2AIaLBZYQ/VusZ3yB5UNgcdXz4
Hsy7zrE0Q4XADfvM0rSbKWQOxJLTrUyrl06rx83hcgTINiiJuOElfUMDxGQPXRCW
F0dg+qCwNmOy7Tj4CEQ4Gt1riWh/bsYWeOcjwSBG+Y8hTt0a+yzA98aS/Tu+D7Oj
4P0iUM65if75yT5jTJSkvHgfFx5Z4uEG880m8aai1pVN/493oVDweEYTio+6CTeE
NnDvTV8xww1+jCvOHsDsdx99WI8vRLnsHZvIBzKm/9RB+Uy9aBAqKtBWagmLC8fC
J3Zigi/IiXJxiViEaaHt1Q==
`protect END_PROTECTED
