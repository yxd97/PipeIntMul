`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJ1OKQrGRFaE60FM+VOL/9L1Ca4aBiEGXo3TjYIyUliZKnvLWczEQXwIA9N8RV9D
rVUnOg7ZfD5d6hxhM5TjsAu3zmJWJmC2pwkUWDv7T6c4VCOtxM0bexzpL1K+2g99
V/GH5OqANbrAlvG4QC7XSzQtKoY61wQSBA5ehYj8x0NK7mlh5T76qEQ+fM3mLqAf
ziyTNLL0YRLARDi2LVClqxvvZ07fZ/qQBhFJf6nas280JNRckrLC/8DgzjpQMQZ1
4HAz91BJ/llfTf6fJFuyGszCTLHXxVEUb7fI+LPFrQ0=
`protect END_PROTECTED
