`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nwbnbjp93sHErFGSNAVT3eyiGXSscW6q2L87D4uxy3GPjZUszKZ2NTvL96pEroN
EeTMg53sChGzxl28U5devYIQH5p62jhBXVqOFlvH9I4Ze5/CgMYggZKlnY/aRnRL
jwdC/UeeWAHcPSmhKeLc8rZk8PqMrwMcfdf7iiif+W7BN+5pWuTyEsw46A0NsmPX
jGqHWhk8yLNUhSy5d2ZpQD8OhkKwYDef/cNe50oPQPm/gwUkpxaAKemK8s/S0BaM
ILMf1GkdZcvnKhnlOZvy/2wEW7lGSuBBryuKoGchOP88Sn3a7v+zHRbzLtSjrlrw
iygwNiuUl3V81jEaBIv5SD6inz3ZFjMVE4z9rIxyraWp0a5RttGtLh+XIEVfzx6q
p6qWtXC8b8Np7LHwp+pipjBPzHwPoWKWe2EQzGRjWgo=
`protect END_PROTECTED
