`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BzF7f1LhU6M6Yl94qdjgNlmPAAsjWa0OsxG9vneGwCnWmB/HDk/m4X/pLasPZbzp
27+vwbrz/xKsBTeIIynMdKtDh2XxjaHDOo68dUJiRtFPFDkiYfYNU93nBOxk2Ran
+N4qofLEkKcDy2AMEeQARko1PYMhtqlswNV2u7AmQL63rOIRJ9BlNKUjtlX7jt08
4Q1F8DeFIT6+arQhfYt6oUlOuMm3vcGm2f4MM/7N1rYn8GAtSTRJuIJP71mXdqT8
2s9uD42AcvVDRMuUr1NZUkKQPFLbYlmUsS1a42h9Al+VY/24cuhHk6R9xbjjx1Fr
EMs94J1MNmgq0zK66w6C7mzPGX/VtbwzmT+SW0PvUZB0qY7yTa+G3TmK0FRgDfIO
Zxm6Je7WJqD1m4oq2tz+DKasUEvZg6ar1JZhzpt82m5KqxjnB1K16hGHIzgYwi99
npWha98hCUddmkO6kDirY7Cw+v6TzYJV9wBVjXNK/CQOY6hb5BiQYsWThiRqDD6L
ltPE8LRlPvCTWjWs+hjOxSPRRksESXs77abcnWhV85Hv0o38nfVwdMA/TneDjiyA
V8fa/jL0mID3mvjm5fTz0OD18jDOAYoCU50FZ8ldkdF9GB0So6fzcHzOMsEj+V60
a/80RHD32A1BovQaa6vM97jfq0XfoyDmm9/VUga/AB8C81/WXWHHOy3EHNVNUN+f
lNy+ASftcF35DjPJd+qeM7l8Xvyw/l5yO16qWaneJcg6j1wkRr1h1ss55L1zbEAz
wxbvxIexLobFXZ2wTZfmY09VV5moCz8ApZ0CDwG0D9xdDqMpviSehEhThk/UUGQy
5xqvDpXJIupjZu8ySlCqc14eEXsAyG1TaMBgZIMqLns7WNcuQ0ZYS5c3ie5UEbyO
4CvY+x20qPvFJh5bMm0YMXeNRLvDZO7Ux9Y0WUOUZu2obuy4Hqn64ZUZ6IReZXCT
mNzP9xqnL8HTV1blA0+aqTotdK0IHXn5ymRAiTiqvRLSNuejrXw7NIQ/HyiwuW/G
2V2lx6TkVWxfGLWp9XL6Qy6oJO1+ya7wn5p9bGASV48osqi3xfPg/0HSb1qBkdwb
HkopNnbRVJnpQC9VZ+FCymKyjoQBfqVx3GZ/GsfQjCC/goDHVKIJvT1R3V9y9lGB
kTFwRWHUB0bP2Zz/KH0kJrXWFs3PRdCVMqXKmnKD36FRAW1c+LI/5Ilkb+/jJRVi
0dOWooQM8XCRqBwjXGTDGkW1QhokSr6LzOyTiQibACgQkmI49JGzWjpB8FgzEhzf
KXmsUnl3UjbUcJhMq6cur/2tfoD0IcoRJzY8wuj83EjH2gc+aiQj+Hn9zd9c43ll
H0tZHGevoPU18us420DcZT8VCFpSBRSVPsty7O5dgJ7Ge5YODZYGHkelq6pNWDXy
531/b7hyXVjERZCxK1vbGeM6xzFdzoVwsuzOUbFJXKuTCH4CABbkx7WY6YOcGtQG
g0BKCbRd3CiDs7UqMSnAh6x8QixDASvmTLgJefEd0q0keAxFPf/I+vQ4O+Y67CcE
Mvkij6OvqtXCd+AOeAJgAe7YF+fhveBcHZ6wquH78Mn6TdXM1qPeO5Zq5EiAPdxv
xG2J0KGzvsf+jRddzeqmJuGyUCkemCWqG9kEp7PYRjpsBpXZdDUSfxSIG7oiELNv
0INjNAZPgd2dMvrlyit3Dpw/OnwdHx7ql/T5WwkGzwWVaM8wEhADCMKbbg9V+PLT
zXIMbt4WQl6Om+tFUoZxdgqXNsXYBc+mlAqdmalhREPk+FTz2X5XLH92iJQvzWOP
7944CtgcYSqE6Hi3lE+BpVYpzybFr3/I9TCYtn3/TYQfyIDSSGwjFEt+hb/S7RB8
ydD+2mM4Nt6BQ5vNq/ZbzjjyByE4CZrMvRtq6v9c5BXoNsLfaLinA8HR/ZHMaZOm
UfeglSisvXltp5o6fXOHhlFwgsX+XiPr66v3mTPXd+U3Z+IAN0LNGT3C8NmLhnfi
GmRfcixXH+6xETAd0OpF9HC3VWidrHfNQJzHUDobWoL5I9c/f3hfkzah0FKlwd3A
CEFLrj/Vt2pt0mR73aXLGxDguge2/avSZU7A0wxWNEd1YTQ1lF4TxXm9PWbDRRSv
uoGj0HEabYJl7iYFgfOEDA==
`protect END_PROTECTED
