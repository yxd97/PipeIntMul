`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkaT4ZYuEG3Eb2OHKZds8fi26ZlAvW7qwx22dcRhcC01q1OlK9mm0Dvo3UBJ1ZCQ
12UBmXzGulZpUjLS3QMdky4br5rHgn7FTL7rD8w4E+mAVN/UT0FNAskvj9xzXQKq
pSNad3ONMEFyWU/+VT/NZvRFotvkf4EwJV2MoPpj6LY5Z2Wbp4Oe1FrzkAOGZizq
G1g78QzZvhCwTHEtHv6cD9jymHmyKytNsJ/pYbhtp4mQZF0ERCkE58qLsMMHlrhA
W5VZYwLiNuR4pE6wTG0nNejzOAbj1PkRBf3T6Z+i4QJtOP4jUKwMw79QVkjkXL1l
6kRIWVLaXfSOpwvx8rxH2gf980hTXs0UWKEShENvK3gK+AeIhYl9m6TDYDi28lka
oAN+dPzIBP5Y6hwiODCWQsAANjJaBOI9rH+4+vJKEyxzFh8aGENFGZ3PQnR1cyFT
tfc/x+uuDnRXM7FeN8c+Yi9Mto9Jml/t3WXoyJjVwChdie2Q4bMmUtsv+iqCdJpQ
/dBJS5XUNNyN6/VzSpw7a3qhQcIJ0J+Aon92VFhHjYAg3hUbH/YtecdzdEaHJhLL
`protect END_PROTECTED
