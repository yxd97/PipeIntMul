`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkC/DJyxkWpqT6LX0j5Tpm2uZsy0oJrkkfiEyeMKXEb/5m9vlQvXGkpeZMJ1rFQ/
NP1AYXXAzPRE/e91g5MvimzckKFNY15jKOPzn8ekQIfy6Bld3Ju6LY1Y6ioCotqv
+JuB0CciGYWLYydrYsXypP76bAnirntWcwzJu2PikoJz5y2legCRiUC7qXdA97eh
r54qO2eg/WuWraM6cChcXLi98eD520mehTreMCx39CwJfF2Y/GXzBa4Oi/GWvp8l
fXrvvbq+bLZeZtenCvqON4AKH9ixgIJKm+6+lRVDmgom2P9UbQk+nAu7ODyl6297
yd19bv4qvLMPv9pkyeEHuoSIrf+aaiWdmHniVINJwexiFGImaWFgfNq6b7JbPcYT
EedRVbojOnARmSA0PWd0xPgjeJ3dtY2TIUroYI+HivjWWLjox9ecsP/iirdi2YVj
etVIQUBo8ppJwup1hWJZuwovgeI8Qi+GQpfj+/qbKjiVM3p4n1Jj4rXp0iOBy0Ag
AN1fkfeVId8zC4Gg5V+yuX3Y4yenelsBOLRqV5vs9Vx4DxA5O3WulDT5UY6LLihg
`protect END_PROTECTED
