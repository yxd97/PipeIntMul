`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HzVfm+agxgbyq6TtLx2E5rw/YF102WdHqFex5xlrqm5PHgO4D9TtxdDcNqqpZsBl
5sKaekyxfqmykC5CbV2yQ6RHbdu0BbHeuq7wSxcqOp3ItqVlkGYms7GfaTVMJyj7
bBaFk3e1URBS7hd2/v567uYEVSE++EI7OkigANJZEe0qCnNzZoAqQEBxSu780HKN
G0RhPAb15nb+drVSAS2HnjzSSODbkGkVjhhD5BIYEJQ9oLMkX0u0gLDruRDe/VBb
2LOaitBMeiL320WfTGs0d6OmZVqleqNzd7/PItTlItIrq2eM98ITk0kE+0TmfGnK
HAWv6ibY34AjIB6iW0dulWSYt/gKCilPcjRESGueGRnV4Gmmbb+/HWGfRRjLeY/F
NSmdYuT39Qs5wqvJEZ39z+2JOmf3Ei7fpotikeidt/FZJTEXS/79/yWgFuO2ppjN
dXVZb1l7WwvS0RdYOnkKfAohVAAcULcxEPTyOgkwQuxAYW0FwRNlFFs5ORV+1Ns5
Vt2Q6yBOcx48dWXAwUmW47vzfVMLmHY1/0bt000yi6BUxH6Yesdy+s5s/GfMMP6D
ciP3EUn1apo4blF2ZxyNn7PkHs0D7QTVVPhfmznFtcyBkDFmaThNkpQF9deb3xyD
`protect END_PROTECTED
