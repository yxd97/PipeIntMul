`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QcIekNGalNDl1l2X+Do5KTU1BcaeBSv99+XRr1vcO+w/nLg/5E4xQ8CrH2utDZZs
w5dipNUY6E+m2wvvlH2mlx8ETgbKdzAdAueml1PSdtpG+NINLZxeEhDWDuyqFoC6
UmeZluCJj2+cHBWllrGQVdiYLIfLo+xOqUcvggE/OIzFY0Bf46qoYJKLazoEu7bO
AWVxoczoSV6xtWPsYX7INdnjBNcIgkt+wuk1cDWUT0M3Ab0NT3YuUGzKj/aKamVG
JPKpiKbrqw/rUyKEq3YfnuMJxTObHqtZpUBCkKb6nSQbgsKKbyPcowXNJDEcCxch
PsInWryrSmsBRTeTPlgGcGBjAP4yEoN59JuIuYS5y+gtkoG1P/b06JHpzv9PSQ5F
2vWOOcApboQE+2dhWMdYadEsW/Jc+yus8EXd7iGHxNKK9GOrLYj5ohzIaf8jqYaU
8hsTuEMdRrq2pcnPINZmz7S25b9YLwkItvbjHGVqCKo=
`protect END_PROTECTED
