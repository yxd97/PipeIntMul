`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIKWhhq/8fnJ8GXOCvw4QOZMjw04667wYWEFSrfe04sxB+XuUfM8cVJQPY+U3+hq
Gt3MzVfJCiWSwvRzf1r+nfBzRQEgEe4nOaQ6dP0JtZk3e+aW5zEkPRkm9ad6gj3l
tOeQwyNZRwb9LWUQUAc2cPRnMtx5lautuN5G0S+7SyIv93k2QGB99eYd3kZKNM3v
M1zzeOqpfwHVwDecuc2+RQ3uYVI7802GRYxol0OAH268hl1Sv+SqyudWAzsk2G+6
3PPHvPHGuSTOt46TnVpuUc8+OJ4u8RCyjPmk5Tf/gn/7mawNTV1g9k9GwcIfHF8L
MT7GG7QTD9DBJR7DaY2dMeunTl83Rj18mAZWHkA2fQ8MSntwm84q6Ouxcfh4elUt
7RiAU0xi9edYqNEQHEUhm62FAubnJxg7Ll2kitbPCG46fs3dc5Tio1GHFlThaqCx
S32UoHNCIOqtRKedeRzZVhNg/QOYD4jWZcpinNihGN1XprHrLxEa2klJufflJ002
JI9cofif2BeBhia9OGxwxZErwwFPUEhATwYA/gkc2rkQjDZYHUwsiE+cs0iSBMIr
N5+0j/Ski8oZO/myiwBKwjZrqktD7PgJ/tn0qdFvrmrrKPTmUZ9acYpr3pmZn9gd
BrpHR2yTV7pCZ6aPXx2TDRhHkMO1Zd1myCdW4qNGwTM5ojbPqen8O/TySL1Efv01
dtcTzfxKX7TEPl3uM3uOsbjndP45QQ19CkveL5SEzVaVgLAmXAgJS0r6z5EgV7v8
JGKxTCm74FoKYE47A4r72Zfie16jfePWvu/zjYuobgMSfASMU+xbxzcSzk0V3OKq
LLVPg94Zbzw8C1OhbrpXUBv/eMhOvmbyoQBetx+87qQ77Aocl4ppbi/ABi5xNg4x
MQhL3WibRHOThicsTCidHp09MG39noB5JeyUYsRNE8VQq+AvPBbT9vaPDU7XkgzZ
`protect END_PROTECTED
