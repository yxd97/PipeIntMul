`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NnYt174uDwCeGQTopv9CE6VdowaUS7+DiG5688SMLbCODQrtthfNUeXvbv8zgchx
Lia8uyQS4pLj46FWqQADhn7hPEiID6Ww9Z7Rqhu9qaSQk4V52iYwkScYS3ub8CKG
rxcbXV8S8+d9Vgm2rnrjKWiHKy2bknqMZPDXUZ6amsjX1XRp9p1hfttZEqjPg755
g4dR8yXQJ6/Op01KoLpamtl/i7z9hVxEXFFVp4hREoEF2U4+lYuAPOxFnJyZOUUN
NAlRE25TbQxW0Ldoou2Nvg==
`protect END_PROTECTED
