`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MCyApnvvrjNBKLWxPgELTVAvdOSNIZCoAZ2KQZK0RBLGj+MT7HHmiIV7Sek+7Tn
+C9aRDKQjjwLBF+B5DT3PCZJkrMSrlrXmMr/pU1hsNVWu60QgVvrTCxBp0o6cPf3
5v/iu7zwzHANVQJwvRDiNfoX9rU8Scc8WIQtYFQvIIJBDTm/rM6MrsArvOMt/4ns
umqQTNNlDdLgQNA+L2f7pYKXMhA65i0sx8gO9bl7lg4+7pW9/gavLrobLoW8YqCt
FkUdfA33m46svPwFJkITFF/Xhcvb0RQqF9+aW+3YIZIUziFUjnfG11QCcxqyx12v
8g3mrMWhdmrnBp6mPbuFCT0zSiipz3itk1LQtUWQVD8+Z/vXK1F9+UIjLjRrU/Gg
Ykxht38Z1kKm25YEkPM84bbT1lZ1CPnu0LN2V1hACy43mOxnGiah0m3h1d+9PZ0l
AYuoYuuWHxV+dZmQTa/5ZDkCf+IkHgHzHupAFjSEjjVzDq7FnjOBvZ/ZNLEQ1bTd
kUzrmc8vXb1zyyPJtdtHQhaJrSoNnkqWHIo8hIK9GuSZatMyaqlPjtKox4a19Vgd
AJH8QvNN9OJVDhttQL0EWPiwOlQ0tmYFVqVNcWM4hyUpgpLewcUfUvnuvWGi2YyW
1wO0Zw2i32H0qrZEFt1NnSVcjkG7fBSCyYJpzg55W9ymaJnjBl+tAjmq91kL9MDO
wbFQi2nlOvmLj31XTme2PJbJmmOwYoxFnO0QPI1nDEQ=
`protect END_PROTECTED
