`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KONeWNL6c98aNd6PCI8PdzKJHm5cmA/NNBUXjwPffejartDCbGxgZELr/e92p/F4
FDAB2KaFbTR/OeXNg8J76QQWerYKm5yeFZf4lKEaRwBYuq8iDJ4p6o8o5Rx4YzV8
iPYlT+Kj3/pLY0u30kZ1L9ksjE746MXCH4FDZvmRpi1uvAlWT52GZmGqUhonHfvb
+bEaG/C00WC4Z+QtFxvr8+xP42pa2EPGxZM0ZKhBtEDJMQXc4p3ZNKucYJzxk2Y3
T9KTxLdMVPlMJk57Xr8hvPOmGCLYjXHPwR5O4YJlKjImXdRrigpBlvrA5Fz9pDAW
5h8G+RfIa3nSQFmNFcMdKuFZP9skPk/a0sxO7zUnk2rtq6BOr9XdZQKOK6YC/75i
8pDd/gJ89XNapOdQaEGugKsDlRfH6qxEZEdWMbb22sZLuNtcagM/R0aKADF7ohr+
+TYGDUcgdllSU0GLLTcxiT4NI/wjtjTJ+K5esh5gf1dk7lyDvvL40TkVYrkpcD2G
`protect END_PROTECTED
