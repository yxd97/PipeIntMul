`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aHDNYjh3fg5g9jrytsRkaRpgAiaOf900PLyUEAspjNvR3W5fsdykg2YOUqHi0Hy7
iuM1s8AwiCLy93x1EUMQ6ZTTJIrOKE5qNpZdY+mYgoEm2h7+rxqQ5pZPuIOVFlIm
IpI9L2AZAtDtKW6XXXpp0TimjuuD00n1BACwYrsjpZKE1SgpL9i6fW5vnCjQpxuO
NSO9y/XRxeu1Nz9Dmv0VLtBlVlaDA95nJfxNqgaVsjmfPBI0OCK/kliRLivZbtCa
uvbd3QrdeTfYKPZhRPpYTL+Wb4yqRYRyfhuZ02GIOZ6X+m9TeSnUiL6Sd+pVhdeQ
DzsJd71Fl1pHPA3JJFRUD38NFIueZm6AjSNZY4ypY4JcWmePmscIK186s3x8/jIe
V5u4KZwO2klVSlGviNvEntARF3lEp1WXv+dQ+AodQLctQhsqrGyenqt/NsB8mtxf
Ggv65Cf6LKLbrAUURcpDfpykrZY+lDEZH2seCWfiVGry4T1Y2nngCNuyCdgwusoU
J7/xozC5XpIvu0qGA1A44ks9nib3Pz3DgvGR/iPfIVoQOMrJ7bMuBS21XM15AWhV
5Y4Qb0RM9Cw0nAsrUFuKbE7NqTHls/ITzMdOb3BUjZ+mawmdDlXxxG1Bvi3WcEXB
Y+k8/MyCPJmnjZejrwrHfbEvr4xmZSIQHngzIInZn11AfZuhFDqexYDTzA/ZKfdV
Io53ZmgyGt6/EbHJCf9W5uXh/+YygvgY/OYlvVnY0QqPOw9so1poSjCfp7TkIYBL
OkUd/SckZqg7UIuDpIeUzlZnDhmKbWjAB3XqdE5TQR9NWyqPJQEQtpGIcTSuR1Jo
7gX1D16S23xNzcfBLTPOWoJ5me5DbpZU6BFK1O94iHNLIeRmA6Hpy631dR6xPlwx
PLI451/32kMYDpMEI3fpCg==
`protect END_PROTECTED
