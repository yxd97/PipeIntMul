`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBV9tLXaRPgBAyPjFBYBqdirP4zYDoACoReC7/a8l0JFrOMLm7LZdi8uK/XtHpbF
DhwHEJjafNOgXL5xi+wJTg4ZIcRtlyXn7S93RwB2TjGr55pEzw4wR4C5PuXiC5g7
eNVRElLlfhY+ypl5PLInoDel5UvUxnzdahg3GU5pzQWtbYSencFrb9odRJv1Pz4A
XqqkP4bGv3zgu+ECHDVGbSIbyHURM5v4GKCfju6sAEdKu/U/3rLLmGyh6wYpTbis
dsYpkOdV/mf2l72FNz6w+TUXwsYtT7gTun0Fqcu2rMODPyBH0Ba8RPTonfmg0jV9
fpcSlau2dpxdqZvxoM4z7toLldEKCdv81KPpcOmdnoRW55DI1nX7H8msRTg67Idk
sne/QGqVi1WnFB/Dbp5u0cNoVxUeacdaFY2QQ0PpdGPP0pofBRoa9mltkJnQz60f
w/PfpIUQyIrzneyNPaFWMm3RMVI09g7JEIld0pUWOT4TARkbsHQfhFshvWjN9wyv
K0A6KVTLrLkrlJwlwlXOEK60bE50HXpc8DiHFe/YeJHwcTIXxa+KoVBizecOPYcF
Hdqo2NgA3/60Q504VmNBeE7MaAXoBQ9j5bTXhRo3g0KY2LjRisrXHACB/iqf6T05
2wfob92ONipoS1OlkI5U+CUKyuuEQ2M2QDR9hl2cb1dLJHfOyKANk2z7FuwI0Jbh
VO4o/13l5a/73uVDUgn/Hf1eFGwpPy99KWHEGlJ7Otg166R8TOoaEQ66T8WrIkqm
t/qvjG3CnhUqo/brCkEJzZxc/JxFMuVVOIv65qWVKbS2njaGRQ3lYorDT8Qrh+AD
KgA/+Q6fntYodhkIwWNXOawjVuH1qU5bqqBoUOkYOZ4usRHqjrJF6BKHMiqQ7mLL
jeXFe4lvNL6WuPc4V2vNBl3zkdCtvIWTlDI/40PkW/4=
`protect END_PROTECTED
