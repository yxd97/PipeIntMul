`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vcraGfsPnLru/Kfy0X85Gpyqgbln46Q5LmqvLsLMncm+rCdGbrz0y7gj2eQG7kJc
auzDtIQdPH1vbORhW8UN9B+NYL88DB5W9eicxAWsumybauHiqrAslVxDSsZIRV8u
+FJOHVJvvD4ItW/a0HJyhXIw5bKWg+bjfg+3bCFWmr5KZwBtg6IqjXOsi3LCY8kM
kyMhZMchfb0V5FnsrW2a9PQIpRyqq21nsmnf/OI+EbVFabkpsOJk81vi/2seBiVq
b2aONQ24reontWyBow3ZAxjFJmPt5wWUxRaBQUPAGZOkevHmH5+wuGAwthedStqj
ay5zxD71GudJuevMmUriXgz0tOog97hY8RqBWNJpeyAwBb/dgeCwI27k8jF8+tIr
jFekLSoDMMxkbG6StYvMymbDBBTLET4UZbBGwUiCZht4f03AK0Ax7ToH9QTRgSd7
pTlELn4oLiKqb3eY4lkPB906NhFX7oVeV31Kc2XWmdLt1dZ4+VHfa0nmnGeB1sUq
HrbX/XqeQtkVYisIeMQj82LiQ3qpkB/P10BwO2rH5S56U2olB9meo57lM5xKZLvo
+lUEEswRf3emvrFqweEYBpZJnvmYnbDWtSqAhQ3jVbi1UwPW40tXeNSxop6KTtPl
XX3znEJ5sSNIrOuwF+g/wQ==
`protect END_PROTECTED
