`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dennJAmRq2b2VF0252vsi3lVXfzc8pJkpWy7lvOSLqfWIm9W8VJ8BpTSHLUcegcE
kkhqs/O45ZOP51v0OajMWhzoGM4dZzjlW+XchjSt3D82Oh4lTHONNHLgffoRFB1z
sa7BwJANCSTV4OcNNf+TvGwUDG40r23XcmPklNgtjodzt0pXdXAfAE0UMqVpBXt0
8zDup9ApCaKj+ooyMTa4aS6+BPb/fE8s8H1wWiuuGwrZ7qy0S9PJvMUCTHdSNw81
LUEJ2CvEmH2HDVobwQA8ijZ3Y86qJaoHXKkYEzxxSA1u9X2Mw36yZdMB7WqpEjuh
xKbyl53dtC2QUxsOYhn+tRwKtNXNYAyHaoYY+iBoWRVDT5tiIT0l+Q5FqaW+D9JG
VPGRQdAm8USOkvmolXc3G5uSDR/ktPFz36o0vCEmgKs=
`protect END_PROTECTED
