`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iXAUKv8u2uTvW/O9+m8w3O9ZaE4BeGXhZHuRfzSU2wF8cnvdotx2gy3+pkgnuJBU
JWistvutOVkjRSC9R+i/ftHS4umHmV4rc4OFurz6LaM7m5NQpFlpHGoyAWBCAXeC
Q2L4ZJW5fpCqtY5Ybi7lVd/X+hl9VEVHhQQmVMFKvPyAzS3U8pvX1NfsnMWxeAbQ
IBxwOlFEp/s+4UaPeS1BLoVMK/gPmXsvsgKU3KeCGg3itAixIgUOibzt3T/8J44M
cGOw8cmCNg7R/Zgw7iWBVM9c9mLBMWaNVgtJawO1DMq4QgA2aZ7xX+89XXPItKfI
/IXOy7wvIUXXnhyy/bPoUBgsgLLA78Fm3QN9wf80p7pSb6UVe1sEQPkHDJa27Zbh
IqFWvudnYnXs06DL1TvuAv64TuUYB1aHZhMLITScXIdrYlYG/5sZ5YC1wa2Z0xxZ
uW/Z4eLWbmx5ajGK2c+z7xTbjqGi77JoVAoQpi2wBHvXkBYhptWnIUUdDJrgTaWl
YWUhuW2st3GbrNKoB2e2geUwjWFU9co9qGK+171zf1Od6+T5W6Tg8FJhdLyrPeH2
EqZY22OF9OlkbJBDOi3NzZV0DS/25TWIr6ozb8Tnqm9jFpVh4JI0UJf0Avt/2tQg
tPGBKgV4hUkY9xdp0iS1HT0Sme5etFSnMRUnnZ5OGZXGuyHXS1I1Pr6D2ZkY/7Go
sxEeu3SyvYJcQgW+ALq0J7FbMGRjN7uzEaUKjIrC1d3Fw8ziWVzQWyAJ38xNCuJx
OLU32FBaf2q2tCM1OhMMDx/4AD0P7ixaLK7mmLKSTdwJ7U6++aCyQanwaZqjG9HY
IK/3vW575T6vNNMG9RyLSKwmHJ8RkJqM1cqOXGmu3OsSEUwJhz6d+oR0fNAnF8H9
2mIUZcEcr53yANGE69Ppey7ATA1n6WT3CJUImv875y0zzZL/xnayxlZ8jBrxdMil
/II/nRlWHrnuToUmcNiB1KN9fAC+VM2Xd9BRAefZqtHUQF/yepj2Ewiq6FTpLc+8
SyYG/eqzsBzhgmMwg8KLqyRJXnQL+PRcjBUq8qwu6Sjpv+DuSbvg+LgvPSLU2zuv
O27VsF14sAyxGOPBdoV4sxUIjfJJAXHq4uV0tlyeAYd3GO36UXJOmr5cKc/fpWR3
xUyBIynzJ+R3aCtOiRSSt2NXwv+8mBjxU28prZTjHGnvfVVj30+gi1f8k9DqyYiq
Cn6UsVnwkk+wSY0/RvSRHgyBu9GzYuqH3SYjPgEWfMv5pmZldgonRZB0UFN0nKcs
APgoDEYyWHF5O9mLSLZy7ixVKtD6L75yT5HAlIHyowX4G8TGTQfORroUsmdKRKel
JcEXhMbUTNURASFosgtaU4MFk2PP0iT6S8xk2BUGCHuuG/c9Ad0kqvWp8IQe5C+m
w2fSXsLZjfwrBx9R0st1VmbV87VXNWF8zU4vC4zogvIQFHpRZnH4ufpUTWEg9UCv
wc9l3LCfopkklPAyKoTdqIqK/bNS2S5/Hg1GO7jpmUU8AJCUf2aUL/5ALMKG7t83
rmfhBaZurPtZeF8cZICD80C7i1E2yRln7P59uyL4HK/r3oAzd6cKwE3WEGtpnZC6
JDsbKuIMxfH1JF1RGY1uzxXBcPNU9lM6nTednK253MbrBgDvZC1oDiTWoSOfLY5S
886hyxTQFvuBg5YWbgijV1+8XqrafLct1GsDXGXKBNdMkt4ad3+1pEv8AVqUQJYa
Q2qMwDY0HLTnZEwiyV64jAwHM+roD8B7YVE2quAoljd78h8SqIthyWM9FL3pnrcK
Z0atJ0wG551mqFMgUI7A7aiwWC8Fct3XKfcIdT/EujiZ0MNnq3C04gTcYLOgWVq/
3AaVF9vjYzPELYDhfuWvgtBT+N+nvhPmUkiLZ8ldNIvxWZUOuTRYJKp8kCwE2tVG
kxFHsJTlNMZgvtHCPvmVL4JhxZG2ZauiNsxVG/ALDTnLrMRaYlnINLVTdPwdebuT
H7Cvua/MRB96N/FEa3bkpNF4hueMrK6oIaI6MvklDpOhs5NG7DKUakKdXuZ3b76P
a5tT3fd8AAaac4f3zrAq6awmvuXokVAevSb5Fj6f/bL9ZWpahCpqNEdhwBGmhduB
Hli3P5LNdQixiGACejrpCR6qZo3N4twX1Kmw/mbdyX8DdVZoi4QZWs6j3q0b0atQ
7HZNcqbqPW2bLIQqixhI9Jg2IQ3l2sRgg99yMYZnU7cFUYN/J6v2b+QpInR4SjTd
ZGfObMVr4nZzHSIhtt4dJL14/wZP9M0Sn3pKNzlFGXufPOYUS2xS0Amhbu1BZtDZ
MaZ8nnJDCPztcdAavC8pHSpLrYqVBzIMitWloTCGioAE5s+ZpUfkQkHLWSX3uC1j
PAoGC3cWKM6Pn8083T7WZ+Xb/iRloat2hVAIdt2TocRrHPdGmpMIZd/RR5FVZRUi
kDF7nRljmdJ7q0KEy/cAiwmWGODDk26eCPBhd/4Smimq2SlWPLWs63pAEY4cJ2DN
YdQlkXHRdiT9Qk5K4CJPZYPwsReauDpF462tGm+CiTCRjrMNRXWqx1FSo4eiJSnP
0g7pDcKCO+ct+1EC8ZyRtkForowPVaWG5OU59eLuxjbqbjGMLMAwZOOLgAigZtT3
ggMSw0LNugsTwXx5z3u2vNLWWpkUB6gIHGXuKRIuLgga2IJ4nUEgpvUVEO520FcV
BVDe8XUgJnZTlzECssRzKEaYMn1CkWHkV73buYmjQQ8GYRVxNXj8470+9dWk2kXS
VGzmoO5SzA2F8ddBEYlzRauHTYELIVmmKGbpxxAm2HBZbd3ROh3h6O5AGHXOfUuD
C+JLfZoFrzxIEzkvx0hmX08a0bf4HUBFqCBG3XKNK7a5S89vMhUXwmbccyxd6P3y
n63Xk2Em1hTQARv16eTvdSy60an1MVJEQsJntrTSmVkbSNGbGMSkl1bbKVZqyZeP
WvKrMAFrv99ORKVbm0azHJ0sUs41rx3f4U3caGkZUtjAvjYcNLjiaNDjpPWEb5dJ
5BLhB6ydsoldnU0tw10OEVzHiLDj/GHAlcb6GS87ew2KwbbeN1taaTfI08kd0xSW
62kqmd82ZRYme4zdKF3msXlZv2TWniSEMLU6/8zFxtahWKLCFkxWYbfbKmTp3yjS
9Pa21SMbn3orT2vnQ9yTdEDtewx81gDywUWOTBYOd6FeTcsXpjIrzf2tK/ndz/RF
KWPTWiv/QR8ud8NysEJICqkgALdnbMt00axCgMpjXNrGL3PSX83ebFqQHOpyHXiz
cEWSbPzBcGBimKNdZ46TGw==
`protect END_PROTECTED
