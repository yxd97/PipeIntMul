`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5orLLqR1VXDfzNkOuvGTSL/DyhmstT3OX9NY+spaTtD3Ev7cR6pzpSHixv4+j0D2
EdaU+/hMxZjjBMp4j0w0MIVH8DqVMfWIJQy3rnam1AreiUj2TbOZioD9d8z8GyCz
EB6byKBIdQxZytood8xTnAzjISqTe+kibApeEolPJ1URmpE4/GzV8Sbo2d1Dr5On
bxJ+nN838AObeYuypvBLpVA2mrCvXwWT4Y+f2HDmROK+lVgGMSwQqga0ezFgDmPt
PzVrbTGHYKW7QJMLK+YZ2yDimHrBcZFffG60g/vom8B0TdFFT+oed+tTZy7CgWXp
lxzCcOy8cheVxona+fL1YQ==
`protect END_PROTECTED
