`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIOIFm8d0hWhcT34spRQGF/cJwwILDnKH0iVJ3B1+9uZHLXrLDu1EHyvSDbjIVSm
MPaIaynRoA+NObWpZAyuE2UnYephMNeUVasVXIHIipcF47L8fG0rbnfYkxsTK9fK
tKt1hwcQ7A2dEMytXeLKQs5BXaQQfcmQlFX9/zl02F92OG2EOOE+C9ULNMM6/Kxy
yzM5MKIbsztyTASgyyWxU4LILO/PigzTqKsWTZU4mNVUz+N8RJr42B6q8OvfbMsv
hYSCZ3A1qTGMhKvCbgcFWsXYjQGSSBtFOshB74/IwAWqZje20rk5QL2wu9zC+FO1
Gzydd7Dsc4856anczg6BL5LXnblv/eEOqBJ5R9JtKrWT5eB/LUuWNoFPNybJt+99
47SqkJvHaZ+3PLrkvj/0Sg==
`protect END_PROTECTED
