`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bUyAlGP5BjtZz5ZaZ/NPATiJDsZsO8sMJSWb4cHPMkeGNVNeQghngcatrCXOfvZL
IB6vrW/h1HYwLTG57QNkD+7I8pgPSZSFemZt7Wm9bib3RJ769cbn4F60SqXMF8dg
GUZU3WIHFi5mINO0Z+RvZWZ+F4L7XB0QZ7lWoobJO1g2etbtQKTdt6r+5MAW4bgw
thhisFvSPT8OjOYWRy2MYjHiWjQDsW8QcoPF2sQI0YH083OBZfrb0vldXYFDmJzx
NHKPcH8b3kEeE7+nixVq8Q==
`protect END_PROTECTED
