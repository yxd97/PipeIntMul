`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meGgC1BS4f8HtRefKjOBQeeVWumvHsr3rAQbAogNO8VFX1zHCFzNxbT9zkpD105w
pz4+zkTocFCjQ+EjUjJXEo1OthlWXV5LBRtWmNGKZEd3cN0+Sb70yyB50oOuEh2n
GhR5lf7K5aj+ZgwwOTGIIYfLD4e/JJSYjzXarTd3gHZOX/tbo1DIaZzuUnvFDDye
V+tiVEIrFh8/q24jkkZ9WsqvPTQWz8M9no1x/q17/Aff2bQ5mFwLn0yaQC5yRcmN
VF2bXjS5UNL6waSVzB6NgdFtE2EAQqVB9lepLJ952NqRfzaGNmn1Wt7iie+iEVDk
dBpMvt2Si2X/8AT0MJJFQV1xumrGOXLQMNJvCuBOJIl/d56+9MxRcJ673mbHxz6h
pYCtyUehDVev8bhgj4HWDR+3B1VzYMwe9HssvBG8nWA23Jh7lui0LvMpIoYOGwfV
eCXfRgHDlE0fnPL6ci+CHxa2LmwGNGalgzYnx0VV3J07b0sVyr4gkYKSu+1UX/A4
`protect END_PROTECTED
