`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdG+9E/sBxCTQTS0Eg9Tae5v/Zon6bL/jEZjF0hNzbfoh5QBFvaSFwt1Wgumt7ZC
LC0WCgGYKmB3IW1DFITIwmmnqmHFumog7mzLSEeCBSX5NR32JV06mAoLnSqL+RVm
UFLpKRjnUySmCzd3ZTtmUdEC40delLer7YwrepKMxpugG722eOogn/UyyzgrL2WL
nBpGg0ljISIPP9sS6boeusj5dWI9EyEDfUVASCIMfeHGoCdz3XBCLX617SMyvM29
U5yybLfK/shwnFb3xFHChYt2z2HBaFKBYY4goKni+GZHWQRefo11QbRpHCKjXvKy
vf2o9teM9L7QrxsJ2vyfRaEwU/mmAdg8VgMYDuCw2kLD1bOEgp2JiXwJ8KM7oL0u
nO8QShmqd+OAjHhFxDtBsqt+ItNeJHEd05SPGo86GKRSkApBuQTgDtdGYdV02SK0
xg8umU0UU51TfoNxHmTcXMFqzf9tXJig9clamLjJoAMPUhdlrDYgyYDPH0ZJodh3
fXm1koI+tDmNoe2rAyEwfBpbBS/x0BLvOsSdvfQqUAQnIOyZ4FOcl4T8TkK16fkU
JBsVrd0tzbKIqxO5IRuM2v8LeHBAZ1Cwnb88zox1OGeLQOHbGVh2UZvCEmA5xrxI
Xw7rQtLMlTVCexTK9juO2MUJz6P090H+DIwgqy+oCfXFNv0WaBBXaGk7X+WYIzTX
aJ9n5HmNixqBsG4as2Zx+tay5jYUtpsnojF1coR/Tl9nR8Uo9YCniY//L6JzhTkr
y2NmYjRxy+T8pUp6eiwJ5Ucr/h8dvVZNxkPmIIqtLgN7sSgzD0g1PQbl9X7atfho
ckpYbj8f/E4VZv7nDzMQVIkkcyPKzFrSCRAXL88ciBcNk0TmanviUfl8L5pT2Mhh
1BXHPvVDDfoujq3ivuz7YwusE9oZ/IeE7CafmVVSnAZQkZQ56cwFO90vzGzUgT/I
`protect END_PROTECTED
