`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3VzIAprfkmDN6Xn3kpsiMqzVphSkMYEp5uiqZNk1MUVGx5v1gTdzFoFGK43FGMGc
f9WMgFZGfry4C4FdRPprZusILy9S+Q1tRbeaka/0Xti5Dw6h1iZqLCy6q8WnkAi3
W3pX3DurjZI5B2SiYNm2T8onUFh12BoVc6QkzKO+jnBbLFhrP6NEZioA8S0oc2z4
/+/svilonO0l0UOmcKR6t87gaV+9hqNLfnCYCqO6sIa8EHtgfNsKCHaLOjJnNzF3
TPyXABKZKfPi/p3H0hnJ5qmbADKB0V0yFAZ3kLivyj/wcbXkMdB9uHcdCo99g2jC
fLtRqhDC8O5GtGWuBdiipQqypjZpsUBStGI+8f6e0UizOnaZqBwnFz6QQox27J1w
J10S+ygvS9TTrzmZXJX2Gg==
`protect END_PROTECTED
