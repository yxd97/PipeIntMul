`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o316P+njFh7MrfDsdSsH1JwcGl/x+6Mr+W7m3YwxfqMj8idD9zYUaHvCHIWDOY+/
ytF/+TPm/KEAosk6CSuik1+8VRU1XNy1b+nGNIYz1G9XyHYACp9SLiWLpWrnmzB4
p1qL2mQvvubW5t0tff2r1Mp0EgzFxl3fIPAmZUoO6bV41ntA9m1lffs5u65mcTDY
tCWIFsUyyQoWm+ZMNOo52GfCnM5w+75E73UT3PYFVqcBPFrcJWqoQn15tRiOAov3
h4Eb13bzAzBFxxcoA7Nn7uWIiWVVMGqY3B3hOnyQ3q7LTU+/EYrdfYD7Vf2WEDQh
SjzG58Vbnipmq/mQwYLyRB+HBVoyisFf/x0QQm6YZ1tl0mO8ruvJGjHeHVTYLtBO
XcR8JDaxeh6ENJhg9LcJZ8SglrvNu7HDqlTSYWuWLXaj7ZZ7+zv5hseiorQm5wKk
yoAGUcBnP4rkQcB3xmFGSVBWWzqIKWdWTHsZ8Izv/2EgmPoPsl9GOz9VpfVeCLfZ
pRkZsi50HYaxnfsMO5HUnHJaOPGcDmzpGQvaR7lNukQsFyeH2YOs1Qif+jLR5iUt
2CyNPFgJRI+4uwOvg0OWUki+eCL/8ibGJLLIT9YpB3gSo1YVG9DQUevdClhFSQz2
T8L5wotCb4BwkZBMlqlsdw==
`protect END_PROTECTED
