`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5nMhsvPoTHLCF6Y0vHd8L7Ixc7FkmX8lsQHQtKxjZ/5xwifRYHCiKFgI9IXjbZA
E6DL5i04d81LtpseEw2vo61bTKz+MdPnYUKanl+VWrsn1SozbWc5hb3uOYa6WGH/
AmuX6G92ki75x4Gb1pZuUAUa1EKDILKb0fMNoItdJTyAd3FUZK7WWtPr6umszld7
9nLyvVTh6rDe87orcSI+6i6lasl4miFUk3MLLBIZEfgr934WwBWm1aQZDNgwU6eY
0yDD3Rf43+Ik/qaAlwuBOeH1FDDZca2tkdT9p9uOycnMGdZlXF+hP+iJdgf/nasO
DjQYi9+qtg9LmZtBhiJnZJRvBHOkupsDCUJEM3vrljzWZOkERxlRaeC3zOSiOhtV
FUq+rsQKaoNldyN8eKJo6c1Gm0JsNAHianiVkbM0Dq20PNuraKeX2gJI9H2xD/Qj
Szz6Hxpzo1DJuUxmW5qca21kWrDK1ZCigEY/2N5fW/ps9gCQnuf6cSp1yFAH/MqX
2gxTeK4SqtOLC2QH9/vwW7YIjs2DXZ/m6CWdaf6Lp0Y=
`protect END_PROTECTED
