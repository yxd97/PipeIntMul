`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Mw19tkUznhvQSpIQ3RGiDM1fqde2O39Xp7/1lTXFAfsaH83oluMTwPCdCMxrxb+
bjRvU8X1yr7VAtncVK5h8vYYEItonZkxds0QsCmDqt4qZYno41KzLYyLf1QbO+G0
es/jAvLjfX1mEmh8q77ynLqmf1nSMtzG+t1d0pVXxlEwGqL8CIJWwfMirYewpc4k
hlJB924qIpeGSjT9nAVM8NXJBDRe/dwxVcEd7z+bpPYtTk8nFROqbqmh9Hi/bR1S
2NfTOtiA3hdRJnF2Iubjhx4CTnwoz9ADA8sKV9flAruMcmBGlb65WyPSuhYHIBrR
OQIuIKnBaoRE7/siaJTMD+N05C0tJW7DCm1i6ErT8IeGEJrW6bfFXCk5+PiVPViQ
ZlQAyDp+5UmrGudctlVdh+xfri1hBSs7X8rD9t7839Y2Usjm8aPFi055tTRQN/Aj
Z8xDlP0UBm5OhCybl8sM4t4vRebKZAL30rn4HdCWF7NSri/jvxxFCbthJVQYLGYu
OA5ncuWfypra7uFPGhO0rHmu/upjUd/HNRqbcds2Tv1XsEu4fQDaLWpCmP4hIrGH
6TAy8IvYiaRrWhRVkbU2h4YnBpoBe6GBvK/ooTZlE8qc48EmGkeYwWPHv2NEGmHO
sKCOBy8x4erbxxq/TWOjBsMvt/jz8gFbeNYbaw8dA950hP6a0JRXI/AYAqkI9ibX
cSUhK1+hJIV0DPIiRc2FFUQxsX7sK85zmgLmiDZGQ0xxbqtCLlbhxycvJtuWxT+W
55dBGfhBVrBGyn2hTgVgMw==
`protect END_PROTECTED
