`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZtn/KdNeHmGaR3RlbNgFbvUKx8xJrKYizmihQaLUXjPe3QkELYU9g+aGmI/093N
JH4h73yIkDnMicKMnRvmLGviNseg3XSLA9O4NtkCdAg15WvlCEW52jR4l2b3VAac
l+V7mMGz13kmmQX/zHhZKyCu8pKiYeHj49syHbuxtKPGlRozyvb5wQT0wu1QD12F
i4lPnGG+AoecC8vPo0nn7eje7yZ56jT8jahzBLYBvUvAdyI4/LNZnBQ3WQep9E4p
RrjxGAFjQGrITugTKmuVaI5d8og5/+VRqBnxK5iUlcoBGEiQ/lXu8o3ww4hOCvrw
fzDPdBxT0xXYPIzN8fckx8Z+/wfGdgga3jdd1LkbIU8=
`protect END_PROTECTED
