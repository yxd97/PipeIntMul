`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
als29PosZjGRU8hueaPZlw3yJ1spdofeKQY4q54XbpixE5LxQ/iUnLucDyRzaSCV
Gm+s8QQWs9xOllvAJuuWQttre+ElbNZ70akYbdJGdgVNdmnZO7A0EUdbhbENAsV8
BEEoCvLZqGIfyMPfPsmBxx2yc79tNjhSR6DfflsAmtRYQlI0aAtLp6eHqlqJSqjh
MP17jOOudqI+UEsulP6US10p0w768N9vXnwWH5luuMuLqFuUUzdBmKMqqeHCr0Ca
DRq39U6tnUsnDZ9TYsmaS/cJEcr1Z1lagP6m7IZz7adcmVnjPSog8Pf8PF8PgduY
0ELQ4r+e6yd06GiJp93Pm5LC9pdtJoDed+1cb4v/Ucv7XT1NmRWaKgaqcRGkfQJp
DjKcYksHXZ359Mlktani5V3DqzDk5YF1MgXN1YzYIa8sDhon0XDkuB2cNLAsGhoi
l68Ki8WlVuLYYxear3lcjtDPlFXJMGNgt4id0V2BFHMa4OQk86QDI5rQ5QQeNJIu
XF3k/4OIDh6ZeKGDzIjiK89pn9KYtOhvFmSuXHTSaEPgaVWOULwTKp0q6UoHeZr4
U3Yq0OL4/3uzhm8peMTARInz52CSb+v6hYSXAuBrMVK6cgluiDhApHtVXw7qgK4O
KwjgitvrhtOpKt2JcDqdf+1q9KwJNEkPC+edfHh+xsdLKWVkxArX9fhnMUT1N+Pu
2SpWjWCxjlpt34rMYC4trjcCeyW7WGD/N1bhZUXayUDnZy7qbwRe4NfrgB5Svzpp
dNM7Y7/5JwolbXpCRaVAqNLiu99j9bdqb5h+AzkIzVPgUrFwhCzrmACpeoB1iZ+b
FtX5rIaZ54YIFmHkK4+FHIxoJ/IhChMH/HAcmFsTBlMPreMr/kJNTR2FJwZlN1cs
JAnHzePL1iZE2ZXoPGGoq31KZOgUQ5YhJVNM/tEfgppmiy2MVZEA2xiQmmUVXMw4
KvB6CyNtedbUYwt+2y4C1FxQxy3VmbVFhwtURGJIQUbZn7GZZ7CoGxu1mqj3+cWp
3kog2CAYy4vt2/X/e8e9h8s9GAJsVDqiwzLD5sfdWwZdmWLqrFj9T5iJ1AQPcWf0
hZOjy+rOLp+ONDNThXzwurN5rrX9fHbb+5nIkq/xhb95NhLamyBmIELTPleUMOeF
pb2OOxq26bf8Zs7W97VCi3k6Lj0z5IuUiGem9JXSALNC6L7c3IGIymJ7tOyzJuNp
Rqy8v+ABEG8aJ41rF/RU64TvXWZSScsqyWQ2T6a0BJMnBUG38S4GxkTer3CiewFC
`protect END_PROTECTED
