`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wk2uyVvfkKRzGrH4CGUGB9lDeW0mdT0ger5hebYHwOso56jnknnbO07mXRNxGr4b
5mcDf4sAEf8Fbznpv4AozpVG4Mbew15V/qsozNY1nYxSK4351mfNZC5HnYsNooUd
Ekgm/evQ8c+CKa/XG0UI1WrCsBFTL4+JbL3s8Tm29R1RApAfDMHhDzmT45FHucja
j/egKdllsKavX3q32NX6pKkG1QTuB3ZgZsmxTjkkwXnIkPHq8q0kbqw617zuDV+q
ad3tYrMp3lgTaZnba247mFQLHDEUo6LYStpXgTQ5VdA5nUqTv4Siaphn3lP1Xhdg
iLCnhwuzWB6IKTBl1Wizxo9FpH++ZYhlFIPR2vTkvuo+hiHYoxzTPLQcvfnpnVYW
z9Rhc6IuFva+5+XQZLyvpeZKk88pP/x6E0u6ShbLkQJycur41isuMcwjCPxmuSVT
3zT8byloL9qcitlv6E3rQQ==
`protect END_PROTECTED
