`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncAYONxCxbTO3D5ebQzMI3KsS1MeD8dKRoO+z0Vbzg48j57NCcPMcvoB++jKU70X
LmlNLhFrnjD1pDhbdfNEEWDIoc5fceBsIjR92Ja3n8ovcT+Q0jqOw6o9KPnwoUfW
bjaEDmzMgAtlS7yEJDUZDrAQnuPcqHMSqCn3tN98JX2AOu9SczpiE9aT56G3Bgbd
/6j4MSxdURyuiDHF93wlWRaqRiC5CrkPrbrF4fiMNk7xnO764pOE2LtqNNi2wEek
b/x5gt9iboXGOOf/kqqKXTyBuBpTYAIuObQ2Cysp63+umURqOotIf/y9Gu/pXjVU
8JTztUgSWGvPrnnWb8/zcnDX4EJ4N9cwB21eHUEIlG5q37glrWCp98CavJwUXGtI
`protect END_PROTECTED
