`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8nnYymOmM+watFPxZZ/6YvTrMJX7k0ChPZUMta0nYIrJeHRjoPgv4R3RAiPZGZA2
uOOA7Omfm8qbyy7NNFzvxtXx3eyzjoQcpMLFvNGpIGUdOM93I1okLYLX67eOt9ML
22ZMY/i54LaBLrljdFuMqaDjfaJ2Sho4iggZbWlDFaLA+ZEJB/A1O2XYwG72GK/Z
8qDeQT6vji98EHvehyzN2DgigCNL0W9sHoRWay8JOg7JLoNNVubXVyH6++zbqo+p
sycVnDfV7hqZuxwxpSnLb/HZsoK1BZmNPOFOhSy2NLc1SpHJeasA99TJEMoTdRxF
i5Zmb5dF4H9+idG1J7RQsw==
`protect END_PROTECTED
