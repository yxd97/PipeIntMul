`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5VOL31oDNM3rGeNAWrtJPy8nqx4wMEYIxoKtCqrEmGHuDTCVLKXlMZ9FsNjrD4ts
/cbiAvuXplRZVlOh6PLZN1JR4BOki2ElgGRVznu3QxP41OLPNrmADC+SAQLm0U4W
oMQBSsg/qJKfS7Cx4A+lB5EX+s9iouhSdY2TvmMUWLWCWyHNg5BpVPaROvv6UzvX
t90EketaQtv+Qi9HlwST9sLIAPyllHJDdBm3ca+vAGQ7nCUNPgdoCkti4oMSoTZ/
QBFRVyT5ZrPwDzgX9sFlXECQaVNQJfRoh+Rg3GEB/73WdQR1+pVLR6snZPxfy3FE
na4G9c5B2ADOl38jh255YODulZSUJ7crf5hnYT41JMRo2bygh2KwevJoXNfIvqRe
FT+oilE9S/itN8y+5CKCdcMFJxwSDaNK6u3S4cBm4GSwJBxeB3izRE5YBIhqoa8Z
GV6ClDuKrfN1ycUqnQ1aMhZwtahDeVhbRyf2GvP0B1wFF2cCu6XrmHlj6O9wCVcg
aRrV65L+20ceiwwvtKDHLC4KsscH/QoDb1PdhQQG5KOPJ3PAmYcMydX1dqYSPFrv
dcbd/8t57uVyBlz35Hcz+C7DFBOkkYHT1KUwr1NFb7pZjKcPQwxu50O8vB2KbczU
9TcfQlsqZz1sJooBNBpf8H9w41SzSIPE/lSeYUv9+EAUlsDBRUtVyVnX8hJbiHny
daFSzwwS0PVgeETAAPrasQF69vmpprhHs5xAUCBpBi34szIt2VkvNI1IgUIJy3LW
52tIOfwuxLI7AfcvyFqyHMnZ/aCrEZlYIikqmExfWlM5au5wJIhXFYCfLxLQrZak
tPbH6/m6uevn4Ri/tBHMrL8lt4vbUnQ/i30HT5CR9VhABj9+2YL7FQ9a7SQ1ssx3
AICRpo54NMZGZSBvPRJ0psOAVKwzuiq7UdIf2qsK+5NdTu16jOxYLLm5Icj3341g
WbdwZYIVKtUIgidcIJ8knV5HIxIuo70l75HNLCG/4WVB3onGsoDaJAHDrgW9JgKO
i4jlpZ9OByPnlb0prQfX4SdqGTghsYBPAbzk54LfZavVeZ0FjMX2KMarWY2eXyXz
cjfS0hSLbfo3/tYi28Ry/Gf7fIbROISd2UfJQfJGl/4Q7SwgiHASpkq+8YVfnTDv
XKMmegUfUOtG2JgcLAOhdaPGd3foWb59j6F5WmVPQvizq0JoKQsI69TjIv94RCfn
/DTp6O/oRi0JXYA3UQMl2iQ4dRAHi8o5284u4VSdl5SZA034k6sTjmWLNfDnaANk
/m26ZBQbf5pDeQIWaCKZD1usJw0Nmddd87ASspX51TJ9XgK9CZgtuW8UwrYxB4Py
Y3jb18dozh8An852AK1trh21co9V4S7KUq7vmQiabgoeAdj098jzRNLf6z6TAUEL
5v/5HfbVR2vFblziVGVu+dd0tHYPU9UESwZ0+hUSeM8o3bMau6LCh0b2GOpRxdxD
TgW8MnAKjlM2JVCmCdQ/L+XH5mdFfXkkD0wVbo9FO4qpyv8z/DBENsfcIWBFx3Q5
g8euqIk4wT6utUXOVVjTi3hIyZBzBX1Q6qD10ArboSBup5xQXhyEfvHrgIp3W2Ge
hA7eiENHQ9muaO+setD14L3dMrKCCd99c9w0WUJBhnEMBAu6H3yeMSBE59PuSXCq
NVpRGRAmNOjzTBJ8ddnCQoGS5tYTUKpo05/EfapoE677+FjVCHrulBxBplq+Qw/W
UrLmQaISOrDd3+hXU+F6Fr2e1ddhkEOSBlmaLJmYLwF1wMVJQBLIPEuSXXnGNQs5
j2W8RLUkr8WBhGMiSwbqF8jsjdNecIgXoGRFSW6cMg/jgsFeXEiLdY30hRl+x1Pn
44O2bAwzHqoGxI732mGm7gQK3jUcYYMp5+N7seAqzwzxAm/Dq+IRFam3bMiQdeUf
NtqOs0XU5UvmRqXCBV1DZrD/hiJYmgxTdd6MMOSzOM3XkYMTRl2xmFTVuEP6i6IW
8lNS8XyYIS0vG7ANkClKgKFC+khSJPPs0DrKnP7DYDqTHJGczMp5GrR2/TlYh40r
/5LTcsAmN8/JXuRtFzFNXJEDTnCJtyG+IN/C5IZav2JjOdv72plKYnCwaEybPZjg
otlAHDlh/4xd+HIzOsnjHKtjovrGcC1p7Q8dzeOObXgERpCwqi+d7ThcEkqx/x7V
rl8ISWWXZDmYB4ONBLEjaPu7YgsCX+Ip9nufLRvRhPsQ2AjnT1XxENGzpYZaytGc
fdDh7DRj7iRxcJx/4jbcn87V4heVB+qNWnULv2blczvy0POQnu3fpAvDRePlf5aU
t3hroJaedOPxyQMEgmsUzByCWMubw7r9N0fngRgS7pRbwByEPOaoshXnwJPPpVFx
JXxpizKN/lKcXnNfKfN16w6bfPfa1HB6JBPtUyxc6NEin6a6Nhw8EYul3U+eVZA1
Nl/pjKV2puj1B1qe1OXj1imymGcTVOFbJ+ZiIAxXUhdF3prI0dF/KDQ4pQ9ZTslp
xgg7DUdymUdcQ/MM4sEC7YZKQ4X1BZJZVvi1gvt74srXcZOrBTnlfd7NGRWDTdFj
NVkYYv2uIFtj2MHAJJZNa4BLzEHOsAI6r9bAbJfyz0WG3NbDi+9z60TtkLXwnQCK
1oBPCedNCljqMl46+PAL+/IMaFqyV9JLOHgGY1mfjruvI2WcqzpeBYlJOE0WQ6Yo
lSElL++nsMEFFDYwKwWyXBqCY4h2I3A14+jwWOlEUUA6JkH6OZ5feE0l1rtxFm5m
paL3tcKvHXEiJZzWlMeE93GsjjnsnwjHlqoH/N1XkIcw4CA5lmjnQ7aB0YdUI+rD
zRZw7PQd2ksaiB2gDKYT8ctr/FO5r53dPQA2R8/EC7gpl+YNtNJNrEFv9euWuIE+
UIWAjrHmJp5OM+51HPZcHlp2Me/p38WqI92y3jbld8aknQKqFfD9tS0xBOrXIaG5
jdG63ZrCLsRj5txVOOSXu027plcz37DxfAp5kPbeQz5iOkJqeO3QTKe4+vum9+7d
QeBkeusVXc8a1/8tyEVDsXEoj7ITxbTJLTA2rtvjSmxWmO39PSFvy3YpsS6TjqQ7
6jr6A1PukXuiAcVknxKjgb3X2Vggu1DqRI2h7d5XHd2Je6qgXPcnGry/cL9FWKBx
T2U4GczbadGTdl4d217I7GprjCPEUYNb8/pEySuf+iEYFzkeba2MvL5Yk1dVE4QW
dz9NPkgckKNd3GHfJYZApX9+T58lMffdaCdL3UgJdQev2IyiVnh8pXFKRw4k7qz3
QRgaYkH/j6FwAqNNIFSbWvyTwYctw4X1rMezAwxC0P/64Sh9AjXJDFzuTtsLDRtc
Y0OBwCWSrRI+Rnup3L1/cFgFlZxVex+MNM2i2Pw5N+hv6Vq4K1g5QQxV0YDqXjaD
c9X26uXqcdZ0o87u3Pwbgyvs8bvkfLTM+p385euL0P19kMeAPgmF+8O9MytCSUj3
RZcf9uBL1EyqgWFQs3yGiOK1XIBOdZez6pz1BqvPAbZzwpyZbXUeLxLCvnlUyii+
CmLpEo53WJeIjGf4evA2dQ/+2fT394hSJTYS2nDbyXO+CcfVjg0OSN+0e4Zkidrb
moxdc3ToFtzq7ZcTvFdzIkO7F0U3a9CJ5S63POdtyxo8f7aMHbvOAPWEMLOL5JBe
H/y7iAoKwmCDMAi6EUnSGdOLQ7ceRbswP1gMcfijdtCuSoKu0f6Gs9XehjvNVEzs
daR+juDgT7odsJrmg4DmdlPzEfnN08z+GEZebdKQUM1kBV3S4JrhC+N1f+ZkqXAp
D7aKb4v1yvqYsuFhwBolyNTKL7N06gngqY2RWdTJmlFl0aP+CBV9o2uEUkfEJsmS
ovsvCDusfIaH5K4W10xTwEZpknYqDgDFg3jCjTzZy+A0Es6/18v3k3zZOLeH3V3j
Gy+g/us9TRFR2mb9+5P8LIc8hqGpTuu5x4MonntUSFHgyQvvkB4zHOCHu+Nfi2cO
vU6lRE6HsU3hr4lxL9T4mugJh/TZ9HfTr4ER2GWBrwluHNihjEV6i8NiQYcA/am0
j5a5Qm8K+dU+m01y3BnEiXCMS/bKVyxO8tivgMbt1GbYHHm/cSsFr0X5X90lZ/uk
ArmFtg7m1zzVke+aiKrsXeL7XUDbuPqSP00Z1agdN6r5zWgyE92EzoMCXEoX8Ncm
ilcvjGNHP8vpuzSxWSo+42BKj9BivcsfaTkvfzBakTflXu3UdOKHxND4P+a6x8Qa
xJ/bTfYeejHJV1P+CkcQvL3QZWC/kliph0JdYd54yg8gntPxSm8NxB+YOrlp2W1z
kgjELqTL9eyqenyMsC2zwR3pOvFsYEt4YKO7PxtMdveBjlAFqqWNlnbJQS99Z0mI
+yVxjlHFU5BFyxM0Ae+o5z53e7W8exTvzE/oYs+jiTwt+rYsUnH+Epg8SpjmOZ/p
RMVJqR0N0EiZAQTaUFikHR3WKNc6Obdhwprsvsjy2kHyWJDmjaZYPYy0cr/HZgab
IX6y1tunup6T6gmg5R/isj+9NiNQb5oZYQoBN57ZBcU6dk3zkQQqd13Swx8yhTDE
Z44Cd5HK/GrC+oyVq4BhYBoG6dz6jlS7thupmG3r0l/zmWxPqk0BKI1ezqYuycQ4
oMa36yWiY8mu55K2fm/yyFkQuO5q6CB18onREmufaJQVdpIcd1Z+55RpAscp1NCN
Zh3BU1ZAx/WfI610zB0iQLuRRyydXyeaLWFtqpOJaIL7kqShH+ZYxWprpnoGhogk
l1IVBuGC1qpxH2dJQ4R+qccY+qPIn7m4qGp6pnaT4Pv9GwZaUL1omLQimfURC6Q7
FsikcG/YJrOmTGIX4oQD5NMRTduBqAVDFGbniExn8VqnxliR+okxBeC+oRqKgaZZ
sA6U/nogV6gG6U4B9JObOx2QFVHntbY4pCUFbXbh0UOy8JF5Uut+DU+MNpeRWgqi
3Vna+xZ7XeId5u3+9r93nz3GxY8aLDlU/1S1LqLD8sDl/N4y/6FCiyJlGRo/415o
FNRxy29foFoxjSONRoxjMD0GhfkcgKdNq+hRvDtelXNWOJD8lmeXEdyu8qg1+7Dc
VgzuFtAyrgLAx5O9uCx14mPw13URMhAIMjvy3KEVnyzh+o0XNkUrEwbo5VzdBgt1
/v/4ZofMWXXiE1HKIXmWqTe2H3Cx618Vr/otBCmqJM8gfbH9ipqCPPrRyjkwcceG
6bS1xLNGe6O6gfclgQAfiVnLqhuPyn2neiX72D8Y797NTAZlXe47fzm5OBmnx7ja
Ay1wTzGNNsQ4lSO/kXqnADIBAsDVGr/DMdp6DOG8nfSywE+n4YKKbKtkD7czwKbo
g48SibKWQsi5Tatpg2N9ijk9uKMQEJ+/dOtIrsynoI/g81iL6FgjCvyFWEUNk3UN
AsdnLtf7UPqs56uXqNCo71mzKP9P2L6tNoERojCHQbsTIW144/jHnkMxpHcsR7JK
HjYrCyDaWXjymED1yOTymvYukBJTDAnkpwCL/PrPQQ++C/7VN3HjfSLmi1OsN8TO
zVVHSBGzlXZh9mvwyOs8eSWenTfdSMc0Z4hOclQhdOuk8xuN+x7G2U8SJF/XTznV
bvkrfeJLO41dsFY7OyoZSHtid3KV7Ec6F7rE+cQBeQPtP2SOAjwmnmX4zlpmOuPS
idYBRh2rp9J1CZtzsrR6KFDpG/9WCATYvcNy7E7LtiTl0uIM1Kei2JZpok1lM9iP
stss0TTSIiwZgPJrIoZajv87J9LtKhcotnIdxh8v1mutfAyFyPVUu4+nreIYreoW
iykZoIZlw7w7HR/xxMcUWZqap8N9ao3bsxB94Sz5Zs66BKxrsj7a18PsM3A0Qat2
eUy4rAOhASfukhDmLEPoPmlfYkgBO4zzEeW0Q7BSLrLSq+A0ZdSHcjOpInsLs7I0
EvfReCl4qTpd9I4G5iNsVeS3ljAeaQnfSholX6z4OWdB07zoko4dUPUcVauKz6ST
3CkiS5IVh+phijkznvUW+YqOcs0Ph5uMMLUGcKstz8PZfQemxZsvdEDX+L+6rt6V
yaX2ByN/6AkgKfr21bAEIcwnlyzyL0l+roRec2SlO3B+EOKW1zMB3jnJIvnKTtAK
bM6W+xh2MO9mTg3vjemZNckqWp8kzRRZsFu0ADOyKHdpHplzN/EhfGY5DAbY3ugf
/cZvMszIHQFoh3ee/CXKuNvR+SpKSUi6nouaZUjBfaBNpAj4U6B/2ehKNaZ0fdrZ
kIr/cOMzKG59lVYnupcuIdBDAOf+iRPnTvS1LtSgBWRXOQPUr9AmbEYmOXeODJwu
yvdypaWwb2C/p20drN+2NezDK48oXlYaqaD4xYjMOUvqJKn2fREZidCCBflSJS0z
MEIGji5rWTSg5B3VE5iiNQFwO3k6ivu8qceU1v7xBh+T3PMD6HXcxpPEcNpK1C3t
6T3YwrVs2yzkwENVFCuZs3uAQCLdQm9S8VU3Gq0jk8U2wGOAhgfwWJedZLgZ8dw1
mqURhQtR/bm0A2A/BowibWu2Vw7/yZzbd3Gi3at0lpfjnfKMvUDD4BOXNrsQESc6
py7qYsOSVT/ajss4Tnet9DGmm9GDnGdkPdjH2QpexiqKx+Ao5cwgbkZ+QAklvPCY
kXKnSqBr1yjnqVYYq37P9yBw9kdQiUKYWRxfKiL0v4B3R4XnsFjxVlNasDU4I1yD
Uj/CAwEXj8b7Nvguz/XASVnnylrw4MUVkgMiD1Bi9FQCFr1lLzYGjBnSvDG5P4H1
Dyp5Jodea0UYlkDYGLvLrg34jta5HBw+3d76m3un9O/8joMsMgLo1TPlhoVEbTL4
/cGIOvGe1Iv6mooZW5Hysia7zhGtlwovLpBYZJLQlFRw7ZUbvwJKlxc74e7y76Mi
m+OI9ogcOwUa4OVyjGNnDG4X9VnlnHjscY/EcTTkYhvXYpNlkEmqQWJ6rEiIJCkp
HxSyy8ZHhPCQScoCnCiqzxX0H8FiPVoO6AJuJErJJpI9GtBWl2zGqWlnqfMu1iUB
DU+RlGyziTtL4W6Cz4fZxpr1Wn3st5dDF2T7ldwPijWoAWOAXrEvg3FygHIQPD4x
M4YCDBcOthPcid5FH25+4jn1k4PK4JZ1m2Zk2OnY6vLvh4cyUHqZvoOQR5LEQnvI
8oFhhVtVq2wR8ZGvneaGycKrjCsbVKuC4xidXwOmZkkHH135MTiCb4f7XD+/zFgm
sPUv0YKmsQMmHuYVodtWM6WYeR1N8n9rnxlkzJB1qXw5BYx2ktmCCr34vrBkXC/o
p8jyiuvjrSbPSQP5WoQRLyTOm2eE+4Q7gQu6IbqMlJrTPAMwBwf/wtmHFCE9zxUZ
4i+e+Wto3QbDoABC7CjfflEGBapJzYBii0PGKqc9SA0BaJ6jZXHC/v+inxeng/Wr
wMFw0HVgNOyfIMI5pTiFbQYPSIywD5wcsy2eekuhvI0yG3gMSsqLT5eorbxpx8Ih
w7vemYzGz0Y75CKUjRwVcolG9WvhCpWqCYJLPTn4GL1zXxTvZZcbImUxmEGFIYfD
htjFuP1Dq9CSdYwPBfxGNiY9baabwV2/Zx/lzyTwWutu3wRaL46JFa+8bDRmwrcF
njh0ZvISLykBb4u5+fEUeJZw8Fl2mFYfTLJ6XjguQosHLEM81boDXm8vOIJLJREY
Mc0qxVGYRgjjZedtNIsWV4h/JBbdKJOJRMzaBVXABf/e46WtqYj7OF+MM3MQP1+L
iCxipHHPQa+pkuLS1JvDVki5nD/jzkCUpGhUwJDpyQN26fEwzYvbkf7hm8ARaZ6m
UIvyQlChoIqYwLZdRJn4Iy1t5QykIeDvS++x5LMdKQEEcMbTvnCM4rHRm1ogA59I
fNew7bnCUQ0Jm1CLMsmEYtRwge2EYUvO2qulgeIjtGL6pENt8bmhsdqZl+9bDsZc
voPoukRpW8QR3/LlMwSQRqq5q6WzpGNGrRxbObx79w+hoXvYfim2hlSucI5+F9rK
vT1FH9klyp7hxxb4ZKZljI+yWGI6zhNfc4AuEdgk4NNq/Lq20ZAFzmq1O/05/8ej
BNgxEePgDw1+aaohN6wgyQRz57LZDjEE3KbGKD8fHXqg2/i3KjkHMqv4mpnkR/rR
Rw+dSMnRBLI7e9Yy+sB1LBLxUNJFFlhji/rMe+60p77wvfvcLD79JXoNcSttNpRA
1I3voA63h09BE5zYE+diDH4hflL315yRfKSm3GbvGbAwVAkvF3IDP8Damrb4zjuP
z5Ujvt/0iZ7u/tkhhIUANIQP7LgLv1PoOZk+2rtbm2aEmOfMSDuH5Voq/v0KhFkW
L+UHgozVjVyI/t90UaADMILqOePfZcnemnvmrcxo/+a+LESs7LpJkVb5rMvqu+Ux
xuv1eamlSguNhSk9MoppTYBGt5xGMx5pYsxnBpNxM0UdST+nzYAMSjzG5pUl4blx
+TmWTS1XBnt0KQLJPdVtwgrnZNTYjA87esCSr4mzXakQ5LrKW3zjuJx2AljveN2a
exOY5li/Kdlr3xlUg3wKWjh6E+/R3BDPnKbMhLkTNXfO7cZBn1S/uttoJCvQSqlb
mtJDPgAI9tIpXXJdVIKvfIGOfPjdCIzkkXr4acyDzkrwynkH5m2ybiIbmIGhysBm
LeV5a1T0tSqXXfggUUArPi/zWAUZg3wb0LYL+Afhb7sG4qHifczx6XCjctChRYYb
CbPInqsZGuv/26VzhyEtC2j9A1MGmEwIdFNkE7ZvV/Nv/DvVwagxMXQyi/YCEyEN
w4YOL3iXztjXP+hE3GqZM+P2xKHkVnLFOkftRINDGW5/ADdFtJpdJ48qzaBARKnx
QtIuAZgeJYdF2iipCAR/s4hQJld0k0EaS5YceC92IP2ey5kwzix6Mgy/UoJvC44E
sF3fvbSGtms/albgrXn0O7zXfqBBSjZDSN+B0Z0lkr86Rx86ZNh4q1NvufN63ZFR
sRLCt6zKsiPdSnncOAy4eV0MmCZd/iAW1VdJg3HQ4VOrFO0ijsupJ/P9yV1GXC7i
wgplhkk7rh6FN0cHnLfOubyKfNsz4GkcIDSkKN64KO1n74AyawpYCJ95EuudyefJ
Ukm/8tHI8xsqMxr3E+wGzbGpltXDsPkVco9CBRytE9oQwlkkEC+UeWgOSkVKYxWi
bNuqqmT9Q1O3EzcJHinsFSEcp+i5xdUg7txuf6dCc8xUykfZWpDgohypHMbVrZFV
/6Jl6Npv2XgLRS3Os5XfyihK6GQIVrrRQ/bQJ1Ph/rLpSo0wFBsjshxVPWk5k3El
ds8oH5oYvvUVZIRQbzQiv2nomEu2qoC48iUB3uvW3HajkbpIjJwxudYrb+hX+bdg
AX4kpayzn9O1KCeqm0KJZPg+LxV+8qvPigRnzvPk8iRGvwJds8GBZPwX9Dv3GtqV
0B5hpjG7V1ZWvorg+7JkxM1iV5AOJlFCTCMQbu03JL4uaICeO51JxI9nuL3dRV4I
f0DwZwMIBAjYBFqcyDaYumdw8jtDcMTQAHHZSRNjeunPa8CRtH1m6CqNKFPMou9h
sLSmZ0mOHbjaTTfYUGTbOM05IdVkJxhSpnPa3fTZlXNQHcpgXUyDbPYAPIBkabUX
9eoAAeLjvlVuBfAC1scRX4HUhc52AaUZMyNkUNv4pFjXyn4f12MZDkWsFe7lS13l
BsS6rAQ+JwKK4gGjPN675NZo0vSqhuxMvXLCcKUgCQTaQc+XcPrTxquLa8zXhuVR
WVnlOD2joPgxqwooOZTAT9aJW/trfF+T7p+zeZbSOa7drl0DJITTDlKwub8F8K/W
qVzBMxSDZbAQnB3bheBLJQ/QBEGPmGNw3q6PIlwZwU/rgRXq6F/2F7d2tno68tSA
Vui5MX4ygYZTPX+vUgRAfEH5iDwo7QVy+ZbSwm5udREtlc6wRrIm+pl9TwDdil70
ziz9Pm0wwc/PqA1voFVVMtKjnsvLSh2UNQa4JX5yVe8utHu0i7cav/LW0RnMJsYg
n9o3llWGO0ORN41byNDtV+xaDQfa+kO87AA/aVXMvO4WfHzaI0qbf5kJ4n7KxBa8
JSRnE6m2vT3hsPRR4efq1NNLyHGONp7Tx9wZ2dkw1igXHb6UjKUOCig0+7BtRsvi
fAdBRWTkEwEwiGCdVwGZ/r+z3c6LzVmLSgw4V1AWnkdFFm/tNDnPc3+596BdqypO
/egLUnUQ5YTlCX95AK8UyY3ABD7oLvzvLsHiPUzHBLBIYqKDQbdV4is47I7mSjxL
L7i8tzZbN/6/1R+6TasdjoV6DbA7rR3nCVtXiC6ge6VkEa+NawnRWMOZIo7zzZ8B
9N7KG865vpFk9lk0B670g19sT+YU4nc6FJlA6AHUF5y8SZVwyTOxuH86kKr+qVFj
9OJ4LRy5id4H/fkvzZM3ed2sBdEeyzNIlVpQGec2tU2DFIDAc9TVOb+iyXGlul1r
7iZyhZ/3cn+6ZCNWgB/ovz1/GJ7jBfJxo7E9+izww/pojN1PUnnWB4v8J/RfTPPs
j+F8DocZtbJ0QlPitp3FRI6NAQJbxl2+h2qQQU3KUDo0VepLwFbDxvw8vtPdjvgI
jTeMcSKYKf8ILVqVgGCr0DhqUqimNFBPVZPnObG7rdcFsv9XtAD3eKfYFvzXIz60
Hul+BsMaCriRBMGVPxXWaeIvjyEDlBBsnh4SQuDQdNCN6maQDEAYcRHnBjySba6P
8JYcOOWmb/t+s4DAZ1QTwY3xQDd6/FPeSAI2ltr0Xd7V9oDQs6ExqYSdPn9I0t5m
wVqYTHBM0rTXEoqmOhE6Fd1mNrljbwcCiqDiAQvLd+JSZ1nmVY3FHr5RKVYUsXlB
bv029H82v0l8uPT+huNpfsqnjEnjH4YrBzsqb1POfV+2EajhN8ZgHxpTVPkN5Hzy
tZNco/iJFpGE4AqKrV7vHkU1ITxhDPXnLA8VRNLd6fJfBD1v6RKBSlfSgYBFE3kx
bShMWuyZAJQjts0SzmJnLe0Z8FJadi1szoz6Y/MEYbtps3a8XD++XJ+7jDmS7p9z
SWmXf4VAvvMZWfvVKB/TjEXZlK8a8A+d/WYFtIvf2qDs70gOvYRg5vQGtWVVDqhP
AjkrsdkTai3NlrZMGqtDzxfr4rGmKWLpb5CirJNCMwl85+7eAPK4jsNkRgeryRBv
M56TZJFfvmqiNJR2uU2vz7QhEfAPgxGvNsg829LW0EYJjW2N3eBGRikp1mgrMkqG
elTiJNGDVkpU7AG+I86nHTV4oIkH5ebXkEc/ebj1g93EPTxaPGJfaRLgom3JszXP
CuRI5Wuj3OvVyHea/6egAhLgjP0Dzn6S4OkcKMD828l5eOynfrzHMnc7oHiIqRXF
FUGbZEiX/6Q361k+/ManOyA1CMCfrAdHYo6m/SUeLoZ+NxvzSRCjhd2acs/Ds6iK
5PLBt+/td0xCdjGBjT5uxowb6G+8RpqqpeUY0m9jCl+Y//TXXoeFpRezHVYd7z7N
apuRXBp1k0PiHUVbqcag4KivnegSKfnPLxU6RUk2w9/XZURqOLVZGW7TepFS1pfA
wR4k7LLUbKU3ttrkMoj5J/4mlDZBJVVZlgbvv6b4STo/8VNzC7XKLTomql4Fuc9p
3LYpHhbBJQ3wzyXC8mlZnM3JiUfyf/W2od4oamAaLM88yVwz2LM0XeXzD1wDFCmS
uMUBsHcwk/KsdwzB4/vMIyJIK3ZhTkcN/cwWJUjFGN5xCSueNXVxipAsu3dHI6Nz
6ObqIjHYxf3fq3HU04o7P17e+O5bqLgzA2wGRYerqLau+hay9kaWDacQoDkiX/Tx
5mZoh4pJXL1IZGjTUlAdpSAJrmaJ1WsTJqDZkAHLYdmkAHd7zYFd8GclHNePQbh/
nF4gtkPxX/xGAWwW9DSNfb243K92I3D23GIUPIsJLpl4LWBltZLbKKZImOkp7j9F
Sqf/evVS1TDu6nchThAGepMLsivT/7V2IHoMd/83G3JPqIDZqMcu1cZ8VSRUiPPP
EQy5nkFVbklM53vDMF1wJx7ds+Ad4u+APN7Et8OClb8n8ZNChT2MSgZuiH+k4Z6E
CBd9APr4iLfzGjXk363wNGJyiQRYG6+IfJXCTJV/C6fP72xmOMGlmv/L1N+0L3ZE
pzinQ0QZqRkoFtjlj3yo72CqKRgTPC24JJTvPE4+xCYpbs0W17U0AHZ6QqyTUTqx
edniy80bBFXoEY9/Lvtj9UDQKooqvOfWV1bJ0topgEexKoAvKugufbMdiGFmIvst
yUssiMiH7qyfg05zOgSLyywBjGNrCDBmbTvU6hI3NGQlWPtqosGfmmB7O8Uj5lTD
IoI0+7O9+5NnN+fRVjgg4TJDPfeRS8LBvPuG0A8AAOOgklstoUK40/2MNMfCqb+S
IxDmR2ZGGIgt1SYv4E7veanVjki4CjVz2YiCvA4al7zVk6M1CWN977O+/rEj7FAq
/L8KQvln6igDQk/WqJ8fQ1a06zT9ReCaSKUo/jtWtRDvEOFBcBQ8u3xyFCGfd/L3
PSU6mDztLvSesJxV0JHUO8nW1KnNv9EtRGN9Mj3IQcM2UpzFSbAcnDXakR3ysGov
6KiuRPGlGqhGG4BMnPlM05d5od0i7IuvDuO0wVSzx2kS+lcCNagvhU3sR2CS+v/f
KbSeMj/J6qBJibUo63rIcb8Qs1cJEZlrCboTS8vIAJk8L/W8hJLJWoeOWR8z2tG5
kzK9MKs9XWb9RY+5t8DxDoRcNHR+0yZUhINZWoFGJEXUnt/eq5wKlSCYimb5sC4M
W/gFRd1s2LPPvGzwDmnmYoewqnWXZksdi3N/ciO/D58jqEBCQR1gprmXnAkZAATf
cAIk5r5iuLFE4xgh8riouLyHM0hyVMpiiDEu464MkzXn9JgI9vL8GPYH5f/EhrfR
qSsehddSVg3F0LWTiYjv/Zla/i16quEtnV2+LyKikrQbJu8GIF9e866gJOuyfo+J
6FA06eakAo3EpEpa3PPVV3kiRebME4Gm/4sLdDrYKFnqUy0NMRrKw+JqwQ9yaC4p
SzAJBrSnqK3HECw+D8XVmgz+pTY7NmrUlre3S4WoL5vcmkQkYjWTILMkNPA+b0h9
874vxIhGeKT6CouZ+TmrPcvLoHBsVT/gDwawacVM0Wr5GifPuUDHVNFrzQn0zWa3
+61OMTomtBHX95oBWJzWAWF+v20m59MkyMegXkkYZFpR65jPcYaiw5/oqg/H0G0F
45F5R49e6XFuOoF7eJXHrf71rDHRx/USC4ZnzX1YmsQuTGGQdw6ukIaxN3SqSX+l
ylIa7P7K2Ih/nfRuG9KGOAicMQKkYLZg1lOxgytUPGvj8KDGCI+WK2Drmj7+jMXs
vvr61u4NhT//pWI4i+5EjPDWWxdtpY0Fwnh+YhA+C68aWnYClbAZLzrwJBWMuzXx
LM5MVlOF4kSPXJdkjMdxDh274cnpyji+8av2Nh28r6svXNrLBEgHUp/hQj6QLXUl
ycRu73of76N0fhmehA1q2CN+FYLrr9dRyahs65xT7bQpWTdVx6bSlPrtWORaiGlH
Klhgps9FEUN3lGi06VXza/uFAbOczZb2eSJtraPMZPEDx5x2tojB87nB69RTqxxc
ySzE7SaBw7lq2CBljp0usUJoG5hy1HwpOlm//H+LfTz8JHZcBk5W7b8ayltgRR4C
aJ86BKP/9fhn4KsOhZ3xVyP62bIa+yy03XZ7oRUAKRelEd0hKiLnRW2nYbPfaW6e
r3sPtftmuxDJLrFyxAg5JZuwcSXqAMjD52w7EPO1UDByMTHS3KRgIDTjB8H5J5K9
u0AFDqMqFeZ8a4jPliGR5TYr2pyIu4rSAmxaP1HdAEyj1Zlu5Lkj+ju/p76cg7MX
CrdZZXRnY1x0ivM9yAy8E1Bqn8gW9/o+PZrTpw/ehGS7KPBmYif1pZrM5UXaSTU1
djUw7mxsYc1hiVmI4Fl2c0zf2whdFmPc02FmBeJuHIVDfJGgZH0Gj2fTwvv0/r8v
4lHGhBSSeQqKxXc99qD+uZDe/u8KpMpnVlIRS680VDxIg0TTk5S87edOxdrjwGHO
bRvFEyAmvOVRXqRsra8RWjWMyak5NsfWDdggP9v7AJVlsv8O6sdeBregnj/aQNe1
JuCkdbZSiwIPOzMzTLEfC0o7M941KXhRTEsD5YiOujExcRVzM95hrCNP7Q1aHy4G
JjJDsi0lOVSnDnqPnQ3RJkiAzbZrNXkeDSS5tIyPTaPff5OxDOWXNnZ4cb7S7ZPy
YojmlwXtNguoK78+lYqnaicXZdHa8w/la010+7UgAYYBU0AMbq5HJao+Ee57boXJ
ISdFNHKPNldHDPKYYG6XM3IB0FXQaM5ae5jK7Ib6eZZFXuMCVtWc4ckzo6Zd/1RM
0p+zV5hTbct+07wTGxJE5HKCzStcYz34O6TxbZhobwBibC6iTchZVQuOVRsqo7co
DZg17w0UlDbyGbI0Pxk76BNXHEp+XKrHk02/Fj7ohdZ6OwNiyBstZy8xUYVVE1N8
3jZlCMzogZlVPL8NfHpwl4bgJLC03oU6gAatfjgSp0Vg8l16trzrjc8PolVnedVo
2g51sSRYF4mTNZPfkJTsOocfvYjbxx2OY7WfUaW0CKNXM+bZCoX3r4C/WVoTq+SX
PzQEhcEeFmLl9JcvE6hCX0MtcVTDf6nEFsF4S8U/t/+M1ryXd/X3O+ItOh+EkUya
zkUJj5ArQy1J3nLfyagmTg==
`protect END_PROTECTED
