`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XSnZ3kG3slPenL4ewfvYTuICjO+fKyyKYpbLEQCFeyakAJ3AXwgeYRhR2YP1Tjp4
flxVHOjweVBPoxpvE6NuVii6+Vtr7m3bL/ESjmK5mKs9W+6+YY1McxoTAryuO9Cs
jVELHIJUokPHChegtmSWUvzgqSM9WhHwXTrNgz7X/JeFXLs6UVPbTMLqwbpom8y5
MHSuEeJS4YSF3D0QzFLYLJ28Nm/o+FUTgXtuHhBv4MwI1+cazhv/DKgpDd82tN8+
y7Hxvcmje6Z2eV1j/trkyN1WfDbWBdpIExfIDYP3SJrE6/6Cfm8qYMdH8GQjaUm8
J8hz+ZxhKxcHoeyDicqeVkCrSYLJktSUqMSEMOX//rDWlQC1HR02hzbePkIbmgm9
`protect END_PROTECTED
