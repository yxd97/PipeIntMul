`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JHimt/fVt8ZO7fNtPvUlhpOxpHjMDl7xHQ5sk8RqbHtU9bwL99g0pRqeWk2x4QI1
51f0JGhKyAWa8/kRMBRLtKi3idqRmlcW7jP+V0jlisGFBHEDgIDzuraBmYnAVbsl
YLWpa9xhrCQ36cAZAvwWBzWHb6YhC1yWQJMUzFF1n5L7EbIo4NxMpPMol60FbAyV
Z4b1/A78NA6lynpr7UXZpuJnMFtmEFYPeu0rwbI1kc5G7Te3+GDFJo+0uGe/LU6d
wJNMw1OQswZt8MOm3x5kuk2NdQLjXQ1i5ANC7qxU9e49wLfMgmeChcTC36z7uHgt
0stj1+WkADTtSAJQqPqvzSWRcmHTmD0FoApa/bZsO76yprei3eePzqNOjOPtfF8p
Qg4481BMFXghUI80c0TpVH/zxpmL+O0b/4Utm8pz8jS3qoDKNDEb00BRBPGUqYjO
eIFJPaHhB1nN/25/YEin03fkb2UlAXK84inIWqe+fNhL1bcJAHfR3+Ki75K2VhQS
CxQoGhocXzWnO2DtveUM6/Peq85ML00HAFyRl64PhS0uFvWDnmXpJbF81wPHvjnq
PFqFX223gSe+sKlZpbSCnymR6XOBtFr6SkFqBN/25c+UiS8T7hMtBX7XjpLQIgpr
FdY58xUIg6HgqFdQe4S7kvVzruL9gjRdh81d+Kp7DgQ/ZB2R62pz8VLZTolJEE8O
rhCS+RvV2UgusFZGXQfOeyGCQ4l3kvbowt5DUvMfjxtb9IG4WLIoHg8lFhp5wwvz
7MEHemTNcf64tIIvbXgStC8+nvChLDppZpvSvNPwZEM=
`protect END_PROTECTED
