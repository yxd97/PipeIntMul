`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0/cDha8UayJ8kJ5HQJTuLP061fcgnrAR9+BVZLzaO360KxFUr3McA44/VEbAYHbJ
REaOXdake1G1OOC0qSynEEj3deGrkIQTfPFX8dzHoUyxf4hqf06jAMPz8dilB9nR
UKpvQ0J77F8/2wIE9CNRjCFu9AHpNaqqKrKfy8OeMk+Fha4iOEPaGxpZ/RFQlqiC
vmr8G7fdNxXnykv3FmBuDo94zq52nq5xuwUU4cN801TiIa+BEa7GOylJEFrdh6p5
ENSKrOy+gwNTqg22b9F4d0k28Uv6G9PAhntuXdwjIgEEVTae/ZNod019Gr4MEnWq
rIBZSU4mjJm2BnBwPWBbunfCnTtq6BIigRMTOdbyh5kT2fdDSpfOJ+kHVj5SRmEb
c97qk3ruY2q/lOLBLRrfzvVd3hzp4XkR+5pIUD/uvU0iVVUTL0Un0+nWWAEYUlWF
7jsDrlPoQz/Egn2/FUBK1Snhs6DWKzM+TIiUYHxDJIQD3YT9LN6qb1Lnkw3FMtkY
Ta9jWEp7eUL/+/15216Xi35I1ijRBVZwLyjOfY9C4abk93l5R/eq0gNlJVr2xiux
DQhv9uOUPzzhMy/bEIu/5hgQGjYrKpk1qYTu/T2QA2yq10wBDjJZzh4/Fmcdwi6N
rJjV3wgRdWb2EP5YjKSvnX/vOR2DZywi/Gn10q/iUFwLLreipJ8BsU0BaPRnQoRV
Ltr7+dkFw90AKtV2uJ2xjbPIwLaMG+zwqcPkq65tAS1a4rk9T4YmStj/NZQ7qfaK
Ca1LLQYN9i5b58QGPUDd7g==
`protect END_PROTECTED
