`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ym86KbnwQCayRTUgDKOmRNp/tvNW+4eh7fZJ/dcvFAw+IFxYgEZJ7UZvPt+w2zTW
5BUiciIUNeMCN7ZSd91vVs+VWK7ezialVlXPJROUQ2FDs/6tg0HU/1Ened2Oj6c3
ouiK1OkpVtkP0ECa6lRd6g7S/qycpZ8HY43jGMEYQ3FN1XhWL2y7hTrtsnMbjOQM
xybJGJh8522zzN/TkvFRGZGzZZYRaikxnhILth0OZlIYU+iKnG47e8vCeTMfg1yh
2anh3uOswiAoMz9pWyk3SFUEvZEV5NhWTUCHviWTc+floBwikHVazmNI0+ykOe+K
VHvihk4e29n8LinENmsHdWz5JwNM6EqU7MiQWeBjd+OnvG6Lyp1f4aglDO1s9sIg
msbCPYZRAWHstvFDB4u127kubNbxn9xoS+U1rPaY0S0ynqBVxAfFxyQS9mnSKmPE
+qFjLQ70a8JAVn4jfYaSMNqtQvUH0sKedYo+oHHxxtZ1QY9PwdFFSwBeKr+SzWU+
rYMO3sPxKbc/U6wqdv+3/YohYb7swaJfgy/sZsL/2UE1Ko+DPJkLSj/AWUhURgCq
4BglENZkY7KtyA7iWCnYwpwcPHOyKVtTaSbbgyZu6hwi3VoB04BGrkEnfM6Je2kN
j2x4QMlC2TfPtGXV3zeX31Azd63Dq/Z0OZO/D8y/nuzrsqzvFMTQGxvuwBwWVtcy
N90f0X2ETNiF0UJ5pAzkkxiyEgTlr0RSdNgb+cL0PQY/V4cLweQ5X5RVdOZXEa0l
3RCERvMxTefe48qfcXNiKAaS+Na/ffbLUGe0JqjW4iv+qwpAwzc7vL13DZaTqxAC
IK7jNjFlZ8dEqhG8nlC+/iDNfTlfHbTWIGQyE2wgTkPDw7JF9uO3ktU0qZurr7kX
E7RP2yquPtrHWhXvnycezxPuBwstUpxErBg0qzAHHlWpy1u3w1KSmF9HZbfSKx+5
5DrhVEQ5phSDfAJxJHcRn8pKpBfPSANjmNFXMOfzcQinYUD+91KxcaIgbDOv/r8T
`protect END_PROTECTED
