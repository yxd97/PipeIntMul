`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0y2C0N0kLsqFD3Rha+8jmPcopMCkFYkgw45bqiHrR10zws4bbfem6Rbo7IIEP1CO
pKDnWkOydcUjPtVjEBhb4fzUhyZ1I5ZCVsmaNTYuCmNNMvfz6iLL9V+rqP5tAqhr
sG2bZ/qhfqs6KeNr9vFEaZ/li8GpL33h6DPGt4XjJswsSMdvTSYmNLeMHvtYY/3K
6M2rMyD3Dwy59RpcX2tDrGXnj3lPURlGldGudxJKplRTUdNRnYSAAejp7BVSF0zs
MHivyZrstwi3/78q2DcdCp3Ys1YhmeqxnEt2OrkHR/5CSgoQ0uC6nIsIPQTUXj5s
qSsr8FxHVgPf0/Kts+HyQ43LOczJKjzhv7r75JZH5agGJRNY9mmBMlpVP3FS1Izo
YBJPDOSX3D6AfcazsM/nonKlNhxmVbyTBHk31k8whAnCxFM0f27fyULu52pZjkcw
AfVNIF3GEbC68UmO+fXOSDWTrHiCBxf+MyUfZswVrn7YVChpRWqA53ODWhaNBgAm
HxnCo/3NjznJptWRncPfPV2hR/1vAEIfNPWIz/0Tl0TDckA+Ra+ndt/HXk/bmLzq
2jOGMz52lOEmbtho1n0dskx6/enZkgH1A1F8mBEvcmN/XIh4A8wgjpIkyWhaXNXO
1cDmDoVUOqVtfe+PgrgHlnUbEJJUNlKUYmAXUXWf1kmtimc5RsiS43/Mty7RlQ8P
uSOmdzAXagh4X4jH6OduovmVxvODtIwyThkJRt9ryMq4Nv2SUp1M9j39l6r+mW/D
9gLSjUvilD0m219n1wuucdBbl3gm50RAyAr2TRltI/Xq/shLB+ml2EoCMf3I8Vxh
+LcQs1MhouM9Bsw4pq7CWu2Fdtua8Vdn3nNxMATveqb8vrDIaMsmLiuiVFNIqOU2
uuPUM+kUdgtZ+B/XW5Cb95G0Zgha0FeeYkoSub7OnnZ94JZ7PBP+gc5cYNjC0EzV
CCUp8ewYlQ5I8AYoG8oubFXzffA1bcpBBmHGpia+lNerl+AAgCg04YJwpdolZR1h
zVFMHUEp6EWTdvczTg3e5t3p/X5MrR0ZTwE2Tw6SVWUh6/39Qi0dDZApSGSexlBH
C/ga+GA7oqUSKqY47+kx08u5fm7OSO9wu1p0yweXzHhsG6eznOKt8gQpOxZwhSxu
BgbDdDywpmqXYbB++w3K0ypuBOi2aDZhZ64gghA3mlxgYX5kXOEMXazSGdAucX8Z
Egj/usDYXuX3/rkVnzktcI4nCknmXKFXbV+0+lvUU2a2p9prB1of1ZD0ucPTw9Yr
TAddF3DB85rRyFO8Ey9285RcnntZ2/ifGiAdfDgD0qeSDPvABr3Es8Sgf92rX+Jm
S62nKUDAROUjpVI6XeQ5O6dPv/cI8ciyc8727JiwR4G7BIwruNG0u0G1EbYn1IkX
A/hyngEX7ZO9xGqp15CtNt9NKnOrctPwk4ByrA/+iDBpx4pxQHMBpWlonugPFe8r
KR6UcIUKawoh8sxU9iPTl9CTnF7KnX/h5TgTGln/xd6112ih5A0V7oU+4rEjAXjH
gkMfHY/MroACSmryKDUjN/1cMH6pF/C0xrUOyyPzN76CyKbCUYxoJC87K99unHon
ncvuSgP7gBvq0eYjifH0f0LwcnzP2Hk8N/cH5tzF34yaFd0wc8SIv6ovHdC07wzN
gyVT5iO7x/EsOQEz16qQwLwgjLMcLtU7nVOLSd48N3aYtlHbAElYMEUFzjPeor0H
4P60J8yz/FcRZftZKfrg/XEY3jjzzfkjtI2wqRtmkxhTrt+LXf9SQ6nO9k3HEOLZ
Tyydol0+UphnABrTzVpwv6lmXf0sZj/jznk/O35h6OSsxFL+/MdQ2/Bskx0jb5+J
Vjx7aEz1/ZAnaiJNwHLk1z+pJ9VA+OcJIFgWd7orwPOfYo22vaPk00v0EgfdcelO
Tk5LoNkAzqFz+FwzW00tswkWas/JwUCZHZZwbQ7j6F1T5VhYrSQ6T5CIQopHdcLE
aLMk1jYiyp66E41X5RBJ0Wfs4EAcAIGYWnEwUfoKh5ocShzTpRsSLYbVBikz0jzo
eQBuXe/WrXvAKHDhqAyWuCVNwANx2vHPfwOn7SvZnQfe88TGLS/50m2ggiqD18H3
565fOZtBQoteV8QPH0qXNToVYhyt6RjtpCNZojVc2C2jyU3VLLpiJ6LKEtIXth3k
R40qrcfb9yCNCJaVfpj2oPWeDlTIZdYMul67DBKtcCXWTyBivl1xkEkB9xtBwhmY
+LECZa3Jzp9h/pv4/5TxmToyGhfhW+SpXCKWHQN1wuasnEniaIPionxEMU+tqKfU
GixRVdBbRsSaGbzCmx+lX2xRn6dmVTHhwgKcrd66Q4q3pJlXL0lcYZeLwNF3Vxyu
3ijbCNDyITQnOdbHSn3ZdHbFZYbBfkEPbt8nIIm1Z+apB609DY2eiWWN5bQJh/M8
QtaGbaesgC6ZKags9hTCbv2GtJ+JAcOS/Oi1hiiCVKCYnvpMMJ3UOPY+xREnigxa
nt6FAsnXe2qfDJKJT2krHxTXfQlUZ4gcewoZ2QhJ48XW2QSGUfr9krlyW+Js9Kdx
0yshSVZppBEfxJelzZ+N02RzEcwgTVHitCgKfgFWOfflXZmKUSsV42PWi8gP5zpM
JmwnARAn/xzSRHxfOVIkgpjuqV8CdgStc66obLk9TmyP1KG5qPD+dPfcMgzw47xZ
CSVOZ8m27+3CCW3rvPYlurkL3BKmLTH3VwDEyuVB3zKhDZvVE4W5NZTLxvl+UMoY
+T+b9UCxr96TMLxDXRwezw==
`protect END_PROTECTED
