`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ewRYTqYFVT93AcZ/BMLlUdUG0TKisr7DpLbLz3Z6qriidpZWgqmbgxlwQm2PmXGG
rg3cF0aY0JPGtnN3/rHLkW3S2EWAejwokyjwAFr9wGQ7TB1RB4/IJHPTLVg2U0pR
3xqgAZyTCagaa9LQejhYvLlSL+NR542P3wQ5sDWqbH9Hhi0Gggh6aeWt7llENA8G
4/e+s79PvfVYoXOznkPga4QRRrsuRpGcuXL1TTioj/9ymKyG5dSyLhEPlvcJIBaR
UstsAA4JcEKitAS6rBAaHtO5HWf0isLGo4Qu3Gdwm/k=
`protect END_PROTECTED
