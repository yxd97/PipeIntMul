`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwTMzkEAZufSmo9q4JX7IHXSyy0GidxAn2lM3TgX3NX7p4RlHnbpBTrUql0VN25y
CcXhMQglS2kH1XL2smDud+ncuxsfn7WdANf8Z6T+0HFcfv7KO4bhx9bnud/HC0Hq
KRn2xLAzlgN2bfhUlwRhmXbL6GlLJre+LahmuwOeUUNeqtVZYQKiOo/0sVrHwYRX
NDXrIYagsITMIVxlnK3J35Pt6cWn2hW5dgOlxA2oDiJuO3RGi8hpnHqI+QMVJb2B
A2L99o5b/kglTCFY1SKVUwjrhvo1vBOaSIR5MgDS6BUeBTK9YOKQUXgra0xDc2qM
Jh821zQdWiJdM+8n+Y5w55LoSP9cq8JS+9lbbkz6cIirh7/QMHAbt/Dj5W2j97hQ
PLAtBrJ/9JBkoQtz9Bie0rR280CxBHS/XDf0ybBnkK3r4dcs3Tm4ljL8DFjC7VTK
AppFRz1Tt3UIY0ptiabmlqAXfdS2FROsmJ7ItxNnnppbErS0tESykVsar0cBDx4w
Yd9XM578eAJ4tNMaEwLOWrrXxyj9wj3cWW4zLb0hMTdtS+W6ibDWiELLqn8enuhL
qkiElfN9kbEOMR1JkQm+/slF8HvzYqKBMnmcUCAUCi3+l83k3kJHDZPrTr/Pske8
P8k7nTl9S6RmjgbHwedet7lE43ExSa2TK5YRROvLHtCTcWos506yOmOH7HKzJ53l
mBMhrv5qJfXCkwO3rHJ67ee5SW3SRkofIu0vCV8JrJOYZ02KyHhdSgUdHFufx+2t
7vQtDB62kLwjItH8mTDngS/dGtOZEEeasKcakDIZ7jUTUa1sLyqU4A5Dtc4G2nTQ
Vs7+qg62vvX1nx+Ah9l6dPeTsi0dbNUm9RtVCXRR+EaVSJ4Ri0tBHC8GOBl9unfr
hCyPLgLURIot/q7Y4pAWNICLSZHpYgyicFsPfcxZ6x5jlTea9h6YKssAuA+B9Wbp
63aW1v3WtMzvs7pu/Mm+VlzSMjKPMDoi1Kh4QgfX/sljHIajU5VDe9uXqO+jmvCH
uPnChgRN03DVh6k+xLNncw==
`protect END_PROTECTED
