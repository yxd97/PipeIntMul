`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VWSwgxx2uCcOBi/Um69M7HJn4J7pahDQzBOjH47g9wd8kGzFsemT+xUolBPuZ4dP
8f+ZneGEGzvxrfPtoqHMqWEdSSfTG0k8OKG4KDmE/W6RoV286EbNAC9mMmuVkS1b
aralRYlfXTilYZ01q71NNc8aqAZ5n8QhUjz+osC8P6iA6LKzhVCwLjQqbUR+qYrZ
8VCH1FKJK0Y4aEZ43i9ky1raKtvmELfo113tryLSlroFuR/c5Ro4sU2gEExES1zO
7OgepUrYZqTQpiq4clM/o4FK8zLASiBayKgVSKAahrd+3b8OnHThOuJYtcV105uj
X6edJQpYvZY4OqhgJN0A7OwKo90thaVu1U8LB88udymO1LJUfZ2MLRXCqfMM8GS2
G7K3eGjp8DmMH1Vf0tYBtxyyWYRXC8qPmPPAMsnqkAVK8yegAIYG4kj205Wcywdd
Bf1AH4beX3i3vU8LBHBc9F6HO1uP9KPv6K+ubHpkmlxOqvMCzja2QL2X/xxdAG0/
ByvPKLoWoV14pE1vCVHpeQDCBUEpPmgD64FcQbq84OhACeJW80sEg1StK1y7W+kY
ypKcf+/Bj+UtRsqZ+JY19VKeiwAb93AmX1LrOBmMXYGc++oJ9BD+T0Y3jplpbIHo
TkPnMQvqKuI6Ej6W0O+7wGHYmJ0MJe962aTWlJkPHdvV13eTi55tQiPadN6Si+Qt
cnZl/JSBTGcTTxn72NvAQ5bU4GkjNFQf18ztQdRH0IySrixiMstZiowGD36/Yt4P
GDwU9bo/5pP1urXwLHajkw==
`protect END_PROTECTED
