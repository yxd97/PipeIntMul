`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3j31EKygKmckoMKorKuES7GWOnR8B9hMgPXtOHt6rY1mIx5dGcwkh9IfBJwsk7pu
34p8WIFYI79QsHZtg3Qv1ON04ho8Jcufa1COfd9tTBjKxv+/YnScfyrp+KJmY64j
S88su/HFDioXJCPZYPTNAZ2Od6rusGBXLqSOabwm9lPiRwGJX3jgwGzfEVxSbeBD
UB/Il6Ezps3vhFB2+B4mZj9eXXJqJFiaWiQsXu9nrnIq0DwgTTE5gWYDqJekGbAw
iJtFW21wS0KbAei+qDWOC2YXkj1WybEuVWOiJ1/oXDZlecx2u3w1I/KgAB9/N/uu
aAZJ+nqj1yAUiToqhduGyTPo/vfUbE5qTIQLTU2/RF/BARk1Ktwc3lE5HMsdbiOM
ly+s584zMV56NPTxJKWIRaVcj1AJ52MSLONituQet+tIHJ5hqLlZNe13D8DyQ6Fk
lGvhK8aspMhyDvefgfCmiE6REWsxn6yDZDAccQCahcSeBq4ksHWkniH4WjnWnzfE
vYV3SAHY3vDvjwm48GewWHYCHVnhJCzgOCDzAMa3GtiSpdVgP8GCAw8yND0fH4ZY
ganqQZD8ywW7yflnRi05w0yik2YmIg4uRW59BwHeo+8rvNTBRMMRSTdXF0VGay0A
d5YgCwZJ0pcfxnz9iMjWbvWwPqntTsp8T5xbrY56mDxIASDiJAK3kZ5hkplIs7Mk
UMVm11iRguthDSMzDkHOq23okwAUbms6rS4vffo6BXU=
`protect END_PROTECTED
