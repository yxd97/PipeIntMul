`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h1c4r/oB0vfSM/oBUoSSa345Gf7492AYhpoFDimT2QUYO4HEfy6TePylamirtDFe
fDChPkKly5ZCc3YypwW3YaSMfCoenFaT3xkVqg0Fcpn4XEXtiujpMzpWNlFnRNHL
H3FxXPwO6ubgd4YEdhl8S+iKAKyG1ibWNAnXLw7SjylStZv0sOdsVQBUW43Md5uu
Ne4wk/OVCSjkPA9MSacLRWo+3RfRQQYFjTggr7yBsDIzMUXpu8dTWZDorxHxgaaT
k1dJ9ON4J8pIjezA1NI+DoONIoftFWEQ90B5zWVmlKls6pwe/d6clFIy01yqwROZ
n5lsizte8K/+8RZdITNStMHwPDinIfyVNgGgK0VyKJDYpXEoC+ggiNdXu32IZMsv
p84mbxWdBjjpjuu0IpS5wCh44AN07id62Z7zc+GSD1UrTUE0pvh/dnHvOt1uuvqZ
uDxyx5WP5G4ZnmfLM2CvciXIYQvyADa4PnKPksIhd7SuJcYE0woKxoR41Dljvu90
fa9/TyIpIC7GQ4JMHDfDprW2LQDNyZIwR8Q0IqjHJW6vY9K24VhFgdlw3U7qxOoh
/VtiZgFZm1//8CixqPhqUAc6SzYSSeErTflV4CXHlEqOqCPzRcZ+aTTEsM2TZ65s
LtQ5mRUm9LmzCAbbKNjv7IMejPebSA9XeVpCZ1pr9AAkY9G8rdB5W63t/McVY35f
1du1YQokg+gWNu3jNHJT8Kwwnlm4Ch8CaFVs12G9X/87AagrTz2NActxVcm2tn6N
1LFbR+8BYV1/719bs2QK0BWLFj16CmfC6F0HtQ/bULTQRLRh0BQ8L89QMkg/d+xp
2aCh5Xqq/3H7wCO1TzV5yOIpaqyb38mPHZx55DkZglDCi3QJsmAJBgED52R9metD
HokJZuDGW+zlYZxwIVFB/LhchE7nvugMx1ZZMDVRTey4zGSoNh2Dzv3X+/XWsuvJ
S54+3kT8pa4dHSSOBnpSs1k/1X9OsgCr7I6KmdiXoa5F5vG/Z/RsmrT3jkmvT+4K
5O0hiATqvwBJerZIN9qRYhAogcACi7Og5eznhKyrMHzDL0mJVmaX1/9s3FsMDO+B
C9vPdUt+UXStaqpIqvuQGQ==
`protect END_PROTECTED
