`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SSj/c1Ym3xiKt88wcUzj9rqJrbp4GcGEdqS7G0XJFN5jgapB3mhoJGwzIr7JZ5vM
dwERzxqrfrEIISpXyfI5rdtnzPOaSwlN2qWcyJ7sKOxajcw/iksCFgqWg6cst0nh
uyUF1G5t/qBL5j7sRqpWiJDpL08BjkXbnxEX9g+8cygwV7UAmf/zZx2ea/cp6zTJ
Ao7gMEgOVKc+ZugehWlCKOCphqgQU4/bRQ6YuWBCz13TfWt+k4+hwJGoxuaimG4w
QctlBL4XcHumgT4XzxLogkUWwAObSO5xOEKjvBYdo65urFcy04jpEmzWVecbsRFo
bCzTaNtRaFFdIaxpR/a3enx9csLnTKF2HBxcZe/GWD8=
`protect END_PROTECTED
