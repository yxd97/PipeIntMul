`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IlksPMKIc9wKTvp2CvwpaFML0wd8YNEmvt54BuJ60CkG+ndss79EIanUxN8lIMFC
ZI10L+L7a5PL2SRoKSdSFbEGJcoXhYCGGp7ZzklRv+AMUHKzA0kuXMT7csm8kNva
DQ3Qu9b/24W7LdNUEMKNk0svnv+iqPl5lh5ystb9TUO6Y6pWjSc04/oFzFThI+hI
Fb6cO96V+OF10d8tQu0gpm8p486I5+AHEejXPM3u1mjkRpcuniKNmoTwzazYYaFo
3ytkhKCAqyh1kFZCW7qRoZTqYumagldm5Ba36l5wsNqpuddUUsZ7+mx1CN32ehdL
VMVfIiZIn97bm2r7Dz1bIq9xP72nM/xlQZ1vOdMnGDijMZQdN5Pdb7Xfp0Ee9hVw
uSa9+dLoDy+nubGXzO3QZjV5af5KBbebK0cp2EDbSC9upGrP/J1vNmNMKmpwwR8z
/Nh3W6NzbBc1VeQQJvNqulxaq49OoYx7TVLh/Fs5pbH6xRRNvskXrPxJ27L1vnB3
`protect END_PROTECTED
