`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xnIFfY6lfNqcOdBSoGPDijlY8nfcFQOfphFgNSKTqNtfaZkkghnJbnIFU7Yg4uCX
MII8xwDy8LgrlQAOCnGII5FKTv5ZG3VX0r05Z+iTcvkPDOp7V6P5F0sXFwyTsJMm
NHRwqVeZG/wkGmy5CcuaXd9RuebiUjHzxlSdMKiBvsESEzRLgelejBObUlDdG0uJ
azMz81l93DKrvALrtwS7/UzLEmg9t5A/aVE0QZcE23Pk9RUkh5RlRx4rNJNlzWMj
wsgkgU2Avf/CWP2bI9e/UUg7rsbJdUNMu4srxKJVZQRhM0cvLI4837r9zSxiJAx9
d5auaUqXLOYtISN5TdxPJvXG2WEC2GtpmHJb8Wc9ObMPMv+KBvVjNwgD4snzcPER
akMvx7sglBOla2uuFUwEEAVyfQyu6kF0QNSp73c8T5R/p8GMMAtwADw7A1CegIjF
GJen6iynwSaFsJ1H/mLe4K6FyEUy+58BSS8oUvCqusSIfMO223P1Xc3jHvcFOeaD
YAyhoxGB87KzTH3ppQVfXBOiUnfM1B4GVDgZmPdm/O28QwlcvJBJQ/ehs1HO2MRp
ScTCglD1QLTbt5dAUuscbsHc3JJhAbRgkmjGoDft2BRxmPPJLC6Hy4Yf2tWN8m7Q
6RANjG7Ui/ZLgJqWhhR2WBlZ+YmVn+SFcGFNDWHYQ2oAd7PmQK/a3wBaNdssCEhL
oNHO+4XhJqQi+w1x+kXB7f7hqZs9D8pKLukuNuf5qPSSVxg5jSvzz5Jg16P30TeO
gm6H/4c2tcbvwF0Z+Lq9ue/6wy+LNGYobGEWSMG+1r618DAcJoAAO6RcCxxgCeFX
vIO/j9WzBwiZIfFMNB82hiOmTx9o9y7T6TKBJ1Lxas5UQTrdpWNCecsUvq/GnfDA
Rf+mLAiF2ZKv3s1WopAUmaItEgUCqXoCUfL2uyNYbRkjyKHesFtqvBChyRiOOhKP
blOELU3MlT8+FufPdaiBXcpXK2E7a4ZyMWCaz1eYgVGlSTg/33cP4A1Sop+KFAYo
2R41KJ2S1tPhkr1fywRzL+zjMN/pzrBbeJn3a38bLjoTJSU2VFdJyM5X1n0KLKPk
NpjRwQzjqQmdWVUHH/iDL4smdacac7HO+1/SsTG8++fBtsaNxMuSWq9WWqpMDtmd
`protect END_PROTECTED
