`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0JGgUYYHiuFE1lhyboB3W3/9SvYaLHSGn5PxRn3gWllFTXG1KVHW88BRzyFDDD5o
x+1XtXlUdfbc2gl2ybBouaeGbNzSI2y568vUwIOlzT7e9LjkYvFShyobKc1QxHrt
Lq1qWWqoQQfJvx26QO6aiWKS93VyAF+d5EvfC5kuRrx41LPMJJMtXl8ionKUbn0e
OPkLfHzrW1oYPOlXtMzyBe8yNXZq2ci0mZchQWooNK+3PdrTuXYdz8e2Lye+6pTP
rJXDfULfU/WXKmVkFpHt6jQvQZvg9N/kshbHV7lrb9xV6p2nOS4YVzncubC1vhMB
lNZ+rMyVrFKlsPX5F6mbU+HdMUk988uIukpemkRmsWPxgLtFuqSnTcEELsWogYsy
HQD9K5mrcV4aFAObamlys2aicNe3Zwn8GpG2NerTh5yXhCAVzN3S2jJa5rc5/caT
YVmy3n8Oq0pR/6sPj0ep8sVz6+NGhzE8FIXkC2KJ+0jAH9jtrINOempEJCifv0MW
zkAIQBgUFhiJv+PHjdmDlqBekj1h5Tw1Y8KOKv7umkBuVCGk69hjM4WaClKK6LxN
hV2QK8baIZHjWXWJU/WQp/glazMeSNe2Oje/mEGC/hcbD0ZMjCxIOSVc4ovofcuv
mRIlsmJ9VujYW2Pbzb/D+BF/SVP0dWaFGk7HweS2O0TBD8KTbQ0l/bJPXfmXYD2E
ku0rzB1xJ2jOUyzgj6SwZ5/vwEkngITJX9A/ZeSU9/es+nl5/woP9rOZ1NQmTZWj
M7rlfIdOP5oZ0SCqlraVNIdLZGl9qlqPMtJL2IArCtyq5rVpSdHxp6tdppzBJsVJ
AcH4lTSNxW4pIuu+465zZhUI7CMFeqskuni7a8AA1lxDmfbKxecjHY27X+zwIwBb
PlbfCk2Sh64YHRxWlpKmLnG+rHBVQm8sMShxZpgf7O79ou19thJCUCAUFUIVDK4I
`protect END_PROTECTED
