`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qgVKTvjlql8Uo6ADsvNwxbkeFX4ne13H13e/3/Jl+Hz/ppwX+UkHEafvvgNVDTb3
5+OCdD8liSZrkA1TQXp19g5+ZA/49JRg26uXoIrlO9LS+pY7ZillrnTD/tQ4JO2z
w7qbqqsRJa2ugBEBfRhITgEQQJAY9J4rQJYL6KGn9OvrRrQah+Ckha++Wo2Sw42t
w648Jf+YTvV0vAHA4uvzwFWkGuyrP7eQkcIs0ZZHuTYzCP5QBRnJ+fjb3OQSa/Oj
wSdj0E5G3gj5OxwfHZGuy2SpVul2NDwXh+kIXNMtXHhXUcFVvYmgO/8yinaSqOdJ
AGaLDK24voPKHGjXHBkzQIa+bj+HMnOb0IIJl4NnTVmdtNLLhFK03WgECSdzf4mB
iKQnjQWovcbRE5O91Ah+rJJNYrKLwqFkM1p/JXL70lLxQcAmAuBC6vUEc7QvQm2s
DrF0ozATYkp5TUN47nfCbA8mLL4LMnawg9X1QA8zVLZLkaTzFGy7DZFEJEM1R31Q
`protect END_PROTECTED
