`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SdWgM5094L5N8ZtfhFz9/JfWfhotfluqNeUiJiRhQgFi4ppQHz9216CtZidXPmzW
K0lGy4RC7W1lr23UGEzH0YQOadyTJH2c3rjM1rXd1YpqzN83eJp8Oaq6kcbLfUgp
v7WquGH/MdoL1C8f2VFpb8eXys8dGLODjgSEIzD7yFczQKIeBR8fKSikWUJ+wx26
AzuEl151ajuK3eYSLOZfC+OIsKqPyaJWYmllfrPyCaP4oxF9QvNwIer/Vv9kGkxM
od+Xr0nynUhTp1MD8uQl4lYfzFpJbPDJ325O4Zme+bAcaa/pE5vV84gBZvX4qFg8
sbsnl8voYZBZYc4ca4TURgcQDYvaVrsQCdAAywG85v211q0SJPskZpupsVEkbZ/9
boN4VmFEybGcoEIPmtOBEPUN2CJywvLz3jRfRFziReBFpaRNpBWQme6Qbf+Qwn3w
2rjQuYy9IhYYEXHoZshM+ucot1IR9agy/oge8gzt78ScGLxm/MQbEF4beZ+KUc6I
0AtWEHNJvkqU4xSNMoAc9bn+aJ/pkcIGlHpUSLcDe/xreLELRVyVUql2ZPiKKD4E
nunaonHyvq1xPYhdRi/WKQ267Fc5XJ2pgVcSOGepEzatIAplbTxglFpBVxgh8StW
yMjlKpjo8wpxGN30rRCLivFQxrlFhj9uD2OVoYhQX7+e6+X1ea1FNUZ39u+WtQ3t
DoisQOMQ3raFXMQNfYavnmgGMqRpJNnbrbYf0V+dShCKiY55ZUz2GVnO3cExermb
WtpmwNZ/hHnxof/UG/CMWw==
`protect END_PROTECTED
