`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
khdIacpzy4NNfZnFZN0nVttexHwBv04QEIpFwKTDz/gAUkLJPuTJSsrBtq0PRmyP
wqUikDWELFJt/bFrg42nOcMGJ4FH8h5Kn/TeN9NRQ/HMKz3+3/iU761gQCs31Hfn
HCLMEa0rkBdUsvx5wkwZsyP9jut4psfiTdwb3dJAqFaIDdRbjv+0B5p5N+bKF6zi
0oB/cAY1j4ElZGV6jLs43Ibm+QD4yJ8+Bs6VVeTu9InxMyUNyv4FUOv/QldTUlG8
Txze6czQE4IoXvjg9yDjx8XCuiOIW/zNNzIHUXMD8U9rjzCCQ8sq7xDyDhhFko6Q
+30RuV11fI6JC7QM9FMY0uSt985iSRrU/W9I53SHTwi4blAfMXyrjN0Yjrl0Nsn+
8126LZIPYp1fPE0KvrLw95yEUOPM3+zW1ig5zMeiojW5LhrkxQ+37ws7JDzSN7/3
HHW2AD9tsFFxCp4G5snWe7Hgi/07M/P3vYB9vFRrVcQ=
`protect END_PROTECTED
