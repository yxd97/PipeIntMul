`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzhCJBhekB0WTX9BG7SA92DvYKd5AsP2MRRu3Xm8oalNLv74IEcBtDwQL9PY7d/I
pvEHtSLUXzJtifAyNjDqLO6NfQLJ9kuxh1VfgxESSH4qwHmfxZ0JouuF3o4dwC7i
598PA3taeRWByGekde7c+Kv051pVxF7Oxe5EXJcGkyzixDE1GJxkJVN+DU7EVL/i
Z+cEg9IsjnbJEO+sso8tD2EfP7wi2p6diH/GcNpGncw05qC+o+7iYj5i8wkmD2L0
Cs525rp3w5x3MagCPglQ6P2dYbDIQfNn0pYQcVxb+zOtIoQ324hjywb/7vcyahIT
h/wvJToWbcOlSFvfMdqoLIxUnoSYC9E0c6XBcbuT8sW/A3knP44d/GYx9ZXRpKDq
8YI88LMu3S73aT2zfxV6isq1onyZFYXdrwQLQBxlLPGy76TonrwHsu0w8AcMBis1
a5wvGyjIfbic3p+nvQMl0bcV+1Rl5a0GWtECHiObV1i62Z/PI1y/KL/Isyf7iGIg
UB9OT6t5/weN63uPhQvX/AVksocNTI5MJCljX/7swMbVHXYrdRUWW23lYImEOGkd
HSDS1d52gy6aAOcMEawbu5a+czcgET8jKOfdBas92fHzV9YPTHjeMYnwPvsTQAbS
KsNlAdtUDXaZcvxEXhkxk/zRLiXN6Os1ZT8FFkcYhBL1r4X6ZbEnPWOhmy8r+eKg
5Z3Fr5RKN1YhK98AZS3C6QLqFAqEi26+B+jTST8LnOAeyT0b3qNPe7Mq78b+CzLB
BzXQS8vTdz9pOYdMWJ3g8mw+gc/2TdHOfd76U7rqL/8JPxIa+xdu+zVppbhjg6cw
c6r+TbLT4xEs9qCYA6m2Jw2SaCxydfbV7MrukIIOM8joEGaGo+f+FgTLlf9mHtP7
jqvVppV1FFG+xlBfU7fsWN9fuLAiEBB+ayhxnytR4LEBrJtKbt7ZsPxwn8rAfEke
`protect END_PROTECTED
