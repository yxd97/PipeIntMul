`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8G6VIjHq29OaKHZdRAzeqsLdjcwFeJKF8ktUl7BF9Uij5Aw6R2TmbaHaAL8STTj
6RmZxlL5JYCa1o6TOv5l4aD+dZGjOjdYtEhevzNaLEpOHUoZ2afnIngatV5tSC4Z
hEtWasw7sXKvVpmzuWzTH7JTMUa3LpzfdxvUGpIkQnOyg8Ig48o21/Z+fwIDOEj8
KIC2li0/qf96MXZh1wKZC93s3CH1PNgJn2NsYFy+ZYCo/j07qbvywk5E2Q/7Yulk
P/My/4dAc1+i+2zFgWM/xPXlGa+QzEGX7TVZ+r6saNpiTQ4g6uE7UuZQ+4uXFRFJ
y4DAZsI01ImbdU5gf6xbdTpoYxIifPXyQQrVzM7NfI3otgDghVE/iBCQpfecbsab
q0Dus9ofspNbLocaPGtFhR0S7tN6N4uHWDbsS6A46xtETzw8pjdTsF5+7L6ckzUj
fBxttMi3ZQlNdPQBDGU5VtDvZtM8P3j9ivWvrELw+GklLIH5e3PCcvDl3oH55xQy
yxq/Hs86uP0FSdVASRwkmRdtrec60y0lMXYEGiYmXzaEP4O1pUAiudvIUwUdF6OP
MNyRQyseE2nGE6NrzaSTSidI431O/x6cF90wLt6uJ9Me9MEAwe2v5btcBuEsShMM
GkYpkWY6gIU/sLvUHbwW/iiyrhSNmEEFTRf4ILvcyEnFJhtDgbtKBNaEQUeVOejd
`protect END_PROTECTED
