`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wEzd559FE5JPt8Cs1NoEVSTso7eSha8Yd4aYa9jfsSWVCiDDuyjWOkMAfdSvTFso
wZZAUUfYrgU9YCyo3js5dpyT7SU3UB0Lwh8XEG/L7w7ebW9yhW/7iCs+MUYR30fS
ugedKiSytiuvO+/AOUBS0WTBBpUvq1Le3L2uaxDHG7H/A89PngwGZMeH955FmaGJ
PsUzg2QuPXrIW+0PNctRUgE24vrA4e4JYNvF+wpBOtZIeCLUQQUvC9hjP3Gl5uIW
u25anT2HiZvuN02ZtuayCucvD3rNDPQ9MB9muquIor3bGbCZ7RwgjjcH0yQd1RtY
9MHtx/0glAVUbuYBhBMQoDVRYUowDhaIJaSRhGgC0isL9n0FdnvpSShscTlXMd9K
47Q0I+ChBhIzPQ9ADaFiBmv70jEFBLk8S+IciYijbrcm9I/wt1Y4GgLumvBwR9RP
pcGusV7v1dvmPqRDbEjd55dhtbZpwBP68Sqs05eENfoi+GuiJYgC4xeR9r+k1Upv
v+5p04gm8txFJkNRWuT3pVIdyTZ9IMLPP4VTmzQzMaAi6xChjj0Cv7WzRua5sM8z
qDQF44F+v/zIxovKwsVXOJJZDPF5XzoKirDVXuRFM2CsyyhX7zAsU+vDKSr6TRKY
wTqt8iOdBFN8PzHHqDHAodbV+0w4xPcaBMjf+cl9U0ysSiMVYyrVG7KeNRvOkC5z
FG04CkcUAuaD9GqCEzo9IkwcdhFSfae0ezhFN7sELa7r8eduxgnp1t6qhj6FyupA
qcLRDaIiD/MybTEF0xBetZ+AzjanToHwcpnSpl5gbG11wnvzvDTJ+mQEeh6+jH3b
/sMuKnqgjra985J1d/tcCkDfgh4U6fUys9/YLYQwZrKKNZnaPss7MHk2gfbbEXwg
gCwqzG370nOhA3S5UGZi3kt1nPQEUNmLnxP9H77eKlTqw2xsz+7lSL88EMizsiOF
W4EEBjeq7fbm87QPuD/pYuPEUhaHSRlEhJediOHxltZxOA0Tmp2dyJq5Hdsuw0d0
1jgNWPib24cUIKnuoPLSTJg83evTGnbIZSA/9FOpNQ3pt4tojVAa8HFJTYYC+rd9
AFm85ur3dOkNG42Lzo8zwCD0t/elAyj1mVeH4TXMc4K2eL9tZb/fHU++PswnlnrX
J+IbYNGcGjB2z1K+X3HnZhJBy7fAUfeaVWTZmaOFGnI8DSQPxtRsHtdLvt/329sW
YWzJ2oiX9/D7DobJi2RtfLJjvpxDIybAYb9WfGIvOMed+gu6AT7oVpqP3uAtxYkE
VCQn1m32d8E5QgDq1jfw5u5hVGF9lSWc5r+b8qi4YZJsD+uW61xU2u5pIZmJW60f
72YrzadYiNAqfF8HSy2vYd/1GRSzPpe5dfK6q+xP/xfG98MvpausYaSkgZCTtgbw
nFaY2XLPAx9S+v1Yfrokaa3vt1J2tQv0bV0z9ibz6sDQrDHInOnpsFjVYa0ba6n/
FSX2lTPAhwLHvYHKK/BiW+GlzLdj47ldpSvYhCMjcH59ugpWEc8MDUSuT0C9hjyp
adcE290sWPwyqQBxnQRveCSoDAv2snnoRflqGyy7PSr96MYuOQ6Ag4CyO3YB9pLl
4QMaZq+mW8JBpYs9WlnI54IXTqdS/8yOY+DmnI7yMJ5pPKKyyoFK4laf2YaFphpE
VKs2opCy8uApQ5x6KGLagKm6RGDxmVJ+mHFJyY37KnrDbBGsYqdBUa43uzqi+evE
q6Q7m5iy3QdlJAWFzmF3iza+a+LqugvhskHwqidgg6wyox2Lm/IS17MEh5pUcCxk
cC048OOYYTYxRFcHClstX/ZfVPZn70jvuAAJe+Zl/ZDyB16I12Oosk7fACC+ltH5
bE5hleIuqNwDoxGUAy/gUF7XRJBcKjG5SYZURoEmKQ2BEn3RRw50GiNNqW6bUgfI
lzwCUSuZGJVo8R9txhMspy4JEGwyTRVQen3hEmnPDQP10wlfFv48AyGenHADjKVo
Z56vPtkWDjagtF8Jwb+Sgj9FHM/PWRVMKXlWaCmZHFV2Cp9XScu/LeKsN9sGnnzP
9VDCIKTs774+Aj17FNjo3uHH/+iJLeXwfuK08y0h23JKp1AIHI3tfPqroWBFBggl
`protect END_PROTECTED
