`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
USyH5H/KS5NE5SUi3+FdlnbWcC2mAou9i5QT6IzJHq86Vi482KH229z7pheQt93Q
pnPdRWZSmG3XcQrIhBvt2NaLf1l0iGwRtz3zfLNqWqhf6dix9evyDTFfCLTUekQO
W5VQzyuXBLoVi6vJGfFLBJpJ/o5CD4uaK1gMIcFRJ7vH0HkTa1LOidxoXRtNKzEh
cD/b3S6tTm3iFAIG1TsAUyiT9T3cBPLtnY/AGTK+uBUwWPotI5uoDzaLDeLIEpBm
Fo0WktpDjwoxjFMqnFPKOZ6ETJEn2d0j5AXtGDceH+6ER4DK68idF0O8dmbk4uo0
cOd0i8lo5pPyuNypg7tuCsA39ukocSp4BP5AkEAIcuP5ONwYJk/coiNk9zH6D3X/
`protect END_PROTECTED
