`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ItWA7aZkrcdQc2jMGBEUd/Isu/K95bl+0UQcgkNDmw8Lze6Of/kY7FgVgxg4zos
w0lvfQd8f/zSpU6t5z7YwJsdmGjQCmajBWgkS8ElPLQ9XTIH5awzRB95cl75zobw
0fIIvOHT513OLhQ/o6vb3BnDXsS0/72LdYAmhG5JshkXtxco/5D09tocstlyQdTf
LG2o2uDUP2cKveTpg/saAvGcx+VAQyjWZZKEdgovulRP78IdcxyTHBToOy2yfW/C
qHWymFR8mhWb0jC/jaAN7sWCSiKUlFPfU6hv+km6Qgv40ZEQ7/SEp9qada55ULcZ
fcBIu0eNgpWQ2PckXNOhNdRCLqIkg5FeNvsGMPaJz2bNcSl/Jvzy8bvT88eEsXBq
02MlRsqxApmYe9N2wQGcig==
`protect END_PROTECTED
