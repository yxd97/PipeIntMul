`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wf+eMFnCrPMaGn1uHXDJj6aSpNVlFyAEYSVQguBxWjmMVcA65JEKUHZ6VZfDbDmu
xo2bQxODO5+P6o3dGwWe65noUHHB1zRHtxLadxIHDiF5MUbxFvveKPKdVYVu4DGw
Lt0BaevE7064ilvVpKVLXw/yG7IzGui2kotvj9994e8hbvKrcPtHRCaugDT3E/Pn
Wnxct7rPjjglesJ5PnnDAF9I4p+Xa1qhswrEvty0NkYV4HFO9njzU90xgtfv43AT
3uGF2EBQvfyZ7XXV/rdpng==
`protect END_PROTECTED
