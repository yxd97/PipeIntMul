`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6i9v3bhyJNXq0QHh+d3tDmReB0oei9pOr1bXLLK+CvdsrKWG8pH5zxx7mRaGnHM
Z3GyUjCPy/aEvkWkWE8UFsz1zKMVI+4SGSGN0FV8xdNrsTUBm6XmaTwxIpEpIGdq
ikjbd0GzQzm3BE2lNPqsa5l4q33c8CCGIZr3PMlyu7K8g80wjVwsTKge++HCuJPm
xEX0ME3oqdswHcc/wVlBljwuWvRTeDRim2HKyYbc1n0LZcSpWErxajmACtBSt0xi
AGdFzkPTNzboR/Iz0xkH8GvdP58zvlmIXYoPtZMfoys/+eWDgD0OuvCgNd6vHlZ8
59fhZTezUtQ1eLb/dootRmufpMUMXK+cIO7o/lFJlNItlwzOWkN/mEkfH/k48BWX
/V5vADHKhVWbh0TtaYZci0VFXlIvAQ7u8aZdsLJkGRHP3F7CtEyiK/gwhCwbblXt
lbKdazG9lIB3jye4PCy0Zw==
`protect END_PROTECTED
