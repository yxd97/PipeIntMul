`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EKrOyx8kqZLEaw8t09ff/yRXujaZ90e7lPbLV7w1XJ/forhu5We4hCpV1XGhO2Ks
NxuNROzYAAKyVd/QUYNquBQC6hUnYKj8Oo0Qm1Fs8V883VO9lEmpSbc/j0ZLJ53o
mxbB/58SsjrqcPrpwRnilhZ7l8d9udZQ43eAUULg1O3pjUSRk6GCT+9ZQYGu6eh2
xjQurUlGH1+arcJiEDtLtxKQ/FtgiyicvXwpu4YvrQ12TrnN35MF9KEXklS2E3Yp
4rxDsQo1HTd2iThT7MaRaQ==
`protect END_PROTECTED
