`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
np+R8V0Ra+BPkYDArJL+Sgk8alEuF9BprrEHG5QTxssgIuSIQFTX0dotNK0ZFbm/
6NqbEcUBd/1xY0MgYFjGmgvxHVVWT8YNRvHFgjjQ8WPROEqHSY//xr+Tm7M3BYek
eKEPe/s43wCTCQwmW3MainopVoThk7PURr46MdlqdIdjYDPd1Brpht362nKx5ZTo
LzDfY4EHol8o+ktALhQs4E49itZW5vVS675ECEeI/oWb3q6t5n9hazW6N9/FC8Q+
Xv5rIXMuCQkYCCpwCeZC9RasG0mO81ritUcGj7f0ESXVeaVy/cN1k06ptZhKXjj3
xffB4PXDlcTkyPsRCs8pzRHebnqZ3plFd1EZP+IaGMAHJsl1sWGQi+mCq85+MX5q
vaUiRNraCDHmr6SAlZavpLwLnx2laL6akQqrY/KfJKrg05LV/leXFG6cizlt1nyM
0IcmhuavVo66N8yUncvifb9AnuZNpqFb0HAX8ACGkHY=
`protect END_PROTECTED
