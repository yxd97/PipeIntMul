`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XcnR8f6Du4cd8g6Qi/rchERDuftO3K4Td7wIAwVbgchDuBvEUJYPmBbG8e+ojiqb
YXhuheiPINDdFzkXT1fFNIZO9RXdMKH05p78K3WwfT3x8r0FWWQfGk28QZMbdqhY
RlvAgvBSer8qE/qTtTAxJ6iZ5lXvIKYbzJwvbuDUkN++nLwj/ICZ4SD5/h1pR1II
xqmXZa5ofiYvbEACkQjx8JjHEsSZZjZRiXSYcAdg9v9ARM1KdylvtPYCM5yKTPKF
gzwzfkF/7USy2OZ8iNTHGB0D/o3ej81kIOo1BGHCvZWeCAiQ2DB9pq6uiomklzFr
L1Rc2ByRZO2tNRqgWCFRrtQaLxbtmzGeCiI3KFEj2Nkqh9G9fM7x/IVgeonnCzUT
0zkf339LuBBJ8VmxoxG6B2UgMCitxeyj8Ul0YgDQGhcww+Iv18qNNPbNrGK2X7fp
1HV0uCBEvx0TXcmV9Fk5gAv0C4dmOA2xmxAo6P2RK/RIUs6/e9gSnmTY5RkWA9K0
Gljm4L7oOHkQw8BOblTdY9Rg8Hinm/DlMhqNyY10jGQ=
`protect END_PROTECTED
