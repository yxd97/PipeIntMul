`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ryuv9dAPpGQPGvg/D5PWCFJ0pVWDLMEgrdmGSB75ozd0FDpfPhb+ya/Rj9uMvO15
PMOpT2lOFFgIdrJ0jlq8Ei38kCHkccgW8tw/0r5ji88fpYgMjCLQquYdPDWZMZDc
SZ5/0zaQ0+eNxr7LQ5dlcMYldoSTC0EHV49P9ERdzBhJLHaB44rv18nk9/Ee12tm
GfAuVjN7AvXKv9sYbg5zI1KLn4/N2kMIKG5ciLcfYOjT3Yc4parWYyUBaIIpXU+/
ynfV/thV/JTC0xtAMQgqjw==
`protect END_PROTECTED
