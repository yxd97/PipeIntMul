`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ff5yQYrPfaWnxv3k7F9pLrZfRx7G73X+t0SN26NYAFhBHw3T+gvR6fvOg4QRFD6y
WBolu6trmsMJpgp5MU0eT8+ohbHjuGmOzCQfTpXbx95xz004tb56dEGIaon9n+xh
HjsiZMSWg+1Hx/yafcjNkitpxnz4i0bXujq0PQtPFFMDSsNm8VfD/Gb3yxLtnHFI
O0y7YKClSEe5Tj+LWLnIOzLzFrGGlmE4Nvbitj+Q3ZQo037ng1AiaZ6Z7V6fFqpx
AzyyoYNJR+B9I9QRm8qBjigubwxM8vfI7XLgm/Ql8pSnSv/UuyD/y3/zkmhjsGeo
CeWVc9i+ROCO3Ud+xqHkpo46vmYkT3p4HpGvEheWkenFSQIsVKvNF3Lu9OxANS1F
KvCqsNw423R9Z05eIKryx6NlwcjKI6IV83ylsTsXzVwf+X/egKzudf3byRTOUYtf
PVRcBqoEpllkEtnCMssMXKYYwjJAxeF5sBu3u6zM5QJnVM/eeHt5cYUaJ8n9JwiH
b2Su2WzxhlYJLSwBgFqMDA==
`protect END_PROTECTED
