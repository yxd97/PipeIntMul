`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+lSYnO6m6NlEK8Ep8x2Yp5iJ1sFK3o6nGtdTom62BgHKntnrmzIaEXyQ9O73eYL7
q7yqKoKEBWpMQPspbitnk+on/xbpYNVZ3Metsl2Nk2/jf9X5NjXCWKZj94AM+EGq
YNO7XmzF0B/+nU+z1anrS2L4VRw2EKGpwoP7jTmIBVxHQe4SrB20znC54eCYKrkw
MM+xnp46LfE2EvF/fYoqAIRwdQhRNyNRLkjer890r7Dq9dGA2O4RwsZMwhfDtfSU
vvrmac/1/TtPK6ZEJHHr1vVUSQ9MgxNNGR7pkfE7GazPICELOFf/K/K+xFU1YQuo
wLVXS56Pzyk5XeLH0SGWziym+L9PA19yE1jQ3Y5U1zaLGVZ098BCHKu9uSvflqu9
7HTV8giczweF5cogLZpUNdwbhjolMNTM8wQ8MnxrxCrV+rVkqWHehKC1Gjg82dup
IcfX0CIDTSnlPe6coYL6FVIVltQ9NABzW2PZ0FnTsl+E10Atp4JwmrgpNEUGOxDm
wtZ6cPsOZX/5aIXRyHIfCv8xvWXZxDSvZCHzojGyUSKXC2JKDgVNW8OAkgkxFxDu
8oFH/ul/8sdR4l3nBIxkktVu9rQm0hGhRv6bh7J+sIw=
`protect END_PROTECTED
