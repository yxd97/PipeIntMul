`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UAuDAqhf39+VyT0Hxx5g/BdkMnDcD/A4f4ON53e0EJgPMeO2Nh8WUq2xskw3V8QQ
90xY4rO6I/A/L6SkFG2PQn141T26Na7C58q5tk+R8zgyZWBI5eM4K+GbUIaH+bnc
eLXfhGGa2L56hcLNMAqfxWxnqPDeV99sqyz4zdo5lUaU74Qpsu1I00+M+EsBdXeU
RoSrSy/smq5Fla0thzFrkztos/yY6ldJ6/asrfaWlTb9WIVfZbLxhIkGUaSvht2p
K14V7DPcjCytoHdZpzGqgQvb4eLQp2XFVuTKBZgRT+WWHTnH/TQ0SukziF5GdtnF
+lvCTbgKRg/NgU74RTk1PCnrNHGBSaouagUpJyrrUiKqXQkw1i4okLt4HJDlJ0/9
eTeKIw01oGX3+mDLrLrHCwOXosir1A15DU6YCTOhIeLrdOtUWq9PvhMwEBZXb8Vq
Kx+dPyS2WHsUlk21JQ3GQFKyUoh78ZN6s4trv84TrHb+MGtDP8Fpy7XzRRPGMH4c
9SfXcOpyq2vhnYye8qjt2Rgp6R2JsNtei8pxvhz9T90=
`protect END_PROTECTED
