`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xl5iGkdByU0xDHQ0+0hiuo9avurSgVpF8/8Kc0GMlSy9HSbytDW1Tgl+q/b/kMG4
xujbX0+iNO9nkHRtQL03jnf6xmuFZHOzyLz2q7MdUQd88CCgn0P72JpScPPkcBL7
4PeKGR8pHZrRiJilyt0T5lp5BrMb92zWbxbgokdEpxpbLY3qr0M0WcDRRVq5G+Kx
5N0vuTcBgW2nUR+4+Bqb2ytTbKJDX3nUPj5ax9A/DGjBOFuZvOmWBizCK0LYGog5
kzXRH7Z8EQwqvoNLswGC0imOHUTbj2WEu5Gaz9JCzXZuyncz36FAX2G9BQrEFCjp
2wAY5Hv/bJA7de4wrubsZgQprIbk25+dNTJ/8tllc69Q62U7nDPmFbJLT8VDcO+D
Pev1KFRrwFL/2aNxv1pPnRfedRtMT59u6HwbBbYA2EdGEv54xXcfXmEjO8UevTYC
G/XXPIrNHCwWcyyBT/z8XtiFRtbHlPwu+aoXQhOzHSlYLZUMBjBgJPD9Rprp0h0G
mVB5kl21qPUKcS0Vy+RdEKhHBlEKSpgvD+LE8G7SU+7A8bHGeZ1mA/+Z7y0ztRRy
74bcOyLJdTFrrSGi7ZS4lznaRR3ElTEmqiayEHWWH20RtmYpDPxSHSPFbLHhNTWr
q+kxFp3ex3T3jSOaFcaSGeti8SqhDbPHWaknJqDzgnGY7+y74MOLYt2MzV8gbXSe
vcF+3EZcGyB5y8AJl6jKc3I1lzU4o8aiZ5ewEVNA03bU5edhc+82t0Ycdsu7FiOG
NBRznL+Mm0USCFbCyy7U5uE4pcpRaPvpbeq+xdoyy4zvx61iGa/Y7f9vs9ddXLlj
cLOW9E7dVZLiNmyd5kHfgB+f2KjOvSCRHp8T9QMEZYgCcEUqxDfv/vBcMx/eebjG
PjXJjaaYDW0cC+uIt4iQ7cpw7k4qznXJsMxixxGNJHzbInrf3Tll/GzudAT14Yhr
2CUfZlos771jn115ag9socRrhIQgBso3KmtZSu4iuoyuCcCD+1joenDHMbacSi5D
VlYG4hN2x1fFK4DMlYOI1E4rLlAeisVhWJR+VYkooO4f2cLiOvVD7P4//uRL7Ydk
a9XUjr8ljlPqugpVzHaSmV1uiRAmZVNzjDBtZVWN7UxkwuX6KnMVAIZeuA1oS/HL
d/qk9ocauqWX2libZPJKIQrBpRNGo2pvcAxDIQb50MIlDR+R0SoEt8mkfvO0fbrm
FY8o0O+fuj59hoIGKJRCDYd71VzGRmIr/U+fvKRvLraxmYuwHLfavCfNYMOUYDks
`protect END_PROTECTED
