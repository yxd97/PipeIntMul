`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jris9iKKTQvuuDAppkaabN/vSBMa0veQHCjUYY4Si4Dz28eduu6eL8VWo48cKoGS
2ZBTbHB8X7p3oRItluje6EAdadWJ7K5gCZ9nXJE572BxJM4DKzqhv91IXeJ0htZC
uLYhxsrOURLZ3V9TfQSFWJkoCxj33T2OVutPsfEGLuFAe7VgUATogwm9g4vvcrIC
mPKOkvj09tMMtUX7V+kTbQmmk6PDOpEHJyQl+RAfedPHemeNvQHDuH1LaH7ICsXu
89aIkhSQMEksvkiRvA6P2eV4XLCt8Ue/pP61Ncb49quwuhZlGdjs4LwgTFq7jySj
5a+Fwd43rQaD0OJ1Qq4ZYYuAxti6STA06mT4XXqwNjJCT8rkN9/oxOlkO+Lt7mlx
`protect END_PROTECTED
