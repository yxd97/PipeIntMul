`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPisMk2krBmYzsHsUOAQOpj4ppd0aF3bXeJXETBZjo9v8bD+cOH/HEzxAxKymCwP
ypSeXLpHY52MqjAlgEx8ZecMwboMReblgjP5wupNNIZmvdmys2tG74cIPLH5Fwst
xaHSyazruXXG+cZ18NlB1g0VXJw84OnU0O855l5qCcK6u9qoAEtXH+DhujdL/cVK
/aU4yqep+QQPmUYPZcADKJjcooIAN2pYa12ozarODSa8XE1rcvew45PpbFezDF0x
qpYrgLBQeOxQkeC5bmt2HiFKOpb4jKaxL+rqU65x34vVJW5knt3NOS0vxD2BbhH8
`protect END_PROTECTED
