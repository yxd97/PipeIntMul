`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXQvZv++iylPNciWNXm7uxKj7AUw5g6KBYZKNnW0YoN78/ksggNDE/i3I5xhljaA
9eLqT1XKnggEEWK3kRPHm9R5yXlM6noVQquBRkYc1JY3iGWmB7QO3M4p8r2/mPwX
Pi1MliIbVC6ywleJ5xffxv+z3/P83GFv4rwRc2qdpqTxRH+PLIUBuiUeNUZP+Awo
afuwIqB4T5ymoe1V0imlYR1+WFrADpLuGaxg4G7wEKmBC94rLFhJMLnrmTV4TR4H
A3NcxuozSfM+I1EiMGzJcn6+f8EsmRk4vtS9nj55Xxj3xkqGgKO7+BMMaEMLgEkX
lH4E7RFhCiII3o+lgzR02lnqDcasECKIKOo+GQG3kny5GL/l7bfblYFKjwDsnNef
L+YPisFoQZTaRH3J/bTI/wL1HHDsyA3HOXdNPqep5fzSzhFhhu7d3vl08uOMmaAF
5IIQCT+stOW4foyneR40HtGfx/1hLTSckzfmhZXZtoHJvmvLKp7N5FT9p//Vi+fn
qeOK0u68n7WXwqxWavVlui3q7nHsDmZ4g2kIbjP7T5YyXtn9LlRm25YWhYceP3kZ
AGibWiSYic8Y8Q4VXvW13mDbEnY1cWsc8HHTq89JeJx4l25AWUHuoY2Jl/z7FSaP
Wli6onVEPIThQ2k4Z/yK//tS+HhdzFPbUUNJVFCK29hXMHPb4RewA2eDkvXMkBgx
cLIf1W6ZhGPM7NLtLkFbruMFy2dsJDmtiZdn9nhSNl1/ZYXpnvPYKtEwsbDc12gy
XjQNGB31+ed4f9T7b2Kyh0Swp1VvwuHnQixjDUAUC7bHDa+Pg/jP89Ebf3w4FmSl
mVK+YW4G5WUbuGSGndg7ms09xun4HLntkPlRQltvyGc26xA75KSDfOyLyZC5+jZF
jqRDDNHb5YKWHUG+5euVgSOpHOL83kFhYjLVlZRwxROhp1cmuu0g6PU5rQSGnesQ
AizoEL0Xq94jeLiidoMfyS+kZSEJOt8DT5RSgA1hi9GLzNHyTAd/eO9pNNILhBFX
unJuUkaU+dUB/oK0MdD/xjxwNxCOdidJlbYQ9kItafYt9gZAnAI6mKMA7VGkBtbb
ZDIZwn22Cv58P3WRMoHezI6LwpiN5tTU9nuDiuYcjoi5uTw+xe1Xdd8m0K40Rktb
tFJ9jWS62PaE81bAAWBAAN0NCAD2zmMOAcPfCx+q8gypxidxoWNkiaAFHvjI3Eqs
8JEoQyMEvgGIADiRKsr/vbXHvwXRAiLR//8DvKRj1wiuLUEGv4BQ++HzVssH+Rid
xjtK1AnfyLXordIswdzTXvwgWE2hew6glmgxX5wOf/eLPKYId4x1vvOmbmWIP9nh
wE0cKtmeVNSDnN65u5ZK4edAt3itidwEhybXiHc9E2e/wnhnXeDHl4YC87e0T5cg
4NccPp3LJgOErr/a8U3nsnA70YoKRXPCCo7fBGRiquZg3CMGgyE8xyW3rmsYozte
36uXvBgQ9GcZD0sXXrEjaA==
`protect END_PROTECTED
