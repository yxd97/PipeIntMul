`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xwrab1EExgjSxTjzlj45+E4DInWzOsNZ/WZkzQXvqyMFmKw2p8DSA8e52jFGpy2X
sSA19dD6bE80UYZ5+hFR/+FTq9IhL9c7o68/z5kDF5EVgQrcGxdGXZx5+F6sAgLF
PpOj9R90hoi9lFx/3wG1FmOvXOoWbI/mr5t3hCkExqJ09LjZeBZR6OyKPbxUN4JV
w36U46qMJ6tgnyPgA9UIQSivcFUYq2d2WHh3yT+ju4CocTpHI5unJjJ5Yzu1fyL6
8PtSjj9BEK6EjDxbFy3e/MBJ3D1ckl+DaQy6SSVAHIGeqizsCIP4Zvn75jgxZrnR
rekgL7ujttb73oslk4NTBLChrzufyBxy6WWkEEnGZDXMnukYvJOvbld2ArcC0Axr
QYERsm9YOa26LywaBoZ7Mcpb33ogzud7JcD8smmiFCQ=
`protect END_PROTECTED
