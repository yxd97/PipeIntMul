`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDQ+s6wFFt2iLZcy/QydM+FRQWERJJV7jzItVbjxdHc3t/jHVbJi4tUv8HlgBkqm
pcbag+q/yiAyT6EriHFjZmiZXiikdS9SZcufpHzOqh40hnZMv8BX9TzM2JrlVejO
N2IUzy9YqQBKtettSe4RNKAhrLjBzS3lxAmzFBXhiVocJJJSNHnQOWLpS8VLTi5n
OWcLKG/lH+ynWe0IUpfacKfyYuK4tNT4XMB4TuLOg1Nd+xTUJWl7BhWrt9cBPloB
pEs8jtKV6kTl7uHGWtaTdX/vJek27KbvH7wyrKWTL3bZjkx+PdKbiYrgZ/DQd+C/
TYzcOArmyz+Bsk60DbzybrLfJXkQOu8c8uF/Xg+a3tleLhZEdhUmjuUqVofo1AgF
sWY04SChPVmYdXneMsrk8zQlAcKRxU+ypXeiZaomZ2/FQoEJVrcvtjOQZKpSlYTd
dHwG0ID97RpBlbqgYloLLryWiHcrJC7P16oBW+TQc/qGV7ihleO6OmxBklwht0NL
8GPJoZ8Dvjg2q7WbAbB6XXIWIbGWILHXLopl8iBVTXcNgFUjlwGifTVWgzKGUsW3
vSMxegfgWcp5y9Ljh2qbLo9e4aNQvdOkjqxOG93HtEq2Si4x46OSfYe0EJy05oVl
6ZvhRDP/O5ZdbPqcjL4qbw8EHJz2eUeZ22Zy/22dCbGrhaoFibJZzBJk3jdPwLdj
BWYdXPSAkbRa9Q0NDytuFxq5OucNtvKOsme6IJd0/CotvIGMF5JeGVXBT663x5/p
LZ4276+XkqMVHcuUsucUZWxbLvghSmNSNiwAP2senF8c4sIbq3F8Vf2liqngWdHh
MIpUtK8rDS96vqXLt2SFmeXJ9JKy1s3ZwGCWRccbAxoLVFESmaf44lq5hyk0cotB
sCKmFKgLq5Rujn0fVszNZt2sDLCczEFg9YzXtHlG+6W0vDC64l6PQbzOXk9+m1C1
LV2+ONB1kp4ACG4aVFhQy5mFa7AdYOo0BXmDwGBI+ZESMWqJwB3VPDvgBJ2IZeIT
DYFCeZ5CU11xrZP+tD+m/lBvAIXHUKDX3FJHZZTdqJAnBUIvhVyKpwWPqDgKQ8Jw
+IHJbMk3+2ZzFe/8Pg0YeXb6A3Yh94+XCnp2iOOsHQpu93v5W23yYr4J6iirv8UL
Ok9iWO4ZvpdnHR+E/grf3b4mP5stlVXN0QBK1Q4XnHO0UjoFYVxY3zh6D/63Xx5c
hOs1X6PGmY8Gp90GMSjLl8RQXLNxl4mV/E22suiBGj4lwebwVo9Ir3+L5Nh67OTx
a+lVuaKuv2eRmtDvO+MxHBzcSHYxYJ1rgXIqkATCAm5XR+0ctqiFM0d/ZEPfvjm8
Qg5stH9YsUcuE7oPbUfDLMAkoVzprb6mPYNE1Z5xvAN4l/yqa76SGhbup13xvUWU
ORd3+CQKB6zeDs/LhcyFf32r90C5VDBKDft1t/1RlrvzH+Ex0HY6utT/k5SPEb/8
7NQZ4lMIhWvTpNtm4S1WWDPzpCc0g/BTTg9JCmbN668ax+A0e2E6T7ooP6tD886x
2fmTu8Yud0qyKXt0QtJNNZJAzPVxvJa6vlk3JC1MdC1OwnS5O2x8kch+UOb2mhZp
i6cdAM4wdqFd1v6dHNsdiiwKH279hs0GEpD7SColjklT5VVqYjNUtmWBId8vvmyt
an2IC6ft2rCSiKZab4Ylbw0QAjrq900NIClCeh+xZYnAqvPJdMTuw7pzydKaJigF
Sk0dJBBXxT94ngXSWOVzboIRvE65OSEdYHoMrOmuFo0PHqG0/R7vrQ/Utfi2NeF/
42Fuoov7wM/qgEaPNx/Uo0gArD2VtUA1P65fJuSbWvu/wQ4TEXl1WFqNQAghsGSM
WiWNiIRmZDOefJlPb8fBiW8pcnP8V7XHWdWb20rBqR/NaVVEhMPMwI1eVGOYrXCI
HWGo/YubE1PCvHdjreRz1PCBGrOOvGkHgcpIxSy/QxzUYq/BJ0dAbtGATYdg8qQP
shux3UddFL5nLyZqvDLuCjueJNO0260gBxP3U6f4VTpBnvcuHzhtNModprPVqJTt
x0ihzmzuBDf00uDO/GKzQ7v0XqRVo7X1e/Znoe4R7WhwZY4QSfDXQPHuWiv/8awz
LSwA/sMojQYhe8DFfh/0pvAKSJBo05tfxtaHUH+MKT15pGs9tsUjo+/fNE4+pauI
H54ELjJwtsyHXZ+74dbEA64GrYNaDO6E5HKjmiaLKqRQYJqMAf4iS5rmwArTjojZ
OvatVELHobAwLghWciZUgNM1N8WaGyx7de6dtGK8kHxyRk66sRH4Po4CLQRm6DK3
SAw3vINWCYctXBLgBTzn6ijii9SMOQIorLTXkxVg7IiMWmakw4DeApZruiMoqXZT
zH0yvaSQt/bPzziyBZjUdLv39W3+9ZlZX7WO3orOimd+a42vBzVJACJLGRT9Z71p
2frA3kQWPflmn8zj3bOVbY4tNwEnusByreS7/MDrO14ABJ4mBN84Hy2nkasoKL/t
QvGU4JHkJX/1Kh2Mv3Sjbp/Oqolc1N5hGqvpE74+Nn566CeAwY0nZnixwNP3xKaz
vemT952OnumHhNvYPmQt2wZ7jwfaNNcH3rie2kmm9EQbGZvr62V1Y70hGrp3Ih0i
Ghz5BTP+rrFd36vXHtB7O5hMCHO0FURCwAGzvQ/xoxlrVDfD4A56QuVwC5/wfiLc
cgQMw7sHPfqgLDp6HRAbITmmDWWlZFZwLoHC9pRGYH5i2CNKsjSfO0dqbB8akiaV
P3y08bfvzzgiD9FmHyD1CSNObE0+syVPi3qHIDZBQNBiYYIff46vODwQTNjMVsbW
wddCSwfZsX0PxNtrSQvErsO+f1AvReoWvqZGrpKDpGRiaxJ4m1XlRKNFKhaXTWKW
d+osuEW/M4i2bCr+PCHmFWjYL2a8ocUaHPtgjh1JRCupjf6TBL2vX5b5c0MLlJmU
t4E1i60ihwFfR6OSeKUoeaQmMx0qukMCAdfV8ZJvuDdCxh+djDED/ROlwTR+RVqi
JjLbC9yMwfyNiHEUYCiBL0PQtF175lLCz5ll/J5Th72YY37+4XO3H9e60Uczf2mR
FHGiYm10jPiQULuBh+weWUZ1VVSR4OQfzeR7oE4gXmS7K/Upu7PIU7u1qUmjqB8j
YPFKCwPvh48CL0EKuhP1B0+n8M2gTfxhK2R+5vDB3OsncV/mZcimoIi51KEDemub
BVLgNcuPVsNJEO2Pr6UOXArUfyEVHxdigz0x1gm2+wVmsH0My4w7hOXPVIQ9/Hb6
oWNwOwxaSuyh2tdPHcqiH85qWc1VVRjys4sgwBnhnjh1uNABHLgeJzjSNJ1RUTPb
zMzn4f6z05cllI9+RV9/cjD78KSDB1LvguxLUJv3KeVCbicC4sw+a2VpYcVmaHCW
SyO1UUbFf6qD+UHhzQTrE8AASkmn7DHrQmxkuR6otuFa9MJ/K52QCP1q3o5/OJgT
JA78LUENjJo7yCtWObikiUiCkah+tZ27uvusJbiDWR3sk9xCBpo850y95kZyqD9C
0CWPZVXTEI5vS4EAcU0oJMCijcgALbcCTMh/voWAiDJLYnydL0NeuvpW0UK9EaIm
WOCwX1D3sAMytGsdwj8or3uet6mzhLZNwDkEzD7dC66iffCWi2NzFgy+MheeMKGF
+AI7trqqGu0c1hS0NpdjPOiWOrlI8EARhGXMav1jOFhpoP9A7tkLVW3oRXF6aceO
etsPCKJ1t8PA8CLI/6jCn836AAvb6SpAs6GtBIPuwV0snuJjGxkg1a6EYgNcuTqZ
cNrprCy/9OxQc63cW1y8OrL1ItYoNAMJJBm2dOTcrqaes++3dZVZ5YD26GGB2TRD
yeBaVnFAYLNjw2QggwdStMk2hXyR3PW9fAn+ItLlw7M8T7XwaplNlfvoqYyZ11nW
+ol7LemH5A6Wf56uOco3RzLODdh4YA5kt5jsuLofBl3/qDkUY+CpPkChBYicz8fm
Uj9Dx7ww4YqUSfpc2CBrdzlFS0synB3OtWkW9tvDOYFcXr6qp2V/xu/KWp6MBu3X
BhKVJWlbt9ksZ1ZaqwguhzwOLwdFFj0Zv8iygUioQafruSLpwFjjHK8WOSsJokic
I+8dCD0jpepy12QwDtx2sFrro5KxIbhplc03yCzM3HyRE35vjSoCoFO0DCWpwNi1
7uQwWL93yT6xHLeGhUyCGNEvZUWOrcOYwvjkgila2xfDiwF7jE+Raxtae/1gzPhT
Zfv8XanIszoOwPtiDbDFI+qR/5Pn8EC+xbHRU2eR+f/15b8P9sIDnscxw0r1n64H
HvAO/GdXNXK8S6i/uvBeXphfCZ0Gd5m3K/pvpOsOfP4U3I80prznsqzZYRSCSsHq
NIGnuqQ/Dsc9SnZZPoDjfWmHnSE024zqWiCp+aF7KyWYcmTPJRDY9cYNAJCGw7i9
Hn9iN6VEX1L1cBwzEtbtbPxKLtdeMy0x3ppeMHnzsGgAUcX4RjKCG0zqlunT8Efp
6b+V8K6GnhcvdyE2+gZFh4y1tjdtLvjGgxN4XEW0OThqv0O/Kizm1qDaX7tKpl3v
YK6JP/ezQ9lJpwkgQFOHcitlCS2fRjcRS6fJHc2wYpD78a8s/aeHMiw29lNP9nnP
EkZNBFBOl8kDJ+0pVonwmR0xb01tDEIjgFiDEf2YEGMjfNQxA2GmiNltXh5SNZs+
Fdl6PsC/ElWcn5LyROGQTtUhYDUWgGjdJNiq9qx5upBObpMqXrnImwZqbl/dLtJK
ZeGPIueOnuHHQ9KFabfnPIrGpUl6Vjk9GLk/AaY7ekz0ynTCf3vNTkCDlb6B8DL7
6hbjxEpwxqaEanDry1tTbdjQ4HMYb7DqxGJoNvnOJZEh0qAAXgU8UNBhuXh9xis5
yy2Rv3DzoWdf5aDai1ZnRq4TTmKYBkk2ZD64DYdCcO13QErjKL7d5OChaPArvoRe
iEI0baNbDmQ+wDoEHaoBVmB5ICtqXeHSyvr010NOIecRjIdVkgZqXqzZJYGhumaf
iQB3/BTiM8r2zqNDWAZU+rY66WJeCSQJZxq+V0BrjABloWytOl9KdSwGAefr9Zry
Zl0uX5UqkM/GRGeKZwhqgLega3KrNP7DltcGR0voidrnI7q59avI84HsGUByv01F
bK1Ys4fVlUaDH2+Qs5Sm8y7EP+yR7oLVhFIFKCSFnjz8Mcr2prcNIdpclBF1M0Ak
VDWnHmXohm1pYgl8PcKIyoDRecbgKW9ihRywc9VB+LhxzSyfm4MMmaRLs37Qwj3E
MKKesRH6aMsPnO3cKioWytcvqwh0weecdXTDFRm98ZU5eP0L0AC+OLW/XO2QiqyW
iCQRIZiSl93w6nD/0ccIoQBmy4lTvnkEG3nIqgba+ly9amL3gtis2t1djhXCD+Ex
UtIYWp+XLxpXQ/uVmgPYYbz5sp0/H6Via62mOw2OPRKWMmR+ONBSX4v/BEADoIKj
HU2BfBoWkefPa2nzHyR8MHxqV19DGEVKlT7jSfjJyI6BYjnveYA1YqspQ5hSPlnX
mXUXiWCDUvEsnQYQbxcDXjizJvBOGV3b4tACIOGq9Y75DZHT/CH+POgbBwCdfxKT
pZd0A08tkjRN45z3T3Aba17Lg2BTwKdxeri8d3bwr2j0aSJhal0GaYV4nxxA3Lxu
Iu1N/vQP34k9GU9WncbiuTTKlXWkNnNuC+0C+E1Mgszfy7hEc48o1TYjBz6Cyvnj
iGp6zbxDvS7mxR9l44HYRK5wF9Z2xezf+nuaS/AccTWONAV0LV+nKQgkU4w4kWBT
0Qa7ELr3NsxH73043o4QKuJtxVXvay593Hvsg35HKGEs+1zWR9gAQzHDI4+9bwRk
PySoZBtlQ6Xw85yviBUf3uRJIMaKtnaMfYVm2lsCDxw40X8rmpaK94ZlA3lb5TWE
pkBMnPEXc6c22DoPmk9b6lKZVZnq7sM2vEkWykVuA1KzxdI9UoUaLyQL1wFPovev
W1x0KufDsxAWczDVi/gjL+K/ZeePw2pczlohHLL1meTMEgw7QMjQGwQ4c5AMWA/q
3D3mjwLK+pRyH65B/rkSYO2q5qXhaEWGFI8ZrVucfcmCHdzo/AgLN7YF3vS1OPqt
btW206IeeFNx5se7Bxo3RL0tKR+3W2mwv0TLxsf4eYhgtU0snps9HaACaMvtAlMH
05ilB209Z/Yv+s2nznVHY/aQtHsoW9UK3gGtGf9kzwSw5bjFl3uvYhFhURTPwGId
ZR4a/cnPoN4ZgWiG0WvEVGkjw5h0Ec9xVNUTA1iQm1Y6Z7TytXz7320RlSEe9hZz
Y6tOrv3KwtGa6hBpzpZIWHvol43+QIawuZS836Wx0erjFDzM9WXfy4yyir86kPuj
45dDEjs8FbcrgHZ6dnJWo4hdrjY8WpKXMzhjIt10VuWtiEXIItqq/U1C9nSI7D/e
ch2VnfF99OPNOSBzXLi1jMdIfLmPLox/Q8waLcda4bVQixyZ8rXdODe3xXLZl2CK
470G01GE2HzlSAdE+m6HVwnFgI8BG5XxrIjl5hhYTa8qHR8dbjhjAH3vT14920OI
f70wG1i6jnEIrkZTjoyqJrO42PW+gWBzhauUPEc6kd6uFcCmjcE84UXvC8+KfZU6
Q7sEM5dSts7Ca3GHN6KVvNEbqOHYmE0Cvaa/sto8EqWgC6FMPXCJzQz38+s2Yq6q
/73o6bY0kvo1nh7Pj2t2RXBXpnJgqJqplU5wX44K878tX69eee9lzwh8JlYWOPr5
9Gxsg7M8d4QYl5ofcPRkIamrQ5ps6m3Tmu6u9ICGpiDAqIAMJdAbAue0fJxv4dfg
8+QpljqlVJeYYaeMvoAjk7247K5LVnX3OW8g25X5qlrn8jAh5Q+qnonoD28H2Rua
VH4YY5HZ2hsRUPB0Rx591MIFI8y0MIkw9WEvrEjQIA56W/A3YLaozfxMtzq8RtwR
f3PqLeh5dKwmgJMGNNLu2xN/hxUNv5062yxCpJkW+1qac5ehdKKMMrHxWng9IJ/A
/hL3v4S7VKrAcr68IhZPMngZoLfxbXaXzfCmEXQ98UH3gxUJe3hchEuGCSyjKudE
R69bVkn9+s3XWs7Vq45qMLhnxQOZns8chmRstL/8OmjafqdzltKCtvVx7B/+aixx
ivcPbFVPC2a6Sgz8TE0OceizsaJ+mmRlm3qKKnmRprtTlsHNDbsklCX9fSadHMKw
mW5FA1nQB36zpV3LT0msOScGqAimURUc/Lu60OlqwBrpI0VK+i9AJR/7zLhoCbDO
eCBqBjHH45jPJceOxiLhxpsXLTsErkJlqQAWXhLLMcmbMtUKm+qbkXzWBzQFcQr2
pNR6FGf/bNjIeIk5KkHRcwY71PLR6E8yEWzPQi0WgDs5+tTkorEz19NeHsvfTeoU
tYrCHAPcF0EwkYhv7g5l7pSr/csQ+CjmVakA29xYdie89n+Z5CPWfaKjq6LJR6cW
+HNrqbg0HXQbxsMKieCR8LyQJLtd4oG9oDVCZ9TZ5rZjF1LTKXC5o0CCRgaCy6pX
hvdJXTc+Yh97pnBPyXuG/LWvXqRRJjSUE/VzI9XCxD7VDHP8Bjc1QuBz0+SMtbvt
8DxW5Kc19nQCKJC86BKNYJctKlcwQPeOrlNas7MPP1exXnktRjbQhVH2B4+QqobN
U2ospUK/6lYP1/9cjqgDCPVyrP8n4Dl3wpwvQknpmOj2zp4CRgtKXmAIQzxO+cau
ZRRT+O1JBl7RKIeI9cyomwBqgDVHVFMJDVW5LDqI348CeOnAF9s53xwozrcxSymB
9tZ2WN/elEW2SRy7FY0KgoPO55hAy9Ri6qrUfX5tYmW7S1EOWM8GhT1GeH1d/KCU
QwAZJQy7Agn59FmR+7R74RQy0Fa9sOfC343vT9y6W7NMwn+AAA/uW9kpVkhPctA2
TlnpP9lbyZN++I0+Qdn7wVTf0AoVWcoQilHbORcI0qKTcwmZhZK5E0iGvVQVS1RY
vTuVtI1MRspgpOChT9kVe02It4ipy3PgVPNqXFQBDjd71iPughypXy1qbiEucdOw
dKlGFSQFcUqi/3JGvqWcUJhaSS9xNzN//6KPfu9nOwM6PhlZ2Q/8naHoyeSmpa7q
2hF4iultNMLQHlr8Tla7xW7Ncb1BtUKwUF4yz0bqBjQeNSTJdPI8C3vrjvVK/2Je
c7cbdoL+s7CP+RMRQUye16y4yXmWcdDdEKUiQbB15MgEs3MvNXcK+1SxykEG3oZC
D5VuEnmXKXG8RXxFEx1tWBePiJ1fv0VnbuUuzpG3Zxr8XcymtyOuYE2E8GcNBygV
zOmPhHDV0HQLGkzlYIZSazpvRwvGCOw2r1nirNg5yk+mv+iAisSfSGxLwX2R+QO+
lv0EXAL6JO9sN72K6tiimIzXt0i7nFZNMMeEqANn15qYYZqGGTl7I7laElY5XicS
ocCY/AUrADTyP6rzzYF0zxF9xAk08uGPI9C6DoQBVI90+gLkGWzs9l7KdQdYMzQM
ftPUyonqZ7V+sC/+fumcJlgXtD448SBfP5iJ0G3TdrnA2bPh9oD2Gts+StcG7vRS
N27c+EYHQa6dFnlo3L5x/GzcDmwBdGB205/B56Onph/CBEh0b3Efxeldk1SwognY
mO9NSp4+CSSxoL31/W6eikJUtWXl1zmuopMPQp6/AxauEtYP75gJxI6LaEs+Vj0F
4uaaJkkm3RmA94DboVO+5ODj3Ye6xmZ7YYwtJ0+FOAFJ2jlMu67DSYTwCV8VakWa
UIS1ey4iJcJCZegE5pVSwtyU95omzSqW3qx/DuFkyTunS6HT63cYJiTVxNIxsjuS
cqiySAJOYc102d9w4XDBM7QgpUUPhAppln6Iy7oY2WCoIuiMITC73g/0yNANDjZb
SpgQFGpw3hhHRr3di0jvA47dkVNb/6hZ85p6O239PBeA9XKbEBjd09Xfu+vuE6pJ
EhrdIsp5BJw2I+HXXh12kTSQAI+ccCaAj6a4F3vRHMKh6eZD2vZazjbLPO6HxK4F
IjbUJuV4QX1M9rAgMm7uxY4WUxS+C9jr8oORZ9A69ncoS4gCvpGYEQy8zfws8CX5
hQfvpwgL2HfTZ4TVPjRAk0S7W7IxSbeIBJChZ0wDolol8UZs3MoAmmE+QKDM4e1e
4vzcyxXvvUJLj+cUO246g98PUmihauVVYx6J+Q0+dQXnpXZC1q7nhQwtglOqMha8
76NB7D7nLTXseURqzmJu9KQ6ABMzlCSAN2JPQiIluPVQV3QRdSU5Ld+Mmk40A1mG
a0qyxoSEFeRtGtIJcy7qBmrmD1AaG2We25WimPWtOf56g5ZO038G2sUmAbA9CUGr
SPpALzGSYk2uKw2HKGJARUr/Mcf+vOip7A7n1d2aaedICDeD8gatZ80v3G9oiiN0
+D+aQO065UEeifsqZ1AYV2DBpXpkdGFsqDzt2kJ5jKEJBWyWKQngd6v/Ilxi5sXA
5OhBW1Tb/A938hDs5m99E0HBt7cLn95++F2EMuy8rusoyU2srTE1ICFaiej1sTBU
a/Ye2Fu0j+XJgARouGcdSHsJZWaiz6SOdxDe+HzsDwF0tohORW/vC4BYlds6syoH
fyNutgH55T8UVVyZ+hlzxjI/yoAPJefDfj7nDMJR9b1YVthhwfwE4nLpfkPjBug4
Oa6ZXnby+6cz60VWo2q7EvlUaoLCYLOmqeinPLBktYLP+BEIM0KFNqeYQxSIHiTL
w6tB00WqKMS+UdIwccfVDM9QbXTvxuclFHuk8vJEHlqfH2Qe962yOPz8IZDVF1pw
rtwtr+EAxpYz5/tbOtWXw1J0aZyVqt4wzNhz/s9IbakORFn9EJdPd4JMLiY3Jw83
6IN/gt9i09DVG2HOxEYEyfj/DU2AO3tFHwsVmDDR8bbnj7jeY4AFg2KpFx3CXG0W
hx6n6JeMUY8ku4RoKaIGbE6kA+jEyCzPTYdU6h0gyRV5QctiEiIpMSjpRXx7HCee
Vw3qALINdctlJYljRa2aXYbjbjSqv8cAGwX+7VkW3Glvq/EJmxNcM2igmx67yHA7
dPfytm1+fColyU9bgp5OQgPt6M+jt00/JPbU2cFm58mU8TERLb2GxNo6CRvGtTlF
gACu0QG6z00tO8d2U0+rMrIPpvoUHnFDw0R6PQLF9sqgvcalZxhMj8jfwFNB6JpL
TOgIsC3x/qXAx4ym3B9xGfcSBs9ynfx3qBc7cjDpz0UOIYAm1R48EStVAp8RXPg8
WzYfBAWTH3D4PdNQZOUlyWcxIDl70SxnDukVNUYqALon5xj4cB3q4rCrWyMo1jeA
WfNPsBjIL+cPUutSvnpYwKT5bFyU6oGimLKTaq3ZqVPKk/RtY4q/hGiN3FHoaeUu
Fon33IXpDFdbydVhdkhIucJQRP9SNfKTtS/dAB6dXCoC9Y7T59Bv5wV4RiqhOZ7o
J+8bCZdP8O46i+B3ofKLnxIbnmDHUXuwSJFFq1FkssWDkmYaVWLFo+WLTyjeiNq/
BEqsXh8GhzHJ1EEvFYYgzExzaNJEA0UdAcG5xQVUV0PtZ9WEYx7cMrK4R5Xy6njj
E9jNFEhJwOfHler9lpxUrg5JDpP4iifjD3dsN0xcZIG3iL4EVGFhIO0Y+loUqnui
9sNgdifXEpZSPYZtww86Q/1JCpiEy90ZtCOIOJNoTdD8jp2bvFtSW/sKzCQaTTtv
YTzd61FlXsfrP1NvmnK+um7tXVzGdb4RH3rglKF+11Jk1kC4gxTEuxF5Zcq2Ypax
sr1veC7BjRE85cIKIW9UaMWBQu5+hOzoShcYCfNanxBz0N/zIzy0JleWDnkK61Ws
w90JYtuI3Nyp/pnng43PumZ6cSdJYaH60V7NSwEHvl0EeFtUpPKjbl84x9gPVKWC
Q3nCBq06ed+miKpyopt+KrUIXSxr72lEMu6rXXEXt6wrcu9Wq5dy21LY8zoLHDNW
glvjfFuunJU+Xn3/fyF9lQt/u8UbQrDVheab+sk6+o2rsVV//xtAtixSQ4s4dkwA
cLjUuplAupRpL4EMGXtAKzSQKeLuivl4vmbCvTZ548cUgoYTRWtDx37p/pWFhJDz
yBqmQhbGatQBma7GQLBJh+8TuaPFgiS0MMb/NMXeWnxInAgztTW8E6UMeLqVGY2Z
Z7vb15Xwp92ok43ZYEM1/we4sEJPW67lafChQQEHNIeGYd1762nYXUwOjSMm0nVu
MVksUbY8TzH4BU4cMtshEq2j3irYRJDVw0KFqb7WbxTbziXYasldOXAjtJu3wRv/
w1OVe0YS+Z+U0fbFx10uXdX67+IeUAUM0mpvpG74PclPW28P47k4SlMYQ7qNRE3S
hdsRQok2KnOjmkPwGF5aAcDyJYlFxIg8XakU1X1bmJMtKQ/q9veHvs/UbFA4wPsn
PPD2fPbBLjqvu3KzhRWesNFgD+K/uEJ+yO7ALQJSrwrXWKTmE9hnljogJdLIGh7K
kLiTbl8sHNyzQQbGqnXhPr3wv2+IrS23DRzW+V5y1CW0m8KyZmID0huZ+XyMtaQC
g2aU5F52v25uRSn6xwEkrZ4tQkMWf/SvlEsYk+b9JMBfxFbGmAw760yXlQkFSRpP
Zs7cRiEPX/oY8QXOK8U7Mzj3u2ReAv1WH329S/FkBghBDLUZiixFDBNmrttdV9FR
W5zG8vCo8FZiUaHALqb/3JdA0EMpCB1P2tqcS0CgRqQSqDhyzt2zGvxVi76yYIZ5
JdpL+d5ucwfaeLRINkmcT9Nvo0QOLE+OKFSjyxAcWg3bWyoyNnMKqpL/Bpgw6NdQ
E3YPYxT+UGNqM28xbn8arOCuEA6NikloNLxcQZtefPSF9aikT6mm1CUzFJiJ7ZE4
Ug1YGcjTx9XAbMJki9DH6RzNqZT2M1Zot8zjLeVZLm1rBazPK+saryVKnhZ26drM
v1zs3gl8/zR1l6ysD/1Y96jNEeD89bfTEgMOGOoT3DMmQFZz4flCaHQ0ggZAss1b
jvNbNtSF/aMB3IXEURrXBU//OcvoIiGAn+enINweVNZw6/pCVnSEfdlhbq2s9WNK
P4/dFaltxmLq52FKPwM9tuvC6KFfhQU7y3MmBBNR+YyjEbtNDr5m55kQnFuVywKE
BqikpjsMD1KC/YIVBVQok/KozujS45DBdxXrdTkQPiigNn+2TDGrNNJ3Fo0G4Qx+
3+JQqClTg/Ugse/uUBMYpjNOR0CNz8c9BQ/O1jUVhWDe34B2HinJB9gdavbf3N2g
H3jSn38xAxIPh6zqGz8qmQ4qZOrzmsiUPYPqjTKXoWJ3oF3e9qyZUKPlrgblBOd+
i2AYXKW6YBgbZnFHa4wz65uGH/mo5rsfw/zR+cg8ZYpAwGBSt7auzDCop6Dcsn7a
7NDrHOfav6FJ/w+5EhQ5Ohibt13DtVJ8N+U5cYZmB8G1IZD6fU3RyzR0BuWVLuQS
fZ9TL7C7oafqpgew3JflZ97zjOxUXAiXli/IC7uBB1BWk8aAwC8/l/OJrsX6CgJS
OYWvzqgTw+JK6ICJgRqBE9X2SrV76vWS/Qtjc+tXp8Z3fiXV/JeynaNM8Rp+KYcg
alipMxedaBx49mM5PSUgFxQIB/JT2JJ9wHHCicrxMN13HWDNZWUeJ6HKPV4CJ+Em
0UkmwZiwJMr/5nqULVxse138LTFu1kujrP58ZEB6piXTynHlQcpF2OokSS4kHcZq
wSeHu/Kw2+pbLC3Kx08UHrbwgpDp13Ri4dZpsgPQ63AhqaW5dQZlGZvxh5cOmPH8
NOe8aRSM7XkigJTcOdy1KzXBCf1eeXDFMoxOppwVPpHChssZOue1PQngATowy6i/
y5CUxVyW0pA1z0Ac0BVGvKt31hUiOGL1NyOZ7S1Q8dUXMC/2JTgaMVo8sdGoAqsx
3Sm0RRA8CXEmL4YunA8yNAYQRS7fAXpUZG98DIQtHUv+xtexniE4X41l6Pp7uc+i
GpUYnhgzVIDAi7lSmpH7K6wXZ1fXjHkuFtjNPCmD6YMu9CG1kVXPi/r7yZmwcnyP
TkN3vtbBgjML6MknwXP/Y3F02soMf+O0AIR7OEZ2uL/qzMc6yCSEZ5qIwcmjlvdT
6N3t9g65sN1ZZmSuPEMwYNeK7paQQK8dm3IfogEJmRNQhvxPvHVR46jvqAxKGZ/6
VitO5EkwHyOPKva25qxRemiiYrndE+1npVRuNE9itB1aWQze8oPIZytYg1Ya0cFr
VwiBVXxU5mYcXe3yVrUVBGyGyitVqxavOXYhxT8rVWCA36Q6Rm/dFD16xDgqHYsO
EzOBeQZxCoqfU18TD81iccRd14U+LlEamdPWCQoz4FEybmxfOPe/BS+V0xG0qMbF
mQUk5rqvwP9o9iOK6MTYhSAWBeBAMNTwUuSR920whJnYbgug3kZloUQptN960HuS
oa0yX6C1mat5BdJNN5f4ngEBH4/HPJUsYIrOHzPg0bJMmdS3UjCWqCLEnmlySWPN
n1N0zuJqylLyjqm2Be6CneC/xGNKI4HdEjbejEcTCR/iQx7r1bBu710PDWKGxhxl
5dq/fvoh59s5c4+34lYf3HMXL+mnKITAzH30AZSlnwnU6rmMJ84pdgd7KQptUj5Q
stLu5Xw6F6I+hNamXl3cl5bOXZzfidQ/27WisPdZUw3VR/9+8amPpBdGUOzYRHiJ
wBhj3dag6DLfPWuVzKEybHzWirQdDqDR346+LkhqIDUMP7H7DryILlO4GDLyZXrE
EEmK2cVS+g3v6n74aITKyxUiyChqdLH/oMDO7YYP6ce9rhwNGkNJ40YmtfNtIf/N
7fXa2Y43Eka95Cy12c2QSogwUrEFobSLMaRldHUjqkk/qrTZ5aqbuATfWW/Mkyg0
MdO1nZymZajILv3WAiYAq2hU4/K2pD7yiWFGc5iSIXtIqiWkETTMn25rBTlLnkC4
lm4jhqdantY4oJV4AWPq7FS5tYZ/0Z8Zu+YdFBohT/yq37wz1a1tAJL+Atg6s6tI
81MErH8/0pD97OR5kBOs6u68JMNfqn7XmA7l9AYJGpb0rAN3rOCMXgEWhmZXSo5X
RQBDLyV0QyiiTa9zmQPXFQs6f185JsmjEmhvilKX/sifEmLHCdtJb6V/4n5IW0lf
z3GrMyC9m5ICzIzbJwo4bhMHsi5Zx2LXWqM+eAepJB8TkIgOJ929VVU9q7182b1N
f9LzzDwIVH0IvPqi+MnjGQ2KS03sQtdydHTclMNIeZjHzk7ziny1XmT7bvhUJvmj
Mp91Egokf8TqWct2wruj1vVCU3SQ1S9UIGYghPS65uiGfbRuvsASOTk7Yqy5XIud
lw2mgVFHRtii0Zhs2ASF+7/ZWFIDgUk516cCmJbyJzb/n0XeJvJ7jUnixzVqnXvr
eHv1RbaTTI8xY8by/yQHVU3iWjPiV2bwq8Sp6kT9cdeTQ3dOdBIBTHn59KSmV7an
46UzPRih9L091uSleURY6XAtniXOOnsDuO92MyGOCG+ebEFuMHt57PtYfW/TdawG
kClTHGr+nKkGfXngmWtBvwsE6LthBc4JBC5NdyBbLm5VGoFezEAkSUqv4nxJcLG5
1jXhsiMPv4gycYI6ZucNEIFe8V+AEHj4ZuUuqXlV3iCIn3tuYjTtHtV1SuohheJ1
PkDLNacUUBuiuM46GsOt5kM9NwgjdwafusW2W4YwBCHb0L238G40PJCgas7gSNmV
/QOUC+OBPvS7dGDANqVgs4JD/LQmomLTeYRE1vlPJuI64ObaMe94PNrTV9Enkoez
T/9g0uDVamsgk1/tfkIlL32bXUWY2bZu6ezNxoqGQxPw0kIeGbp1SghDCXynTlR6
von5f04P+4eq4IYER6UMulQj9+tbqPkgKfOIqqlv73/30X7WbALUN/VSw5CseW4V
q0ELW4UclT8mojhHUQsq+vtWmb4U1DJJz7+0fH5kf5bzgVy2lrN/0FSiWyQmWzWs
JPw7AhpuIf1jHtwZtKs7fjXTtj+QCbtGW9ADeAapd0QVqNNDYQiFitGJfGXc6NC1
Aqkzuu09nlOCzSNgJcJDPUbYMwbZAvTGKJawMj7isJAQ7N6S63eW2T5BhZXOfq5S
xIzLox5jD7mCv9La9L70wEC7vJWVk44w2N9zrtqWaYdP3WkYGaDUbhxAS00XBx6P
G9smULpFGKznF5G0L/Uhmx/Z4Oxd2bLtgheLuJrT8DkA4cUWnkuqcxqBfuqhtJ3F
RFFmz2WOXiCXLoKTSiAMShK6uswDOgfroqLj3DvCITM8dsQWayw8FXvZuo5g70q4
CYV5SLGXuQ/FKaOTg+FvoZ/XQU9Xntm28/83rSMvpCTeibmBZPhCMNuNq5xwCZ32
WoG94Er8ase+/1NdIGUAsmI0mFgelHdvZzhThBBrmDjwFrFF4fpQoCfIIKH2NBq2
+VQebupn99r8U40aAPfB8M9pdHrGtGrBhHiJUIQi2EiCdSyds9gv4atMsc2/p4dN
K92pS0Oo7Cm8uRvSg+oxbgdHqiMfn575qEetxGsNwP6caJWEQqqKjm4ZVa6HHVfg
+/3rT10GmFqO78W9R2U3qjpikKtfxRQviMRvuPALZXLwhSkz8gxswgjWUYE944uE
gSSFbJZ3CP9QrbZSwBiiC17SM0Le6GMmMkP6jsDPbY49tsl8JSNTz96Iyv/n0yOb
2Mk3EssopOSgEYURhx+xs7N/VnxX5tpzfiXYcyJ9qGPuoTy0SGc2AqcJBJ6mJjAp
IPWXeYnEidzhTSWoVVOzN7pAc5A07pcwHj6YdxjVDGR3cOn726yBYDRyl+ESTqoy
UCI5SkXE7YzJ8A4ZhHzhaAtDt4iNxt9Ghx1271YKnF/9JGlnCpcBgwy2aiHhB0B+
MNBcJSHCEVtIjv5o6YWxZkXyWJc6Ix2Zrm+VHtXkLYS1IkAHXoPJQLjNSSHfXX/J
tQVGsDJQ4Yp3dRSe3l0eHqz2exoML6s472ZRqsln6pz7sQvsj4vS7XETsF7ukMrn
+dnYdfSCA2l2JsLCCHlXzBQj2vRw7vGvEsVvPIxhzVGGwaK8lue5/2RF01z38qZW
7AJHdfMTM68/fuEVF4Tunai/Kz5fn0IJHI+TnESJ+taUZnGAimBTVI2OQBP7yGoj
ZZTi8YVPSQnUf3M2VCvJ4bKS0vkEIJQtIZuHS6+YApdVO+D0w6yNS6kfaxYUu9Gv
Gr0eAmkVQK30ES2NTliOXhC9zpB2VOymXHYqLPUKhN84B7V7ukbqnoAdrPkVsBUw
bhGKPC1paSjC0sRAfodWUh1W8OyvPzgkotggjgxy9RnZ8b35XL1YXix81K+UWNiE
FhAYjCop47KfseqSreoQxNDfNDYaGl+aLcHk10GK0/fa6pzcGxBfjI4KfYLyHm6Z
pREBuvdDAPBXXvVyzexv7bfoEkOi6hVxN665T7mJgVcT4IX7P4Lid4p2Nd9pGhAE
zX/HGLW9myhGRn4pgx1ERkmC15Hk1XEUMKKVbnYnxbTU7Go7cEPTgB7UOe+dcWvF
7ykTcGX2nDtrpq49TJZoz/dW8uL0w5FSPgptvo+qiDL+dsdTXj6MIqFG5G3bU0gq
AuUXhIeKeXRqXebERNHnsxhHy3CZBFkErEJ3ty95M0UYHskyOAyCPxccmPwQVZwD
zmJBR7+gP8jdyZDkkyS9MCkfiDRjpvB79p1DzDNxIgEnuITfW/JU9huZKZGFr5En
TGzUEfwCJ2r+Wvc5Xd/C5h8O5CvTN+c5V6jNP0bvAMeHxZHjrhd8rm2sN2+57t/Y
rq9bVOt3yrTetLDyncydxPN8QWc4MdvKszy33A4QAHeJhT/4Q+rDp8ZKRqRlFE7N
ZyDgPYgGnxDvnDyWb9ish17JsLxa3OUpkNAFUmoEMwCU87D7k06FDtIYCFnrd86q
cC3CwxrfbhArYkcsdXc9GYDunaiSjv4VqIw+sfCgTHGjJIb284daD7tz87RZ+Yz2
dx85MTlTqsyqgG6YcUZ6nD0LDyk9lZ0pjxWP7BRWF80XYlSbP/tjuzg6MeaL2vMD
bTiDqwxfw85HrvnI0YuJqHd6fF0HOhx0tPY+g57IzhrpARKU4V+Mj3huDEAzl97B
Pp4blnsHIunJtVlHnxJ/FOCsFnpUswt5t14hdvwQPD6iUlrVLj4DJqoAwddo2l9O
MO28RydK2WRcEUJn1hnixE3Wm5rcexyNqQ2XUI5kAvI4neJvBGqgeuH0xhDkxHdE
SC4vxoZc/2AGi3HzOTj6K5ieWZmzPCPnBrD1wvomLDb2pCY6L0ltClvqtrrb/Y+/
g6wdqf3w+zkHgxdADPebUP3KVew294NrVq4AoNNjoaHyD/1WUzai/crIrd0pNhSd
Ke6kWus/YP6OEGpZfo72GpVyRDlN3EUHiJcreFCc9noYrAeUlNykVhceLfwn2Vv5
3hz6sdELK71Wb8WGjuIJJJO/YxUggGqRrot9u+SFtWwNyCQ6TtOCrqnmeFneZd80
3hKL9sdD24Lvip0Y+KS7m2aa0PsjaDh6y/9tInD71JIR9siVENMygH5HIDKBf7Kd
UMyvsVHp+T08mhA2zinxi/WkQt5wKInYvx5GnzLXkC4R7ymyRRNgyIuSWSwXuxno
7nPE3Ht+8DJqIrIzZYKafbFm2YqCpnkRclGGzltEGReyhl1xYe73gQN/r9+zqZL4
eaoD5jhsCMvgHUDsDNvuqyuafHJtfmk9SHuGJw8B4yyhGnsmUQnkPspVgEl5UqxV
laNgfLW0kJwDTtkGvp3mwlLnS2aikwWGgrGeby5YvkEz/xj4ulIv88yheHvivmcg
JCU0Kmmv5+v4r85Ona+Ui9x3pa5AMIwg+oyqQjag+jAbkUdc25vwzfd8DX429D3y
lpQGGSEbYFxquD6PO4tKh0h2c/Go88aqbhjQ+UOkyHMm6l9paK29va1gzpanTacW
6FWEWWqAMV8KX4rmpEkaxvovDCGUhOIfyQpQK5nwG8PjbscOFxKotZ64cKKoCFTz
K1WQnmELKN3n7JUHvFzNmUusW6caDEUj9n3qWKFMDIG9hKJzN/NWkW3NqjplYw+4
BMt2eLJP+tJgfaS2qYZvIE+Wc0fJnJbBzUpF7v933Gq6dgQGwUPfggwL9gw9xxq0
OGHgro/LttjOBCqE+6Y8NiEDIoDQx+dHrsDKZK8C2m6B8y27Gj+uqybYIMi4/QXz
DniBJ/+Fwr9qQFn2ZiSFeP5wYFXkZts+ygH4/d6ylw28Rul9UKc0tCRoTWDU6Lf+
kqiPIh+EK3PMv9mP1E29kdtzkMqXfTTZj1Q/HIQK2nPZhJT2vbLqTSuOrNAXmTfb
79KbVhn5CNBviTWG17fSxfqMxDkDDfOKmsMq2D8KEZJMpXhr5peDA2fEuJcz/O9i
oChTJjahoCw2GMkYtH2XCyiHVAnzwleDjRsHzzluL47JwOAWt0LI+AgqIOqbjrBw
OTFXCYgp1UzVKQAj/RzcjDvlnwUL2frVbL/RWVx6dFKS2snGxaN9Pdht/YU/ziUp
WOxY2eZCpFZpDmQnDY3MjknzickuDlyc24tiPVmGqiqn27kUQ5kZP2uIzAJvv6fZ
jTc8tWUgXC/TimS/mXbiOFGsRKmRBx2r4myUgUBo07YKB6k3G2HyqaV8Gb9BuauO
Fwztq5J1zBxDXvCk66FTZ8Q/1czJd15c+8yGTVIPLatrj67TgZWoFKOiTTNdpx1p
WYHG9A7giLlZ+I1LpxDJtjqRLoY9ueeQT7/br6zN4NKO6n5dL0L3+fUbU3wJy8ap
G5WveJuWJwegt0gLeLcjjZRU0ph4SiwjnogyZEKH4hqcYvZ4ZtQ3NcxShIzKXfhY
0Wfzd4AFKOfSHsmbUHgJqj4FRGpLgt46gAKUqoOFSgSPuD/6bczil7ST4ZO10YE9
MQx59MQA1414B7DUkpq5zb61X01Ps0ibAJNSEIW/Y26qpx535WqahQzTPa5+keBw
EitBojvRQrfNnSUKUwzKRgWXZrNUctvtLBUf6a6b0WQ/rSxh2w/NcOgvQHCBXhJP
4B6Weh3sZUzvGXJP0ISAD4nXQeAlYEME6fxh3O9hTeS8OgSQTjVkqIlyK5Brusus
QsHlRJzUMN47fDx2SvrPILMhMx/0iwMqyc3nv+kKbq9Q8MP+d8oxBuBXuFNhUb8v
8gRpvmvZMRdlLjX7PHWoE6bsXd6Y08j/89yNFR1SUN7QxjFvo0HH30ox8lx1bKHX
b0zXxhP4YmwYHomg1/svCV+9FhKCH2apiw2NtT2RyvHiw81t0txFcmHTzB6J3uPi
mXeq/P3X+AjJ7axy4Eo+rCVcHTu7+6gnSkcBbPP1s6vbQ66qV8o87Hl4pDDeTukm
qlEJZw6bujbo+3kOS3xGXFfasW3ur8ZGXrj+zBO78hg8mXZQi10ldZzYCKj7+Duv
4Tk/Gw3IMzTPkD7DAudOGWqOgEgqw75SUjojEEclawwG0cl19ghA3VSjOqEwNpqs
ioeqi2ROMPfZWziabppFn+7gy9yY7Buoy9Mrd8lz3XBBHR8UEgIk2ncRWBpD1yWy
XFasojSXd0FtTfakdXgXAPmYkYz5yIHyvtCqZZryYIS4C6TKNI3uEcm78W8Fs0H+
M0r4AnCpnFBxPQrLMWJr9ER09+PcVB53tcuZLARg/s+shJ3mPIIuZx/C2m4iJ4wx
JyUwmK7CAImwXyOrGipNHAsJwLLPTJhPgV9CezykoNHoL7v3OUlUgMwQxhi+wSm3
pxk3qqoxGNgkTal1oOsyyW+XxGtu7jev6y2vo3rfmoKh//zR8YH/yFSZ0TA81r4B
6XKHZdtF4gGqFyl8rtVdGQ43s3w5vtWVw6G0OhJRE06AfEo0jjmam0VvJSbvCadS
Mmx2q2bjjSNaeZlPImoRkih1yLFMPv9EGm9ZTt9i+dyIIjdg4ZCuQCAYL1uufUti
qmp6RuUbGqPPeuwK9dBdbfaGm4XwGTKulY5PVAhHWcDSMbNLbV8wZQwebf1sqgIn
xtXxdtG+TSuZJEUHz4Uh4253GZy2SJ9oZ2QRrtHxrFTuua1OUTXrur0/DB8EdSWn
Ko9r0QkZKVbNSzdc5t4Cw+GSGIHrf7syiWIuNySeGduoPLb32+4SuHwfj4E/Luxc
EPN6XQH+j+LHrOApXqEchDk44WbUZs41BeOBUB+LEb9+WBxny8KWkwzxATc7I6Nu
WeLlzqMcGx+2yr7yiV96bZrkK2wd/c12Autx1it7zp3RW0W0GoEQAFU5PBS4EwOt
dmD6EbcpyPkRvrOuffKUl+Jal2a+8hOk6RUSpE8AjG8hIRyzQThY5OQIvZcQ/f9X
dVz0x9w7+Vhi8vPjYoQV+XqlS0uB3HBaRPAav2sPzVUXK9O86Q1qtqZWpBFoyZLd
sGI0I4ihq+oQAk6onUPN3UFWadDMqC5inaBAdgHpBGVn7InzSnv+ZNcWK3aQHMpw
syJ7CNysQJmfVGSBdpD2I/CTwyb60I9AKC5T0MKZTHzlsdwjIK94d5XXsLRkzwv8
oct1SNijg/XPDiI63mEEsa/hnHvzEe0D0u3wnhWymdVmNAQHP/0Fdmqt8aPrPxRm
JIkgfzW/Yt5ZcIkGpalFPML4EZop9Jv9bx0w+vWalTS5BbZAhDiKI2WS/vGTQFR8
ri0t9H8G+lDeIJYtCHxatgeIQDFrnGZ57b6O4GpuSPyB6LBrgYEAS4l2YA/LT0sm
0tjmmLLExETueyKas0z3UJe0p8mfHEPS1Ega5dVz/MR/Oj8I8YRLNcMcGRWQc6dq
0laiuJd+CnpNNH3+lkXVPQMIqzRkN4xicixDfVEYIlJr32H7aO0RmjG3ZhDqwMui
Zz4UdWSmPnspPe79DSE9zjyH7Kp4Nfamch5uYp1rgNDXRMSJjYx7ZdiN7H7+sW+9
K2l8Fsopd2whsix/99QY/dStRT7hFCOp3o2T4XREAOf8ip6cOERMD5aMumPOX1Nn
h8Z6I8TqfG5AiBuaeb/NxbyazN18smLUbaUMgFX5DSN11iWuu6XqO+NeLDVk2UOe
FoRT4EV+gTnqqwNpU3lbUYxX2E9x+IR8d66beun+TGSf6uXSOZbEjFa5hnzVMygx
ubJIuaJwi563wK4mrguJ09AkPMNNN+YBTLnMsmhXf+Aqs954fXNB2SAqydyT+o4Y
eJsuQXQf2J4rnedV6tcxGzj4qZY6bMZ8dojUbWFwvCPx/XSylKAjh3tSo7qYUu0S
2snXaw20Rfx0aSZtVAHKGYy1qU+355ItD4tL1G6IQJreqdZVbVIBN8Ac3EZz0X9q
kcmGOaO1i2mnQMghY01Xc2yFpus7LRN2wF6Nd6H5FA0uZIPDa7/OI/DFwAKvK3Qi
dEAlPcHDvbK20T+NKpERxXEHRzoj1lEMLNfUbvvwJJ8vNkKv6xeaf1VpgbAQAQ+j
5um+Kno1KtZkkq+mB21ibBnD1w0eIIQvT1kxPUonm9Xe0TGJYagEsmAJYrWW0Zap
xZ5pYQdhjr6+VBnB61nPcqEUWLk8dx7j4j3nF/dQCFwV/oiMnC+c4r2LlaFgO/Ae
/UO5zsvvuEo96JplKxf5KDjLLb0Gny8rsgW0lwd+b14O6c9iuQIqLfB2v3/B+1QX
jK4WetMv5IniqPkXa/kPvQcXyhv3wA41aiHQ47Zza7LHiW85eMYStEcwd/uP72+t
9LoYSTQ9BT61+ItW3iN1BOdkcPtTERp9Wo2YGuL6SPDu793Ozp09KKVt49xkulaL
zFKJFAxvyaMFKLU9uevdY9aevDda6BzNimrDDsxk7BlbQM1/yguyB3EV0tgdYICi
5Nl3c3Gv45bGr+sh6o60iwuxq1rgQW4VtnKtDY7Ej9fYVZkXl0MevAW2wOW42ruU
DlPg2CClUhQ1SxP3NaMcX5jFtnm4TZ3mK2rPSzFPa7vZUjyPKAFoaiBfgSrF/2Ng
+sOCX4+9vl5IpyXlWHYbI+aIPPpalwV7W813BFSzOIqm5+O4by7n2NgiQrM72D38
ADd9A7/i1jsA4CJye9fdL5Be/h39t4ya5pso37YmIy8oSY3x/12uT0FU8rRXT3EY
mm8jdO+e/gc3NImMML3LmoHFESONjPe2eyGjeV2S6EZbqiDhyT7herc8p637RPdp
nJ0W+cXyLj6kgx7cz1MaZppn+ZUbs5pzYrQLIKQFUwMWYIL9co0W/eIG50LnGDqT
Ag7TeFTKociOEZSeefJicB49tbMr+0TjWN2E6kFczir3zfhKTTFRRWjRbJmTrdKF
yX9PJUBwhT0LzPQAsAB+QYk1c/omw5Nm4ajb9KJw2wI37DnMWrzDqgLL35O5uHAW
E+jg7kJlU9ABsJcmCx9Tphdkt4QdJzc9r7Gsq1fxxFy6XxUcc5OIkPgX775A2wGt
TtOFjZf7T/HmVuA7L5j4IjDY4hzPEGVJutBNKNYSbhLxYjw5mWBcIPrcKbOgKGXA
mVa4OLR4uFbPRT0JrU+szxFQe5uSFCzSq1nEM4axKTNXE+iqJjUvJCP1POncdn+K
JVvcwlD91Heph+KOcf+HHQ9zrE+jJX+gBEJaLnQcC4bgipiEhwRVhsCD0l3Yzp7y
ak0UsW2knQJzkQHwfick2KqVdTb8eX8t5q/F9JwIXdsVF49qd0rrOuoaDJkJVRYV
WwyciSomE3QuzX5HaKi7QHBdl0ZGP2pQB/dPrXued6nellV4Kdnt8gnM6SgUWdD6
dEreCLkyYHNnIdGeyYdgAo1k0WlsXTMAUpp4Y0S2coWpvpzWn+Ymf6+CicopwM8P
p9mTsJTHEnO0IRhnIW4dMhOQSo/88nFX+81fG7b5yTtWrZFYhNPuKdK8/TonXAi1
JvE6/GX8MHS+ARnrXJCc3IoGpyzIO0V4Sj+NPNIA+Lb36pDfaKeayCtWJRY33me5
e5/KcXo5LFuen7ifccpe+qPOTe5wKE0BT0LMVa5zvQf5N6vQ2Jy+GXWm/5a/0tOa
ISEXFkFgRRAJ7Ykl2K0zRY+ApQwEJomO6WzoxtN1Qk+WhYCEe42xFJQlwySjxUj8
pDcTRtt3e1Go/4x9XpztyVTctokzoaDLVkIu80kiwbunXJsQ9/N9HxixvxhCQgwG
pMbgsBnamToUaZyJ8wyRAvngasyRGLPLLALAq4OsX6Me6i4bv+jmrfAbC0X1o/zt
sQ/DmC/r1+ymi0lEj/4Sh2ONNGM/0QEB+sCTA1kqPChd0foPy8gCrZzkqki7rwM8
Edt3IWZDah2yzi9LTzkihz5C2si97br+opDOkyXA7UOIzUcFmFPOjlhbu9Q59MRI
2xErpFFTUqX537ex7Fvizy4Xej3bATwcee0Aw4bc7NhlZjvrPtRtwMMJy8gY1XCQ
DiWjgxcdsw5OlHTY1WslW1y3+6aQPom3XIbRek5SHXOPfJRdeBXvCkH75GPRhW3W
5D+0P6matyFRd2umt7X15eQB9yxTRph0eUjF710cHe3tabx5yNoTnKZpasq0X7Av
M9QVUoS5Jnu7LCB2wiJfcSgL4zoJ2/xHJNLAwoStqhuAn0KPcd5W7IBAeye7GGd8
M5Fl+RFnRtOduQhDD7akNWa6jnVCNVveqjX9S5C1ToI8rBYrZbDFYjT6TdGw5jz6
pXy1G9Xv8QKfrHuB13MpaMy5HS4+e3ByzL/qzDLzRA/kPu0DjNQonk5ykOjlYG2X
BBQVSXFPmnGN8jSnYwx+bK84EjMFYmZzN2etPg22SWjiCMLenswQxxkMHjkvTgFh
sWS1kS+rEtuKiotCRQQHXZfOgA2ExgIl95elENugI0AR0Y0fMSEDGKhtM4Mb6Dw5
EtwsNBAv0O4R+tyjFOTyxaNG7PWRlk1j++OXLMxsT7Cncg+fVQfIV43eXwIDQoQY
/AmwYxNK16A8EhZSUU4M2E6tUMAlDKe7iFlxFFrvr+bHBsY0GvGT2SwGpYLTnF9p
3W7s/XjYIccl5UduaHkQbMHYFJQT1CjHnpX/sEhlFhrn/CmlR8A9Xa3tqU+LRTrt
aztGwcPqXId+F8oIkItW9u61HWq/I2ySqvPm1YqZtIDsN3/BXq0F806MSIvKBrIx
MNsjsFhUuV8p94bnvDCAUEyWebiTDP7brhbMv8kpJktW2IT1LhXDI70PqdbKW0FT
STY6r+iRhT26msUn10eozD1+5/UDzByNbnBdQC1B0PnO8L8TgHbePM34AU9hVLVX
vaV+FtYXn0KG2xs01yHqQtO5fXyaBvT8WKxcEV3zap/rSYeSnFnF53DnthE+jgIQ
KCXj3NMBhnXAVGlDUGKZjE2WkclYQL9OKxTVw1ivAkq4CN6yDw1i/j1lusfXaEvF
8j2D5uq3rYuqaAb3UZ1Whz0LKB9OxtC9+F+58mKRGzyTcOM9sXktBklb8FPrWP+R
l8AkroPB7Dma2v/LqsVPtnq00J6tEV2idkzqDSDRKvA=
`protect END_PROTECTED
