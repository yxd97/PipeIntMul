`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uC+CXbSYBNOvqa3G+qa5cuiwvmcFYR2mceVLTYNfdQfNPoNUhXs/e4AaBCP+Cu9n
Nf4S/sDoTOMoBEJ+72TuU79cCiouL93T1Obef9vXwKL4MBtiisRBltAZdQjAmssV
xTcx/8gK0V1+Xzl9c0b5ZVMsscCdHCNWJONGnqgsQC706J8iUD+BECFd07SHhAC9
0NwpdhluNoGK/jIy6Q0hx3Zi/ESrSnycmNOYuU+UACRS/Xi6RwhT5ZP1ONuekOi6
e3CkYJwM9s2DZhNQEE7KeLWkzZguXDWGQqXfJ57sM+h1vqYsZoxfHR+/tVaF6XPY
2HnSjTGfPYbXHzeBe1KtuzwTgU6g69x3f/7yRioVB1lhiIHGBQp1ZiQw0JF+RuRs
OXky6BG86up3aY1H3YtySZVbCSGImA5y/OKLR9js5mdesbARJ4ZI6bn6UD4bC3mU
5QAoXS52aFAuIxXtu5/gwu9Z4XCY3/lTQgtAZlcUV7H+fdEgEiusVd1qYcy/cz+Y
`protect END_PROTECTED
