`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W0xprD2csFMvZDXV6Jy/LyP+cF7fRTsHODwPGMCRVtefwEwMxHxhnfGb5KV6NJBF
uGcDeo3tG8E6DL03Xc6vgPv+FekNu1yzuh2++Qvp0tvjG7BI+z/Ofn2Vt/bZxodF
yIdVKR+HQ6FoDzFtlTQnhQ40TGtZ7QdtLhrp86tZqsZqCfOjkeMkESTxE+daSDrZ
/03NEp7yWb9INPnPokkrD7FIlcOW+aONt48vmQBVk9Hl6LDBrwOGMn+HqabyvT+j
qNrh6392BhIK1NB4ZIDQHXisITiv9mkEEWV/7H33vinsLUVHzEsGgX/nasVanKid
cft+Je3RZ+L0pi/nFBX7SkbBa5cm9pGACm+0VW1SgyQjjgEzGlahP5PI875L99M8
zVc1g1BTfafA61noXrLihNfQ7Hil0QxqpmmmoDHVXWY=
`protect END_PROTECTED
