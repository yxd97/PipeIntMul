`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJa8DAB+sW5nXOlcwfnUtSCToAsh0WeHvzTps40FfWRF3UK3Q6gfPnGVIAcaoqMG
HCEIcVZ/r/PvzpqBvM5w2IsJ/ucEYhLKptNTlCZyjGKlPfVlEfhkI57Vzcq4pPGH
OkmfgoP+V1NoeKNhl/3WhWy3lOfwhB/QXRbSXKPCWZnq2oBAiFQ7lnY3DC4TdFbE
+DU6Q5ZpXNH2G8MPkFsw0EbAy3M6OX1jPr+dSOndy9ZAIQ524z3mBo9eAxo2aHSN
XXimSyOx/N1qYs/VWOMdYoGGweFT2mYNN7SeMjHL4vc25TTB8p9+aVAR/r2iiwqb
b8P46jpXEOORSmNrn8+zckurtiw+mZLQcl6MYiFYArmf6u+pbMlqo/tzj1XInuE3
C7qmud5YiV9LsYPNydRsIH3QLH/tIY0Se65nOf1vrXZVtC+l1jCy2aaxfE4xg1RV
w9CWxtBjuV6NyNKecUI3FYajxgaFD719Ml6uN5jS3+1OT5AARuTACF7EdukrhQSO
cY0T/KMUzgrmvlp6ZsgpwVSgUDGsDkosDEpUWPDIL6X+HYHMMoeTpWrZBFscLS6r
NVXJ+OVCdBEi/Sa0ltdvRBvSu/LTHj0pw2jyPepbHYP2UbQ3CwVKBafhOwxHdxMf
AbYFUn6mTB0p+JO8t0Qded4q/1pLDwHuF8WBOl7/flgtTLCtoBR8lrOeeLs8a2H6
ifX8VKVt3vYDIOF9ojkoAWzJ/x35mL/OzZoPP1xmN6E=
`protect END_PROTECTED
