`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Or0pU7bwc1YJBNYlrxUYn6lG1H6WXh4nSSa8VBqSAsu2BVafUk5tw/YD+Sf8UPYs
PyObDo3qKUEmH+P1knNbDlGmN1RFsTaagCoP1LemvpH5WosyS84stUOOCDy9HuNN
2gUyvWMLLlci2aJIQskgQYw479UiPtQszo5D16gHjMUwINqbSPKvz7VNpSD56LJL
OUPgJp2ztPSJeXj0upruYkZN4hF1GRiXd26p5blTxKv977H2nj3IOuRv7+HAdUKg
P0EchM7QiOfnYN2bxMi+Wo1eCzmFT1XPnUDJtEWTWXOl7eGAZxETStutyS9mchlo
`protect END_PROTECTED
