`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYpOLvx7MQ0JdNMCJ5UYzl4AAgyOYVbHNP1+mVydWeBhK1vER8/ZE4AALXNvaZZ+
6lpffqsr63icytluvwVhcPVADpHxmB4IuX9Lfp/PeppGKb6xK3pyS0cqmxaf+1wB
ifs19Cm3zsetv3ncsQv+YGK3/l1KR+IZRzpI+kIpGzY3qL5A5x4Yw45wQ6Tp8wxs
56gYSsVwm3utH0ecDwhUDOiK/p6z9tra/0klb1IZxL0D0047qrNCY5HVEev+5PDr
2oILeTEiHfSYqpdRAwU4n70JK9ahS0LV11fHkffcd7YCSSdBEZK01u/h5m9FHgg6
084zzYYZuCRAv32o5CYmaXkQdowtbMl8nJSovbP8REj4ob3bty2vbDpJc/HCELot
x0GYtAQyMWYUYqVCKc0E/D9km8rj+g5mzzHbHuoB3G+uA6FRd4VNGuW3RAxF6FpS
qjz4laG8ZyUC+POIuYaM/xy6pHKJ/GKyJuLMfBowM1r/E1c1216dn68Aiy/BokLG
pycFyK09f6+jSe0xmxqXm6D1rEmM2p5zBvgNealq6li63Butso48/Wkxgkeek5xY
FuMaVaP75L+H5WS3UGDvjZTSr6cHR7rVox95VoQBkr87HKLoxjKLgi1F+9h4yHRt
mn2j3D8zaRxTFwSO6WPh7jKR/jS/4KHNRfms8LjM6Oz3tYgYhTip5IX9lk/BCpcc
2fbuxt3tswsO/yZF1gOE0eM8s9u2DiK1my/qbX57Tb+3vv47QQ72wQuahYXVzM9H
L9fyBSGARwDKklPGWuMVkvGbEbWlcpuUDxFG9ELXfv2q+vxALoV23m5SxisMJBWc
UcD2MGtU8BaiU5UPsgoVkA==
`protect END_PROTECTED
