`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zqa9+6y+WJklh0F/P+HXuT03sHbH/2ena28ObWF6sn9GiDLQ29fs6N+xo0bYUK/F
5INCCdZlNM68aYAwQeWa6jGJkioK9mfm80UWEHBm+741xhoQkKFkIB8258/V7AzR
T8lrHu6Zry31vssZcSiRfcRKZOGxtIMFlpshJNbHxIw1b3Wcu4tmKsPURTpLUztC
DjNmTlFq1MAUDGnJbYMsMdNiIoqgOhzlmJxKCU786WbBrXurNNr14+/STRT4xS76
eKAwjeU4tmA/C7oC7B6J4uCJQzd2QlBILP8PEjUKANSiCr1eC56TqWk638jZGRYj
WGX0SgCPb0zvTjXt3k22zxDMFMmPk+ZaiEhoHEj7eEXdHNN8/zLLRUloRfNVWNZI
eAA9TE/JwOvORYg4vgrXFQ==
`protect END_PROTECTED
