`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnaMnIqYxHKkm8LldCZ1/BjxS1bEdKOzyNsStQyC0UC8QKj38RLeYU+2tki8urcz
6MB+BpKUyxZsPj5kLY7vdQN8ZdCatPms1eDJu121+JGu/DWUedFwSzYI0rStSHxb
wsW5VWwDusHnDCEONzVqmkmyo7n/OaO0XIw5WvksCYBtJLG0AP4PXTEm4d7zOix3
nakzJTdjzEZaHu1tOxo0EbXl6rgX2okqZ5plMHnxrwCAwALmPzfIjSMPZBUt9tpE
aSE6Q6fk18EcNop9IA2IiGWaCZrXeQhFPcolFPz+OzyS+NV9Thf9vLfHYgEtfN9M
t1k+JJBerEEtmUXgpMJauo4AyK4oKrXS97KGCnYwmaoitHhaG3bmdS4YEJO46wGh
bYIbdRf3Cv205UblgtabEuUho9QsbhcsSyj2lFyAq/3pGm1in2qkp3zFOPYpagjX
`protect END_PROTECTED
