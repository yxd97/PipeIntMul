`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYso/OWvac9SaNLend3mdscB3Rc88P9KVPNCFEhwYgvBjy6FVyd+s2w+4KZTbg+C
/PXYCEVRTaCbu2BJHvXPx/MbIrvri9/ocVTCkT33SnLyke6zB52j+DErCN/Y3UvM
DZMW6Rb/uBMv3R/J/01FJWcY43U32PFuGAmRfUZkvhtiuxxSsw7Vh+OVniHSUI5G
Nn1cZVQVdL17wgUmTTzqDmQ0gs353tNxiRbY4AHikCmEbsPYwmWzm5B3rgqCSQTT
6DFgK3FoFzS64nky0DV4u25F/dCQRuCi0puB9SUhsJHSU6s+O9UNVvRpAwjChitz
FyX4bdSSf/NuGTvxhVbIwfSgMM4A8cEXql5u3BnBzztXrlw3IHzX9JDEfA5OF+DG
O5eucQ/Kza4xhX+lnapTWArMWLhqBR9ye2r7a/jM3VZLfMwyAvCLKP91eatLBEA/
3pQvTFkSgSW/5QiZWcDBe/EpGL0BrX9n1UIjVmpocc2pfI/28tXSGb7WERwTfsdw
tAvdAZgfXUssUNIxJg38uCj3fe2nrIq7So58/9jlhX9CN2awRgb7UiwfzZL7/Sez
ic6HaGIkBaBZWnil3A/bCo1RXav6QA4TQAiZ7HXjtdci9TdonQFkYaiRM7GmeJTI
fXFL9lUURzj+n6AKo3z1gNb3+8B1XJ7KUs87cvskEFu195+688VZfA8ntF4WlRiq
uU/qDby4fQrCR/+TAiypygJeicAmbUUwkeDjNJSeUfD4BsGvmyf/fN8oIdG6IhvX
T04nXlCoDbQBhjJb1holWjJLQErTTMYo3ouxcJqv1N3SzNjG4+0UtKqMSVKALoCs
GHhoMWc+zjurMPmaR1GXJi0JF342VZwjY6ebTmw+/0DyMwYDoOxYmDDSn0k3XhHR
UKhTIaIxaF++SXTrt/E/CefLgly5BLjtKChhW7xPOoW0P4RJbIIviAPQ7QtoAzUq
f+GXmTvgkOwwN2H5AHDdWkcms+CDerQNbjuw5O11jgzeVCXDgztezM3mKFz0zjlu
1Kd3aD5tYRQxiUipykJ7GXqL/quUOYb+luxhF8t4hSmvDIz8g+x7sZmsoaQcI9B/
G3thqE5zh0IO1mx+u9esLkfYlJL7b0fhnc+Ekvoo1G/OqD0XkfB/xWw0FWETug3T
EHtJ2W673jUYclZ6P8nnXTSQuE1+l50dEEruUnU3I/t61Aqmubr40dqcdll2C9CK
kbbhDsG9UP4jDWEtD7MrtMNVq5dNYbtvjCQyMd0K4Bwiyg0Ri8kaDvncIKGxXhfv
IlldC/aWIDJXkqzMkG7KIy7oYX2wnTBwInaIMJw48NdpVWlxrxvhacob5PaCbDke
5YVDzTjGtb8qsb5IPwflFCH7WyTnH1y3nNv95i5aziMLTNVNRbriB1VOBcjKrL47
2gUZzBtGH6wlymCBLBMD7PFKbYtLdmHdTSPHLw9SZqVsDg43Wp76gg1NvzhAuVBP
boPXNhJxwY2wpwF7/MNSNfYGoXH0v9cx43dk74lABzVqPR/1QGUo66DFBqXd35sk
6HEq6YGBFvG0lEiaZUSOKpxTwqeJMiPlm6avnRTaYgx6UEHe8x7auxkPP/BV+26r
uXwWtpgwcVJOcjySkSGakZyFRx+H7k8r8C+L4b0HSAkZepn18wXriE5udi3kANdy
NTdP1ESSGnTnuZvoa/89LGUwW0ktMySEVrXlh/hnWc4NLwqzxQ4tC0jswbNLjbYt
FJPDyBLuF7A49U+WfvClt6Ayl31CB5dYGNYGEeKweUhSO/oDkoROb0sxM+BYV1v8
MU0MnsZPSvlqU8TZWT5gEyb+tNGM2ydwFZIwk6fVC56pvrmVzp8Csz9FagL815Ys
CM2+qHSxiW3puRvRZFyfC04RvySPMM7WTe0MIdjiNyt77kRRGFzbI2Hogxg/bi/D
kO93Gaa97NvTqC4IGEPTyMnLs9SOgTIvKE/20hP+lNGVl+sK8PjzlBZqm+dNJmp4
l8TNa4gCCGWi3KSpTahI0VX/8bg94nma7geHX6+BThp2OJXgKjtujKip5Zo6A9Fm
oLW5T3mlHS5rQx6WIQ+fP4J8U8B9753/3GL8pp68yV6CNTWkXa1Cl8t6cdB7bz2F
eP0f3y05PHkfs1O3R75ou59e/w55BkAhnVrNNNVpObvk4G2RZQJFefvgFh6HHt4H
rjk5Untwq0KeflOYEUWDIK8T3PUCypLrJp6Otypj3Aod7asKX1QWV6FRT2eFRYC+
pX2YK1TojPJkPZUNW6cIKHgZAiDa+L/DjJqGy2V/xLoDfp06FbiW4VnUajrRXpgH
9zdVgKclvUD3WxwcAQuF9jCMb8wb5s3eF2lNT4IGkdYeta+lX8/Gf5KcYEG+2F0/
Yg8BT4PP2zLKfbk1/vMPvMo/mzTR52CckcNwviL26oO04hqigyua9CyMTwzcVlpK
VRX7LF01I7upPgw54bgCkh3yEH7xxYWw/BgvDzOkntGeTD2KhLMXLY7rCcgqQPPH
m3o7hIyT7fjz7ZO5nTYOctIl4m+qrPFtOP7vvPTavgqY5cbY+0pRxU3zqTpZz2jY
yMwrJqugbBY62H7FvOWaDOGjK7XTGNxCLnf4P9xwTuljziftM2+m7M/DslbEy3Ks
Kk8xNwoK0EBOXCfy1RSWe9xkD61TFoMx8OcGqWAVOMM/7E6T4QuFmwXcq3HJkOX2
kqk5AQSGAxCLqHzK/xYHGmf3d9sFRnp9iJQtRx/wosQLP+kGmBLwg83xl4L33uQm
yqnhUC2/AYdyC7MeRCVlgYV1fTmjJlXjMbIuJCGF4ECSPKfWfGrRlySyp1j4N0bF
BIU7geNbWYektrBm9BHIo+LVi6lrbPbylxFrc1e9pBeixWAWDSKCU5Ar+vyZXcDn
Zu54S62IkBupnLg7Dj+vJapzAyPwDubP5Cj0sW0oY0tVe8iVfpuH6F6EX/ts2DLo
oPfeDMkLi0+hX+Y/RyQeTIRjPzfnB799IdynEgBi3/Mp+1rhlO0A/81vbmlkt1Xc
XVLOgPI9fxIms4BkO6lxrQvIosJHjcpxHL/V1uzND67GNJbK6TwD0Ziy8Jt+EgJz
AhwUDRoK7KVJ5L5hOJoZreD3MCd6DTpc1kxS+b/1ccoOIXbzXIr2CI9zTuxmuwFr
1Ee4qVhAiAjrznbHrOyyy3wtDBHxdwUbAcQ9o8/8Eh4VQc2QIDXLkXmeCw20Q/58
kqiRzBmKoCa6QeW54ChyZjrLybIyoWemaP9R077CCwKpGPgxDma4LxQqLqA6B4Wz
UAmG8YBhS0kjk1fwWuc0A2gPqap6T5n6bEdfU171BOOrVMX9u7PXo1EnSAUmBtGE
oTNVm4LguZL+YscJAn1gARV8+m+cxzOamfk2ocHIivBc+JfHDIf3LhORi8mZMPd2
W3O96V/TbemL27YteQuJsfbRiCmIEDxxZIVxPlj/04+6I+BDOOfQLHmyTz2RDGJi
l2nBpuxfIfqcG3a+itfdOnM0B4KPdduYNwSW3rZQdQzCpijAnKJ2oCsRe3RjvknQ
7aveFFY/ZA70mhUX+zzT0UwTFx2ucE06nBBuEXxnBi+d83Sp5IS9gTLwosix2hme
Zmw+y4sAYKYj6JVBXRkCOEbpyHTXT+6CzayEjO2k9BgzZvQlwNX0V6oOSBa7DkHF
52++F2fZR7wyqQu0A+JN+HokFjOh8pAtPP+qq7nfsT2m7uKhEwjJXNKHe68EnIX+
z/t44S3IFjQI97KEtsGv3ZemIg9AAsVBf+kXu16bLXPsBh/6o/WHlS2IBftGkM2e
CnJK9LixmM1+ExXnP8fuf/1ofvcXwIQLqoMhGymg3O4aZgV3D5ZsSg+aiQr/Vi75
2cu4xocUGGriwdI6iW+2T3q45iLUzl6gLTbFy06az1Wl6qPhtpWk4WZUaLQ6Mbye
8ufxmBldEMNTtVijD4vUgPDuvdb/lQcNrO2RXXcOghEjA72rL0xgaPhjIO+mpn2D
4yQ5o9Uk6LZVa65j9nP1/m4+1+uA2fc9QUgf2688UvUQ9aRp5KA0LkDfGbmNlF0S
bfYGrsNXsZgT8h0q59VRFq2Q4NXseXSjV+fnahoN3/thgJ30CT9crUr9pj6nEoUj
5Xaaf5YuEbSPVtwVECCTyJX804g2dmj9AJnqG/LOGGvxm4LPb11Fxq83O21XIhBp
kmk4ng2UDgUEIOMY1u3vUJkr7tT8f68eFSLFJCxTA+Zj5DtttVV+FRjD+6T8mOH2
9I9XrGa1dvK1nzb+M3VgPjXFkb73oJqilObdfH8WZYwyO0oBy9g+Djax67dvcluG
w3krjDqA9JSfMLePlUwjqirMOkLllDxyeiTZGdE7f0eIXgGI6y/UL1cTgqEvAzVx
6m0VO4eqE0jCYG7zN9fzzwFubsTd5YpBiCyOenFXf4pHjrkje9QTWkLGgfi6G78A
o9nCC/aWTiQVi7DX0+pZdvfTQYV5dxsf72BRB4jHFWlue0mQsB3cebEUtwhgFzJP
DbA+9rGfQk2jjG+fvFPxz0ef9D1b9q/J8cSOYoYP8pu0AjghSxLqAFiWjYwwqNpd
yT/k6Yh0jRCdayChdeg9tVf6S75RBuiLOau4n7Ghetu2mXdfwwOGNcUlOjU7tYB4
y54JchHsgYu2p8UMF41X8xOChcMnwktSeImtrpyWQ+WICcfkcg7naSUz7fb+wQp+
kJG0/9+Ks0snHdJpFuveSqeISOnYoD38K6Knq7/rBK5+0J7srU+J1ceftcaxOix2
SQXcTx8xjXevx52jTR/i0xdm16Iu6rRSaB2js8fm7kpVuj9SuvZJwIDVBDD/uqYO
`protect END_PROTECTED
