`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L8V8hS9hpXP5hr0udZDOeS9ANBBQgRCkU7le4JLxkCq9+BHihNwSsTveDUzDyc8B
iCVlq0dAI4bTyhDcf7N1UwUDerK19175lCCxv/lAddGFHm5GweBuW8e74Lu8fufB
xihIXMSEMj8Xh5zZ1J2+KwrbzvEFd/g/nQllwz7F/BDYVm4/vVIp46e3qQD+uk4W
WnFRjf/7xgMirAZfhVlZaF0MtQ6ymlqj4mJavog9WZQA6/HXfvdPjUg7U8m77qbr
UJ6qHpCauphzFdF/zK+2cFJskftmGqiCtYz+IvchUj0bL8P0g2fmm1csqcXfvp+J
oUulGwQMmYw6dCFVJwoaVTBAOwApEVKHIKSfBL9FAIIy+RcaGptEloukTJyyj+Ze
NLsq/TQqrSvEdtqrrdFdtl5HWiP5+0yE67ZkSsbB8Uu7LvNAEtr1SMnv9VotenKU
EBVGHZ6ClyFWkxG84icbN93Ffd+Cw7iuOoqi4kczcdXZo7Oegu+f1aTTU0K2lHNs
YKHipx0+683bOGJXFSl+4JBfx2uVCmRxQ7Jrv41JS2MoH++0LZKUPfqMVbnU7I4t
IUEX3aLK8vQiPuj83b/lXTKe6dQjyLooHPHRCh0M3LQgN2PRJhFY9JRmTfU36E4I
fPmk3oxqzfmi7D5Utqe55AJUDueHDRqkQFleY7PaYmzUH3o5UQoSjuAO98hbzaej
MrBdoF9IOlpicrWBqykvB3cIPGm/wD514o5TILwdAQ1QbkyOFnMfjK7OeA7p40P6
ozNWsyqI6Jx9YW/B7UJjfgdHN6tXOL/j29yJTnw6bX8GooJTlcyuebUwMGvA4eZN
OtG+dwQOlDchN9LlHjVdsE7ydqZpAel2oZe4dH5U8F2orq9Utv+/anovUNwOKU/E
0Zrc/Jy2aF59PdGd3Z0GDevqBaSgLrEj1r+p7NyOWe5Hn0GwftWvmNgcHCRoA83U
`protect END_PROTECTED
