`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KAsb35lxhO+H8pnJvVD73HoVmUWPs7kjiSY6+gGzwJiyLIkfNX8hPSDB59O+yB7U
MRi+jV9AFeKah+kxGBmYWPOheGJPeOc9nUF4Mosti0SXvwbcTd+BjhO3R0YMIjSZ
g79aZYcDKYtwIhGRsyuAnz0aPsIQJV2dJNCLtWnFJEo+LekxGBoQ93fT3zU56rf7
VT8xDILDvYI6/pUozx3lu9EFFUsChu9vkQZJHhBAL+bCcsvy7aOYaVYwmgsrSOCK
AfV7eUKDqZUPixkQX5+3A9tyN3T2XSLRBHMx88xZ1Dakmk9fZcW+FJnqicxXZVsO
0sOKcE1+Bb+16o/TB6iJOZ630RbCFhei1n41clQLsktOzK4Xn6Hnh8Azf/GZRxNS
U04jfLk6yD6lODAplj2BHEcUn6Nn24D2ezTun1ljA2JqofEwN3wAhSyKIUFO90X2
j2UmOslQLx/9uwAe3PIRiV32fxoj1ZqJ6CuYM3TAg384G+1j6GWZSi39skHLzjpR
DJGPJZ5TctlKxDmWPnqnUNAm4g/6e4ohihAo/ZPa6HLXVcd2Tvnli1PcwD3vG86Q
Y/ougRkRMUbV/usKhiGm6UpUOOANA1W7t/euZ9J/01CeSQSgWsCQueohV1OB9QaU
4nQmeGCSovzDTN7hQwU5aocJ2tz6OqZUsqmnAtW7E5a4rK9lH+geNjW/GJreuwdZ
fPtJcpvo4EZn5TbMgpPSGkLdGD6Gubs5C1EOzD7z9jHO5zXMw4xQTAe3FpyrBO4y
Z1Tvb5r6xyI6VxkQGGP3Zfw90J8TVQPy4+Y4/fFXn4BNQQzAZUzcrVmVT19mORGG
zjPmWHF6HoB7rtfP9+NVWzEseykw2a4m3BqMXz3CMx5MG93IVlHkCzWres8tel3D
5sNElfZdAw+4UkjRakt20LRLZNGP/KZDLtF56vmY6W68LuL01ZGi0Jm/xz48M0Vl
zkwM6HiT8MWd6nNnQQtUHZH4VvoV+8WJcvWZGmvZam7vwaVY7OSpGwoW/0K101c/
BPL2N9lo/o69Ud0oAunTsCQ+GyjAz20gfnYxA1gGkfrBTfC7YaB3yt8eutvuT0gf
hQuHQCeK8na3xG63fbWY+Kv/lVsk98Ao4loDoJ/kk5l13TU3GA+PqhwgXgsSh/GR
YMvSzaF2ra+7cN292Gev9/rusbFRxueOyspuh1G5/WSvLi56lwwORxq789YhkeaT
3HWwwDTZbxH2YI96003B+oWBT3vaujJMp9222t77w4HYtZ3qCqr2VVYynlbPw51h
idceNttjzNg+PdAEO6t2NvjZ7EYuoaIMSLK6psiNdsDuZvSViu4Hy9kxpdPkuOBb
lyAWMyq7ThquHDXch0ThfXUmZVSGsqVRuvL7k3jfhb/9UKJFNiqskwToAbiD/4c6
cGhe9ll4hd8wpy8ocIAduArvHCvmGd9S03BYdE/ynPn2gIn33oP74gAkKxMDk46/
DI2NAegqlE3xjH6VyJcrufK/5/9pAXssELzRcVZt9fsuLcGUOxDOIQ/dDDnQWlWv
n5kqg7iWpb3kOtaSBHoOXw6WoD+L/sCutGvOLcPxR4/cH1NmIb5EffqsobVN0xLq
gc8MBvjYVbaXntOpWOzF93W8czNN4x5yhHEa4MCO4wAo78de1kb+mhfr7jlI/8VV
urna8cnydho9Z3fKRBnzw2oTmieL5z4+Bkyryk7VpOgCGrzJo6sWiM0fXvDHnnOh
Jmsv10Lx9ce5u2UYbbKFKDKnrQwLJ186Uy4HjfMKGdeXNi1tIP/aGF0GP1oWdHdM
AFqQRnbGZgIKh775lSwzBYw1E/uMVQUa0iBWP6WpVXseuG60AQE2qOjJuFJk4MEP
2xTFmaMoVi+6eUbTkJep8AACyqrUuMEdQdKVqPllmYmVoyazaa2pk2ZBgmw8lhBN
h+BblhR8T+nN2YCR4ird4i2Q9y0bHFeAFTJbquIQuCS9cpxqJRb6HuBrbDMhMEVi
pozZa1jkvuTO3Hgq5fSFd9Sx2JgttwZP49/aEQ3MK/4mLcMAtgQo6hsSdlixRNlV
cKZm6mW4D2xMo0eDbd2HZ6dWr2YzevkGDdSseZXCrqxEjhR0qN1vlluyMflsc4P3
jngqu4oqYs4U7W8Z2f/7uDeAC52UoSgBpbeOIxCEgAiNC1n7WBTiWWIbN0p0fVZ4
Wzc94uOGZNXgfEfVjdhjF6lpbWH1tVu0Gg33Ut/FiVs=
`protect END_PROTECTED
