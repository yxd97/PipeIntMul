`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqg+5YIrkpfh5mEQpQVPosMlz491zdSYOZC7zBKZqJlOeT8XTf1NHATm7pELGj+C
nna0nzEXzl+LUFwL3vdOXa17ZPZGKx6dO7Om8LtZ3Zeg6J4wZQ+6blcJAeLjWIX+
6Xua+2SyhN8Y6E/yJF1/i+rIzhjgr5Eis1LoSxyG1OgaPLHF31T8sxuk8YMW43Tl
2cjr75X6emLOCk80nIiwTss1wGTnRAHAHnt7g9rlBr+wmCLm/Bf3DY+njKLiSXBY
sJxkseDZ3lLITc97mHJLr8d4YzRlbrVdmJbIdNFRn7N/BM5Aw53jsQdlTHKwoZmh
jxhzBmJjBSSwQi8sYAn8McaQ4WLhKcjfHVjbita+2By5mLW38lvQpSoiRbIp1gZs
TpzSbZvtIUj1rh7eCaN6/i+RoCm6rabXHidrgHZeQgcRvGwulfMDEAAonVERdFwg
O+JmCFA41ImTgR2df8SxqyyAsGxIqyvFRF2Lxe3W8qHDCsL75zTbPhSeFRkcdloD
pNJ6dEEkqA2B7ZJe8XNSV1goHcgmDojSEDCfmCDbs5ztXy7Pt6MYPL+INRmU6SI7
PhtUELova6AttJU4xrIbuLxkMhCYorBsgwmuddD5IO9ZTv510ezFl8FggbYAe4u5
`protect END_PROTECTED
