`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MxDQYMa86RsiS9Qkv8AmDyLh6pt3kCxvi46KRoaZDetWRlILdpKQrsE1WjPOYxYH
p960A4DZSj6OXrGxqzxQWBL+0XSlg/4TkKpZEtMlTNffAUxxes5irB4+e59re89T
lhJiTFtIAr62/YVUPbHkhoshGgOeKVMDMXF5oFl+zeqyCP7pfW+hhYzsnb0Z2W4Y
CmnqD+BIpfRD/x9BuHsuSHT73d6fdPU2G6X5Zy5ZujagMYnPyOVWiuAgLDDqkSCR
`protect END_PROTECTED
