`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SH/g0kPoD7PVblYPa1ExOq5LfADi7HBsOtzjWzsh7CojBI2qvXbzYppH0valhyLu
gtA5swk5SprvdtbZWGEFoTljkYw5PVumb2dgaYgFsIWNvgm3ehvF4dgEgu7IDFeG
lAWr7Mz2WWUaGXnBjl6HgryyCiUWyJ2gkmg/YLLzSrkAQNP5RLIaMs1wxIKfy7ie
tIdpEU4oLRYdCDAWZLgcryQkQZvZsgCfZENN7nC41zCqVW4fjwXjTrCEhHakr5UO
Oh6xDVFXLAtLxAFgAnhapWgQzj5G/xXlhE1+mUdmAkIDMsMCrJXRFj37zZuBcdX/
v4JgvRNb1tolFhXVjK4Mzc/SKQOB67t4m0cid883dgSmGlhI9yxGl817009ksgT3
oHy3DDsx54bwT1E4iB20pkZjdEglKuNwK7CTahe/spq9xP6fUJZsHz31shpQ6caj
RVEo1gUS7os1D8qmNwsj6ypfENshPYPA0zpIkIE5SQZARB/NQGenMkUmRvAwYSwc
l/+yfWiOO+fmFrchdabZZ4jtJyWME8PUzfwmw8smlgS9HyaoOWtZM0NxQR1+FtjT
reVD39KYX2aldygQHNHV/hB/89cBE5z/JSpYLS2X7h0PD6Q2l40Q0h0lXKPRHshu
PaycwDxE1wD87sbF5eufkCUBOfZp8WAd2orEASMxoyw=
`protect END_PROTECTED
