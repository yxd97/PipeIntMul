`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2rTGzE8YqvxrNkzXYUkB4Hcc4ZyEULR8ko8finVdUA1k0x5zlBQZDNwb2La4XQ+
yUmy21rHO2W9MGCqWvw0Vj2jm/itohQPfybZsUCN3dBO3XlJ+7god3/GxsKPY0St
S/FXFpmrKON5RSM6p224qxCSmGjdXVH8LiogkGzMOSniCxIUZhXdCn5ZYyUzjg2J
6HFElE7xplAaTk76pRi6mKbBTuW4cB7WDFuXt36dfagRP79m3YogbSILezrB+xg9
OG5kJU1HG6Nao1A10XVXJIy7H1I87pUxpxFGmTmG2+XZOTckd8oIvjXQ/iJ6HIiP
doKgctMJFHxe4YIXP5ki3ib0L+ME7xoac3Qwxbknh1htCw+wf2km0dKvz2TNgSnA
QpCAaUFsfQ/taoGoZ/4xYSy6C93u0bbYaq7YzWjpf54=
`protect END_PROTECTED
