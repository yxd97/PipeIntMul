`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S9jkREqiB7zXHIzhBjKvRMEbAKGqpAZeQdkDvFwuYLGbGoHv97dilnx57Z6su20X
Hqy/Fu5WH7DqNxVOEj2B9NIKaQcjgeqj+mr305V193T+1/onp2jcckjU2EJdsLLl
ngA5GIlMwA8yNGEu/Mbn1hkS2vfKIQUXNdP4LNcurHpODVO3MiguK6F8Goo4//u9
FAbXrKfr+ia+YLF4iHwCYWkDWjDPs2kNSXGKR2K2w/Kr0IuCio+CYgKBGygA+DTr
eb8mRKe90Yj+gDamtrWlu/OJyMaxmHRu2HxdB2HQI/CEpqk6sQGfB9fPb9BiTYGh
4B/LVTG0FiAw4jbnr5UgUXTC1vZLiZ/WhD90KmgGfSABe5d9zSDhoY610vJXIAe3
l3khIc+BdsM4RREGB4OlyVhvhAhAjxJI5K1jnshjgRLtyqTa2zSWY/EjJbu1WsM2
365tc246bX7PmgFj2IZ3cecGij2cq1AeO/EBVhoVlrwjHDZoT8qTPeWGpjiLZmzG
sI+YkxNU5Fw02KfLkNO/xdE0sd4d6t9memppGPsXlfbUXjO0ncJ7xugZ+hmfdzkv
UZUiUHoRDRJi4ZIhl+FQeMiqvyFLX2A7oBimjWx5lMG5R+pARWcD5cE7benshth4
WJMSCgWdXc7IaOLL6p3RI34E+Kn2B343+iZvcpuMGNH/EYdSsD3yfkarq0ylrNDC
H9lc/oNgm/EoMkOdbvKaLBkogyb++NR09O7wYlv9rWW26apERPj4jXU/Njlwv19s
kW/kFJtvv2jDoH/27nC13XaEoL6Kh+8TEvvrN2OrDCbDxCNreNdq4OFSNTvQeaGv
ocTkoRJFCDB2AVirRDU1Voheu17qrmi1KzIT7g0TRpJoAqPT+2tLUi36TSdt19g6
Tl078o2vE4BmAXALVI+Gbr9TLxO6XDT0nWt3vRpV12FoddSellK+92ZozBv6CJCX
WZF52EsI9F0JHhWbfFHO6PVvFD7Vyo2pYiWiBYnzh+Nxix9XCo54PDe4pfKgXVKt
SvIthdmUjS+nyr89zvF4SzZwY9VCRlPlACxb/XqawTmhv6OwaT/fvML5BrGL3gdR
s0YXhjRDUT1EcuNP2IqrBGLBYT6OKX9taZnbrx/fF1bwfXSQ/zTusqVCVfPppWm+
`protect END_PROTECTED
