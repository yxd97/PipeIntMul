`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmeDC3mRsgg5zBpjx2VJuuniDxyUP4kmGujhZ0R0kk73nPJi7DClMyjF6XmdcE7K
4UkGgvyJmm9LRn999rDpYFPRrfNhJBw5B7MZpz0dNF761z8fbg4oEZbJC00PCryY
HM4aEsnCUVs99mknZZpotKu9ymbQ97iagUVul5DLsmT1rK6+wQfZxhjWUDFFTCDl
lK1O1s7qu2XI8K8UpQjNoHXckIGpeX0IQ7U4kAjq3ECvqRbuIsBya0+y7IDv0dYl
pKbOWoi8M29ZgyFaJ291hX/pEEYH3lWwEfl/JCcV+6qS1YnWJmzD/akV9i9dtXnr
r4Tf0FEmmqNSFrmJW3XQAQ6ZkRAPZESuKsb/bT8eHP8dG7QZ/jR8ysuZtyQjiQ+A
rXtDjZoCHo8a59eXmjkDBg==
`protect END_PROTECTED
