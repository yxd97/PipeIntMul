`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eJn7KcKw8Y6oWx2yWXFrae1FqDfL0o0xr/anjB81U0pNcixvnP1WjMET/L3c5Qs5
We/4Ss/lkSWYSGkMPuoG1vQjl91jn+Tzjh23g3xrIvCF+RLUskSYklbiZ4qF9k9f
N4dpvL0OkvPBnFNaWTSQ0JlNQaIH1WKrqsHoBSQsgaFi5EBky6hSEWJr82DRMWzT
4k6nIOqTf2sDXq9APDF6EUYSO102JPlw8IbONXdmaeymb3kyWhqFn7sONgJDvDx5
AVNZF7u+nLeaSl0OA9sW7ZuD+dtHCJoq9E6I2Yuh6oZls6bWjvOCWcVcw4FIpzRq
X7JRTDHQrPHeMS3/8AeW2nIiqUQ3ARrizPfSY1HBWeaTgeKL3GPTzz40dR7DgHC6
dTMyaKzfuOjI5JoLN4mbMogV0eZq92jZtsh94G55RTxMtaowq973IHg5o4rq7uo1
0EmiDUu8G62s715IKq+aN+RjkYqiuRDhgw6LBAJMlTyuLeFk8+OLQTqZ27gSu1Xi
`protect END_PROTECTED
