`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
49Z5j3TBqqC+2NolzGvBkxKdxrmeXnmvUWC+/zmAYvJYVVgvqa2TfHRWWRF2iQbS
YcDL88Pgc1Rd7XdMwweze5ekGZloCjtLaiFDrX7q0wY95MiRDcvqKWOWjEYaWG5y
Q4YkwqOueb/6ymB44u3Cn0XXPlI4x7TUSRBCbVCqGeo/qxPK0kBLmECZSaGYT7wO
k9YQRXcfPPNr7/+LIcJ1+Mo33HovsYFmJHYFTYmwP4SthbzVCyV0tfJh7PTmrcCh
aLnkVofisQ0/G+MhEnIJMT6syLzTsuAJgnSl/Bf+z9MIMCLCG7z8ZYmvl0Coyuht
vVVX8Cs4r/4agR0l1+bL7OVfrY1OgL5HiLaXCAqeK4/Qg3nuI6cCl0GSCU4Ii4Mb
/VZMm6Cmj4RVMqJKeq7ANYKoVW2TAC9apLIGlssFFQS4FZsyUNINmhPp/hwVojs+
2vW86NNSoIuXvI5fOK2gFcsJ0vjf6JSP3UOLhUbmk0bmVjNa/jfdaIel5kWYCSV/
`protect END_PROTECTED
