`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+GkgHIfw5WrWBgNz7PsGhFwuqoRs8w/9POQ35KienSstetOfv93zd+/KHLc5tDM
7ud42NeH/bLoeZiufxSshqWY/wwL1uHjfmI9lFvvfXLSopRLwXL+Y+KisXTVHGyn
4vEK5svYws1aHr3/UB9n1iVRzOO0WqxZXtl9LS3VnuqXVc1UmlvInzVRi5LpadWw
I5AlOtHqAcUrr9xG6lEq+2N1rRfm25vzmhLAqyE5zI1Bh2iOlLUFZSvh4/NXN2Eb
lJY7bvh8e7D/+1Yp1kyD9bINGE66Q9Czf6Rx/WWVzWPyLiB+WQProEc7MSJ0jskg
QT+h27EBTjSaVXbF81yDCNA8b23rL/sKg2E9IXLrEIHMQysZAkiKLz7/klMLFQK6
s8jyMIkJdrXEg8gFsnDrRibatU4WtEB8+Qf20QCaMvLZnyKA0SuVwEdblq6CqNBx
G/CeEQCJs0Ql7Jbh9ISa8nJUPvS04JAVCig3jDh7SD3pg+SOtXBT6dahifiCu2wu
`protect END_PROTECTED
