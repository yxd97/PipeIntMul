`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zrjEWpyiuxxY8+Ec/c87lA9RG3bZrRbXjXScljUT1wfYu0tE2cT3ajzjUGLAAB3R
ye0H2YL5P3jqR6kTBMm9GHxBlDiA05F6efMECwwKHoZQEhiUqQuJ//hd4qus+ua6
nwOK8UAxyiyt/awVkeWOFbW4psHIHwezkHjuG2+HWv6ltRS+zJpsZAfbQSj1Pezv
8iQmMelhDBbB2ATBqF7wWNfJ5M6Wq5boTOrI7ZFGGgIfsxETAcg1oEHB+yZDoIQn
Fvh83uEzG9SEbf64mVSx/8i5nL+qXeZUj/6yN5lnojPUiXX1+doTXKkRvIwfG/LD
UjcPsqdc2+ZntJMJBAOeyszoDZedFoF8cRt2L60bME44xflUBMd7d/SjXGy8EhGV
VXSGK6S8hlf5BNGD8vqkYTjDLngOYn6fnBo/5zDB1mwMicOzh/fjSMY69Bhowx/a
`protect END_PROTECTED
