`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYvmc/oXJyrD7Bq45kTcV9i0xNyt34VHfbg6O6L3JKQXT1nVYu/lLqD6A8NUi9TS
ndAH+YrS2LjD8Zf7Rdqc3tfkmkeYhcY2bJP4ewhLBplERDQi36iUcrrZ1ELgvCdN
64qb3g9jgHjKftPCcYT9UCkj3F97yrd+z7hgYCx3xIYYAsJHBB3BfZSGtO/NRuSq
dD3Da4a+nEomhTXAU5icg1YwVnfY1xbOHuRvNqCOsYdoO70dw4Ag9mW2v5gVZMI1
0MTZq9JOLGCO8hQw3fO4vYKXe8HMQes5fsHIpaYVzJtesg5urq9qgx0BgJTa8dMU
U6GofeGTHjCPuhuJv/qBbFWRYZ2Ci9aFP5hkDpbFmZkZ+tCgBJZSRR3BsR10FA6+
BAfz0fRQ4QDyTEWQFbTEE5wiwTsbWr47g/rz3sS3JU0WpiJLJ40tNg/rxqqIFOAb
ra2HRVgXWPgg2poKN2VtqgX4KGh8O+A9ekbUUcjb2PjK+gJ2jxpV1Mvpv9FM7yKB
/xTv0NiIlHBZYQkE4Vntyi0j67htywW+pKnTMms8rXYSjX1fRYdacxErmcthqHCy
yyrIQECGxidLL/PVJHt8vP9acxCDsU6owU69wSuHLQ3f5mtfRZ6CIjd++kC78Nti
VFx+CX4TaoIxkbbfmBjpNMGm3NsVZjcfp0FArznsaoV3JzhbRHJcz9SLX56C8H4S
nDZz7n9XilloR3T+4KO8Tw==
`protect END_PROTECTED
