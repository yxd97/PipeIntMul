`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xO1Z/koVTFUgmq9OgyzJiXmnKJogj/BEq6xPskO5ad0xu5pEWFjVexPr1QghkFlQ
Sv17KKly77jTbERMJ/x11MbkG4W4yxE0gCQ+iYMakjSkzrQGtnVCDyHvFhUa3oHl
MqA3ZpqBrzOXPLbeUUJAFtw0V/7CYOoJzSspovdXAgXHqQ79EfrL/1F8tNT/0HsR
eHSRrBPalYJa/OSXfFnG75qN+feRu9Yjqh/oqqlIiJNtwSPC7Aq3F0TVT2he6axM
YBxDi5BJDIn4KmJF3Xqb6Oxa4cFVx/91d+Z+iMndh2HRi05PedF7LAP8kqgNsp65
bYT+to7L7WGqTW2yhkv9xnYTmy4qLMk8m49BvZ+iQs9lcFkugUBhNbl9IoxpTUUk
fDr3rrAFU0UK5Kt9XkeXSVL7Km3HZnQuAvaOicFSxPUuNcVUdUxKBY1RHkq9WC/A
fySXaX0hi+D7CUWytjXHkgZFn2NYMXrZbexcNTkopfaRL93MkVyUXoyX1aPv7riN
31fQGM3OvsLo5yDMxJd/9uiUL2x7zOZfVTFDDbBko5xRg85vyz60hFLL7q64b+uI
PklHRBtPCuWcBg4t5nttIS4idybgrHt1felbOl6vKaDjL3h6Sdser+fxuLeT8aiX
6u0v6Cn3DhZz2PpJp9X7r7f9VDG3Wcc1PWYuAXVvz6vvJqyly3aq2lqurZCBrfY7
`protect END_PROTECTED
