`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPKVlJrwENe9l5AXww5ko89YnG3WUW+QSVyOiWu7wvfT+icHFo8OKTrP3of7vNo1
YlGEzCEm6XbXHm7qK9VzKyGWPr53dJMAPxi+uAvuqVep/EQl2UtwdCofa0TYcAMy
iN+Z/8VdbaPsSInxIg9d5hbtz9rdiCOx2USMCrRfqn1bYTDCNxMT5OeAS8/a1txu
In1rwJGG4UMQ2m+cyx8J0KabCygRT+5hjRLIuVzbCGTkj6HueXeNLIHp16hN3gFe
chJ+4QzjaseLusBCXHZbxduoxq+jRUSFXfyTDLe8phboXvBw4IDICPAaRrgJDhuJ
qQgqXDDnfcB95fngFRLm8C1+grb5xE/QdsRbTSPxS+QFSqgvqdMl2GXITbANLtOz
0YKF/P0jQec0Zd0MLB9qcM6ksBDwj8iCbI3SV0Do23W27liznab2uoENEJME5Ecl
LbfJ8xqHlK9hg/O/e7ExCWoU5kXFwKu+jbLFj8fDDKFa4FkaKWwUOaeymI9VIYDg
bjV8ZH1Q/rqnr/iDaxr+1aKgpu6NhP13luU+NiNlg96/KYNPokY/joqcecDE9YoH
`protect END_PROTECTED
