`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDR6aXKxI8agAD3hI7BjFWXwptMO4k1GQhuLe0NoCao5Q4Pfn7NqHk8e0It5cRcL
ACuReDMZVNkr2EET6Rkulhi26KecM4QEgsrTlqOppLeMR5w3dzcOPd2BFHsmOrTT
xvXC9mA00rkPMSAABuUIPkRxffDku2IIeEkhoDYAawRcHrZyhkLBYotSVz8mjQIK
cY8n7WsTFREu7udhwnsREOqsy6Fag/avteFlRu1MCO5VWHuLXIG9DQW+/9K4HtrL
oDca7GTW8Ro4CGJqSoxGJSlrSJ9Nz+cYrTVKpTuiLrn0MB1l88XG/QGyTzoL2NSx
Fgi6w8RFyCjsGj09VVWzn87KhOl8vQoUJ7EnrL/hvFhRLa/zdJEx+OBiMOA6Lshf
Sa4/UELE4kqeI1eFX1AsGWSrU+KLz8QXEYqDDJhvbz6IVSqk2GOYZiEmp3VzYA92
NYbwk8Bs3WG+69jgmxO/t1GwqPJG2jTx9qkEmsNuhjlvApNpahTC5y1/Gfz43KpY
quFNHg+oexBcB0Enf02YPROJuIbY08BAc5xSronDNcZL8JsL8leTzyAscWqXMKsI
o4c/MHwDsF9mwDlRJZV1lGVy8/feffjq2Zkh3cSMgPzUMDog/EIroqGjgpm1QeoI
OUwdK19S2el2JBTW2/unty1rDkHjigpaclTh+S7VUaXsJ9d3Bj57/IsW5+K6NCM+
ispBdtbjt3x+uCPLykBLwt8+Wi4xKQd41kidb/nWb+6TR4DN8TVKFw/qwu1bwjHp
KFEkUnSMc5Hzsj2NLPZp0gSgVVQWoJUcij7phZ3K82YqrDxMvTFMqbpFC0/MjDIh
HyS/yCf41ScpyKBQQ1RoXA==
`protect END_PROTECTED
