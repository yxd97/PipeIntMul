`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
amifuogQDhILm7Op3rcXsKR3c2mATbR/rIZK2kM8sAyGqgp/Qjfv0Mpn+Nv+wvaB
kSQ45E6BhYYen2f1CtoMI/rlFjQFyw8V+QB4UQfhPGjmb2T5FQLHOkgOwNnp3Clu
QmfyP3WpDI5Ir/HUDVNI25OV+JN9nfEdOZhgPs1rj64GdOPMkK94KiYrj+GkNSFe
kBuWlvvibWuz0GWwAVhUazAGSJRvCuj9rmqCW2rjz8XcSCBG8NHygT4OEu3/6UhO
hiysrGzQPteJvcnea0VyuQg+Z8LK+77BCeQYs4MC/OF7aAsgHGYZyiVeBlHUH9WO
ZecZnyL2Y/ITFKvPilOgKNBHCS51JjNG1bjDtz60xEpZKiCrLIvtwb56NcJzoA4M
`protect END_PROTECTED
