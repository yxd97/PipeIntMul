`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tTDALhep0bYx5Biopabz+/C0xuv4LGWJWp95HmpTHAVS/zCK93oG/yey/nHCs9jx
MJ4KcBk3kbY+HzmrEH6lD/o4t1Mi9uqTYvxqMzanJlE157r2/7BCq1VGeXcvvneq
EuaeIlrRRR4BAVbjSaPi4VM/qvIqtJNStplhX+uWYmKcD8WJWqAs7aAVzO8jAdS5
8IubEQmE5Dr3I+ciW6Bk9r67Eh8/lrza4jPKar9r2srB3nmNK0gDr81fLUOp1d83
ULO0oyy8FYDvUkve+ajKR9WkHFUUw8QjsqKKHv0msBrZT0hrH4gve9JawJknjt6x
r9NzavJY6a9E5LkZVNNKDwg7314lsTQxi9ZmmE2ZTQo9PFEf/M++g2Thn5ccd0My
HdK3GiacIrLv1f60eZaOSq4XiTPOESTgJUkQ2Qe62qSwGkgoSfwhzzJgz6NTp5AP
QvnNza3P8z8Ju59u1iUl722+OZM7SG2BMIMDqhv4Mrq3MMeFrUf4W8+zogCXqzTr
3Ofvyjjdmzh3si7alA4sl33RvizytIv4hHDB8NVNVIk4mWgIPgPaAtpf1MzzBSGp
rAjuZ2lJWL1zBGNkCNvtltWE5Eb7dK6MrPrUYGrj45ZlaAUxYvoEEcWaJrwldtfe
aAcf8+JZ+Xk7hrgdnNOzYvmCmVOgcXUIgKl+R+pi9Tq36VY68t6bJkRWwNiq9gnR
Jha9e7au55zgf8E0jjTxu3umbrGY6IyBkvCZrgciyGEp3q3YaaZLSG58KadzpYYT
cTD3GPe1E56U12ds/pXlSAqV6vh7ysvG0zVGb3b3idJI14HWFfug3CzF3j9c67oL
d88XgjlAZqO4cJ7vXh4lGnuImA/qsvexpup1xkGakY6fScjok1vOuGoDorE9D2Do
JHmt2li/U5tu3Q6Pd5i6bCuDzDny7cs9bjamzjJBt4fcagHrVXyNIbxP1efeDUUI
dSdcIFF0BfSmpPXTYiCF9vl/axTqE8sC1pJy9x1fkXxutUZZggvN/H+yqM7cpoCS
EoW3L2zcdkugZx3Kj4ae0IqxnfdjTZsPv8STVO+WlzXBJUPmYH6UUY2HRVxS3CLH
YMcQLmJNLGZ9SgWaTiU7xbF5QPoI6BgJzHVn1tHYTBcKeD0y/LWrIVaGYv3o3Qpt
BiBKpNNUIs+Hl3ybCGI8CxPesNqwPjS1byXLWoKpxeRSHXF8OLR9TyvbewqYyP+n
eIM3zycvsMMLuG4ftj1+4vcatkQqJ1ZbLkwvvuDy34PChJ6asTVtKEiEIoL/zlY3
uXT5Az8m51uzJ9b6vjWCU3BM3pVlJqwx1Lc76Fv8Q1xD+wAUM8Zi30iNhPcVe3FV
V5doIXan2ohWQc8p/WZBFI6Gt/jH85mX4f4luefuL5JI73qe3fHNRw7oL4SDh2sT
yl+7soLQcSun08mqGsrkH2B7l3vt2lg5AZIEl96qFtYPbE23yw58T1tpiIRCbG14
XRzSJSPnBtNBErDg/7rJGCist+XkeNoDvrlJntroWJ/ONGWRXpre4YrhptL+dYED
VF7Omg/De0E8ZbZUCZYN7IcBcRCzF4ZLFd3GsgLShvTVybFDbps23Z3F6p2JJ4gB
8JTsCSRLJJi9q/Z107LnL60w99kvciz/Vwh+mcIB5ndDCcVEmsijfkGdC87VBG0Y
giTmkDjyrRnUmpWLkq8/bIr6F4/clfqlcI0434rgGcH2Df2l781X3o0VQy0rhAzO
+7ncDDDnrFk2shQ7CtsNheljtl86PQsDeSuLAB9JpU9frmkijtRXpVnczw+pX1OR
jFg8fjUi0Fcd4/wGXG+pn4VeUOYqFCehIH2qLniZjOh25u6ZBKkwNWINYPJhxndJ
bBegS5GxlfOibFx1SIpEIqkxJtTg6q1STWDV4gf+6pQGgHJ8SF7iQmkwUcLexYbq
Yap7RbEHMxYU/xphPc4Bx7J4HYtRLlrcoCEDQHw9a9daEg6dbdNnLheiT2DCPGyX
wG+s4Xm3WgvyzJJF0mU8sTFVMg/Ib5JSWbqj/GDhZNj/84nnKP9WTiyLhJN9a1CO
PZLW1eVlh3qMhyk/3lPMOrg/lkJiPr4y61fb5ESSFyp57vvZ3LuRKbMVNhE7fj24
NkE6ZyV8VeLveOVE1A7SvAgEZDeYFhRPheMZFbPl4+0Hs4EMXBHYIq5VRINM0LVA
Zug8HtRQKIB/WNViLl3yj92FFPUcpfXuTJzRv66odKfHBVZFTijwWr6NMH4vJvhu
VQtunt0Cul2uRTxwVilj11j5iPskrFiTKphMnNcvj07GvVM2kxm2KAZ9HS0o8HkJ
lz/UPJes6BczvezmYsw6ELcQ3IWu9q8oqz4Zz6MnTI/WyTgBlSSkzjO+rr49B9y7
aMfAkdBGht5NvSOE35vRKkUK/dCBP6InhBQvcEVloSVMz+yfMfwCb4tb/GTiLpHW
p2nXinZZorR1UHsq+pT3vXBTlIbM+5/0GiofVUql8MxQ4g6ai568TKT6cw302XbV
3MuwSUwAQwqh0XoKLLrdQFiVbIQ+JYYcgu5e2BoZGBQzSmQto+w6x6SdKGZmRmaK
JIx3g6kWDhgfoLcetQ6np8RAr1LbZqcO+Tbrygb7OIN70s31JjbLkxzn+7ky3/Bp
z3Y65ZXzo0nYXYdGhhcOlGZc5ql9X258A0bHL5cIeMkALyxLyL18xe3zwfKR6K21
tueCauDFDiKj/qM1gf51fHrG8W99gsWERtNVO+HW9DJ5bOJy1S603pt/PwJm10v6
EbDYu9x/JyOE3mRzVWf6JtPSkd0Wtq8Z1CUaoo4TvCJe3Uml88eeyeOXwzZ1DvBu
6uR09fKBaoF4FywkiJp9dCACsljYLgM3ortItlcwkcI4rBQrzeK/mVUtnrB+Sk8E
2sU45W/harx0e6vuU4zxZmafF/yE0Na5SuHqEbqg6+CqyOvCu7xd4Xyh10NJ/B0R
ZusfJTHcybhNmMEyzetQcHB+mmQA9xclbHRsZEmx15TqWBIIvysJihATsK6gqBdH
DETYda9+gq5KlaVZS7D2XzfHvhrOQTL0a70MEcZxturZF1xWngBmULkQ8MBQQ/dh
1h/2k7giy37MEo+Q96Nm5Ua1qLE7u+ZfkUxTdcJO+d/5ObEqLAysz642cKg0Nphb
b8mHhJUWt0C5DTTAydsyzRHjJmj84eFZw+km6oDgyCGG65Blrkg7DK7zoSEETebX
dtl+H9VSARaGLrtM96Yaw5ttCC8Yokhl9VRe3wD+bXKMjtDjq5LJy7UKkpNPQVx6
0qzTTqxASfxlvHLdb4UY6O12NGa3Bo40/LIakRe8Z4ZQLP+h0bm64cYg0p/5IkQL
8TB2c2i5es53tYt5a33ci/4pFdGzHWqK6oik/KDIwi6AGfGC/+spYlRCDXz3mSGl
potd7ZSXYVZTmMM+XON4W2gmNGsTj83IJCG1mIRy5QfA2IW1ikKmppkJFVruypsg
xiY15WfphdrMp1L8keit12vtOclfUPyfe8VIch77QtU/KrJnVsAbjSYIkwv+idxa
u86KsAH1/djJ0clHUqNi9B6ZQNbynkMGgnIl6UNTIrZWxf0taUZdD3w0rWAUq05a
WBksL68iJStPQHgLjgTXXxj+1cmZ1nxn8rldbIR139F9PXgJkGJuj0CAlA3czkwe
cMRGCGpXsxIkngpGOTswcadtjL7RjhUcX30/nfXHCC7Fsjqtxmj7wLH2C4AcfSil
0KK5SWigylZm5tDeTTLprRrJinomkHMq/c78JRbpLmIzI7LjPOQ9os4qhecMFErL
ssTUGdcDLx6frfdBedOM8a1oUMtIWk+ZrHNil70oebciuZTk16Bct/RFljtS3no+
c426SJwEa0qH+a8LNGno/z/pXZZebdb2oGh3JAw0Pkxdt5DmKqTiXos7oGFXuM5t
9biw+u6+s2x/3EB847s/DXZUEG8VudvLvHtP3VHumSb4UMoROBZ2E+/gYpdt2ruk
AtefMwElrFNqa3mpXl7JdH7D027Tdz2eNERG2tqwYbJfkCW77T8ufY9DD992X+66
OHlYKA3dsCoy/orZP20pm5IAsaicJppdfp5WolI0kLg+bZbF8/ZL6dODc0F1Aaki
s3tOi+rzwrAlCVLhSqnJbtE0/REDjV31+KfA4Dc2+eWUjDgwB8HkrZwaHglAYFdS
HtwCJKO2VryImfLGDpySWGTV7aGEiQmTrG5XlQVn36EvFsq14Xwf4Ug2TZm1Gg/3
9vJRlEu8eWcx1/803NweFINwFYZWrw4gKXEtGGERmAqXKFldmPmRbW3neIBq2MZX
REhdrQnNXUN+XYqlLnRyPAJIxbvrWkbhSRUDET5Kn2/0Etggq5lipaSU3oVYAJ77
RER9DdK3rvYxLGu9HDCostxjf4PkLxzgfH5rFtyo6PWaoWyEzG5/Y+RpsDSXmTe+
AO0kyiee25lYEMIIvv2gsifFgxYVQ1nM0XT5xIUzqZeqE8+nT5mUjoENhPLA/rJK
JCjcylPY8dbKLUkh0abAfeRvHrYL9o8b9Zm53LQi1riUmWel6fFDh8H68oBS9nZz
n/nEbCHtX0k+0YPP1/XVU92okc5dJzNxuuGwSOeUrTup9DTlw8RnTeW+D+gsNojq
5WHoPC3KSL/E1MvwmpFPXrQeaOuC+RgilTeTcDfM0Y09ykqZen8cC/F6+OJnkMsI
MDdGD8Wtyk727YXxwzZIBbv5LJ+H8gPpyRE+R7HJ/zkxw7pXWUgCDKoHYBUYx5WT
HLQRk69IlgLkfXmxTIswaE3aTdNnnfKPWfFgRTEUvefp/JzBjF8c/FXcRwXotXZk
ZJ9EFzuxlXegIfgbsak45YFk5BWF9BhlLvEI0lHXBzVyIJ7J66ub+pX7I6g3APTi
nQWEmwckC9DyrdsGNZUu4CqhE/qak4oFoL/IAVSR1a2jI/ADfEZA3UPUmb6aeW6D
1P5CqGDqSOh2qL2LVWg3Gi5zjLEcIrOI1jRzJtpT+kG2ORLjBv5D5SBXBi6P5BSi
eyNyWTCrqGCao5Jql8OEH58uYr2FmR3YGyjwFBUT/JlWKo1YKfDlC+sZW5/TkhT9
VI8cRj20w0qgV1E+rNDCX8cWddB8Rx6F4L5nB2sV7ugApyIQfsaskuaVR4dzxJ6c
bCleebGA904AqOp4Z7IRgqHDmRQZCj9RWrspk7wEaul9CIM/JUPHOY+lnmJSlbfy
IxmyNoOO1uajdi6B/Pkm1+lkroAtG38rFRZS4bFAVenBf/LgBsE8BCkow66KRKpn
ZT9CaecTrCwDbMy7kZMTWPPiif4CfAIS5rrJy4A/dcLE+GkUCf3jviTd+HyJo0ib
uDLCnwa469mLV0torcaD+or9DCo8/AaDnhyeAl0SE08DxmFkctnXOdka0LxKTnPx
haelTNuEKJyp6bB8XMgIROIsLBQ/bmnAV4Xg6kjFZ1RZQ06sr/tAYQuHdY5N0q7s
PJMikw8XeuDlF2feusPRnFXh0zcTFOzM6lulezwA9HNpXO+D/vqoG04ylqIcvin9
kfBUsUu9/Sm5YBGfPJleyVTCSy37CMrH0B/R2ljlcK6OxzemwO0gMoIW0jkXmEVc
mTH1bTMvltqNTTMGYL7xKoXDXM6vh5wbW6ZgCi+dsduUh5K6O19eJI/DClyQVD5s
JhWqITkPfyuDwe2bDdHZ4+K4TFC9P8Ld3deeJXFrCEQF7amyv0CZ6Cr6uuVUCLWB
qNqe8CfQwS336dcaVxgMRfYhlondzJkuMOhrI5xv7uva/2aLgG7e48gOLQxZqZKG
AtLufiAUxVsXXBQu2gWhe6CVE1ZcSPGF88JmFSnk7CU2vHvOQF0ni4ZZxsCBkFgz
U9tSYzvDHGCDrqYxLB2kjk4dB2CO1FUm0e1TeyN7byDFz+BhhiaLyCUz3EVf4CRg
sTLhHFVbPSYwjoJBrFhDhPB8m9bvpdNh8/Hzz5JCebkMa1+u0lBFCKiyhibrlZ+n
itEPr7uemFB4j+y1JaccOFqTZhrOCcHjO/qzW8pab5BXTFtmvnfObMoVW0kuoDSy
a/JDJqvtuWvC/kvBlIJr139/UPmsQUTFFVOZul2jQkOfbl2UrgntIzwfXoj/CleD
SUmMOhirpfQrkls6wOoyLBOayIh+8vHGHUpGkOmg/0k0yaddLyDyIuUap1QASqB/
32/BDm+8vyaVsugaNVi9Pcnes7IopJ6JFNFejZ5S6CJ0NJkMIbuiZIcyndHZmzNh
GqFA67dWorfgfjxYGX6CrT9vq5o9PwBtoentOyC4izmeHHXXqp6PRMap11QV8Bc1
YT0UG1Sc5xCZgZfDg19zz0rk/WRhkgVeDKHbBuRU7HYF3OB24x5csJbjtY8yjHRb
IklERhyqTc4bGvbT2VPwPr4d1tC89wlXBl4FDAsjAXzWpfJ9WZuwQHxldxN5iL9O
jrHZFds4FBZuS2sWEnPxfU7dvO534sGhuUqcfmz2yZWo35XGeWWw8ujaGn9+5Bur
1gnZmsTY8MkP1/88yeIGZHD9K+G5afjkRuXQaQRhU1BfMI2HYoId9dQie8WGyqNH
MvUVkKbFwPSJJ5Hfl9mjgaDuaGQ1eun0D9tzQeuP5HsXD638Txzl7qHmJfe8EyO0
P3EAxm9APjHL/lURrbrCLDeMBiibNqeFANr5ChfMYgIY6a9w4DeDJHKdk4VnzpAp
mTkVDuI9YL0KHUxiArTnd4IrTr+Du+M9yvIkXAIAEzDD5QtVGGuetzXU14rFy71k
G5H/xnte1GRKWMi4hWMvYflFdABoI8GXBL5N3sVf0a1s7aKmTedyLtvj2u0+BlTM
iLEWi+IyEdqpZhsfbwVDNHzQCxdePaoBlnb6HEwJHwzhaFPEuhQ8Qh2QM1UKHXyy
b1srMAhPZGArhxF9HlqpNqmh6YKGy+EHDn26FfXW2tk7yEoTQHz/Q4A/wKNCWVnY
oqNMjewxCgIUeoETUT/hnzTT+2FZxjFfuC5sY7qn4wOp8Q3d2NR/btNaTOKuSGjL
LhAc/Btp6PGAaKtlFu7bSPQBtvFyRTnGa8NrWlb02Lsr+dThSItagA4JbCOwPzIm
phM0E0lIKEkKu1G/ZxD9J9dEseu4M2fV6LRYY5sQSbsPV89wwZsPY3WiELQVuPHd
/QOrI4EKOE/pfsHUSPvyk6V7NLl0b0yfIPrNbTZP7VaETA+7t45NPTMi2CWDhbfW
jYlYNvpZ4xIZIay2L467yGrvIZgTqpeTWgbjiyJY3jJKFLpO4LdC6DSq8CYCUiSB
LFXGChWSgb2920Y5phcd+TJzjM79vLIE7tIB8QuipbJi3jDZRthN7bc2vQSzfoGs
0Yw3pVeNpeFfO3oKVVxj0DYmeXOAUg73eT5EbXQ1DayNFa0zvX1nzPQJ9N2wS5cl
2kO7evk2Q4xuvrBoZ2xMHmDxxvMkaqpCeqnk10cFoYeJYpCl0mlrJH7N5vlQXL1Y
uZN83x0A5664xJGn2JMIWdD7FCdohTKE6lIjF2SOsO4XY7r0uNh8geHmLaOd8kTH
rBhgRZZD1xUaiqCRxqyI1enjlG1mkxfVrKWJxLBiWXE3RU0MQ0bineR7PKU3wmec
3PK7VENuw0xsrAA0X73z3zNVuJ4uJvgJIGZkz0nMa2mRKDvAoqrJsWRA52MFyl7q
jhFgLzRk9KTRMu9fbVvHbNeF2ZG5Q4f1iZ/KZ9oKWOH+34DRaqduy4Yi8wucHLNd
/NpWY8Bpw+ivMamoLs4Y2ErYtsIZJ+1BSEc9hyrvTFs0dJaA3SPgxq33zxy18fDM
oYeNxJtBYJf2J1x45YgVSW87Z066CxxHVYrdTxNeWYGZk8xXaP/yFnclb+vqUtpK
E+g92K6BNG2Z2XlwkfpFSC1nD+wzOgjOU2yNpasIWx7ChG56KP0/qSbyWfyY4bK7
In6tMY5BKrIGLvHm9/oOV72wo3a9f2dOWH7ITtsqWFbqkkDIhdFpgY8EugCsgcKz
q4O94O7qm6/xEwgy12wvhNwJlYuQR8B0R7Hg1d9D+J5xBBhsTt4GSOrWdJ6DULBR
6ztnzAr1SCZ8nYK/iRUDXdGa9kzSKaDpskU/Ye7p17f8YFLF1aOdiI0A1QpBOxZA
XJ2Ghd7uofGCHN+Crm/kWukYMITUOwJ/yK0Nm5Efz9Gnh6nonOeAQB9kQv2zNgcK
KSGlXFLgaaVizgzjrEHUQhaJ1OqZRR6qhwdNYQAeg6isGt7mSA2AURLbk1VcMyEH
nBtyhZ1BJZALRvgI5PMCPtlQMGcz1P9ofgoJVuxBDj8mFxAte47nvjvr6jjUXVy9
AET53S3iTtnxCpy7EAchLFxdMN6rihKnVQpuQDAOnsb94J9xNpMYyIjCy6SK/pAJ
Mn20Jh8LWa5rbpRWbcLg2BcSN48/pLTTblx9R+h8m4fcC1b4XooHHHuy26rsR5e0
N6VU4eGxgEe3cHEECniBLgWxkP5MV++p4A/OMdqamLHJTCosAMZiRPpwfNsdSrYX
XEBgbeyWdyQCP9r5LE0iEkckaBT7Vi3geumQf7guflf6Ru2NrDY/Xs6Cq7wQyrqo
5BqnR7AdNVwWInmWD6rjQdx5rU1X6BTSfK/UewQSYzvfxhwIX+z8fnl8C0c8TQPO
mvpsjdT8ez7LIUHpJF06ICv68Q2UIzDwh9Y4URYGrEkeHrdlYjhZmj+I4ae02Wmc
UCH3zelwW1wQwLV7/Gwn9TsnA0l9aEXJefWul0hswIbq5W5i55peYnXF7UBJnnB7
ciwWZQtuPGcAY/HO4E6JMSs15AoGC0KeqL8QSxBvR+os3wgUYcjyJP/UBprP3gnN
HkUNYRWo3dlUnhgJeHPbHbRLIjT4VkooDqA4jLVqCI/7vgykYl3VBYDhktPfYW2i
MidLVEwMtWz//bNgCbUZR3EZSev3DiVOmwvcHlEGsO/Nyk+gDMVZWaQodu6CGjqG
DSgqJmB9xdWyxS+V/yteRjKSFMLtuQByp6YxuHHRpvPPda68Oa+qMnQB2nICMBnP
SmXidQhyHZNBtSf0PTAcdeuZX9mm74dnO6HJdcTTxrv4IcNoIrXk53aZk02K4O5p
Vjjvvqn5WH/nQ7WEglQ2kTJ9obriteWajYJ2q1EcA2u23uBm2GK1DWsELREgDVvN
ClqxOGumh+EEhLHe+0oVNzqWSZj36FX9hQ691DI/GObboWV1GrfUGmn+b+gF51yr
st0D40AnL75WnlKtslPhFZfXWedQcki2igETOv0qkrNC+4qN558sultCLGlMKGXR
AJIo1Q29bEJkAJV29Fm6b48D1Yn8a9zm/eQeXADcd3N4cL3jsaeLqh7Mpn0RW6f6
M4N9yWn54fTr9ZZCeJla65xyhfOQsQ9T9n0pb+o+MvKu49qssDrZHwUYjzi3ZObG
J1FPuwuSbbYNB3Ie6JSZ05cixJkmO1o7hBT5k3GUktp13+/kW3qgSSa+obb4Bh/n
84K9fceaO6OkKCkY2nlnqIOwqRcvX8ouhYkSuCNJs4F8TWp8lQgggtzJAY+rA5y1
xlbuXhVP1nF/167xtwYL3ORessRpoMjFSIw/+AsuEX7yNqSiRsLKWC8TFgwcx2Ba
MH7tj+TFEoOVk9MJV/ErtCLM47RO/7Xn0Mbq2Hg//JBeQczNE31wAYV+/gR0eDaF
Ri1G8P3UK4FBrLJ7WfdZX+AjVMWiqLqKQkWd6Oo0yWrVtgAa09vT9K9YsahSxJ1K
VfiryWb0ZvK7DDyKJ8HtCX3YRblQD/lmWReqAz9hiUvuA51DBlpL69SfQrkzHy9u
X56hfTdiukowxK6jQdtfqZXKvky+vh4o0LEumPMNcTQGoOoSh+OT203swvwJ7IBG
ZGC/0LXRBMsBcbJcgvXUY48dgFRSLdNrkTBnIYDDarHxx5ENKECbPIX9Qbolakbn
Z+dadiWFKbfi8MWj2eZBwxEvDPmGrs/hSXmkbF1rW+5Sa+NLz4jD7Yddr+TMxMzj
WRwG9SpOG6VHetKawGwnR2rEGfeSYnHd7BVPd00AjHpIp0fQzMtBHXOYF/pioT6d
Nzy93awTY7CI3xHoZVAyP/6LXotTpXU4lLLXdK/8DWiHqspLT4CmLmC47acaJj3s
QRcFIzLg+HJU9OCqMaUftuucmBs9L4qompBPtmiD+XTZu9MPk7r94chn40Px+EyG
QjvVWiVBdmL2dfCXgRKJCNkQ2ajhIHqNBdvmatVS4fTH2jjYw+IfV84oQIZWawpz
qdT9IRP42x3JHPCGnCh4WME0beepF64X2NgDtM7v/VPQDDUvfLxfxWDfAib4QEVd
5XYYRmbqGFe4DToey/TMt+PJl8d7RViJh7Y5QSrwXeArNPvlYGuliLwxrsF++L8h
sDnIpWUbWl4CUtwTM1tf5EQ9yGGZiJc6/NtTxgBLDJ0h8Agxu5IaW5zj4uSUB32B
bt/odDk9N2okc2zvyXIcGutL1kz3D80eU4eT4G4x/Tou8FtQSR1xLqxXUKEI77bD
6NB3XoWBw3KhrLga02BIQnSvwtjrLSsQgZm0qDdnEuacv/stPJJncZI5E4H1/Dm1
IccZfEkXlGx6oAf8PCKXpCBUGDNCCbx52gfcSSpyvhpVGi1mvvf29D9SgYQQs1Kk
fzgPzFsaslbrGZpplwXF2zoblJ18bh+paFESog1dNj7jG2usCnzEKIe7bfJqmbcz
3HSv41k62bpBLjFsXV74dQD5RnJ+lAV5A5Ms6U2TIH96Jm9QHeDOPYpGRPnmdkDt
ejz+TUEgDZqvD8xiULjUsfou6B3+COQrrKaCnV1DK1eTHbbmSN5xrsxp2aAFpOts
om89CvgoRXIjbpFkGlEQWSdSWMllOe36oY8ZWnreYjbNeMQKfD0UnJwcxMEn1HJ8
D+uPQLVQNYnwpRGPXkQQpbHmiJIUy770172a2fPJFlsgbFfkyq2fnkoopQLdxh62
CXEDBGGY1gWVBaJi/JaY8ku9Ct7lW/aPFMW4StV+hDjt9P4xpWXMUBUb8Av+DncQ
Ooh+QdpgtiTdXYab+gxhpSGhtGvyA5MjOlj0/oxxBwc55YGjHW4GZTRtoG+I62Mt
xizD9mkFIZm1XCaI2X2MOTMrJevkW2LorSLRWPcFL+GVo4dmrl8x/DWlZL14Ozwi
/mfkpEQCi0J9N7lWaSew4QCBpxW4j2jixQFBUa4sYLluEArb+dBFmuq7TjhH4dkN
dXqAT2gu5DZro1nKLxdjbA6IjbFLEYAEBu+e/5rJrkuGRByeMlDTbtLRb2B1e+nY
khs4VO8R5B7QADO+XxFQH5Yt9JhLZUOnNcqZwhfZxlM7KKRoKl2xAyXlzIjr1VUp
IzkGyISW7KwnfGPvys7bXtiQq8Nn9tF47Z84Tew0zRydkg8T81d5oxQHjrVToDj1
vTDU3VuUciW+YFLkx4MzvwnBMrfaszE8uLAb+NG9nrykbOUz3SBvIpBDMthVYRVi
6LSmOg/+49dDyIzPkG7vz8qmq2QfJX0TkZlQFyawWtDIRR6Yd+QJ/lSM9HffbMss
tHXM0f6tv589mkWaW7oQHplhxw2KZ6WS8+/0qfkujmU6R6Pxr2O4LpGIM/jC9BGx
U9g7Yfc9zzeKIeLsxqJeFyneP2gl5hh1gbSULlIhnOBXfeAByoisBBoRoC6tAdR9
reV0JdTiwUDRiG5k00xU1CiyKOItaZUNWy/YdCrPUyi+F67EFeb5wrYpWcWGBK7r
lSOuLINWkVqPSF9h2QvYgAnuevaYOdnrnBvTcOJ5zlCnxm2zmxEk+wUphxbni3qn
PnlTlOlYgs6PRKZXRvuaFav93e9KZntGRHQLHpN59L7DOa5+DowGfklxWfjpgf4X
6Rl8jgvdRZgkEUH+wco2fpvSyvbAR+nAYi0qrIxfvbJ/t0Hxz01qJSGJEW5dth7K
02in1s2+5umR2hkFQiFZ2r2WXg22V6ycK7fcv2fMw9x0Q/kVTndDegfNvMDRXPk+
m46dZyUKfMLZKIs0SUZudIbvaKhlb8J5U/Utjz40VWzFJrjtQEadBgV90g2dcKUp
Qg+bVbukgDdkCW9iYhIH+ytsJNSAlhVs+BKKhVd4tRwzvN7tIWZcizcyaj6ZbwY4
oAsP4zQ/PsNhmFpfFdzrAtItYJC3lS1155cbsbpQ2py9e0gURu8/imHvz63ZWKbj
DBzZSQLgrR8JR5RYQuyJNqQWTne3EMIGRP6HzJvD/YlU+QTf4h1rcZ1Q0s0ywM/I
uIkyLgG/agI+42Bd+xCxT6Y7V7fG2tfCVlns8hUYP+Jwy+9ZRIu9y+/fNmJkhote
nzwLAUZuL+y/P5ZPoVL3+rcTUnh8OPEXVICPG9H0QgJvVyS/lwMr2K6JFYHGywy+
JM41+t0z6S53T5QWDQpOqJyH5IrEFyAfk+piuV28cho+3Nc+bpcBMopm/6d9vIQN
ajZ0N0pVnqFvTnhWTt9Wy+b5lZPBELYOEohDMhLZ/sl2oX0f1ej3lV2aoaMTVq99
9Exlg73PDfUFXFy/YPHVPpQkpZd0s0X0xM1bjx5OpPWLkR/YLT7S618RhIANUdBA
89s/qrFVIlWs6a9jBjWS8bKYXbqhRM3C4E+nL16Znoy3aRLzjnLvKEjItPZPtSiU
IxRyytBFzyXsTDL97nwAATgfpeKYVhUWZJdvGuL3h5Uv9W6C7YHFXL/cfrg95EW2
smzT//NH+yOAPkNM+mJsBPSpTv3jMMQAvTS56+rlHK4XZk7VPMKmtekXvV+Yhsjl
0fYxMzV/6ArSUXl/jcrLl1d0N1avOxz/32qkj6Vy+GbvQOK9Hjcvdo3+9GaiXeFX
+nT8kHN/yl9SFYgIS1HoFalRoDt1BzbhhrnRUaO5AIkemlwmFOGimQQVLY+z3GDi
t3Quce5gzKxXM04KjLAa7DX6iL7YeZj/+YpY+UkwxJJtX+ooJ5Vj5yoQ5wnjIDO7
ZeUwD51b3O34dvuDBiywFckCjJ3KA8X4r9yOabeKddjukDsOLvanYs0fmxvDWzYZ
gl9Z5ZsVi6hBKkMOZWeHUzfZtGSSH0IQMMo5YshsCmKJdJQ4e6pgybdujhBjKWzx
D+jR917d1NuwwD6Ip4ox/nLYrsjIetEsDgAQ0L+lB+peir9hmI1nHGOc2uUQNVv/
p64QMr3pOqBAi+P7MI9uIBCimQQjXVnZsom0XRXdhS6coJUDBmaQ/Z5LEdn0TsCQ
V4vMx5RZn9AbYKl4/cQDOb2tFw8l3lt/muXAwwjNKNNo4lRWJbs/l0L16owm91J0
NiCSuUNC38lqa3dbiLrlIWsiczJmUCn62Y5on00KFSRc8AdqfnjtRL48i84e3xaa
4XL9hpaKhdTHfTbwENw6mSgp4Gw8HdpqDiRVeyJ/8rVKthweZg8AuVRlEzj6MZEf
5ejxsVMxAbfIQ4Ht9EHWrws6h/MqzF7DNCwnKi+mpiE9t3eqex7rBuYuAeuGUUVZ
4ZEg+jeiKkhKFAtQHbVxMSXQhAylCnFUVv25DQmUFCGA1dFcidaeOccbDBIWFmWK
0uMdpiutZGpxAAn7kcw4WKyr/VFkAXAi2TcFJowTQ+hqh2ejmCQnoqV0J1xUrfKJ
4mq3aPyuew3YqsYdDTJEH0H9mkXYRC9hBbgX2z0q4gjB6YYcLHdRvM/su0nyPfKo
e8BHEtatBh5KOEMurae8/XLCsxSWtgDMrwIj5eqCQuu0cdHhdolowOBB3T3bdcjj
NZgS0L2j3BcMoti2baMiq7+UKw/un+vss86b65rCUB0xFKD2qatkDIUufaGfJ1yZ
mX2LSVtlBX0FNzHkaVcS2T2ur1WAlsijHZBaJvtgMGelQwVXMH9S6u/9JetxKtkr
dwAc2gEBlKY9DMyXTUzDZG+qIut7rzkC/94fX5804hYStqMqPIsZrVaPn4dtwpZz
+VY6R2mFqgLrHmnId0Bl+QNBTh54mQCxCEidxBQdJxkiVVOlBg/B95fXelVbDMoV
Wyagcy+j2CGYLM9+ZyCdQSCKyso3a8QbfPnFBLEPzaq1Y63A8Hl10ikVphk8/mLI
oLJycL3dbBW1PvK2X3SJ+Z0ExX8fkev2hhl3++kepEZ6rloaATPMXSvCCL5UoroF
oW7PTEShw1QU0Ztbg173LPYG7Hgbb8fFXDfaaJ9Cf98ytczcsQ8l4hVV9C8j3AMI
aazv0gL+qkJkYLVar9SMlHo3i0mBR8K5c5eoIe5xkveh1BLlgiQIpBquPo8ZGBqq
2+w9xiAfdVzLWv4O5N6Oozx3WmZbSjWDHfWDLudOC8FUwlxqaedrcayUxuXIXJNV
8FIf3DhlE6ZYhDQc7CnycTudM49AurwwbU7CFJyeWdmzHBSkekSTOTMHMeZafQFb
ok9EGc/+aeC6Fhyf7W9vgUIW63gs2dsCaudMnszJotrBmyNe3Gpuibp57vY0gFKF
pQL1L2W4RLDC1X+Jrn3q8g==
`protect END_PROTECTED
