`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xj8syrEiTQXPVrHrWm5sIVBCc9JsUqXc+SeFGOGtqTmAsu20C+E/wiffc2mVcgPF
tM02vIAIrmGotYoZ5V86fUrF5IainkyDBNZOHTkLwn0XYq7+BX1t8pBpqGXZm7vm
AJMEk/1oEqNmH4sFNTdao46r8aYb+0yms0ysuvwqE/8wQ5p9wJVI7og0F/Qe+llj
8LZ+vowe1WrVjr9WhyZlcU43ecQVuXfwoo/ev1EgaUOfZsMQ+rW3kHapGrQVI+DF
1XM5CUe/T/VTi9Vk1Q161+YxvWU9eCTgLd0qPUY/c4Qs17MvI3SXZNeF1HoBCc22
`protect END_PROTECTED
