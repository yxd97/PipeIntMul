`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jzeZc0udH31+9h6vB/deXcnH/Qvu8FVo16id7xjxma6Q7DXvxmQiYoPAEvidzS/F
pXhARjxwR/H4oCA2BIA6+W0o300GqpBfiX3yHVvLZkD+RLHJ0j1Vp1WhsSAEIecD
te+RuCFjY2xqUc4p1KvPVoqrmtwc7eYp1nSP64n/EfnvCZxwM1cen25l9cFVeo8i
uC1MKuxn4hlzNVBRUpfVuCC3FqcqmeR5q7/PSJ38ix4jCdGluD5AR7CFjB8prrd6
9ocLXP3VqpmHsgsKlPd1V+gPyKAlv3p0qfvBZs8j1heJg3iazqGEI5GAVx5ZWnp8
t32Ci31GAtrkn8KQM1gAI4l5PmjgCfm9Cv0q92Z+exdJS/cD84PklnWbnNqFHeG8
Vts9cK9qXlNcFUUN6Ld34ewLyAKCdax++5WUVFAWoDaAc9JgxlT6Tt+ZbwfActfF
QzRIoJ1j71U/E8uN/c5c5WTMIbvPuYfcXHE3NsvVlvb4GbtBIw7Z5f1g2Qc0a21v
`protect END_PROTECTED
