`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXEmj92qRgrZMDko3qJg2aU/0l2Hb+qz6gPBVqojYzk/GCRRO/AQUgLS83EOaC/J
uNMyR+EUAsVvTnwR2z4e/PRlk5RSz6S1z6u6uc4kSubi5Wnk0NsO6x1ZCHdr92p2
Ux6q69WlvHfMdPlsTsLgFQW5kGX5FkFzQRmjPI4vowYL5ypbYYYsf3AAO1TXKg7N
yf5Dv7HpYK62RYlzToon27aaTKrzq10/5LGXOJSev94hq2jXZakBeVvyL7CR8g3n
QvsjhfBNAszX+CJQzcwnZjTZ2dEqLas/KGKuQYjAVt5Gh3bfjDoi9R1Y1v2AXGCa
9C5wojsRm3du4w0cm9lCiMq7fwC/uCZcE+h8JXcULl37RNWo8mWmOkzAxspWhMCj
BPJqbmUg0+GEcNOzl1fIXyTXedwRYBppx3YKxlHPBgoLX7tC1D5L56ZNkL5tG3NK
yZATkbFs/fDnbPGFwReBTmg1WNfVAYM6aagMgIPkJG4XY5Y614WJjcdFAmbgWbt7
978zg0BHPaX/jGLgfo+wNXyGv6S5hrW76q9S2AmrlHRknL/HI5GZdFdA9iEfNB85
qLOB9KpKlN0RwebpwrL5kBU+7fQoD5UyR4GE0He3oP/Td5gE/vH5PdlsHRxT9dAs
Kz2GtUqm9NWOkG/2oBkeMirTSn8xDVKzrYhoUcEvx2EEYRXtu4dqsgYETFp1Cu+h
41ojp58Roi4eCytL1sLWXbn3++7A+EWHFZX85/PvuX+DhhOK5nM8Ri3Qlte7rT8D
YxexjM3QZ+Nh5Ol5hPRsi+Aurhf6iXjFSfTqXE2tWRxKScYO+V03ssdUUHUiiT36
fJ7s1QDMFN3QqBjuu7d1TeWuy9H79arSXxKoNe3ikccDKMfvbVwOA2iDsmkjCChO
Gb3iDhPu9318wR2CPO5OpvuJRzf5oNRogClRBGLs64GatLT9uti0pYc3OFIMWvkt
`protect END_PROTECTED
