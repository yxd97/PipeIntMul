`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXiZrGTNM8dYqlCGI1gB30YJa/Zb7yTNskXJ7Nt7BEiDXH/W+v9llf4Hj8osUh9g
XhVGn+Ijz5l5LnaiaIQK8otMHQNASyaRalNWnEtRDB8yjx7fbBQMr3B0eyGLqlWa
lEzLHxf73ZvQhkq+nJAtjmqfnAF1dIwSkE5YOVC8QxGkt7Pd5HEAw4iIyJWFj++Y
nupETypoiUZyTCHSjuG691oM/RWJpG9IEjx3fD8bSdInXxcTDt3/pgSGZDB7+9u/
gC017QIRpxEZMzd1JYakJ7+YSLBsNDHK6Ptulkk/UDxCm60zFgmr0MqvvFvQ1lvH
vkTEsxZKQieTSf7W5I8ylJaYOo6WHi2tgupmDQC3arMxRQXcHFyZ4QuV2wehOjX7
`protect END_PROTECTED
