`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CM9jTYBVZU403ZpLH/qq9FhfHjh5+yXs1smZKmkBVoHFFHzyrESscoqFizkw4Z9P
NxYJ/4SrYvyZCHC+KK0yJLztYObK8v/NhlfRRSxr85Uja9WD8V8wuyMxu9FuunTN
ao3NNrDrvCk6AaJXgpoFVKFcdl0Csoj5diCw9rBi63AWCdvo9HixrvDKs67Rsj3E
7O09sYeCqpF/W6nQEycbzUnPJFzHb/QVHuRVy/a7Yo2BJYphVnHzVO8k2mEJs1vG
5gD9ZqjJ5AQlWtJYXUsHxOxow5Tn5fnAGm7fkcytnn6FWvDnGRKJH+DM858awcOp
z4mDXlOU+BnV/WJQzWFgREhYH31m8XgnyYrKCfia9XRKeREN8pNEJ+2RxW5/gmar
THej8wAMkRXDH5To1PwGQBYXYckaZu2RYTyK2zWMd6W1lXHrRS6muzlY0N9QTkyd
53RJY5AgU0ntNbW3dWCci2xOf4qAIDWNNCAmo8C0yRFZP9V9oXpVKczy1ZHmn9rD
XePPU3b9JFKfLxkUxkFIcw==
`protect END_PROTECTED
