`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xs99Y7jSuOyF90C0D/hin43fSKSd4yexOn98YUu3PgF2/cXkeYEU5s2UrLRyPG8O
VaFFf8NTNXKeUlSkJm5Lfoh0IBrkjGQOcSsJUvLCmTa9ShkNJegFUT9JXb0J6wsD
KTm0jT1uBWk6Pqg8u5FVWVSYzaZ+7CtkweI3J2uWawlj5aS3g8PIKA6hhrxD8Qak
r40QJgn1sadFAziqC9IVDaatIBQcJf9SZn8O88zakCaB9t8hLD2/im8uJHC4R4oh
IywqMQh+pprRMLcdnzUN9GaH2YNmBU766K5x37ZzBYO+GgQWzIYHdF9lY6pn+BuB
1jfNEyMDhCm4kYe6oja+8w==
`protect END_PROTECTED
