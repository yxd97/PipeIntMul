`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjfZhBvgv3RV8UDt3FZHUMaEKIHzTXit+Hsyu9K2nrGWM4njlZBGdDWOiThQ7eJ9
qyVCv4h1hsSsw1W5Je7DffqiHGnB14RfQtS+egm6jBJhNBAZK4vJIMb7MsJ99QSh
k5vCe2MnqroPJ7e5ehFm2trmIbNUV5ZIriGXaFAk5M88frnZNeNjDkY8rcpu5FvL
WjSn2yBBnJmU54yI4TC6fxIVNgIUIWZwTe0UyViZKXgOrEoz1I8ytNjrI4AvKA2e
lEB3kkjAjghpsFctV7hhVfBl5l7Xjd/Fv8osb6VQNax9IwNGsLwXj8yMlWmLpWbP
R24lButKrAZvpuwl2GP82VzDcGDYQaewZS80SU7eBPqJ5VhWbprbeKrRbVdJ6DMz
2YiglW7lChlCHKcVETar7Fa2vvxEUjdKJgVTaVXL36X08T+ynyCW/7VecZi1ChtH
`protect END_PROTECTED
