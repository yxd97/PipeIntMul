`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ymFaMHm7eEVeJAm6L8PQUs1AZg+YCB/e9DjRbNyhG4Er0BvbV6Opm1iIqa0HpDrg
Y9mgqF5iGZTe4cPIlyeMOtuiYT7/CBupUUt+v+rtzTfNLwbA4GQbj7Rj/4xpeRTT
wOgsDQ4rpi/VSRVvAy5bVbfIW01ms5llORr92lDQBEZlQx3l3rWZXQUXpDbTkSmU
SnbftQVXwl0YtAuve18qKje8M750cPKQoywCBA/KBw4AX8b6tx8H9KQvxoVgqEIy
jz5INU+5vIU8UM3CRkJ6wMNLkkdhBCJzgRc854RJ+fzNYqZz+dYdZGaurjjSl5cn
cS3p4KNvPZ/eHwsOlcijO3vZsCed5BXoE1M7lriT+jDWBL0aka6R5UiTL3rKxIPM
OCSrdwWthvh4wk8skraAgchKdXx/ZkoEPtuBuhV2mvyjA5FudjMcC640dE6wEJsM
P1DeDAiDvqhQtV/4cO4USze5rHlkS/7YqU7xe4A/dM4Dfu8z2EvvVVYfhy7Y+f3A
S5VXyEiwLQzc0GI1U4XFKltr8wIcKWl9W60y8eLewnX81saJ8lCti8RTV5RjgyXA
o76X4uLi3GwVZKbzxUBHjYMZpsTdawshrtfWp6e/dT5l2oQh/SbPGmbjfLipsgSs
lvNm4fmfp+jFZFAs0NQUYFhbLbIG0ErKrqpVeagHQQc=
`protect END_PROTECTED
