`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IWsTMvtM36gLW+D1Aqxs7CHA1pNkUp3aMT3XtXmcumA/C6IO6VKY/O4/UKwCwao0
TvoP7/BhskZwm0V3QMVV3E8tMUujSKywmLk7w6DUOMhpZYCFDDvDnRBM1P2O/oOh
n8ppGpbBOGZvaZBrthtUfSvAVV6nBjmACWYVU7hwOX/nt0uKkvCpBQfziNSoHglr
lw9bfP8LUcUWYMiPk/xvXDYbonRYVCguyuFAzyxwOYrUavAeUgHJCs5ovtsMzvA0
GSuDpfVuvCxRpDe2zMcPfrUZMHvT2UzdfSw9wQiLdmOycHEFREsDK+ulk2LuAkB4
778pB2GSUJPsb/KZo1EuKFzpMot/KZKnxE4PZSk4LcfGrHFMa9WhiDWuIXhm/feb
YOG8lMpFs5Pf5qvW0FVOBkdDXInaGXUI51aP/p2RQIA6b2f/1kslRotYL6UnqEaA
4ZYFRDbEb6psLjNnKOQ7991tPevsP0nopb35MEt246sN0bFoE21Bfand2ZUVkplM
JvOV3bM6ulfI1bViRPrOiXBZXSBXt7cVwInX6C6CJQ0ca1GIs2T+Wfvx72eGtmtp
//Wz3eXjlh8jCCtbjKKbWAiZSeqamalD84HhpyGMIzFMIbhsWHH/1RQgkT4OcfBh
xyNxEKf3SqCUI8flmalwS6e1oFq9ty/8M/bu2DAudtNVitFYBjZE3F/f9/rqfCPF
yyfyCxVwbrqy+doSLjWQ7BF6C6DFeF5a3/HVf3DYowzkplem8eF8m18lgi2u3PBh
G+H1aGNrkWTGhDYJCbEm4H5Zka8cNCTpWPaK9wH/W76pHwRW1Ne8o6+A4boO/xXb
q8lnDYUFcmtIb+ZG/p7ttP8E7l55DV5VqvGdeP0dFkPWMQp6UmnSukkb4AgavgTF
v67Bl1f4BTIV46flbM/NJwrpTrCMWsjjH9rkWTkH01HGP/m9m5sOmuwmIScyoxAE
7XlNa/hSliY5tbeLUhlh++mm7Gbx9UvwuHKkJf4o5YaeGhW9JPrA3/ATyyzm9n/l
7jwG86yQyEHdQiL4rVYCG/oZkhz9wSUKqXkTVTKoyh01GuoeDL7vlIjIY1lB2Ozo
7DDcGQwej/1hCGSukHYZa2I4UXD3DwPVMfQaSoOeviMCWKw47C04BI9LQhkJ5+nq
eKfHKEs36PWl/zVrfqeXtAfFsvOh+Vs3p/eZTfQaHbs=
`protect END_PROTECTED
