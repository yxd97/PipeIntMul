`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ry0esqrX2y64MaoLvQ6S5ftsBecf+OsjyxcnuVvscjlIc7GRMyZNim7yRUuXpprr
AGeEIgG/cV0zpebu8iorRQUwVzmXb7lzYQ9ndp+Hp3DunoknFHKEFl52sM3Xxgi4
WUluAxQwZXEKApaVVyNlIuGmhbHdb/A1+j9aXGzAUHULQMCs6vN7KxFMcqpIy0uk
YsYCYB89xgD6K5iPOlXM9clIA2FFKpPFAH6eRqo3cgJ485mp/4Eb9AJ4ETo6sUj7
TuxcvhrHjY8Szm06iq4avLkXcYl1wU6nWOUXHdKD9cXrW25gfCLvD9VWshWJVsQG
tAKAFrr8OJuHiUo5JqaNCLiOsrROFq8ApbWxZ68swMcHHKez9pUQrNBr/mW6n26a
HjBRzw0Frp8FcF8yE8btuirzyIlzQpsgeRgeQLZvmK4xcBIv27G5nL1i3oH83n6Y
6BRULICilF4oa3vKLk4FLqZdmzmHbp14HqJUfjhsvEbUM7BJhayGa3gjEYQUJuhy
/Cq90UyS3gPxScNf34GkGbQK8o/fX82iuDdj9a6TMxZiKqzS6mrxOUnoJeBo50Nj
o8/YvDPY9rZijtnGRxR/7hZQ0QPAd5Qb0IJPzLLCRSyyxnnP/yFBZQIoWtsV0z0Y
zllVZHO+nQ3anfnJayg122JXbG6I3Cm+JhF2eACFzAtEty6WYLa3/9Ub8iQJgsUW
hxovxiwVJSu0eVb18BdI+qPITzkUGBilZMF3N2Xs3pGrFqA2eBRPNYqdC4l30ecm
xoXHh6VZTNKNCZcqESmeST0aZ9b44DSKgfHIpWUyWMVP3tGlRBg/Je/SFI5CJsMR
DyR2aUzR7UfUt9zexndFdZPPnaonKMaGJyVggoRfAB6KUjy5aoMHEPPh6hR4oXR5
DBmN6R15fJIhFKwLX5tr5kjoha6wLw9Xo/9ote9iMVXdphiE1jy6Cbk3mPGUiC/H
FEjUzt+Qsfi1H3gEj3AVUoJnGPuQ0hevoXpxUIh6A5LjvgDOLpPUnnWPWpnCAZr9
zXZLEui+yBWdcfv5JW5lZuyRvr5mj8cNg9zIpC/vqQHV5Wq45F7yuDrnKILOWCNs
LsWRNP8WM/XoLTtTdvryRY/gy0w/MlzntWKLE0KM79twJeXwgoCCjZ7P94HKgjer
YpSy+eujh9U+0AWpj/T5K8Dm431i04weJH+ixum3EbzKruLM08ufgccaNJ1E0Hw2
/dSrAfY6v1gXFg6U3FnL5TsMTiXvU1eypUOkvwjqAAtqscQC/x5Z4LzJ+R2bsiLn
7a0JijhOYbKjrqQ85LQ/i1yhkVaCTu+NpvjOAgkRSdV4Vx3eLvEzzK3UftEJTtmR
g895DISdkGRMA+DhSuw+WYsD5CjdGTXq5skFpnWV5SGn8nZWrtNDPJzj60MfGRWa
GXiKw9FbnE6lltNZs+gtEiC8EfVA966BXm1pJC1mtnSJullBJ6Rskhd/B+3R4EoS
oJ/cBDWTL1etoPYlZWseD/WqPkQfsL8FWn3mCHWZozWQNkSuSLqBL9cei3ezbfzZ
4rZblKz9RUq6WEPpCU4/zu8tpi4tAeWoUHo7WtGnof7Gj9RkxZY4dc2P8NMZdjQR
+uM+mTAXzKTNsbZgYv6w4xKyXyG36iemcbwbzIZq7jRsW+Cl4dMrWHRW/FwwomCu
D9lj9RBil3T+k2wiR8TJFs5TyUoq7fmUr2ojCkUb3ZuvP8KhvOM6m/W7jL3/I9tp
KibkHdi+X1adfXzmryrjXsqk9Essjfr2xxYSIJN+Ny1KxqUmX7qaylUEp6VgPnk5
2gVZgNtASPJAMk9eOLUnJsaTlIX0/9aJaEaYbjPKeSvLyk1/whk+Pzt0WqwIkAp3
Nk+gHF9TmBgGdz4jARt+jqFYfIp405s4Q/7aFzNU0PFV92e13I4zToOUr098EAXt
uk7wyJAihfa1KgAYTRNJ9N1TYyWtMmChgUcDW2hKGGfHTK2aKDcLui2H1aYtWMoV
0jbiPJeMgH5Hr/2co4AcsKwlz3x9DNn4S14Y+XaA6hsdMVg757LhWdsgeALL0gTG
lrpJn+QuE6eB5U2H/kvtqAc5d6nv9OYhZDFlImr/DmWGPSjfW8isMn11EwjOvtDF
xAb4FU4iBkxiEZFpLe7nb2Xqat9CMjDIuZzHQB5/0LoGyUuvis6Pj0pbcBUSLYms
teBxSzRfkIhhp9oDmzdSlu09OZgjW80DdY3UcP1nX6YklpuJeGZK+wiuXE2lH4qU
LJEtLcnMHXmyKL+l83Z9J+oWjYcmF5UfpJqk1r6hqsJEl3+EUpZixZohVwA2FEfe
P+OXW17RSiPrMTZuNdiVPxKZ6ATQS9njb4yuSZGEGlnggqxbF2BhcpnRhq1itm5h
pZCc3xAMZHPAhVHKtjI7zDS2FlGesPzZB2CYG7ZiC7N3mEnbKkvWmpqJlhbxINjN
8AelsnbOWWAzqXZka+M7ktpg1xv6KA2hJ9mvDnYR+9yXVxx/wNdnDpHfHWqOureM
OxNcWwz9WEpsoBO6E6egFObveWwvuFSemwOWcPZT5jHJ7yJYFWfZPPewjo+b2Eo+
7rN+dXA/zB0hcgSaMb+NNRhccdQx8UyA+UquAWCV/7oQukdZtR2b5EYhI3ekPdbM
I+3IXFNeOZa6VrJNgl645CylZlxjx6jVzN30vOJMHxseFjpUEk4EXcQ0XrlXQ5HW
UZc0gNXxThh+1n8Imqiz1UuKUE7Xh66DGcRVEYKNFKbnjs6ihY5E8hvB9cqpehOc
8FpzaDCtnZG0NxRyWYGGuSZVl7s+G/2cHDa/wm2Bwzau9n05DQTZTWVmSs50Fb6y
QCtkHXYqlef4zQahKEQWRP5QeTPHxZcIhilPvJl5lc15X+v76iEiFHlFhezFzcS+
tCmaFFM4MZWoF3N3kzCm/tovOh6b4A9+NiGVhd27Gg0nDhruNv+j4+eshkxGbgGw
0JHtTcgY11VZfsyae5GjlV2d3v2sK2AFo6SqUPf1RlHyKCt43444LFw5XarS7Rba
a6KRKDT8k3lAVDwTG6n8DKru04E0RVG9gLKRL9x00+Ztyb2ViG/g0IkvzwUJk3hE
cZ+eFfRphnTWstopKezSj9gRbzIcKxBAw09nsy/I6fmcZD/lCzvl7b86w6Ogd2yO
upBqDuAhy09aoLiwmirgkSuBbYUHV7zNvPhndU9JPJHPzp85kQdDM2v4YrSbt49l
hghLhcnBztWIMmYqYx+pPA==
`protect END_PROTECTED
