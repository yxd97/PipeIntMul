`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwtmPIE7u7Ku/+W4wKEnxtjm8R5r9kwjE5a3hXnoOTYCF4udi/pXb6wwTTIdAwyP
08IGD51novV6ghU5uCQEw9DJtGox0pEpN4MXs/eggfHd23aOqUDbGcwe3BROC7/v
tXMsNsykvsy7ulajjGEZ4k0HNSPSyliJILa2lInoIKjhd+RQGCh/oVyh3GcaVJqR
Sx1QzVRomhzAtD14oiVugwSWm9IxVtyu2tjTL0mrQO++R9EElv3Zjngq7tSn8jdP
+zEZ6zgrAvK62khvbuZOsDuXv5WcV2U9aHYD3tiWSDL/7UIL3qQcqY0AhIdBKzBF
vhkqjzyl7dHAgxfsz1ZNnW91YAep31SDpNSBQ3Z8ojf0wIZGWlsXq6xFUNYmWU93
8Y1drsiUQt1kpXX8Rhet2k8F+5WBEq/ZY9Ko2EmLqw/JdneqyvkYphV0nimLcYmJ
88GVKO9ry5kxH1hpuHCsge4dTyHP4YKGcLfCz+qfCYdKUFfGk17vvNhg7YpHCJj7
o9N1SztJmxRf/JzXU23T8GFVXfAgCt7bigtAmvE1rG5a+FYpkYIrsUdxVyY/sc1v
57vcXnekOGwLwZOSeBUpVdHAOrg6pobTxzHPPDWPT2N9wMZ7sS01vT0cgz+onMDx
xCA2MmrKSaAVtvWx/pnIv7qo2+nEYftOZxeuRgPNByKt6WXIKZJTjd6mayWh/2J4
QbUr25GYAThewscJz0vIM5TZ8AM4qVz1LAhp8fi8O/4KaM9MvR2VYc38vgB9KpbE
bkCzniiISKjwZkCA6eZP5lgourLtiatu3VnnPUMf40AuGYkda9pjvfDcUU7lpbKC
ep2mNuMi5B3HdPV9g4rZ6nCiOYjkPg9gh3djorSzeNukFb3f/xIWQ0+int69dQ8j
ub6OqY/WOVll14++NyJgcA==
`protect END_PROTECTED
