`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jk5tk5GUhdTDg6LaZEaru5ChuJmoNtzSXqbovnpSn0MvGd9adxcPem3r5mvnIdXW
fvqyWxiVXGpVtM+NguEDMlWOkudnZy4PrTm9V2fLxpT4ETeGIyiDya2JSbKiwn8t
BsXp+VQaHFR3NV4YDMf/lDDSOmNb8PE3yCn5aMMzOx73aD4OqX5tZZuFVUYF9LXu
BfrD9IVeTTux6mMJ6k4CmyMTnUmxWl+5FdjBMHt26aHzJAf+0uQvYJhToUpFpFqn
Iu03/JjYtS3Dl/69w62GaQO1EmaSplOCbXJ9bpzEOald38toG/gnxm1pRMXREXKh
qTR9cWb1wkAX5AWMoaFaUsFZWXowd9GfNGC2GPJ00plwIrWxiu87PSgL7BjekPRo
/4Op9tkvuiE7hTbnjLQOn83S0kFf2MaDH9zN67AgRLiYtJSZ90pjI2bAM6AnYMk2
PEdI+jcm0umKFtUSvRsd5HsbgHhTvwzZXANXflTtw7seJ4B6iT4T/8nfMfUCOppb
CkSqT+PwNgt8IbDVUNF5gUJjcTGKvs7n49fDRYMmb8Go6BF36KbrcY+/mUllRdGj
QvaXm0nXV6+Ap0dOLAeG//yGJF1hVgdoIWYecPzBwZ3HXY370ta59u6mcmMh3NRO
ZjLhJjdaPHRhoSFisdgHgXeOgkuNHUlUkDHnlpnqTaUxtLS3a/paV7kTeMJCSWml
3eyDoCvvxHGbbE2sWnVBJzP1mRBi3eagy36/NkYvB0iQ965pnSuwomFvdtoWAKhm
w6qZdcPntX3U7QupOXWXktP88qgCdE/4jMHAhhka3fIUgIYjpuOItE9dvI14LB8R
VGaXNCoReEDO0fr53PcmShkJrQ25Ft5zbLwpzt/Pf0ltBRDAwENcFZ5jENIbOGNR
EOmhbuSBDNGfWVRLCyX3mBazuJOmoFs8EiGyWPxqFn6MWJ+00dUFrzuVZpbuSc9C
foeAsfCbNidGUl2KeesNqWQ8bxj34fteWC4ap6Xlh9bmNT1/26waILiz5Cghq9QO
XppUSOvl7b3/MKpuUNLPevagFtbLkJV2VCg+l+ZSaN12sGUG3PZ9kLaasmDYi4R0
0C11SMlzC1KgZNYTBVa5i4HlSsi/U/xIn6pKNjLA4C2cZ0Bwk0lqkOKnrTb+zj3o
eyiFHCHkdRfKLxh8/xyVaoErBnP8QjYZ5/DSujisWxfVFgdT9dqCP8Rkj/ohsYBf
suoOMFxw9mUBJ8HelyPS+hCFL6CNop5B9t6jb6XHFNIr4a4zEdrhKXLBG9WxHfgx
PmCP0VssnkqIi1hCYaaqG1oFkSjUCA546MfwqSssl/VlAGkrDF/VX5M4LqLHUwIf
aeGXNpceTztvoC378Ia9HKU/NdlRCpiqlqui2Sz/9O1HQpN4YrbIJvHFd+O6LwWh
9pevP/Q0J/8o1VLOfTsZSEVqza2c8hLc7CLx6H8RYNlxLU48x0Eo5VP/bP6wzOe+
zCyPPqmCdo77vRFgZSOmKQ5FZFPcWE1Ftwat3II3gl5BzKIgGTzhjJvN2BouXe3x
IqHI8qRGJ6PxV6sLD3dIJ7gM1B86rhEF9mHi1K4ydZMvyXajokwGvpH6SQSwP5FA
yGobT9fbqhpTGBBlXFdrOGCOz2Q/44As41avYC2dcaShq7vHfgpchOq1GMn4Nkmx
mcQzbCwcD5zCPGBj0kJzFnJQE8H7i9iLrsIOfVzUOPpZn7wopOjW0YJY7fI+TO+a
al5eqcxEAJ2SQ+Pd6V7SDgP4DB8y+8mMrzYpAqY+RkCp9/Qj/yHf5D752NrBGxgl
2VlXVA6l0txM32rJRe0kSEmeQZXwUvyqAUpHQJ43w5ExCgNCT8k2WLHryHtiqneE
wZqOneE/Qo6bWW4cpiNSgkGvoozDGWJLb8pxorb/cgzajsS9x1H3TH6IbZgfc2K/
+tGuOMAm+zSPmZ8JMBadQYG1yq2W4D1Jd+3XE30CKscJOIyPVAOvJnQCK/NDkiMB
OKGqTUNh+vVdGIMlQLrZkq0+kb/09qquKVMWX9OuAEYrwcXI66pXtLTu6q0Mskq+
6lvLKz2HPGH+mIjZLDRjNa2Kew4Dse4iaiLnMRDpM4bmdsKmaLybee7+wdn2GeeF
VPCN9wNVZjfDm4Vq9zB1T/3CNA3/M5hvksjfWa30AveN5UrxabkUVfoNvUAiadUB
LZNALEokG8ixa5GLRGc1YQj5Q80SpdqL69UXF8ZzVB4Gwt0vlJaELMtoZEF8tRAz
NC9nY5TwTFbJBDVT/Jdyx+HV4+DhX6CeY2vaSqjqzzhPTRz+EC/XcoU+W+NwH36c
xUOr5H7BnDUcxZZGNw6yWZVyUBKXkxlc+RopoSdAXXvgRpIOKoFaU5fsZ7mO5zwf
hZI+sTsrlkfJ5MdvEX2yA3btcrGI9xxWd/thLQQL06RwtmoFcHYiIUUzf26ZoY5b
7ZtvPCx1zGqJCL39OMrdLSRLp9mHwP8hzQ1DA72t2wwIOMBT+qXuNx8JYROGxq71
G/ESYyvAzBlmh+Bo8WmDTvAAyF5gp+GBKvERat5ZMnXoSsdcVFNTdaJRJsjxBTVV
8mDHeWl+I2GWrJgYgk8SVV6ZzDrGakcLZZ2w5IIS5FQcapOmvv5d3Q6/suAX71Fz
UfYErW88envv/dQnP0FXs29+kCl1RcZnH1lEynsq/7H7gfU8sagB1xBf6q0K/YAi
14zhSCw8brxE0UHendjy3sCFJ+zkF4ByBdLl9SZdeGCZVlMKUtJnQH782flo2iq2
EUBgqizeCQ+F3O/A/+jArBAW7JpqVKYskWYjQxeYzT8VtJ/dtcSOs8ue2JjPNZtm
YYStBn5eHkEpalvOPAP8vRMpmaGeufK/d7J4Bt1rbZOG3wZ8LAoe6Utw0/P6ySDj
mZMcX/7TObHOpOj1BMATL78c6m1M/aqe1exHhqguKn1vB19eKpu57zKqiYI1ffQ3
RUex68hiT07xSTDlhQXjKhesP6RlUK5sMhw/PSKoNd+JCpyi7lPPiEp7pe4+JJod
ET+UuNGg9aWQra6viKuZVIP1H08v1LYEKjPd56cVrdaPRV1++tz0gEKKFg+/Ri7u
+G5OuKrlkigHV0A/kpw5h1qqCT4S6wnewKczLG/CCWqwjn/igRe1ODXOjsTMDC4t
+54Gpl1IjGQFYA80pZk2coPQI3Xr84AlYdCnzd/sMDvroLU+pW8i9TRI/YKim1NF
aW5OL/CgwyOwk97i5oEY8LB1L4wXOtNzrm6B8S8wKUxPjhdNEUa44xaKTInAHvQD
KsNVNClwFJvmWpBsElUmllV3/P0TkWNJhtPYPbyQ4uKPua5zfYDxyrCZR0UrVJp1
2fUynL3PX9EgqtywbjCfimpVGpbHAy5iGlY3M5Tc36YtIQaEJuoZJDR974iPhPWA
iApWlJ+45ltLmB2qfEdCemul5rCWGZvLlSUx0/oaGlMoaiYPC5EtQ1JQ1ibiaexg
Dt3N1ruTNBsp9jsbkZk1XAVUXqg2m+C7727iP6Z3LwcFQ7BAK758hqxTdCB2hSSj
Xcof7Pe9ciz2c2hKXxBhgYI+qBOONPur+Gu9czifTf/ccbZ8omZrAtG6wwfezu9F
T8/mTrxtbaXTX321P1/zUCYKwjGC7vT5TJ6Va4bH/vpZoXO+Zn/gLSbAw9W2hth9
cb0Ao+8QCqg981ct9ETpftcUqJqR/GkmALyomGGvWPpitPcsAIo3zGFg/Ut7LBxB
U+Nz/KI551EUg9MXyUjCqvbq90ZFQAWkxbhfDaPvVGQ9bT91V3Ntdyi5ck4YChKQ
lirMKY2I+Uop7GPWVaUOhk9VqeRvfOigI5rZSMB2XFoOn7DHhyiUIA/NDnceEsRP
Vte1gtvijEbMq20b2nJZ9NKiW8RpLKBw+SOZHJU+HMst4PQzVkrp2TdhsL8YftN/
g3IEsqbJJ3hIuiQgM1qg7CAJVUv1PDOBvGWC1BH62k9axlFmdZw2VaDaMuLYEWUI
u588fnGdefisi+quVMJPb+5GqjebOt2prWbblu/JRVKxi8aXW73PgJfurO5wDT6z
ClhmASymFXOPGT2LGyK9xqFpm0ecl8ZpU9CiQvbR5TbZQ1lui8e+Vib6BG6+bsrP
PQKjOP5wuc6tBmboqcuG0rOQxXS3dPq+fZhm6LnE50m0KYatcQixddk4sXn/ceA+
gyu971ilcaieMFmcSAdxDrlXsZ8KviPIU/i1LeDF6Jbq3LIJRVQVZ6i3AqERuIdF
8aUf07XvLN0Yh109BJaWHU/tX1FyUxdvY02yQEXOMHzJdke+usNHAZmvzFHkqFGF
fc17/6Z8Lmykmebd/ugN/3VysF3gHsL9R8eX/X2c6/YxB6WBu6vIKJOzS0oXqboA
WAv/nTmxj5vlQdqDltO0TUEcQU45hNvZHvOCtwcd+64vSYR6/hh7vAGzruV8bPSw
Wm+I36lp6NHcf8Ro30qTs0RArX9JxRMO7AWOhcXQhitAWc2x83AK1uk2iCJRWKji
/ANGABkL5t330PTCBK13qHbz2K30S5sFMfBPoHApVYGCMkTUeUNPPbiBbGPQ8Oo/
kwkiIzKLRWylELf+L1PDnllV+98CEBidcFRSVmJ8FrqXxRkHTx9IZNIYS+SJ6Zbh
0JiUCIfTBbDn+1RyITcQWl2ug2OJ7vRAaE0CvDCYTUv4QMpje+BLUpDIc33OrVSV
DMoZw9r+2l+z5ezYVY/svHdkpwxyLxgmVMny5b9KWAmqKXyBA/0scVk0okhXlLX0
o2Ypm5XO+ThpBiwQ66C18tIcegUzjjV4fu5mZTMMHgraKptsBmtQqCZ75F9TAoDp
AqGhAPq+kZ0nUBZcLoOMNUswcV68g8pOqWc2DJnLWGPAkK/ZNEh3lTgGUZQoP678
ZS1QaqNIipzICukzlFuiKbSQwfCvVbzvAIQJPPTEu2ON5ihyYzgBDR6NjDTu4lDT
H29/W14N44gWLReUAwp1B1CU1u/a1g3JR/hc8WuLdtGRSJ1gMtpJSGrDKlrH3pgi
wWCf9qoecmJ/aF0YQgtZPyUGZkOw4wtYr+WtVaRNJBA4Hl4l4444eNksxTYAsnfn
fHBG7Hz36z8vWpnEg2x+EWGq8kNoJ1fz+bsUOBlEOyGDMZOAirLm2O/+P7E4k8zZ
Gsj8gOI+uz6BmwUhbRlT7wQ7fBqJ9OFOVr6V5CAKt35IjO/lKxLxotrgY47EMdNV
VlNXIavZRi0+gG/JHAgQ3m9EE+pLN0mu3f6rwuZaBpRY1r40h+kndiSC0TPKP6qQ
QoMeplOd3GI0wcXQL8Bm3XDB+vbki8yXR2q5U7PYTvTT0VSfmML4hBYNh4ABq2im
2/IoVev0eWX+F4bj322lbk/XK8guAcczOPU5WrTHfPH/n3/El3k4RvGN5b/3kmml
LkENPnN2CnJyZCshQNnxD3HxZz9JJ6Rc8nVf0cyUcvmXImQj7mt4b1Yc0v3HYGtt
7HUZq0cqEkfQOP8aLiAN3G0lAJcpwzoYkdRKJoroI8lNHlA+1lyURTjCJpj+kgfD
0m3xWtsXC0gd5udS7Xt+q+sykl+cRzN9cPgxCMS4/gBS33Scyyra5o1WxV+swLof
89L+MXVgogL4MEfzsTP51BAEJWGPVsq+ToCV930MyByP8C7blRidIodnI9qUBxsw
jAEt6fVGgfZCiVx06BC2qG1K/qlKm8LQpJcnZQ2iySYPyw1Xxw//kmIK66OpYxxq
WrMpC2sV60ZVHPWArecY3kpaNHhDDc2uApT+I8WpYohpk2GdxUgAp2Hnl3srxXWM
QMbcbkaSHGVKliEp7lzGPpIknT+d2YmeVNpmCjOZq6QTeyyDfGL61vmJ68Ur7DnN
mbQ+x2rdPkRGyDx/uPN/IjBwTD0KFHTi2C5zzX6HP58NYj+n38pcpXImbQL7vihV
+4jX8Sd9KImFkyLx4yByJBbj/11UFUBP+d1/Ycsu8IN9sLEk8gSv2Gs8caFQAgq5
iIatvUU+NA2jMa9gT02hZo9bcI6CR4Dj6aTDGedMuHcZ11diZxk+7He5bv2IQx4M
1AmPeO3fjK702LLwyInUgtQZyTx1jGR/YEgzBIgCFRFZ0kAmT547rMS9RfUlV9ct
5U/xZD39GOahPjuxQWGKKW38kM3flb5Xep65TAtlQH909WptwUs7Nf4MArNki0mS
6viIoIdHrNj1DgZgsFSs9ma7kWOZYTbcLMYB5tyuh31PUn4Vte2MZYAZH13Oc+uQ
Gg+8vmYuqxrbob9yCseekMTYvu1hRnzFaKHRtFxoySkjGow8u43X+DewUJSL887w
HfI9YfO16TcyriWfsjl/C/qxCXhzEeLGx1XSpjWF4JKZ54keJmwyuUPlQH5Mt21B
XRRCTCFpAaBpqs6wK2gknpA9YAVvjp66ErGL8fjmHftrs7D7reWSRVWD56g3t4ft
hUi+C9xbHQWhv/Etl055ZR748h1JQdlaJ3D2n8h2OEQSW/HhxXgcs5yODCe6M66w
nMhcDvRIQJLth4mJTxOOx4jXuuxhk8fcABDEV544eFHWCMBfaMEG5ybWIyJPLDtJ
5Dhmj/r0FjVJtaVQiTA4lodN6hhYwC64d+seCGtyPlNijwTA+Z+W530OgwEUVA+b
gBuFqzSfVkYdzO7S0HqSNBENoDU91KdZvM10VtrXtszzyQa4aTP5F2Euo4syX7dq
iPSrxwOU+Ri5USXUWQE29LUfuHiGZKFfhOiVX4yI6iMlMLoHjr8fkZE8gTd1VK6m
a/rCqUFNSCnP0VMQfV+PUDrUCIHupbwQuwLTMcB/UsgSroA8vjLUFAXLwZe2kzgx
mN6DHAR0fhC5YWp5ZZX/Jy6Gh+SMrXFMXIaWessBrkH3g2zyaF5M4w0Jn84pdTAp
LnH9LpNpuZE6IOkjpVEUhBWpo2mzez5FKgKY1KodufrWlJpUnFR8ZmWD3D9se65d
2DZTF9qFLa3m+8/K5sQJx2R1ApC+tcnh+VjERzwDC3aYKdAoyYdI/znKViUQkWBB
5QFzeEpk5w7ecJbjJ4oB5urG/T+b2+uQe2+2FiS3B6uO6pQxx3pKu38n7VMvgpfG
u/4xc+HPkmuho5sP2ZFWZTphvU/AsdoGrgLflqNFbIKxn+fbBEsrMEBmInsbQpxh
W9NETueG+qDoCz3BmV4dl83R/D5SfaCp9crRE1LEBctES2YDdjQq/P9tyjj9bLxY
7Z/jAwel6rL0DVRH4AiNPxiO7hnxP6OnpC8azJO/gkZmo6DO2Qfn0kpVaT09Xa9t
KJdeLCEq7MrngJaYK3xHWUTS4lXRgF8LBqkgBCiDq563UVsqwuwjyh9xibHDGznm
VxVUqkwWD6fneBriZefspHldIaDzy0uBq9zm8i5NP+Bbt0Zsm4ug9IgM3RQBS96W
hbUMSwh9ywhtoTiQg1baew6hQmo9+wGyYMtVScrKykIO5WpE/Hw9GEDGCvRwYDn6
GLOnqop7f/FbkGZD8J36EyqCpKmvnB0Y93LiK70bf8Q/cjdZ8hCTHRIgPwe7j97H
SoY7Fh63M/Tl4+i11HuCmC0bgp+y5RI6VUcHZF8TsTIqDNW0mW9LSjjZenUPE5Kh
d/4IzqVBZurgoOMsIFpeJr/1Nx+Fgp/iQvg0MZLcjWKjvXu+FQ6Jel6erNYXWMiZ
ahijg32JOjVH1jYnzaOK65jnbbwLH31H8iFpo6hlRajM0XZmSHIBCEbadG3smxV0
us4z6b5El5WOVPXP01qyApTT3WbvV2+2ccYIxfN3GVN/l5cRSOWyBEto9HTSEeQG
rrDSYxukUY7HgMH3w4h37OZx2d6TJaffojvqNhEfdOnspiSTqmhuhfz/PofK3BhY
8VTeATlFqlPfZrZM7DpR5SH0g9Kclgw1SNa2zwd5fxsWMNQ2vpMF6QtF5b9rWlut
iK07RdhlYAXaG61EznU7n8mCWb7q03wbKUVVDdE7cy5nStJ+C5Pip1+GMRScikzo
mvNCFCMRe9XGg7y1lAZFqUBEBLidm3J0V45plTWapHX1tBGJvShy7PuTRScnQ0if
OCfyGhVZ08hiIbfqwvYgyKOp1lqe6+AGlhx6F49xmslY2E1Xqo7v1l5rVjtKXtFK
fahkGPGTx9hBh4DqdH/FLFLbCP40GpyAZ34ied3zBSa0ZAuRad5h+0/xB01UktP0
YvjdnJ1dRFZIBIdpbCUnan3sIWogzw7TfYDLCpnZdwtmbse6lM2o/hp+YrU0T5BL
tKOChc/+B+E2mdHCAFnwOt5lIuL1azcIxLh8UmYLmkXojVuBG8AixjBimANHhHf5
vLkudJCbAr/6YdH/24AB+ZypCwVAHP7+OfvTioAV/fZ31NkDl2wkQPCSnjzo16NN
09yqXNdmI9/HPZj1Dju8awKpnqXrpCb0ZVu5vSa1jS7Hur9+KlK+mtOt0USak0h6
j5AIdxuMrDwxIj4OSCw9BqpJFwSLbsGPYUb5mh84FnSQ5Jzr3/gogLVt6UutLZVt
NeTk64zLUNe+mN3U0KDZk3qNVsNilXpxJW6eALt7QtUMeiCnrkDee3Vj7sP9bLYy
AcC089wfZ23tzJDWLezWG7DRKgJRtUxqRSORUTvhC+4Bjg2BW4ZX9AkmX8GD1z6L
Re4HQU11R1LuJIZa2R/3w34675slEnUxmi0cHx2R7h5OG5D/IG3V5eysljnBrWlP
oqpDZ8CCH9M5prrrSteQlKfI715mhDT2IThFv/sen+NfA6ydmsakeRQaGLfs9L5y
lloJ35xi+0mj2vFsmr/SvI2SWBo7bkXr5LrXbvZPdTnE4ySQOtt8e9Q8dJKc4A1m
H+llBFiubfLYbINCyBvJw3QzANAXb+XUznKPkHJ8wz2Zp2F7s6lplHnXQyqbMT+H
8R8VJj38owQ31qBeBzirmv8anMPWOr1U4VVS1UDlbiD+WPCff4dekQI4/AdWMv6r
aeX+PtqacrrJk3Zh5oGk7f3lppn08vxuOb9Aur5CkVAcIjptPChOwLvNHHU0eajq
FM9nyCxt7xjs8yDP1fuwqOs4Ke+ZXPOc5ZNqlbk716J107TA+tBWDwxUnIfFSLPC
4QgYgxCpE/qh0urbjxcF5Lxlo3cudKOw6rXxbBn8l1BbDXv68pruIbZPRnT4cS68
vuY0Jo5rRj09VNspUYfw9xjzHLO7kzedpLyzXJWeSMASj6JU726Vvl1Fhw22LZRQ
3VmW/o4m+OtHfiEx63ocxQJOL0v0wjE8H1QNqFQggy1hGO3aojJfmTSpQxfW6hdK
aYGGib/LjEiA1Tl5AwZKHYXCsptV7L7nGRSsVve4erwBp8K0evyFjOdQVfd9l1GZ
lKDQZBH2uYhrl7bZOt8VoYgOeGnlB6MbWDSGyD7ZXtmvoUr4SKx8RFhHNhcBIfLI
rB8REYs2Xp1iD9NmgZ72500CeucZwT4zRR6nSs+X7XNi0G5unrHmUVlG0BT6UDOu
iGQPUd2PTmvPFMW5Cam5qmT4M3PfYBctIErAOynx8KICKM5WCkTixhNpUPa7sVwd
xUVab1L5ckE0hgMhBuNuDQ/HDELBy3iYCByc7INpzqNJ1MxYdCIdTzBbqeRC31DZ
vVK3yfvSVCDhV3aTGWO7AJqH4/OeXSQj/W95v/+/gDFzAw6Bv6LxrBXTdjWMzCPn
W8W5DgYLz7PfUCk3ciklpvoBTtY8dS7Y1wSok+zmgeY7UcfkmfuMN6DcJmclLLSq
bsjvE1MAkdn/q6cW1WvLnGAhfcjo+SOk3pzUl3IRw4wCpsJit9uflD/pZeBPqmYA
8+chysppF6/KbGrtvylDZdE6AE9Z9zdAZ8ZwQDsvQ5ilf6f9OgVyPd35n532cOPb
1EYw1qAkD/YbvoYcuwE46FLdB85CGdPQV1nDP+J0tWj3OWWLQbPtWvoLXFmS5tRx
V5fS0H1VNEgKKOCd3u3hAwk2VAyt34lJXlzLvknJIzR5A/ARLjnwvRv2XLn/Y/Ad
HJ2yt0AIcnSQBoUeJNR2stBAQfSMXK3geRIS+VWQcdrHKaIHp7wK2niw2uz9P3Z4
nY88OFMU754MWAfdU+iU7gEByO6T998ciemwuSNv5cow4YnWXZyEs81H4m93hPP4
wSt0W/FzY9hbUeSRrRiuYr4jdP5/zuxZLaySTxk5fT5pM8uCFOBWQDpPhyUReu38
unVe0gTckpJBd8ffF2szLlCIE1GDJ5p1PuAJRwX7+CxINqLcpICuo1RCYor0/BI4
wyro12vQfilCfHbjOrBQerS1VqHVRL4hgCosFzAS43Y12CAMSznZyL8xAn1C+Z6t
Rx3cKrNJlSG47OZLPSi5e82lDcQTxYVs+utNKoYo53Q0mUkheNJ8yZEawplRSZDe
ebZsmZczTzP7oz+rbqFrBAa8x9iVMxsYVcpAYVntMhebHOBqx2wxAbxRhsJR3s9i
/avpEmLmLZQU03emzzCB8h9wLBix48hx3cUdnYIMCdXm69AqNvP0RWt106jDeZLV
TcU+G/6cDseZHvESSe/sSiB4IO5SGG89bRC8xrYNTkH3+XYhGleUDEaKHY17fW2p
FL+MBEqTC/+HaZjQF7VIgfgDgYHcVM9Xo5TCLCVuVurtv4mzZzYug5T39quiax1O
lEeaBcJq5rZtVNm5W+la0L6wR6hI5c4riFtfeIZXy83W++GBiO+Sox+qrr87q6Ol
EWByBrpHaj8MC6hVdcfYhDXZg1G5mQEzkOSSpzyBZK2VE6tENXz/AXcZGnIhOnej
ziiJ1VVLuxpGDYq+GghgU8RoyS++Y5NdXTln25uilJn8J1WbTWt5fVjQKNgRHi/4
n1rxreDyFEL34xhIl8KgTNiCCsRH7wZWepnGE0Wn6UUcwFKeuDGVJGuRv0TRuJTp
iCnWcvvhzJHInOeclI7MhE8nxPo/xVA5K16yuZ0yFYJgGBA/AYGfhEBPGDcAFzvH
C60dipGS+TeeZsWN6au+5zYHV6YPgMscF6u8RWpHMjr2PqTCdSVQQ7ekkOcgIUbK
FuBo3D8Wcw45y1rSUG0AyvLA76k5XlnWZ5diEUy/OCTIOnR42ha1UiQkHJWH2xrJ
gxCcc726lTifvJOdca4UXm0RRtryT64+LJf8o11WFCsYgepkTX4JpIpWkG5SjPGN
ucmLHliOoYwv8+gSHLig+FU7ERSXYEpDMefHNHwonJ5YSpcaSAMrjDZWBqYFXElC
Hur4Sf1eKB+lnX/414nEeizQv9hn0OEhBYsckQMIUoR/puHqbTDtcj4aIdG5iY99
CpNF5aPdfgBbprWSvNBI6SKNGvK9oC1Z5TR9hrUEW9XVFsWOcVvuG89IXNm/61+W
vfQJmlcmyjcjqKcJhHvVCO4evz9rJBw3SImgKkTyMN78J+3xhJhyAMVJSbJhXb96
VDarlxluA70HuiIbQbuZ6qAK4EABZ2KELDS3RHJiHvoZ9F+X0J26hCJJ8NDbe7OG
umx4TGDBb4bGQN/31OpvO3xhycIVp3qAzg204BPy9twUjWUOPmuekBqRga0X7Vxs
zUzBS4lZufN/vwocoHGsAZnPxpg+RPoOf03iTt61sM3a23nP1DbV7oZ6Lau45r2N
fk5qxNIyz4SVl2zxeNHdJxf974Kvjbo7leFyT1ZnVwTSpQqCo/CkUJfZnmoovpr8
aUgImen0kFBdfodEROaZv7M6KCiPlH+YMM0FP02D5LHSi6vqOqQ8wpsCZtW3e9CN
NMzlmK0HHEJXm74aM/FNeoBoj4ca2d6tsChFjz17m1VQJxNDtyWvC1XdxeN/tQw8
fTnAd65hjF7+wisgrOaxqmJHWKdVjyuuf7oweN/vZSU9R/eknfzCCLi+QT/AUadU
9ynyJARfVPwRCfim3d9wkz5yxwjELCj4ToDQRCA6ICp0Oje6Y1mme3fWSsXS8vxl
CC52u4GDIwtWyOxGabRU0Zu0EMfzCRL0dbwYgDsNA/UboQHgMj56jT8B7mDa37Wh
/bSBB6Fzp356jw0NNuzKeLS/71rtT2tgcVJ7zHYkQXLochcn6d1qoIe+QVd1IEgL
QzqwVO54f5hR2hTopGmSMLLp9YhwA8QwIW9AOFp+gBPyc7GcF/NtlJfdS4Hpqf8F
IkXQiO5lHuZJd33sfWz7nu2i5VXFLeNbKykFe/doh6pyLGYrX4RIqyd28jNLDIR2
j6rjnREZXjAug+dLPBC+y96E0NRJG/3jzHu8h5xQeBvORcMEPzKtBoEwCUeYFD3r
uGQqmSLeaQDO+yK6KSNmSo8NhDpUuem6C1vxYaGVTvmt2A+NHCIAR2w+tKc+eB5f
u3wtfzg70Tmhqj3jqmbvT+1ooAgK2JDOpqJtedNg/ftkptS/PWOcG/EybIx2tA4F
BBMDCN/Mw+kpf7wl8P39PXLLa7RjivITDWbnCoFAXLmStWIP1k8+hW3+lRQyw4XW
7Ct1NfbDTfcz39xJRgEeIGJGri+hFzqP11WUiCHDglPfIIOjuZYUzrIHqdv6mKqI
kzKaTaDQ3HygGUYaLoqfRDfs5hwS0BWIeOH/LCyIE3KK2FyzVF8l5x5C/fz72qrR
DDEZNDPMhmUiGYMLCASXp+ZwRVHE8IK41uJ74EHR9T3wKPgTT9CWA28tY7Ob8O3y
NOLKgOpaAT+thyGQoXLK4SBpWf/am4GX2HaNOcLcf8+eOgZsPEFy11APBxpNbDZZ
LlhOFCUATzixC0BUJOz/O3Wy0MchefjKCihXFXSoSv24aPXgwujoyHeKCHXt5Iq0
Dp+f8I9lVobpL9FymaVAvs/WbtInoEIp7vcF2jJCu20ihk5p5pAsI+UvkJyduZ+X
9U3Ctk+4EGRGFGz5TIzKe0QNSj/A2h08WWhSk4+0rGfxCY/rwbhjveRv9PbdbmkV
V+ISDnbmREsBDLGdpGadmULlIIuW+V6cjz29v6et/q56R8nyDd/hSxgSedNOMZkO
knBpQ+t7+PFnUUA+SYmAoqi0F+XWmQ4zp2x3GF56josVTh4NMb37TOfPsDVTD48t
jyVtqtD63qMp/egM6Nf+fvkwdq+YkhXbAzxvgsRvkwFiBaPdZZpbLoWNOX0gqLTM
TWaQ9EuL+UHUPjAhnLVWc7AFqDqqMkChTDYKwPU9OICD2tdjt8BhwSGOWo2zLj/7
K9q4MdIlJBgfE8nvLq+FWJUo+CDzxUidR8rfHot8DD0eqvyH0Q+yOaujFDnBjn8j
0P3aP1w/LkUbT5u+V2M/1DAR5H+ROVkdvd+4UiSSaZm5KuelLGcNWxyYJY0VoN3w
weuDCpXutoWKZkWMGth2kjxDDLjkTjI1n0SU3ewXyx8Fz0j1qcvxYdGGKrqk1Rd4
7Q7LVtR4iMDTF5OrTSg8qtqCQCkwka9hLFCwnIt5jQykshslVpERQiWhaEUuLbiI
Ce2z8lLJdPztuYrYHpqG0Klhm+q65OcrMfdhjUOywnEnM8AMmEucuQO0nI9aY/gK
akwD6ni7yMYLk/FRV2c5tvfafDVsSz7H3Mhwe8dwtr7Cll7b5ynxS+VZXdrnhNmr
xQlavoey7cQRw/IUJVKLZ4eiI5+JzRKTrQBe9rupBUG4E3ArA5YSEOjsoxr5/Nw/
sXvv23FquXe2Uwr7geoU20DXv0HPlEC0ccbrZJ79Fjud8/AClH+ENQpTOpcZeRSh
tnj3LQGfmFfnVwVkkj4/g4ZqFavraLB5rqT6yszw1xW/H2UzkCoVHyPrF/m+hI+q
ffVVvo1YtyIkvaNlsmAjop3i09ILNjdKfrEmTCduB32dyNCsT81WCghO8DOMPqPy
Gk8Nef9AQlGpOmhWo2nIXR18CGvn3sgH82Tu/KVFAErvUjCwk7JZ1aGerIpa6GDo
/xnTgNqhkMsKdGbgQz3XVTe49LamLqxCASUFenbOYUg8ht/9bQg7HgqQng52oEK7
TgNMfjCptcxkf1qiG7qxn8MCamuE3SnoWlj0vVd5pNDyvg1JgorqayJ05GtrBJwu
KprIoI05dV9NByJoBHFY+8VoFVyYqAectSKgGDaNmNQbxDmbeC5vqmCBISz8g1uH
e/8AKpf6DjDu/f9JcesFo5YpK8Q752x2yU8w1CQA71p319XFnBTuMqO1CjPNfW2/
nRzuAT5x1ZYlAIUiYU7Hd1vJgWipKP4+bcPoJEZnf69Bmj7yRJjHUQynhmbApcms
MJ19EnzH/HnOxuGFoi4UHWWiTvkO2QTTjtSmxDWv9uXAvmjw/c1uj5w28uqB2NMV
fRo/KaQQWdmxD8m/ho1f1YAYMzcdwCud4mqVWsm+Iv8I/iECoHzzVUG/Le4ISvlw
mMGZ/5LVn4OEA47wnalBdgIOnrZD58tVGrAxOPNjAdRlFti6G3hoOYPQbquzDtg3
kgqkSqvKc8xti99nwpULxeZ1SsN2oyDOgH2jbIpBsRCspm+j/Qll+NH6v2LGgpIN
EUfCZidwLI9zZYWImCJ3lSMXpaTVZ4nuYg403q9OB9tVtAopxnUSYkCN+C6w9WZk
DRCMgz8lL9LY6xNLqP8d9a6/c3ELuLyIQsvglFU/sm8tWrQ6w8fAgRya7QTOXfqJ
ypIacoKtqUPDOVltTMo2/NSem98J1oyyTqolu6YI/qt/leGAqTXNu7CcN+qehLrB
D36sPUFeuUs4QCi+IDvYiEVe82M++nZO+GUtekHn27rJD3FBvQ16MNYIC9q3q9ka
WnhMS8Brnx06E9dec1mU1LUvlJy89Lppbe3lv7TmRdlOmdc5EpLZNNrSFZ3Z79zZ
r4jA++v+BGe5rGDwFBrhZvzifZRRR5MR9LPEoMXKZS/cr2Hqrj9f20xhQgxedCnI
kGw5p9BRJzCRUVIg/XzBMlE5RDHhhbcPy/RhDpBZFWiOpW9LQ+K6CtQ/Ws825Ryn
76lnqQnjab/5Hmev/866DHXGa5y7rOwfO937+Drz8UppXkdpmJxrx51g9r2jexpM
GzAiy05yz481VuWBKAgsgxhHNygPwucX9oL3Krgd5VdmWlsAe0etZJvuwIZOG/eS
hnAjhnV/9IKz9IQYxwaL0pfWETxtRstb4w3GtaQ7ITPokGrvycDr2Q7a0w1bY321
Vy1ULufbTh1QzTEe9AeMb5zd/wmZPFHKIt305cyumlsVBRznFJyEBYXkE3GUXqbN
4sP1D5sG/iNFpGm3SGFPbX/0SL0z5JFXDw7z4TDqG5+ndu00aMKRSvkf98d2RKbK
CmNdqdZhN6A+4fiE+HHiOZY77pBySKrZ81Rb1RwZlXIZWjF2xCMSEA9kjImYlwSz
zBRSIUX02S/yiqbRIjkcPeCQECiwNFd7IHDnsnRgE3pTQENkOUzphB5uf0V4PwG7
ozeLvlnzctVhNCoqnHA3tNNSKiVTT4pudmvfdea7pFNMp65zllHTAi4hcfeW/T0E
PxVesFBUKeGe1nUWTIHw7pG/vF11tQxsMWmrHke0M9jKYKgUdKPAzScByPH+pGD4
SCzQO2iUVlmXjtkUIgjBGrh3vvYGf1nRZ41RTi3vcGuhhwLlHCXwxB4gCV58jIUo
/9A7QyuEQsiuQJX18gY6bgs3coxSdYxt1F5C5P4VTexmA5MN0WzTGb33BzE0ll6F
gVfV0sM0zI2NvR6+yAHVEweulJJVOTKR/Osm9lUZo6OyCvV5TIhQs3EvnTGZFN0O
6SPlnxZ20qrwgKPuEC5XLDCKHw71jsiJJ4myFEp9KGKFMYdBGTZZjJduyiAD/PK0
hEm61JKamSK1cM/vk5jbeR5HCJzdv+KEdbPTDPk7C5zWYojmr7N0U5m+U2RvrezJ
brqG5OxkNkSKsG7uquUM0A6CuMmNiQq77OjDWrEUwVW2h+cs2I+m5BS7qKfvyW/p
/q6OM8paOJcb/gzbv99PHDGpLWozbiZIoB/wARBnfNjWngMa3lTXNVjcizEAw5rN
kchnJD44ai2nEQuwkpj9QrYyeCOSVkJxKyJKlLvZQzOP5lNhbaqRyxswPkYTPAHz
jw6wbdjn1W4FXq+3g/As/SMecdaANsdo/AwKRlVamxyl3VK+i5xuQMtfeq1ogHiz
W9sqqroVnlARN6Q/fva7gADbPbVleitw1WyCQXwxybAWgdJh3KKpYPI4ERU4ZKeD
Cy06LcAs98SwgNRzlL2RWQ6wemKSXFkqQ5AZB61XO/CUAynkBX4CNnV6XyJQHCpm
ZERUKdEjXRSkBLjtKnDuTRzCD3CUTegsBXMRd/8jbLl8XxctfknDjLb1iFfys7nE
fuQ9aSLygdPma7IxPwLOgAsXZkzeowxYkduBD3TbBAHEfdpUfVnTIyBV0NNscN2x
do9TgIH7jb84RQRrY0V2OCAFDL4+MUhHsCEK+SPHw3KSaT4N14xGXgY5fm2pWOT4
pJYFbG9EYVmTxt6S/+x16YxO7DD2EOGP+fEb8TEUtRmBHKEV839HoKccbcsJiefI
2n2abES1vBD3zFLlzmydILEWRjHVYAIxCqfNWK7Fdwley6sfUJlr0Z9Vr5GWiqcZ
3gQJk18HMUEoB5OXulsE7A1vM31Fffk3JnjN0/a06C8sQ0uZjlONlYkpMTGhaQS8
m0IiE+e1a/KhwCXPOv+S0sOf3w30FJS4UQVJ5kQOWtTZkuj7iAsnIUxH+7g7L9OM
7NA+XepqDXcweqFG1bg60823nfwuCJ8M/DQe/sCNbw4iansOh6S/b998soH2Zq8Z
dXOm+kFUIuV4rJrAVABjNbjWT4H4O6UZNx5hqVHyrrm8I6sD8jswOqTTqycqfMq8
K9CDM5CHWvIAYlSMmUqG3tsM09N7TpNraoMkbOyoyr+Y/qSZEAZvVJDikXKC0hWB
5lg5afe41FO0Tosi97UgvM+hy2Db5RDFyYX/IspL5a0iqVI20W6gtBYLyqwTPstN
xv8HZSH5hbdGHW8NM3ehgF0x1iao4K+avq88X8TeLH/eJzbT4KUHYTsrYJrKL4h6
NI/h+2fcQTRDM98BCCm055cnTXH/OiWe9ujyGytzOBLOAmAaLMgAOCZNXabBEN+I
f5I0QbtpnThq6SN4Q2vLdp2LY4D/8cmeX6oQh2gpj525yMuxinkJjP7d2VQxHN0X
vYDEchKyyuHijJnFLTzqB3kHIeHlzegGc7VB8k1+7BqaZqzsziHsGtCbT7SoeOsY
ksT1mzAqesvFboD07Gsrk1nphkmRm2wGVyyInX4U1jXevxHHIHsc30ns8HHBOily
TZ9hKfCA2u1KyDOB892Z6+PhCBoPcbKriApcnGSk+G4lMM4DXlS8XJ27JKdInKE5
PjGdifmGxDMv3owHLkUZMU1lAHY1GL499iiXnbal2CmAx1l+lZ19QLSC1OsCBDvl
Dy4s5USJh2L9869kfBiT2Fa1ew8fjcdRZifEVHeg8i+6qe+uAoKRBrf/WGh4rkyT
bIAV/3mZ13A1eTjs/5JbvtKLpROarbKdHuzbfKQWDTdMRmOtcQ36hHle/tuid/9e
PI8bj2h1hC2qf77+JuYdNSk08Uok8hDfgpQXSsWVC8y7SkTty+MX4Q8uFF194rpF
WJTrbCg8RXR1gUdwLLJeBHa1mmBgRDqOfDRBS4IVeaX7ZKcPwskkactAv0UXWUDu
gCGFvy73RRfVzf8prGeX0Xo4Hpo6BkFyTgCpegi5VoD6jfeAC9jR3C0QkRwj5+on
FVc32PM0QWxOxNRJYmH3fGbY2aA4N77TlRcrC4WmS2DAhjBvFQgFtqYiQsq7G7q7
Hs2lxvJ604T8HbVNeIMIjJBMwSIGNRdW2qNgtEbpxWsosmXpt94UsdFYQeb/wM4x
iMN6+YI8//Ae2wkIjOeKswtFiDWOWX1tfR6jRl4Ow1OakiYTgwzuMIX6lp+oiujw
s2Hn/1wb4lX7tUlH233HYa6UwRz2oz30uMvb+tBJnH7jlu03aYWkZpVm75AImCKi
8TTKNORsTa0hK2q++0hcQlCuU/5WwpFVhmll1BvHXumMPObmajM9Tl7kejNgYrd1
+8u/kkjYcFkCiejxIhXCD6ffypqbZnKObl7HHa4bB9EcoPPN9GRnoxoglT4jnQ/f
4D9t4qETyJO5/l/6GIAlMZqnfpaN2C3zZ3MCRqeYGFqNmZV7HiQZIOY6p8x/gyTl
x5Ry5ihu3RYiJkaEKEDryrGlJg3DAvkZ6pu46hWgWsvLfvaD7SC8jK9jm3skIWdl
Oaf1Gwql9xni6yzUCnMoLrx5afVibi4VHuT+ChcCkGDuYfIbPxz9lmCKGBgrjmdQ
t2TZWU4++Imnm7Gbz/RCI/NBdyylf9R0AOJcPFiG/ghdo7sKXOACv+cLIEQCewbq
ygVhhivH+4pukF4oPjoAa5McYvnTkJ943/ZxKkpqCtq8D/6NYKWsQyPMMPlaCGnu
UR+8vHFqzhizgRecWZrcxHacSfd4aaMTvNPE4NwmT//C5ILY1UbJ0wix33Q67a1s
jBmdgHshMslyv3p54siOG33fFT8sT6U/ttEGT1oNcZu8Nb2T/jmD8B+aX7AQmz0R
ckrRaff9RKnkXua+1dEMiaJ1lI7Grg6UIjpmMeH8Tk1IXvlDjKeH22eUOM/i6C6T
ZCbb18rT2g+uo8SCr/rpEGYqYv+9wv43MDEtsilWq2wOD5n2MaH195myUlvVcIXI
CExi1IHcoWAO/IalelDyTfY6Kzu2F8B7pZBKOm+V6Jfm0tIea+qWADRdvA/sjBIu
3xTCW0BjleevcWk4IvT/gvTHLisgm54W4XEHdTC9VfDkQR8V/y1utYEXm0QkXcDw
94jmZlGsYunsq7wgCsfC8FYfTwoL6VHDevmVKLLuStSyQbR8b3Uqsc+kmn0hOfYp
XQxpE4ozCgGRpWBmFxv1IEiePbWnn5x7s8yYI3qjYAWjsBPJCMJ5u4pSMaKM+k/D
h6YCvuqjpGkfSHt63hf+XnU2uPdR96PLw+wMzYdtq4GwJuzKjrxXrAVQCotRBFTm
/R0z2r5jfMCX+Dt2LFc+t0OfO6JUKC215KCQzwBF0HjmotSiY98M0DeKagyaqSkU
98S31bmhKYbuvOZHeHQ1C9/kBouSz/wm4NMvEaAToPZuQbnmkMbkgEbwa0C7PUQH
bSy4Quo67vkzwcBNCSaYNskj3xy2tsKIEUhsXcUyWCiewHUHOH34aY7rTMOWFlcv
LwuaKuV2ZnGR5EEo38C6QX7x6Wu4HrTaLUjeAsN9Zqu2HYG2YhpzukIhT+1Chuf7
KOEMnS9rIo0mbA8/Yv8/ycMKKfF/ZTxrsLnvGeJBaFxIvsa6v1+dD3ZMij3yda5X
w7wMXkBkfJKk7sX0O7X90Im+T0WMdWBjrHjup0kX9g1SrVLxxsh+qYe9Gm2coo2V
oPRcG187ChakbUZbYkEzVPlOlEHYDoJLiVZ5dEANeijkqWNylD0VjfJbH/yONRYB
39t9J5FmrhabeNIC9M/raFKhA/h3viUAZ70axDQjvQz9wcVpBAGL1y3ex6DDG9pW
VLFfbFpJMGE2GD5GqVt+OI3eZS5S1+5lJTM6M541RGTn98Deiu4ac/RoULuNs9L/
x0Qboz+jDcKr84BVogC9ghPRYtzxv76+V/Dk1R7RXEkux22S9ljveJj6nP8ZsaAK
D0k3a64Cb734JGYzgpXPRqcp/he+4J6o0F6ZHAEjAIgd8yCN6/rIVUUrCFg3r22k
s3wjuzZ6mpL+t/1JkjfR41dtkTRIIRncbeTkatOgvYTmuIGr7QBriE9lBokdoWyt
mSyBKS32+J4DQkjufDx2rzlZ/JTAiPB/V19WqL1GsjQQlpXk0qDtm1V1PLOb9ngS
/E3vF1Bkkqo4T83Rpv9fONgZg7a8Gt+3abKMGPTEWQlMsmWQPSlKGo8QfnLJtyYZ
S2i+pjTtzIGu6PoTGgwT6GTRyONy4Dh7ObPb5xho6izx4A7Tp4Tqm/GE4zLVOAvj
KwP/NAcFIShcBDz+fztRs/qskYcjAbx85jWSSiTbpXYuAzkUrSsfB86hReEuHa3g
G781IkmTtTdLgRV2f2Ibz0n388ikXwyPLWBV4CTEVE4baw6bFwSe4iwJHgAzInju
3C/3d03D8Sx/mwHwCvnf/NyotdAptReO6kh8GhhGnoX7uBMsXYwwoB0k5RvQYNEU
L1Np+vpqXBNDHtANfrXs+9f99ALIvzF4DzWgKbY5cs5DDpqjJ5UyE/aDrmUH6IXM
mwYGLwqXS6emJpkzQObCqV3My1WOioWwpOXwlcP7aaQxTuxQ0D0nIr9msCt0vT1C
NBvwdOcckizRa4EbK1VnrWiLDMmUnMDmrmYi9LPAZgdXEXCWmwxv+OIILD0i47Rs
m41wQN4ch52wnit3MivbHleH48E3BJV2F2oLdomlR4zwT6ZihW32m5hbaXEIlPhY
3LT3gqyhixeM2ZdWi/atv4mr+pRiv4i6Vgb7/cqfdvIZCq3VlqCsSnhLqssld4Wk
/6WUQ3tHUG8iGWysPZF+pVls9AgSEqkN9i3VO47sVwvN75TfKHeeZ5IisvAygJsn
yG7dhtZdr9mylN7akHvq0rOt2ap7Vcz6iPdgL4Ep+cJcoyx3uPoPcmRBOao2zpqz
DN9xFB+qxiVj6HjYSostMM0O23rWBvA/pR7BFwznCv/QbnkhK04uFY0coJraMX4z
SOINN74jBf9d+J+AiRCVyErRAHQtKbPdm/p5TflEPQYC7gYDk3hfLv4h2mNDzZa1
5n/sslg28yo2gSuLYMRn+G+kgzECH9j90PD5d3knvHQ+MWEvpCFoS0Pr1qFcDg48
FX5/6mUJbgCrZ9yy8Mhz7ixxE6MSNO5BVpqrR7FkChKCRnZSGL/UlHTm6r2JJMA7
1yTOi3wfrlPHPI6GG1Vndw8Lxc6aembwralZh+rHaN2YUlWC8lH0cyOnzIdoxS2+
HnIBPg9XCm9MUbj3AU9OcTVK/jquYbq5pZSWamd5oF4MpWdsTg9VICcmRxhXalUn
s7uUbH2lKQ5Ij0E0VMwuIUIGvQtV47EjGalK8GDTeIZZ9mu9ocmrhSjHsAqqNsp2
PFDY5BhM6wawgtd4wcWeHKHQLAbOi2pcggjh27kcXjhJ0y6xEiwmvyy3eB9D4be8
GyQNkwQABcneqhyyYImtZL0InF6w+XKX8uBSyY5kjHCwp/6uckbxIEj5o9+2t1wG
CYva+ADAUFMDHJOdwcm1Q6w4SjxdcC9Zm4fIp7YEColONZW08kb/sXV4Haykjsfa
Oi/n0IpsUVLwho2m7n4eIcNvBrbprJXqpYRr1wpK3peVh9StB5bULcT6rXeK9+t6
54HN+gst0nplOuVEqoZEfWaj369oN9K1qDQ5gZ91JnQXZWNFAhLBkIIlISMAh2EZ
Iku43FksS/wDXsLFgW34YG+SZ60IcFYvRTJoSz0I/7M4kNtmwxsnROtD4rJ6S/RQ
G8wrtG5r6aUDWWdzK3PZJUkhsHQbma/4BzvE8m2BQHxeXKGSu9il1cqwheI//1a2
337XTZXbPh9s+b9QfD1fD1b5u8+Pvvww4bE3y4BJ4ilke0MSiwF3jn3+XpYaN2E8
m9ZOXsaePdaBLbF0kt+Mi67CuL4GOKRXuLok0CCIrDKA+G6QyQXXJguFZHJ/GWCH
SxDYg6gq1n86bmMFD1npnJBNs9nTTKTRPVZHE8FFhIVRnuOnzDSXv1gmrSSG3CjP
dMsdzUz7HI78zmyD8VEdqIswNT8Uv4kNA7ucK0MShHVmvjm5FmpTCYkLGu+Uzjxd
PC1zuxzwSic601XVeUCblp7WWAaBmCxZdoFXAqXobb/36B83cQzVInm2Jj2xmoz8
yuL36JyEvIyvI2RRk3bUU9bJ2XrVSSzgv+ayTY13Kd+45BEgJLAb1P2G95O612WW
xP9lEiDdDijWvgxpmwX5k62PpjOnAAybQn23SLUPqq3RuPrGn4H1WrqdTW9sxBud
PdbbzbgKBhDISwlk3fevL6+7aZIp3tE/Xr0cXUP4e+MM4qNT2cYb6LQDYv2va9bt
jX1tntF77Tf+9K587C+6+ket9ddiygBQZBwBpJ90OIar9IqCJZhaVAZQq+GqKmeV
V9ovTEET9u0aY+5iemWVvF4XcT2q7+NreMZUvBntNHHiv2Jj+jiAwYBdW6WIqjDW
o4FGruO5XxI924sbHZTWG3IP+4W5BTVebE5mj32qHHvavZkSB9vatMev85k7Kjli
K3VB+d9JLVbvpf9wDy65JMz3/DrO3/Z6QQBb/akcjHHzmJQOGWb5BoBYK5BsdQIR
qwVZAtNf4CNLNfEcb5GRL+klBzGDJ545C18EDQGUfKJ+T4SF7/qJkoWxa5SX+D5l
YHbW2nxw5u/zRJfKbrvlu6mLcRGFSdYaigCN2VLzpoKQa8pPuRR/aKKoUIooq8FD
kkq8wAWEasb+VOTPgbvgjgHAbmL/p47Izk7oA8puP4BR0fl2F2/ADonSyyrziKmr
CmpweAyUzheMh+e9GoomQdkPx9/uMqRm9COe3umQkW1JazaBPQY8An4qKW69qhjs
ZmmILrfQ1+AyCpid/8AcJM6xAvvxIJNTs1tSYHnZDIaSGwGgwJ6cE0ywMojd154m
pJ9+s485aWitFtRDqXAoSi9HQskA17w3QruZFApikhX2iFCclqwqdOP2HUtepHiL
4UBPqZOcA9bjnS15wRaLU1i3Y0JYchArHmt83s3oXlpWAWg9SrdiocSAtG70e14H
oCgypLpiY96iCt1DiUPv4D8rMMumFwV3suGqzZpy+5ox1tDSuHME4O0nBYtGd/Qr
A/6BXtKX4E1caVcBODt7ffNdmzKZ1vYh0ZVqvA5LEXZnrzzK0Pa187N7M0T0MaON
kN+sNg2RIxZ5/B4zWt958LgR8ZY+MTaOMc2AYRQHdOgMJCKUciVjHC5CYinVzC+d
jr9g5AXMBzR9xUCL4LWAScZw43k2yoa5vTE6oG5oyNiyJLkY5MGq9I1fEo5cWbll
HSNAvb96PsxJ1tk2JwGxj7QecFLNegyW2b/aDnH5sBUtxYyJkCYwh6eNzOPz+bvx
jtVZdYqaVSf8c+zP8lFvfZrNfkWdu0w+TGxn2f4KrWWHRPQAU+ZO3fZxMyNDsc5m
o0faxAcf9s7NGrQhnJnkxNvxEdP/wASNX5fRhWWR7K4BplxmzK0c09kp8GWxrwvD
wzv5a6DCqqNHaeTjPSXVd9Os3IyejIjjXQ3dC9LOk3kflEvL3mHxDjYqnVPDh1yC
Q3rhWNUdPY/edl/LHPp1AJGHCDbKiWXFio/hAOZOubVSmHb32dNEYZOKaJGxUjkv
OwIMcdnQMlq3QkPO05bk1uU88Vf/LdqO5xbQGaxhY0LrvoqcYJFYlkNaCv7ezMjT
VVmroS698v2om4sdZ1YEaWcD2lSz7VHucwRL6vuSwvKK2/dhVagrZxVdO35muR+g
6esaO2i+ZtHDSX5yae73sEz41uJQtaPUepeXcFojRSx6qGx/WqMoD78ueXkTqVLd
s3pYV4tqQngdhl4CNivgM+EKnwVUbYGIthrXwZqlfRPHKTiOmgA2e0eFY34WRTAZ
Ovr8/rTMOB/F0kYTDCjrWblCZ6ZhBRMjfnJb6Tv+eilQFWUPIy8YP2UqQIt67AmD
WYn8Cw5axUCgv0/gIetjtf4AnzWzMY9x2LOETh/aBh1Bzgmq+XNNh6RUtTaWgz78
c58vPGLDfAJsATM5X3b5iTrlzOR2VjqY3saUr9NpL1K9zip9LjPKuI7b4WJqq/jo
Kn6+TlU0BmAgTtHqqIbKnl0mKxcuMv2t5P8p9/SJYZGbna3SENcSOHuRQVOM+Fgl
Ss1fOCH8tgDgbLuioRvnrgqhF5v2NQuu9dDy+IoG/aLgzAg4uI4nn02k6yh7yYlg
pxsBJI8TDeFaeLlFe2amXUycU+UpG+oyYkQqnK6crNL4aVfi7v904bu/g07eDk23
8oIz1IU/xPgBIvrguHjo/R3u7C7XS7OnVlglU5gmrNWCZhmZep8CUnmto8MxlHrL
Cl9t8xkXbUGIQrc7NkRbLHuveM4d6xK829VF7NlwAuMfmyLg6gx2C/Tduwz4JGSn
uvfVXzdSs1mEOFI6QyNeNM9snvFCPEFPY5ghOQXa80w8s4kndc4+XpRMBAse/52K
C9DcgYwjuQNMOq/stRC+w+vprlhZtOqOJRa0RLdEcAODpVRw4l6wh0gsYlItmT8X
0dcfC5CwBhI3FGNMQDxszOJLR3GftmGwysJ7+rTY+Pho9YVIi+3OXQvrKZzN4hyF
Rbx1msGwZHDJTU8Zr+NyybHzdvNZGZOT6FuQ3Tras2Bv1hw9chBhl3i73x1lmU/D
cYYMlokBtCcUQZAG3xYry8MW8aXupc4kNV3ID/BLRuUkzDoUou4+YRTHqrPYDs7V
u71+oFWTMfudER0xh9cxQMdAMTu1TqI6P2ufWCVFXvxwhsV6FkW864a9yvbZz8OF
VHO5WbeD+Ouqvg1+Z4YlvHABTwRcDgZmelQfEzhO4ctjlV1REDYF9780Ivr6gRoG
oSE0Ojv92gn7aUhI19x1sIlz9RCyCctaVhlGEEQ/SKJ1cY902x2PQepR3LTPTAUL
ZI+CLlwZH11eNUKxjYrFIuk3etU97ilDFWBrLOKwYmeydaM07f6Cl4Kl50u32fHK
/fm2stlD9BziUP49zMun8uIVe9EJ1UxnZeb8/FaJ3inrL+KOHklSLMnU6+7oaNJ+
NN/0m2VleNnePdI+WA10V5PDOzmr8eVXnrwmrWKkNAiYcXXFtbk5gFQ01NP6f2NM
A3XtN37Tb6yFd06Z4sTLcyXLvK5vRalF5lhaYS6Nf5AKKhOsqXTDoWFxRjEARQcX
EjSIm6SmdbZBqb5gz/E6AJJrvaImV2XEQ4Q2eewKhP0zVyyL0M8nFeCxQhOuTA1/
3vcPpc10yj4cYfwQvDiIqrTrjgttUORiSzreneuMEHHhU+6wKX5ci6h0OoRCjgHP
PRuUnt8Qqj5+XW3cOI0EK8JZBdrypTSnYJoTH0mlY4MzlSR4EDCh4qS8ncb1GWA/
2AXGgZQZYkTOOcnz00zgjsUwuIo9wWktqsIH+u2VTfsUfipSfLktaBZt4aD/Gu0v
30JRWTFIDSSIJM1hhapqHwyKBzhgcgeth3t3BTGEmOj3tRaj8kGLzYloBY5WGUZT
JTbldQQaOuZD4l5u7oTsuuqcjq6CBp6pdwzelWfH41v6tnOHrKZWiGI9Sxj4/Y3S
2jjFtTod2sorOHM6ahMMxfJHJqhZlkvcBus+sCX7RNdymPknTPUql62ztGqkwTlV
q2TO3ZrHXQ2nSKYmtU28mwCZbZIyLPlZyw0kYWo4LDT6QLsHb7EW7c6u0wq7llSy
9Mhi5aGxkBGu81p1S85PAH5YCEsqWnSkc9sLS/MgC25ckpGVjfAhwyoyTpqy+Dx2
7uoDvNA8wMDTxO+BZhcBKB6fJUpz9Md+7SwWmr1FZMPo2Vq6+EZfQk4xcwmiWohc
hSE15xiOwCgmlwCgu1nUHym9uYg5/bCV1thGi9opXpXNhvy8tDMTiwqNvAqRSkkg
yrv7HPD+PTBocqqL1RxRiKR5nqLqKMy5tfFRrslKWeWXyovDP6d0MGwxRuhMmXZG
tHzBlrYlumkjGyWZeQB3j8zjRNlerZbiewM36sjeVRhXkt+XesMZpNPbrKsiTrEy
mMlVfapLzYBCildl2jIehTg0MuPQHoscSbh34QsIveIrUTuA+hJji7OSREuec3+d
gr6k+yu3EhSfCVm1rCPRRXVYwgVmSRCSuotAtKGibOKLRPdwAoxdulDiwJGvp/oY
CP/ro6wwFWC4E0xOf16fZ6IU5/WJBCrLUZAAsov63FjYU9MN/0XCVHgRoC3OAsxv
AFsc1wlSQ2zJls9DKHzz3W+WrgXB7IJCAgNue057MbO3KdVBK7uMblpN1BkN68xP
Cuz8V1Beo8ecXNWkBacthajOQRK4rdnXwuhOJDkBpFaxNO3BN2nH2bYSv3czpOom
/y/3d7EjA+GurGYU4ojOrKpFd1+7C8yE3x2T6vYjk/FzKLktTRXblK7IeI9FpXqC
tv6qjlfipTiYTPW5OqRgrUgTgDHPMIG7BAOCz22yw3s6JI9fvkXbVf9TD8mCKVtb
oyxZDM7CIeJJJhXxCq4xFh8pjPrFMCRnvGt3yx2gb8FB5SkAKerFVFpjaxqB8CUF
aZkjYsCF8588HQ/ZMtb0XJTknnpqXF8UHaWuzkvLSsXrbM/NrJ1UDgT2l+eVrWDE
2nUTFENQe7zqn5fWIDr6v6IXPOAlWL77148zxeZbK3DdBQwk3fgs31M7T4Nm+WhE
pLZfVqGXp9YJ7Rd7nkEQmmResBEuZ0EGHEYSxlprdghoOoVSB1SfMZOOfo5D3KKA
1X2dfRVnFBxW7UHW9Xl7Z/ei++/K1T8YcwnyhNdcb6wG1R0hLGJipgxs+0eA/v8U
wFWQBTk9kQpma5ZtuUPigZBydGkUyMwbH5kunFSip47K9hB12cHnQjvimCQtnEmz
YoSVadi8CRhE0lN4Wk8YkrvXEML9cpC4MUcvOCJOethFcsypHSyhVvp+thtj6ExM
Zv5+XBo7FRRcdjYGLZS3BiY5RzlDbwPpQo6NuieyCGl6VEwJ+YIZ8HabRKd3Q4eX
ISu7kOZOVjbxPF4JtMG42JWCkDC8Mt5SshxjlmIs+kLaNZRibn4LC0NwSRYeJUOc
bT+7xpXW4nRUGTAENFVSp/M23ROO+EfTXM+yuvtS022hhQrM6KH8p8Wv90HomMYj
Qh1PuRpqm4fcV8s2PRUrwAt924vZHjUEaIiUQHQmq39vchuSDkYfyzIsDeZBHvpP
d6h7eucP/GUJ6aTeEjDuL60+ZK5q3PXWNaD1Z9TqnIgVY4sbrXW+3vbvq1qn/8QK
NV0X7NIY5VfKaKOBPEruNCYRpJqEEuw4fyM0QmkgLRXmOPno8hoT/A4OKklY2G29
dA92YCQjDic2L8oY55Fb29lGjXsMCZIGiVL5uQKj+zhaTlwjjdogOUGsEgFCKR36
MyLsPvNQ/G9Ife2IirEaOWn0LrO2BX7tjhOi3ZW91zKCaJ/WA7p3j50hhvH5gckC
pqGOTw9D9VCoSMlISRhar4T20JIRCiGVVwSnv5Y8NPuniD5OsZ6/N8vNT6YogAt1
HsIXumWpypiccm5jRXPuLYMUcNyQVI3AdrHNKZARQUhIRjpLs/TdMtfs79UEd133
8XWETT29IzOsahjy8aoUjCZYZezGPfYcywG5UkUKpUUGhAZ68yQWLoPBz3MyMVBb
pPfsmfa3LLJAUdE1mVDCrJCnWAcBfSubJbcWs16n+BvDoQX5fRJgAHYseSvZefdW
dSGw5xyym/vuuP8xgafN+z8lv/mMTNG0jbYwB+EcFvZy/rWzQVtNK9HqR7GaY0xZ
zYVUarE+0LwyF+mnOijUXzsqs71+Fk8hchzBK2bhzaGWP/Up1KVqp758YOIeT0Pg
a/WdPH1hQBfy9pvfYWW7Wr05lFXAJwGqvRax3/jcGKN6ROPnJaJ4GSL1yzCm9JsQ
22qf5nQA2LIlhm1VuHXoap1c6JkRaZC9qkYoVJFjXGgMgATcKotIs5qJqDSonq9n
IjRJvFW+nC3TJ87lDV56U8Tti68HSwsWQPZkhsJy7d/5HTDpTp5UEvIiIUNCQErc
htvaEzzfrBB+jR3vrfzRJSHxgsqu4a8V+bdwsWhTL2G+wkzk9YMuu6LW3Ji6/CjD
Qzg51C0NGL70imZdMBXoyw5lvYI7YDsQfTYBY11yNNfX3NCB/WLGz/1264DNkT0W
JiU8YvlvOUIusWOc+Fqo/j/sKmWK6WaCdauFpj7tJB26trs0neLYz7HrJLsQw/mr
ozdIt43+N3yLnTiYUz9NMd211yw3ir8MM9ABcwhYqAW/LYb3H+pW92AwMRTrtcY7
ffeEP+v0PilA+mj6Fd9avmRNJ06H6CMeUsQPVptD87+zdLFEiOQxk6D4G7lmjQPS
iTpu9lbdZgdBTYySdQFwZNhtBfqa1BAj928x+QFnoBnTTTEenAwcLoYwCKRzgvSP
XWyM77gPZgfj68PQoRkO73Vq0qJJePtfi4mg8htvW/sBcWyzyCtKBEwY7aaCp7Mk
DiZx4Su4dfvvvqGzpeNFPTnCIA8Up66qCFF4vkIr7WyKpXxOfLBhEP9Ij9oblWSP
has0/dYHQYqyYX2yqMNjFB5MGq7F4zuPHPdqnm8LlEYca+p7bvAWsxt2Txh3VYu1
hmrl7oUpVxsUiM4Gyh0t2VcvdtNwvysNshH/0IiPVySZowZ4QW0rZ+7woMYvRlPB
t0fokeIKFEVuVBin+3fS5Q8ctlEYpUkBjTUX1ctHWOs9XNqpY5bkt8l72A5eS72S
dahLsrBRyiFxr/5cxTPFcnwPkyVr3sj5vtDBFjEwDKPBfDDi1pDaA623qbbm0fN5
uAP7cCaEPv3IX6Vcqxa76mz7sc5H2F6QjqTsPR67PF7ZFO4Dmmgy6SlDEY0JLWDi
znOlXKTPnc/EsmAlXlSoLzDaumB3c1pz0P4zwMJy1GTIbdNkqpiyjjDTp7156akv
/H9nReUrdEXmdiGsJxWWTbGAljcH1c/FmP5NjU226R6irczQz/YGpxkwAto0j2k9
6LNgLA6pm8MmvaBW+zadpls8OHTojEpsMNECyG/Qgw6tdFO0DslVPp7utCrJKK0P
cXDYvgDHTOKg/f51joLqIMAyCLYPKejBpziVlxcoEjNpav+pDFqjWGMGVMZ/Y58p
UPcbAiyBjLEE7Ey7ajBx2AqMPArx8lJbkgxDzjlavbXMJ21U2iUe0abhB+/XAN8V
yLOQU3Y3HDYWitW9pU6vqCg1vO611KVQsuZ7doF8xgFfcWqc4hscCKsTPX1twPYb
zh8KgtjD/pOuTC3BkTyhwjKw8W03Y1EPjpF0mDjyzXLOZSDLTXlKLZWd2xm0bN2J
tqyOxiginp/a44vw1OJb4iT8JlB+gwvO+UGw2ONTOFDy6rX3nP0CucUkJEMW4tP3
42aa0+cutS+jXWKyQHmUzcZQULHo1+wmypHz8NQhgji+TFBYKnrPcfQ24U6smY0Z
r6IF6wSD5TS7ocqlmrrk/+Moh1irV8B8cLnXLvtrTfomz0S7x3px3+ubn8E6BjR3
SM/hcOgCBMvYkcQHVB3fYH1zoovAFThYjYDTOm6NKRv2LhwIzYNpelY/fK74okSY
6lYbhHbjUExDNsz+iCt97wAq6bPnDn4S2iqbsH5LVf1ZXTcRb8QS+6szst3fQJbZ
zQ8F+MGIsf16Ia/iHrxkAL3VVE26BSwA754/5SXpkhaJZI75hI5fath7Fr05TkYs
o0ZaNOmoWO9sX6hJ0tKRdc4rqDSS1fdcP8lpDkf2c5yETlIO6eHAvckosc1eo6jV
tu+ILK29d3DaXnz88XUDyrPOsSzi5W4v/pa3tfANlR/80sFDkJ28P4WZ/jaACDMg
i3CpKnsi2K1eLvxvWk2xw6Ida0nDBRT9V5q6PFsvfb/l50ewDyvYPC3oBNLrUr8G
RgvjQfz8TugkGwKsCLT3zoHgLyhkVMbfFx9/vkkgfqU555XtuTWRhI8LiFUQxNJ1
1ktwpjbu36niFSP/3qJgDLMywve70HwGXRPUQjUJ0sX6ubqxW1EfiT0jzIoTCoM7
asFFNKqyKZvcor/7lISo5aGzeCPyKbkVreGeFzLptRvF9cxmNVkpp96OvgqrOZbp
h/S0ODYatpoPyRJ4IRSqVKQGOdRROruHaX65Qp0i/NtekFWsYnzE5np6ZRt5Mf0Q
7WuJ3jVSKFBnl5/7p+bBblGFkxfYqYG95tjumtqkD4Bt1Qcg0mYTIkue42vtpioe
o9pnYZaPmHr3AfK9PxIYZy+GxLDzN2VLBnH62lSZs3P6Bo4pdIa+agw+Jy9ajsEg
OHmye4YnG37VAW2buefqTxakZAOBE+rOOmwMV+5CXm4VzioCd270pG2DZN/eVzxE
EHo5r6clhyh1khQiE1ugXnYUsCE4hOeF2JAorIOAutV4fy+dmNrrpDQCFFuCybaQ
QzNo4eZzengjOT6cenJ/5blZlQStaAxPwM9BqhXUFYizxnlVn+q5KBuGcpvQQJPx
DY3irervY9aNIrgiz8AjpoBbvGmLxU1LYyWFpK+y5aUk6dk8ymJqrw/L17thWrwJ
wS4K+RbiSQIqgmvjcpwOqMYqPat5AaAK+UMU0UzUXBP3aZzLPGBAr9ZSe9swFvaY
Z2v7d9f1LMBkIrox7AJRXp6aGEUZTzjeLGglppPJvL0Rp0aRH7fy0OQ/sEPuV7rB
0kc2orxslmnUk+8XCmwLb/evuNRPe7Rt2pSUeYWrvstmoz/J6ipPJGXJzEuwIj3X
rjcBBCi7Duj2Go8swzwIPXqiVStOdXjQmP2e98alMrJ5J25SNL7XFF+PQH6SKDQB
eXStU/9xUeb13CMb3Bf7thC25rGdbFSxbHiBppWgO78eiWzboTVlk2jZlY7DhXCk
5LmCdDIdK53ocm9JRseqJEKXIArnEvK+GBOjYs2WVLBIAXMxNjT2ERIkFHPXFt7b
n4qh6rn95zC0BzZilsnuuoI5D/GC4JWt5s1alJEMS86dNvXvURvdUVDbDIAl4uup
SK6TRXOURtIBmcx+2oec1JlLoca3ABJt7QHGQ0wrgw5fvM1QDPbYYRz9dh2xXq3d
SCfkuw9edWrl5lZMB1EybUrGNmW2bWNGCAX3q9IrlZslkGHOyP8s5ynd3+Nbe51I
J/yMs1G2kLOQSsrzrsnjQOFjMgepOWfyedzobpjkAvr2gR+RPobt1k31jnr0sXZ9
n55REmOHhXsx5qRgWe7p7XnnhWu6anYCXuoxhjE0JMatjbIElgIDvz25nfXGi6P9
73ZX49WIc/Wyfluefr0BWnv80T9Ru74nC0otQL5IqYpfHYcwS9ytvx7b+EcFwZKZ
ZGKwJcfEIaW0k8vMYeBT9of5lUIf5viFs6sqtdpFnzrcaTQdlZHJxnudwqLUrz1Z
ttoqQNmLftHcwzl+e4MsgCzyojjz67Sdw/JpoEOD8R7eTqXxgiizXISjhBlt0ut2
txI63aDnfQRAykVWTpYDWhqL9tnMM92Kmk9xkj7aJm1Bt3I1EyObFiDaQLoFW8qo
7D5qma1BRpjkDU3kYofPE3l9FHRtrSINsUqUjS90V0bmucwHmo5/w8OBDsmQjpZV
XFav71FIbAfM64TToKXwPTHyf5stiQW/rweyZpC1uMZ3G5gslNL1N54zxDpMa1Sm
MXVjsNTbxXUywRUU1zDcm7ESiRKHvzKk+g/y7/E3fgocEyIdNKLGzxxxFzR5tEm7
ooZTh/2c5e7nGWZo6DdZYNMnAtbTHC+KJA1J0pbbSHUMbjXnCBnz4i1VeinhB+qS
Y+Bc21LSqnIId88PjMhri2oWkIjdSq8x6QKhkGtmUOxIvb8D9Wk2SCTW4rRIGGKG
2N/m/niqW+VCObWHmPzhuK/e+jBZIKQ7gOUlSV1Ni11B//XugLuqAhY9GchEWlJP
ylFS7ByyK/9K6d4bTJ1Qjy5cvyE18uDDOXQdKO3fgtmaD7ygu/rk/obB9cya7DiT
BqOraJV0k071ReWdXp2ptK9q5BBTkj4g33ftLZhH7HBKRZBIHx5JZtO2IqocJOB/
almjbjeMCJmNJCXZC6svBfqrp2wC9v6FUpOSWofLGaPR2t+iKN9vLpqqEN2mMpVn
p7lk8v75GSEAo/uJvosk06ObgCfVO44dcuK1XWox7eYiRJI3XP9ZPjgk0z/Jfhrw
hG1eAqV4DYGiHSQR6ihWZSfwmwbx+9Yzw/izxk8AcGyEHOg9P+FwBtvKpsRrxJQW
61gu6dq1NWgMVZedGSG+ZfT40FTzdwyGhMJb/j+dANnaGBlMLZWxyrszcpgItPT0
dKngeFB/5WmdzClopcny71p71vPnfF4VmQXzfm7zSlyt/xLEeOUo11/jfrOiQ+uR
+0ryLu+opTPOSChYtzdcGO4kNRLVK2o5rxmTF8utUNheqM+VwIKYU7W7UQdyWynQ
EKzADLbh7jWPknSN1IyDeT4AVf0L+wJ2WXMAoDQ5KIUJntoo08UWun3o7tNu3ChM
GB6nT/3KX7ERX0uMpckoHhNxSa8TMsUcUrgQog+KOcY/6qr673LecaSAyzJ7qevT
SnlfMKP3LLOGggFJS6LovB90KGkEfdbtlw+fbbiQGiUTDHWdF/bRrVPR/2aDN3o7
ni5ict36/iDOyhaxpzNJRx/YDpOBt0thzeqRIqPmXJf/SBWludCNJvrRlCi4zyR9
`protect END_PROTECTED
