`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gI1LMDRshg73n7W9QatHuTMkcGKat0685TCd5es/l4IrRD4iqS0gxVwfkVyoZR9
QuqcoDt6X7Qsiypj4lC5HyTQVTkdOOOpuJB+s+m0B/3wnMF1/yG5Rk0+ezPOOvjA
44mSdNMsuA7D2CGU6HSn9lVhfwe7ixIWg8J33PyziIrSbcjoOE5tvM2mlHfINHfy
3Jk5bvIwUUz3KmlB06wIpE6YOUHixAxggMea9Gk7fq8YMFwAwPI2jRVcTia6ATOI
F63zm553FZCFNcqKbzr/jhTkE8Xn68AYOf9nBZoi6meg79tOL+ftzFEUAv8eRPb8
iulEi42QettTsC4MTIYS9f5tU7yEUbBw0prgl4Hu0eTOgyl/gMG26GuFOWOpoOvi
hwSa8TrfsbWo+NWWUG8oix7ZotGwhzWCItZbcKZGyGeFRNyrQ1V0nvigu8DbeOWB
0oI+o23TR1HclodWLWyntdtC/xJFmmPNmBp2Ulo+K4AlFEPKGE2s6zVo/IwU4CXD
p6SCC6j1oM7GsfxtS3CfGBXF+Azx1FmGdn1abeTBPlwxf5ocs9B62c+Vkh+sjiq5
SOssWQgok36awcq26EEWNqchsm4vYLVteADK0xT4R0QakyYRsTjcbJwJjUNVWVRH
KX/gPlvAhKREld4ZAC1BEmQtoIe7+4s2VRm1EAVkE8UMH++RyIuxoVHDgWP0yFE4
2ob57KR64YHomVCN3rguZnkqpL94sv4A42GDTiJmEWxiD0urEEwr+pylh0dWddd+
HbrXWFoFgHOuSGO94PzwUqmsn2gIbW1nRBlhE1gNe1x5FrA/rLUYd879DrUXEVj5
EPIcUK1QIUE2d18JIi0nmCFUmjHQWnO+/kcpU5oY1aBQTVUtVI3Nuv/2OLKTvocm
sqkzRxSXxKs6B7T9tL55V60KFs+neLfdnRZFXSlKwSb/ZohHKgMcC9rwoNNZOu/z
ptzynsHl6W2vphzk9GpJtsCKaFAM/mCYOn86TX3IZPyU2kdhSzgAs5pdNkkeVrAU
DdaifoK+RSkAbfKE+qJhfe9CWQjkNfNlek8M1HtREV0FISYsrTuvj15lJ4yl1u/l
Id3AaKG5rdFir+mMQ4Dvpug4cAM5pKvrtJQW+9npNEUbAnCQalhZVFoZ+1b2Oeuh
hJl4PTZkGY10gPO9kHOJdxFRIdHmNeOWvg6cWy41cp5S6VBUlfWF/Q+518kqJ/By
/y+AVTgYcSA9h4EbSp8osD7kv+HobKDFpKdXl/PsjiDeqsaE5CmjrmFQRanOTRnn
GQVJGYZNYA+9+ESgXbXYSyqxupG9Ys5dhrM8IX6Id7vBGKUzo37f9frDk7YkA+eu
OEgDi/geeOk8PqI5ORU7pWgw6HHMR6+RoBj8KOaX2nTWUCE4KpY7R/TgFydAIu8P
ffAlU+DENWuoFSBJwuvFdT46N/KbHpO1p/XH2eWIrUtvipO6ADNQ/9MY8V8sykWY
KltkfhGyNkxq54O36wPUfMCE/Kr5M4UvpBx++hNSbqqYhmO/iJ5zGT8Se1VCv/je
qrEmDJ+PnEb8RcWHd3rUYxu+4iZmdiaNnOvDGUIccc9JREfNpWAtHXyPH8vsmBpL
RTOZmgitcN78RcOFA/LIgQg+LME1bWh+hhCYVXTt26VJZj/tG4OGNKM2UrR0OkmX
2JgOsXMzWyx0qoP0Sg1dxQ1WuibL4JlNpekeuEO6MM1a8wb31R/ZVKGlTGu9K1SK
oaBHPAHwJrifyS8crL4jDk9vFcFfmKs88z1lGUXKsy9pZ9IWlrHDxRgnAFTywjGk
k/6VoylRk0eg7ol/IPAkMysMjs8fmMZO2nPZuX1Mn+IqHhWuO9jecoWVUoOZ3TrE
760nwSFBRAasSX9/m7DPej3dPxwF/1LzdifMs4uIkj5MdJ79/WTsyRLQkBUyRZtM
OPjyaWztCbS+l1RLgxih+fP00aLmvFjZtFpp1ZH+87rYOHUDhluPeqx8ZXG/FBcY
QCeIkR8CIQr5c+jNuog5Ao16bFV6Wxf6lJaetf6+k3dqMW3rFm1hIMznYgacCw4+
4Bq8jbVcPYNQl9+AGPDzMlMJqi5v883zHLC2zRH8x/rOnF5Teksh4yHXgtEuFQkK
JRC0KxhtJq/f1jgqaJS8pmMgNUx5ltFPNzpf0bB+/97EeM/ndoZB2OoE6p/mbCZQ
Y57Tgq5tzTQc8UEP7KJwa0myl1eW6Rw4ADnVLsUbJ946gD9xcx4ZIDd5uLnfO1SX
qF0g7KowJ6FFYvzkOUwAn+etT3PB5Sp76hLSqJrpUcK5kkCxwf7aTbiwiidks9UJ
mQ9fYUa2Rk9dIgQNao0l+Y03E+eFiRMxHHwwGAH/1BouQ7OjjXBjcCqfa9Esgm9f
KQ+OtYwS1yY6G5T+qDVKA6zPxiDScHqENlaQfsFxtUNVf4CrdJRuiA99H8rJlvUB
aYFD/kd3/IEtyliOpZ7nKTENZN7NVIzu+C2EJPSuhKwOCimVSEtjxbFraLEhH8s7
ZdxFyZZEifhtngLyYynMaYSJobMQ93NbtOb8TDHpwMzC31OG1Uhfa5Cxsq5xAjQ+
oiDiygj8Pd2vmBXp9w2Pqi06BX0SA8IkiQ7rkg8l3FKN3rNjUL50OEHDW8Ev/jTY
IjS+71q7sSP3lLe7yE3RqoEacrSMh3TPx/qMg2+0sfpIBHDlgkjklx1Vrt/8cuL5
E8r+DascmXlKK8HQ75v6HczwNzvhaqeIGpXHneOARuzIvNmw7QTzz9L5z/I2y8HE
AUEojKc1KwQWwYbxazbD5tMCr/tPErmuoheIrQC0CIsWHQ27Cuh11E/Tv+CffKI2
i7T8MS0aCftAdNatPndpTklWqfvlzczHmWtIPMemDdt1UtVPousq5hpWbSU61Q9V
h2INaPCWDAG8qhhFTx3O9p1D/5mfrPCx/83V5y4iDe9YgMeDDpfvVl7c3Z4k5Az5
L0G3UZqjhA9czLrGyBC4YAcR5rXEwE+Cvsnu71Cl7x+c6pzKWbBdSxAohNPkv4d3
mktEf0qSwxCpiX+IDlECZJ5OG0MbumesOLpv1dxqxY72VCOIQTP3eLq7aBKfirZ0
CIgiL3GVLrrnvEGrf4irec/h/pB9JquL7DSocEiIokt9Sg5lRlxTCU0RCcN/TMeg
Ka7QyfPPmormZoadziXYGXEcyanhKa07/gcwFnLLzj0DtCSshj2q5DJ6MkIE07A0
DjDSBRlAvdbZaBnMCII+CJsZ2Gl0u+6VcojQ3SCQCpJ0f+bbjLPc3J3DATXWGyJ1
PPiPIJqFNMu9cXR+TJDo9lDZ1s9I/QGRRUjt4fAQbEXJ3ZuHXCwVWF0BLqTXew9E
jo5KYzAAJj7ECcaGUosOP55OyGpqI966SYyzUyo4YNvrP6Es23nBVRvhvJYMv/fx
C+Qyr1UuqfEoqHol9NSIv+upZxfEYH34Mx93A9piugBRaZHRDHPMIG4tmheIlSwM
XyEQvAm/KumCLCoXauCzW7/JWFQFrvmlkpuO1Amk4yAcobeP081m5AH4gCNueQPU
BmtuvU8j5wxU0zWYNxuY9iAymv7OS6dfH49CYjwk9hEvtAQ+Hv5nXok4GYRXKZxI
XK8eQhB/j2TDi7rZ0Q0mXNMYUYWJclV1LbGfH0CA/DPbDO+Jdk2njX85FtwYQrXw
aUBdg9HwGDnhufSz4C2i5f5B+mR0f/JAcJR9BZug3pUvsfEsYs46dUDsAQRC5EnS
eLE7JrERd6cPdlipizntNUxExwl0tzQuFEi6mfFmXsVc0SfguexRaCQ0opXR19qG
MQnwIBVC4Bv0t3Pj1dcrlD+rukVZC/0eQnkAihIgB4V3ssdBxpiDdjWhBkz7TPwM
Sj7YVU3mXbflaXJ5tbXyx92XEF71jn3pG1IVcQYCwyAkY3O+xJJ2DxgUbrkMXb9+
Brp/vZH5AtdI/XG6ctlj1M7zPKe7JaUdX5FNMw1ahaIZpxNB15B7fBshax4SFuYl
PCRUlwij1Ohq0vmLJfceNp6V/EEv1MiD3ERgR+ywPgLsJZ0W4DeP/5AEKhKqEf94
V/2gGNtKNxjsrvC6VKT7iS7Wmv+hPMinY/99L0jz2KdxvQqzWZGbtZu/wqY5+xJl
nGeKSZJge6ym/wXzt52qiPQ5yxLl1NUEv6BUW6fEZerzCwxDUzRDsOQKETd2FLye
5gqrJhyajhGZhGH+5F+B/sesGo/sRZnhkz/shHmIPzHgwIZLZWvaC+JA8WNfwXGo
1kb/n2sCfeCoQZA6cqTi2km1E5L8rOmN177W5HYKrFjGeHr9eyKSZse52elFE6KN
gMARkJhVva9oIVHHrlp16zBR1v3Uc35HgMiBBZ74tUOw1mvV2RUlEHQHPOMZLHHb
6jiGzTWZLAystJe1SSrd1tJ/cEV0elBtl93v4mGhMvyx00SgREkLY+LLAFVrIQWj
4DdGsYLqMceMaqWlKQZGptqoWupzZp3VcOnCYJO0JY+/BBitpUWWPzq6GfyrB52G
FPOH701wnb0ejTaQFDdPnwR1DPMMyfUFe2GRvq5XdKprKxVW4O8RV26DKdMMrBm9
v/mCo+2ADz5dIwvz5wNnmV67xuTjbJT7PFAK5FBoywrULFjmPWY0eR7ECl4zZXcj
IW7F73ZuuJtHXMFpT+Gh+qGih5jzIiMNUbgjl/2o7/LeJhK4Mb2FzyBsubP1k6kQ
C3fCQxKUjSRfR89pq6y5mmj7gNNJt/NmcSCYVM3oGdwDruJPQr02U6jY8voUxy4V
5VkQgw15FMM5TFwRkbn8EKXYxqwm79T6jSn3BIZIPU5aLrnyTWdqS+5bfI3butJL
qYpNbro4fgtRAst0+9gtuvB1Ifz5LYqGIB+g/PLFRK4QnYUYsTSH6Q7mO9SkWZHM
uxXWUIBF0gQIIPxColEYa4AUDemQAbnzsOD16dVTqpA0Yfityz4gN+pT69F3bihQ
FR3Ao7MmQ/aqsWTtT6GhxLDbGbMXmXMrfefNJdzE2CKFmMRanH5BBFXisaT5aVyZ
Wk6owT8jb1wjqtVnSpKdZQlY4wAXR53vo/8edlE7HE41i/imWO3x8Kb13TQlbsa5
ub862BSeUy6FGvfgsmWxomuslgttPhRwfYD9p+YaP0NLClok9uQapX3PRyoQKauw
PuCkihMVN/JshgYvDsYzqRynmj5LN/Tr7U04v2MeVBTn/pxfVU26Epkn5MPaGWYb
UwUvXR8p3d4Vdx+dz/O5vap8+SjGnYrNZs4FBioLPNAa0+aRV/qxm+GdNN2adQ2X
1dWaOsCJwBloq8ClGUxIvZqy/AoLtZAiwVZvqLpyd3tXVrQzjP3eOAIlDSlSEJgN
mNq71YSBGowazCVET0d3c0fIvIw2Pib93OBGu3ABkWNVgMbu7chbtW1xCA2vcMI/
GURoFbUwuZaTpzlacz/fb2vF+PXh3wkNi5k8a+De3gAR29SaRwDG0QHPY3AHWZul
jsxN6TCQuQpxfrIZji1FKiHyN8jlvZt7oJ/Ch+B5s/QS70436Qmzszhz2nsnlr68
`protect END_PROTECTED
