`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+OVu5QkLucQ51N41uh8y3UiQrGomMXR5J1MjeYutdfV+CL4hINYeQ5cKYYam8BdS
Q/Vcp6Ny66OM0sF/i4OXQxvgDmZEi5fylquqs5J3LIcmQyIB0yPRHKicCdaLhPVW
neJ58VA9ekRVMI17fXW/eOPlCHfJKebCFj4Nvb6Cmc8Rxcz8+RIXzkqXvq3drzdW
9ILvVC8jIXC1mZgtdeXfTDiA+AZTCdUXIMLMViRYMKSDaeNbAXX9h1GbwIvWKhCT
iMtf8tpk6htvqenu4fKYmWVM4mgVS813LTpb2HSo0Cz7m4cOb/c2gzYFhuYSxen7
Fic+4rT6ixI81Ar0oHBobs4zmtaOIFBsyun36gIQyaiZ/GSA+eFwekivj41iY9PB
1CnLBcaLnpx6j6d8tbTTZ1KgbFxgusKXpMewXMFOYxHsmc3phHig8duv29PmWE49
1OnLjOrJzpOYM4SztMQKC1GEZg/4hqbUHmWJR+pOd3tbYDbKYeoLLHf97Pbn+4bQ
a24kNtvsjs/z2GaIVbynP2mTjMgEf0bOEuKYn2iMl37WFDLRZ+PpS0plS5Rdb324
IhQe066jVt/CG6y1ePOYTg==
`protect END_PROTECTED
