`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0slxHwJvmDgfJ3txPe5czTgoZ2U7+aPpPsPBdUpoEE9R+2o6Gy7etBVcF5DUh6L
jLEdlVsTrI5H/1Ga04StYciEbfladf9/Cjrevi/tRBNP0zN4bpgvWXMGnkKLE/YV
IT3BUKUY9rGKKZ5YnLr/XR+K0pFhJOk78t4iE91tFR6y9QZkERVPrlwQU/WUVhmZ
Aby1PSSG6tP034bAs1Sm0ANwaUowXM3Jef6A+TpG8G1P9Qp7bK+FCW8ErdYJAphe
CopQGovtVYu6sJ1f1nVFY/Chll3npg3p7hbbGRhGQoTwlMK5kyH6AZqQQnuhpGsl
xvZV5QnapsQjXUuf+MJgFB0aoZR/O2ePejtJQwkiYTRMEKU1zkZmbtvtnFuH0HaS
XYs0vmzI4wlTEWURFP3F495/xDC4FwJDZiFxAXeVyKMy3dyDgxqTfFVTz9KZ9S7e
OrQWN4+0f7gV1LXAqustAuSJxXI8TQSjD097jhD2VLujd/iDGNzaabMtXxCpdNFE
VUeQwyH8ST/VK0DW0KBmi/6Q6ra1H53P4lVjmf9iX/NLybwFm3Pam3HBZdNY0BSE
Pp0HQp+LoiE7yT/9h//EoQ6H3Th5P75vIRloFwlvT9U=
`protect END_PROTECTED
