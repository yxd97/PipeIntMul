`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgMmK5gENLMhoR6ZrceBLEpQfIXJ9ivSr1taOWlx/cnvS4UUA2J0J3qtGWsK0fzg
9Mm8PXy3H3QVK69NdiQsjxPlgW8EYl4kMhv1PXOvIiTLhQJ4XlQ7hMX6KUtZ5h4c
zN3AymhCY7ASJsX9m7ZZuGmM8MO1cKKwg1awTrzSu6HgN1n5RY40NOVY6mtdTsCr
53JPvUNuO0oVmdKRSX6aHNdYY5gFJZ7vMqMK+Ugq+TQVl5rXdU4mttqpKlYBwTmW
+nye71N4FmmtgVDxXF/pyybGHjnZMIyyXjNTlCGG3+Txs2LYv37+HMXHfF7nUu35
I2Ug7pCr9BSCKMu4uag9jLfEVmCmG0Z9YWjOv8Fz71DDmNTzJ1WaQvhoraKpvQ3A
`protect END_PROTECTED
