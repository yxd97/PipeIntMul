`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ztw0gjhc/BbjQ3V3qZZJwaS8ePZUFyZU6+tLThvd1o35gaUaTp142bE+NGG08Z3n
PUjRPEqbhY4sWZdhNfkz/aq4yoTApzE2qYsxNKPKjbCrZp5oHEaFJv/FuhnXNl+J
c7BDhtyur153zws/xxUGu69XPV0eGvjtHq9Hu8//vL2NfAZ5aJsa33WzCsbq2lPj
wTocu3NRJIOCyry5+qZxDPkOaGg/CoGXPSZ72+18s14avHRNAFFllnusA2axyrjm
wD9biW2F+EJcEcJUZmpZBdrD3ft5D87nQkQj3fDXJms5i4sLaJEnbgDLfkaiRtnO
p0mSd6hzQiov18n6ropB3lFitSUOJOLWRiUQurDL/qM+VpmIzr3ehwHsZ2WJuFsT
lNelCkXA+o7IgyVvmPmvFIXKvUg9w3TlTsv1WxR3Bg7VsnuI0JHrJBI6tbFHUzPi
6UJ4uH+OVYzPenMNapUZkTfXBDMQyztGjydR/QW1qE0Kd3DbUKcX7u7nszHxmw8U
mHovcuqbxqpEtjleKNyv/gayeV4fY1WBmBDTAkP4tWqrRHMEpxpR5DCHtEZ3B6Px
wYUI75qcKJVRbimHo/il2jP2SexhKG/s0+w0gSNsg/qIvULDi5Cjv5ombB4ifGUq
7qVBOMXu9VAs8P62VFgMoubGhevoaoipJcSzN2EUac/hkHSZIuPn0IdCKTi0HZY4
gJzPPprRRXC29o4jbvThQfWKBevZ227PuolRbUOD3vmNMRelIYUW0+3pZ/liHGA5
h0rIvSdXVMgQDEzrbLlmw8U6yFFdm/hJpAR5vpJSHKuGZX+4CB2vqhu5+at0yE/n
Yhi/8fF6W+iSybG16REtMA==
`protect END_PROTECTED
