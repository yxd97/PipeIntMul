`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
01wwqhZVsSt3kANy/GL/wpH6tvQ66eat08WjoYRTAv+zSX7GFQpyjZarAXAylXen
2dpZUAJvi5+K3jksa/EfxENasFnZKyrkQOoS/Tzan3pWHTc6w917AUdSyy+9PMHK
ZTttQt6EfX+u3+NFPtwX9o1DSIZgvK2sq3CIYyhEk6r5L7dzKT1yvaZrYJPeXHSM
xy7Ou5uqEIvpe+xY7tm/Q0nDwjCEXNHrfKSUvu1ltmibrMGdatr3pGmSPWD2rTgf
WhmP4eY5k0fIkEeW/ElqT4fpsdVHmEYEufTsIf3Bu6xwKzuMFVSyAzKvyBO/XMfu
0pnek2+34HYFf8JtdGvr5ax65zKUcaQ1SPpb/Pmw4+W1Y5IyCCFBaYF7Q1IcwglH
EUzNOFzoXiLt9BjNaA0uu/rLG5Z68QqbhWol047/lfo09P9aOnDXU2bKW6nvO8LP
PzVp/USOU5S6F0wJwhSrxGkYMMfHhUrj1NrwH6RdHXDHSvHebD/aqSnPMKLYoXKW
DjfWeNFEs4LfuWIK6wVDrtJ1/v/iBOG21DNsJcRMvI2H92lIWM8Hsu+njtLnqACn
`protect END_PROTECTED
