`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1k+aBGcPHur7tBHBDKWlSrCnLe6aFe69Ua0GVuOcyijVIsVlzsH7MPv4aie1Xo+
Uwws//gnYZJKlggbNgjZ45cxwZfCdPOrACAcMXMq72/ydyWTdUzqAcKQH2WFsjkM
5gZgftRxPn2tH731rg+n92CXCnpH7I4CL/QYb2dWYgBN5+uC5vPZvyNnvpEI8mZ8
BTRr2DgQH7c1xeLU4ydGTumepd/zlrDwTQLsLgVOZIrj6ACLWzYRaCHxl6PsGz3d
TgPuNpPm7HvMpXCWlHnwU7nLUmGx3cX8wXElJs5szJhb/ha9BxpTiH8nDUhgybIX
uiONTm1NNG6kh4YaDGDTwhiwwEuMqHr/8rDhL8/SFHnyh1ZBgVSEAdknOo8BssrY
yyVg/BIkcO4VA54GOrmkZzWxEb4ImTG4tkQhBTd9xg14yLR65KVhVJhTm4v6mHCP
`protect END_PROTECTED
