`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9awdeuFh2C1rIuPGE0Yw6ebuGgWECFsXfWre3s1K7daftsQODLGg+QMBj1I6zud
UECrPdtCX39qbe1jPXoeZAUHMLLF99A4MODBoLj8Rc1sEetHq4hsr1M0X9xjsyuZ
MAp1s3KlnggBUs9h1lhIfOGnXPAGefhMnU0bMg/Yb59CGJYYqOm/u6gCwSbT0akM
a9dmyPxtPJbRzlhghSSbv5x5AzN81sYb6MANL/KeAeLvFwoPEXjmgxDlhHHRUz/b
NL3Yb6p7hU/rM4yXvCBwD3YCyFG3O2lDYt1TyxdV3x0MMpiMbjAl4BkQU7pjHazq
JaLf1K0qe382Gqs3DCmuZlrysJJRyOaWWAINRx4afsAniC/4X2boD5cNC9g0nYtY
f17HczTwmBHIPSJzsF02wsyKqC9aYsu6N743ZmdsiYqwFutS5ljsjv/fnLxFYTJp
Oh8FVjHxKPRbiX5PfvQ+tIehdWKkcuQTjbRS0vAvNTBszAnWIppiFGhfiO58KzQF
tTMEU5LfiCnEYO96y/bvAtLB0kYYZ0c8GjPZv+M5JG+q8gTqYU/ZgSDhY0K6ibTD
l/eB3RtoeXIaFt/QkPWX923d5GSn5wjNkHfmXiZjpau2vJrsnlNYj+x9FCBwKqNw
P6cFsAJgOO3U98trloNvJpUCjbo11ewSkc+DfW8WGIZS7rVoJBVVqG/lPGZEpkZl
IECmpz/3zdirzVNM+EB/CcFq/f6Bh4aADKeRQX4amRTws30vWz3Sb8gmPws78XqD
YNcjznFgaJ0vtmf2FnxZ1sKf7u2A33Mw7VTXqMmtmLkD9y/y4cliKwUc1AtcUlZp
FNeOhzTpB6/rAG2qYlhnpY2c7cL2f9OVh64Pu7vZRs38xCYQ74AeQI953tTdA7+5
wKFl/zEAH3AnVoMWZ4diKB6HCup98lqk4SAuD0PEOGXM9WjJMToAFy8GDjUvTMhb
N9ZdOXa8KN7LLqhTCn1poYJrXmEQGcUFtriY3OhOUIlcpFcGT+PRi0IjeX2EAE6Y
9/3jD8EyWoyuzvq6fUGrSg==
`protect END_PROTECTED
