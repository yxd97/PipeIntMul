`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6HBuESlXiqtxCsrgohSLZhe69E4XXEjoyA4sAvBE4gO+2lk93YNTq1T2jWWRtXG
SLPc9Dod2B3CJjMSVAzGDrHh4bqRq81fv66MwSPmfFEMK54UEe4HIhq/9azKR+jD
A5IYYDgVgEeSXu+eNORmMJCzpemjcfkTkc38aIM2WXxpi28oZTZAKlkIRGsf5cDE
ozG01KKACgA6bG03AFdCH/opOFYqGU8SpBvZxznPSWiEhjvsgteWEktMouEmF/az
6Pu4ZlQiV51mvb3eZl8TPEqWR7SGVRnyi++ME7e1XPpBt1clWgmKm/WW0hThfBpu
PFvfREnlnADCuz3JG1qXOkpgVMCOEzMECokACeeGp3rBuiv1Y0e1gaUiB2sinnl6
cfM4u4pzkLXCVD9WkM17iTYYQTs4BRh0cbGEvzAwCHf2nLXqhS6qWM3CGdkiSf35
27f3SBSm/y6gvKzj+mP83nkhdLg6F7GNoOMgUCy2Sl/31aLWeyk4doGKJ3evI4Hk
ESktwKpOkf6JRQnG8qOEfZB8bWARghbNislmi9+1WYpUyNPTJT6h9h3+GLvybWRC
XlAAdpFXd6gcflsS9JNm+us2/YUHCSk/c/xlh8KLiWCKLNjbDWpNweGBXe4addJn
iVyYOlpajHosGqAk6rZSzVQBytUbPhuoCEM+pKh9poIX2L8Rn4IOSNLWCeHWoJ6l
SXW8b5ir19PNiLI6l+bJYwSMk6xFtx2/0paZLF/Z8WGIlfThU7sGDA7cy8YOtEzd
THIkORRDTNfkFcUCoBeKRn7TxkX7+mGVPYEc3ez/f81E2C4IEebUuK3kMVonU3te
wtF5dFDGzL1yH3ADjGjy4DzJXSRc5/QcFQ/Xr0V94JHWXisAynVEIUp/PWhTOpfV
/5axzBx80JRQ+RMBNWU/B3MOKB6H4iCQovmxfg65YggAGYkMJxcoFjDvB3fiHnw6
PLDaNfB2i0AIr6wzgX2+24Set+y6zZBh6SLUy7dMaa5HWujPPBHsOYn2TXSDjcN/
M3ni+rVS3TwfzAhBlNApBG+OOlEmNhByrUxd1pCAPtYt0BTZE9GPo7ixsC3C746S
uS8Rii7hVk+GnGNA6XEdz+XQ6akffAGDtg8d4I3ggVEJT030R4kk+Eo2zW3Hj5hg
oKMJH09lKqXZk/dVLUS1TmUqqgMTNOSBJAg3E4rXcKIRnjTgvjUZeSEG08OshBHb
UojIGlYpAOegW1UxofthlJrsI9ZbFAmMM8CXVBzLnYwJ2AHNv0i+a/YL1uA28dTm
UBGkG+fIAkU/U6y81NiVMzhbBgiWpOXwAKjFxbfQqWetuj11bCTdn06eVvPON5Qv
VMxGETq2h/OKxFqjrx/DyXEBjH9t8RHEo3aWs36gIhH4bL75+EM1ehfZJtrTYRIg
a75MIy9arwR+ZzwsIz9G/r0uC4/Jn4BesOPnjiZagroFho6ERw1fAaUNl+JHAaR5
odF8EiEOmxJEiaoZumP95AMVktBS0McEFzvJUSMw8lxItxxOW9veIDfzr9VzxQgs
Anqx6wD/LEorvXyDZr75qQa/Dd6F3O5rSpTP9GZxOdZzINpTZwUpCV0pzatbf75o
NAjMXUjsG02E3ZZ2eifAMd9hyv58pCRpysVk4ax7pqiKyWg8HsqeWjHLEWNLl/ZO
VrIVzOmdF026/ICyvfyiQ8gBwPeRGTywOt5MkRdpzAlFSkHKSyPxubs3n1L0Bhz0
AxoDgiWQmotPcX6tXPCZ3wj9Zs3pcy+vwp1BQ+qw0vQpf/VWv4wxfUB2mWni2j+f
cIrIdZfK5jChXuBt86S1BjeqBKAhsDmsJ0WogP0KP+8Tu+5jPNLHd83+XBXrMol2
brvqpQykD2kKLAXsUhSNnvsKnMNgqNZz+B5vIsJvHe26gbQkdvuvI8o3/XWX6fgQ
x8vczZ3FkWfx1tBng/jXWNMInYlPrxi7IgjDlVaC1b+31YV0zeY0x5Sd5NH/BhiJ
Aef/V2pR89DEBrcUzlzvy2fTcqChSEX6aLyKMI9ZRypZt0ltOIrVpUjac8bxkkyC
nRb1gBSIciWEwmYXP6sp2K0Oe6nrUABvu7oYBHO6W2G2qu+pxZJgEVd5PPvXrmpA
wD0vf7FOWzJ94ks3fsJsX8To04uT/HOCy588Fa5pNlu/AzsbREXtUC5YcTtAEAgD
ZMVnQHzFCRpm+vhsP4F3jc5cJfiCDBwA2dht/BRjVgM0BAFqfY/AFBz5czsBtBPD
128o13+GCi/Hk4iBSfcWtFfV5Lu/SFwHywvB2RSt4Yy7/7OKk2huv1sWs0fo5Bbv
OivErhc0a3v6HX6LKoH4FMX0xmRnAV0kZsFUAJ8YM7AaoMroVrPW85XxsumteTee
kJ6mROPzCweupAbRhRMP6mIbIzolDYRELBDkW5EFhmSex4/LVDvJlKpWBUPibTn9
kopaqZc5gsxXD0rP8CBpwMbsMyFkoa0sQr6hj//SU4MHaYLqNHm0dEAefKZXJ6iR
tAtZyW8utC4UbbbhL0xxgVzp9qYRZM5aUz97eWa1O8pPjeWsGI5yO6sZOFoLe9gq
ndpiT0Eb8teyBkwUgbJQvFN7OE0LGzF3Ot/wtX53XcIsAgj1F2NYkKsXZH5F4IEv
cN7ppgNnt1YFMvpVUgOosP1wFZ6ZIcBUXPQbsKkGv8yWvSJZfQFQCW9b3Q8ji/ke
tiEhc77fBR2QCj4GJFUkcqQ+aiSPKWSVEfK8UdgjNZ3OkILoDbmUCULjh6Ncp11X
nWf2o1anWfKBxmwnGUWTzJpu+Qdes6uNlzvx0IaDiHzko8eB8qQYCwmpNHNXcjyy
ee4scC5SAdtMeQpyyoZ5bInI38uOArOtqtn4ZKjQvO/JhOLlOwpc5FS5iVBhol59
rRbGJiQFBBP0k+JAQLJTpR4YxoGXtvGXctkPKYhRXs0QuryTxg++WBLkExUnqSB0
+AkLG+TiNqnTno7Irqrs/rwYJBpuymfDk3ek6Opa9J+TJVA4CedWnWDlfc5Q4Bov
GN68v+tDH87P9rEq0nAH7cYrsbuTOoNmd05ig8FY4vvdQLG9oth6yyp/i2uSiLK/
PGRe79/PiOkDFMI+7a64lUNCGkGybjK2QiNuq4tm/b9hQ7rybsNtDLGMrGKG6NW5
GO+Nu5V3lh5st5zqhp8Gcb35JWkJP8vqwPP50Yc4yMKV3OJlSbjE3bmPuOYZMrjx
`protect END_PROTECTED
