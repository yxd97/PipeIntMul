`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+4KgzuVDAFuXpUxKfqq0an/v6etJChzvyyIF19/9tmsJyLNb09Y6H49V8bON3TD
JN1EeSn9EGrPpaq0sPckSq0zY9gKrZEA3XD2iA4RDDO4tVEOKQ/FTOrD+sRUhZKs
8TUKl4sTgrEqm51EggrUK2rWi+EbOKVuteChxjwkOLYiaX+xGFfx7/ptAoM8f1bZ
EABFA50GPiKunRBFn08Gq5TetLmL2tsQbZOBBHfpFToaOzVwNrDnEDJAqKuzeVXG
XOv7GjGTGnf+PoPi06DbzQwdmtsEZhpnqrON9yhUBkGpl0P1rV1IKXJKcg+ryBDR
ZEOFYXIyIG/DqgOOWjvvbfDfZO45Je2vHcZX9TrAgjwtx5ef9gXWORqzp5/UurLZ
LGPPpc2pao0Cdeq3xqsgR08yAD65kbC+k2MHtVYxlOHSWMzK9mvPgSh0KYwvCsms
VS+QYYybRYUYE2eDf7foJEYDWZ1GvZQGzdjQnDLPGKIaybDp53fDo2GOCfzZqUBI
uksJvibSTArSlUuFYDOoSERRjzv4yf4JYY/r3ggzNj3Oe9dEZ+0uTnJYsjAjvTsK
`protect END_PROTECTED
