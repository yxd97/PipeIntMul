`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MMPVc6h1/RKEOgi3+Uht478lC8hPBKE2f6vGApAFIXGlTZgjIIHKj/FTiATCIyfi
5uLZ9KHRgwSExtKKGaYkdt6WlYPNKfBv76LbwjrcsYyt5in9Pmr9epNlEQbKRlIa
XWfwV0GmNeOrv8KeJoaL9R0Ik47GzMKVOWPUsp8dyT9aXj1CnYSO9QTMGdqljhr7
cgRJl42Azg2BCOd7uduuYwNDEIJLG8dMHRK/EOZ9F0p6R40FYxTdnnc4dK9FuFel
2F+A4gteDV4ipEWZKFTage5cWqMRU3dTpHfN0dxS4YaKE3WeNBlc/RlczKYur1co
xGOve+oxi4VhFqBOI/5UjYuopOpJfJi6xR13fEC+js0Cksnu8ADimOUcuS5PXjex
M79WSfHPTAh6tdmCndta/eLNmbiksp/ijmRC6Ngs01ELlg14qMXuXi4REALgzhQG
t38DqlHf3Y7CyScFLpMuppQgG6qeiw+LFiOboWVDSL6ALH+w2q0OHZadrec8tlsv
/Mh4GIlh1kEDVCcFpTE+Ebrrw9Fyqc7YLF4lX0sbo72Y/Nhv65XlJOTQaBNGMAb1
+0DeAPgBUjOrtBreAlyrl6idENQRpLcjtPRtYmE4rUDrnHGPqy9xocn+jthM+LNT
cIHp9AnLvmszg1boc3xencfx6s+7mmAMyzITB0z++8KU2Tc/y3ubDXSKuSy8WQRQ
z9QQ9hDZp3cOErzsnL25fuPjnX8KrqG9azg4Jf1Nauk80W/xCop1JSzuNW/xzOle
U2Jbh9hstETU1YxILbyMlQujRRTgaf1SO7wLvbIXDQtYJHxcnbkIhKla2oK+J1BQ
GC63YoZvCB9Cfb4XCrHhWdS2vMG8nyzz6bUI0+oMmZ07Ip6k7D565KYGViYaWBmD
`protect END_PROTECTED
