`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b9acGd3b0pAkTE3e93BsADDMdV4QHRkfOHOwegnyQdq8Rk8HkxrZKxyC09N81v2B
WXwgddXLT27ew0Dz9c8nLviAWJ3g3LZhFjWtqRs2KLH1uCD7uT60jb3U3eo0udaK
a5kPsT3i+yxluGuXNFOGcHE8oskIGoE2FM4I2AWwpicG3g8oULQd4Cs32XXAIprf
GGWBwvtcZP9fKHjoi+lisl3gy+tmXeZdGs2briMRLLffJYZgH0XQJHJtaZoQOY6F
e2jWKoXC2aK7r7CuTUQajlRv6SDss3am+kmN5FysCOi3D+NOT9jdlykV63IcMfPs
h2Y2vK3vsfYFrVEdm1Ing/jM2AdrRMsJ8LvMLEInqsxexYkNoP+VX86YvTk550N9
XILIvLXoDwp9l6lG6l1hNEp9TgoZvlLd7uPDEhEpmQSJpoZPKNtW8yGaPrBT0C/h
I33LKCr5R2Y1ui0sakly4M6QkQI6zb/osQHUe7Ij2mCD5FSUx+nWs3jK6cm8m82K
UOhtD89Y7vr8Qc20I0B0yh8gZR66KBZ7TpAX7Ih4SFBC60SYx8XTJfP4rALzKPeh
WTCPaTwAAFZRsVK2zXzAYDMr/JI5MKMH6ixJpPX5L4i+BjslDfMiRQDHTS6xSP5o
g5/8xghTONTrl0wCnM2ouA==
`protect END_PROTECTED
