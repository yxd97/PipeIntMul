`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XvlRT23FXRnjzmggOg8cWNWHS0UQEizVbEnzrWRJHno1pIjxnW8ivY5Kw3tGgYfQ
rs2OjXqyTbebnt1jmlNRRjrhsIRfGwV4+5ynRVvdj3JYqutawIuGUepBMTHzB+sV
gt+WGb/8YYN6bgpdpOAcZCXflAqHAtZ/e9aTTJfTk//WvwaV5zBHwCREefT6//Fc
WBYXHcfp1eVZiu+kmApKfFgH+MUQ/IfV4k6muYY0WolfYCqHk35oFzbt7ktzcned
qroUJmyaUzeUDDFEyTLWMUckoKDIFGOu4/BrTS9qucwQsUhALUnhuYmrdMSKKTOl
st6AC+irAPbDW5lPUvVlyFqHWw7A2MCisstDi04Thym4e9RZ2gAghZZypXjGF6yl
GaeGT99vlmkjL5V6KNOrgElcdStIOJb1eCFF1C7iB2VwTZtlfpY3i8qRT1Bcppup
BoZJN1IJJP8IQ4pIVZX9Wk4frtHdoPwQDoLbGI3UeM+27CHUahaGbMdcBPmuHgfc
l728f/OlpIaI82pqdIx0SWGDGrHquHgxrCuZmIRIMWxh9GC5tPI2YQ2bllrscD7e
iVYgPn+J+yOmQX8hYWiyyW2rmF4Im3eL2jAacFPMRb5Q9KDd4HhkUHP85CKd+Fsz
mCcSK+Qh5VsFwXKyBzQdvXygrIpPOq6TQDSUgSbk06ahDXk1VG2eGwDPlzdluHjL
/3dVs1UXt442lItzTOl+u5GdB6fiLS+AfM4KXd941yVT8NK3Kyz7tYaFpIVLtS6v
90m6acdzm1grysD4OnhP85jfRqyc4WdwhDGs2wFlmKDEG315wXm72SB34F4WeCxj
SK9Pi8uGZ5lPgtBj/vqI+GVt94SHrS0ELXo822hadBMJ5dGjxArtt2Um0y9fJAi8
aByKZoBOnhADxBl5Kdd9u7olaWBMrWcP4ltP6lmHeiYa4Ru7171drzdvvvAnZw9l
`protect END_PROTECTED
