`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KxrBO3+VbKzpc1hV4MfaMWUTNB4sxnpr1NsVLbcJDG609w7ZotlKFCm7TmeqDO2c
8MfhX9zulKtrsGiQscfU/RIhhKSNLJZUG25jOOeNY4QZguYuVc2dmutZkn2jlllt
Tmrjl/wVDGraFlZbkqBCfVseVCdXaljPWlL2DsdBZyMOQsMlOKez2zSdSqCcGT8/
/rtoQZeR911rVNTxAr/IhTReePdI/Nj3y6ymZzIGQBBeQO2eBDHrrf/7nGlhcLe7
9RMcT2fHsdk6/0eTjLoH9E1holekvEU+2sRoeN6EDbfAYjY7s6Szq5toWtl+asyI
8cn4MqB1zq4za6Awh4dO9LR18/N04thIMXSJyHoC5f4eudhuuNecMedUSuXsNlhz
w7+tB72f6zH3t5FRFG0HvVA2qd//Xgg3zRNTczaBmcaqxky/If3Aac/lftCfk57B
GJVy493+DAUIH1GKygz0i9qkOyODj+Rwzwbyrm+ii+sJfMJSttLXQJ1EITIbDfTv
C3/O3SXcugQmEE8fwIUy4yJKIiaDeqKZkAE0lx1Yts0qbeSDi0neRSOBpvoeekak
rljr0P1LVJ1o1kyb0DdwLEcX3C7QwwBOOLVl5z6kicfQBb9gWmp/0xToHWib83yT
FSQZs3vTZ9JJTmdJ8p8lrv8LLg+0hbYaUF2d/iXQo1sKAZ6Tyg6XLULP80U5ddCG
zYXg+fqdjLbmfx01D3Wu0vaYBKqWvu4I9jbqpyZsGongGURfO0nQuHjMkSzCq6kw
XdiZ40cHeFnYuLc9QGnngK4XuNrznZnhkVc/MKnwq5IMizFpkO6O/XLw4IvWgUO8
fXQGnpUZg3zUiQ5ev9+VfVcvgl/7Luwg47K0a9FonUCxqMcWdSM889mF2RBVsREr
YCqp+gOXUG+dmpqAQ1vESXFuZqJ4iKqEFeHDgeHqogVvpTeLp9iEjBkwqufZmT4h
3S56YJNhdf6SeljLt/74Ng8MPX8iHhE3tfAJbuexlLjmZy8zMzuTMMuCPbeWqwI7
QKa607JLwxskU9W6kDJjpjMkOcq1Bl8BrJZaGsHU+d6ytC3stlUUplD1h1DtDGt4
7qxcJWZxN1rZ6HVt1GNrNo6xOAGRnfM3VIDa/9zxB4Q2XLp4k/OLttX/rBd0v/+K
bLPIP22T/S3+MbjZbVp6XE/ZMieX9KApl6Zt3n+VtmA=
`protect END_PROTECTED
