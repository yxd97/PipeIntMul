`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AohGXsEnfFdsc56jJfctvfc6OZoPkShUDo0KcSPph+2rYCa9mwh1y5lmlPeqsN5b
qW16+4RqWV+SD6Y5fBjNI2khUae/nbTjLnEljTMgZ/ciYJWwnX/QJ+q7EVbpu2Jx
QknwVREchXjQUTiR1IpO0bxE34TIwO5ZIaKw5B93LnixJ6nbd8SbPf1F4VpQVVL2
S04RNJjziC6DtBGtZblm0+86jbo5zLuRovyoWkmPBkx5bxYsQK2yeOZ6yCUhs7RQ
FyLclVIoJCWVjTSwl1HlhxQ14aPd/34EsHAbJSU/cyEJ9GT4iSnRYk1QXouD/Bs0
NiUPDx1osKpZlbk3YKk8O/TmO+MLcysoB8K0XcZWJ0gQEBJIhvtqLdawb9Q1WtX6
fI7Hf3lCgz0SFbROsQJyyc9yYYF3IIg97YB8Y5nrIRE13xb1tTEamM8Gzqi2pgfN
o6fWnECSD9wmokiYXNQsGwplAehAMxHJt/g8Kyk852Tqo4UvPf4UyiI9cyT06UAj
ZgY9v1aXJ6qfsmanhaRAuwjKg/8Lx2o91LkdhR/gHdEUcB4bxelQCkYI+7fx/VPz
ds1Z66kEtxBi9pivZCV6SUSNwMupPniUwAaX2q5ZmEC3VXU+7IN6PGJaVwu1mV3W
g7ba6j/aKBhDsJ5nkJL4DRJkK7GkjnUcK0b6jBDk67BQeBnmCKxZsOqJnZEsD7Aw
fwSxzmXoPKeT+zFCqjCzoc3qMGjQJLjqgsLTR7CdPLmGj6kpAwlL6NAI2aywd3AF
yFZ6OS5I+xvDg5uYBsbRHkYiL0lQhR0wLv1Ewa2MpZbCLCQTiKBS49C6cu0P2/oA
U0ojQFJ5TV65jpYWwSjeC5RylPuuC+9ObrehhuCXEPQ=
`protect END_PROTECTED
