`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lyqyVI8fAU036V7o6qfS9u3zS1yJEWpjY68yhn729McJ9HEyS0Aj7v6R+rKCF+4s
olMOq0AIi91Vdi3OEj7jZKWqZaSu5jN9+Wy4s9iGeablJw5T3g8IpJRtjvido5be
Art6ECqdciHaD0t2SO0e6myfQjLMkHT6d6E/ePwEtE/B2oLxlMaCkbBdqd1l532f
z53RJTX8rmpnUlhgjuXiaPCiRdpDqUJ363ki8Kx4ACtz0P95x29q8uPbaE3cXJLk
RjNnMWi+76kOFPPNB29XSEHrfEg+ZZLSHys8Xu4yb7L//tbdGiNMFEpnLCeeTcPu
wvGoU4og1cu83mZY5vJfHoSILcVICcRYDhYZAg/qdLSkyG9aMfRbTUNGdRe1+zpp
t9L0SjbatItJR4LPnfwfkaVVcwq4ZbRFjeBsE1sKpyR5IOPY9jzqs8Tpgch6TniK
+OrqWw4wzx1FIqsDE7S6XiuU6fQr2klyV25yITzwTgvy2FHdhy8Q0+Pipq0Chga1
YJZiw7QKrHup/RiS+F4WkRZp5ahlSD4DZR6XMKJZrOBl5jGCs3g72+paiBa23Y5B
4q3H5xGUqBwg0SKexvhkacWag21ZYPkU1LNtzq38NxwP23lhYrq6zDEVUL6o13/0
qvEV9lqWTlrUDQjdsKgsYSS8EmZnPD3yXK6hq+qg+YOOEINvOGN9IZG41MkugWR4
Dnu1ILarw35bd9HnuohM/2cqZ1pGbxv3L0PMYDvZy15e4Amdh0tXocGXb1kMRg9z
EPOAHzH345i7X+PvJkACdG+oMm3k0k6BKsfO9rwfi9VcIx/VGw90J4KtBkvHcXvI
PkwcoeZs3EV84uVXYCYYKOSsVB74ZabDgYVZwM1m1Tw=
`protect END_PROTECTED
