`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7PQofFYyaZoKlgiIf4MZ2fe90avGxhnx+R53wJiterDT6E7UIRkIEaga54A+Xyhx
D8NC6HO2j38MZpz6x09fu3zSbTmcVAWoLZlS1nI1ZdnzJHXAEfu2g00KhZXMtaYo
l4NdmbeOCeCaun85gRriYEUWbu49MZRCV6Tb6nIoNZp/ML7LB6W/Epm4zeRCseLS
Sk0hNCuuHh2F7KqALOSOIoe62coEIX2zhip8YC5xMR/mEPRFM3F6WQyuAS1G/ATF
E1K5NumGzy4y1M6h43kRHjb80CCTtzD2csDEbtl27TaW3geSXVE/bN83wOxhdtMa
WuhzjDP7AEzWn/pvE6jLWSfqJZVJSEr9AGy5bQcsnOLiEH//CXWQvvvINWKxNVos
1z6aCY1VtHZo4umwMa14igTCTG0siflPU2eKLevTAVwNHtFOPsmgF+Ykefig5D5O
02yeVYVeI7v/yirNWfGOgB/CLh3a2sDE9ryR/Ax6mKz/EgzAnOPlrKWD9v+0Npq7
X51ggNNJSD2UuVirIqEGf0OeIdp/9lx39ydiktdvokZkPRJkW37p7f7HEDxjhfC7
yHGt6Kof17x+4tA+YWk/vStC1w+wl3SPmxht1x6Fkl8=
`protect END_PROTECTED
