`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5/SjyF628xyRJRkY8GO3f/ke4iDn8AGAsY1137D5G+K6PGePRIXOZ2aLV/I5Z1E
K2Bqa67j6Ov6ZGz6vlpiasbbyWhcGoqivMczrNa3M1wMC6GWWlBdcACP2IZL/xQa
jtWRConQY+V0cdIhy4ChrF5Rkrkx6kFgmI2Wi1TmYMidk+zMeyaXSrvIoMA9ZGGp
n4GS02Uuw85uehaJIViE+sQLzkbm4AnDo8BERL3zazfXpHjoE44NkwRfELyDQdts
M+NOmuQoK1k2epNnptUgr92yWDZoo9jLUvbXA38EHE14gdMySXYeKLm9EZ3IJKI7
44UgDzpIrQd8fYGAIZRKOQ/xphtT+RhbNR/BePC4P5PAxUkQ2U57ljt0DYFyQ7kf
yQv4xSrfjskde+opCgDGVNuUTqMMO6IjKUsMHRdwI5CpikG4aJ2Lh5iZU+o/X0Bg
d+sEX0jtl9t9Vl41DEACgdy3ekqgianZW46zxLPrIDzjwOHgJAvg2QThp4kZ4PUT
j1cpbjc0YedTXS0DAprY3rCN7jx8nA7xS+CKBr3nkAp18rpZZIqIHgemPozeNdqZ
zMZNJ4uoM5q7Q6lLD9Q2clvEjMrqbR8ACraanEX7zAoLVSWxo9l67g5GeG4U2yfc
L93hvmbe6XOyY9Mwn4nzBp8x8bOVABFUvjJRl634p6ibsrsCNgsR2AqFyLNnJQh0
5xHUR+D8zoF9SzHD4nDxYOmwfF9PLuC8KG/ae+jE+WiS73hZabcrFNzV7o1TtF4q
q646+kL6MAEEvAzrJ+r2f2MNpSxP115uNMS1HlZfwZge4HLqorD+vTzNJvpFhKMG
bREisRrB1SPiZF8jXHn6RGbZXwFbS/sttvjXgp60Vpdz61LAf/rPk1ss/RlYXRzl
C3ELzEbFokokiceSD8jiXoyp2XsdEki5RF8fCptvPTHsFRCkJkq3CWRFIdVCiYuF
FqCFkdY1dIE0Cfm+AJUGDpmTEQ5mf6QS7ZLGPQkjrw9vuq7b6VkKT71tcs69PcYv
wYLSHdDGkpM7CpZlyIFmUsFFXylwQvuQJoR4/gdDAgaXbuBUQZZyUXZ+A0oeYJRX
nrFrJP8U4uMh+i/83tf/tiyGQP9wT9F2D3+WACw8NaZt5zx+8MwleWdJLGC6fP3B
3DdUQ31+tDF23oNJ3vw5HTm84NiPxNwvNAwWiZvOStgaKWioEKMmUNdpK8HmHT/n
hKRDdtBrYSKw2qzLF4zseHi6Ym6uq+vPl3ydkPjDGvGwMcTBHI8GRoapDQ0J086c
/8zbkc5B3+UlWsTjMHzMu94wNBxDYiI/9mTFMTNyfmo9O2eP5uAU1k577SrVhyvk
OK4zzQX1lNEn/jjBZsnOrxe3SBcSoGw7v3/0BkMM02CDHu5KR18jvifhIFNNg5iQ
YdIh0wjNz19Er6gu0FwaY0f9I3mttZvyh3/9msFKAQe01N2y77v+w+mV2v+3LUDT
VrRSxFIaTLKR8yut4GFy7KmD5s+4SkifstjD6miR6Dnll0qjoQaxfoSS7TeEu9Nn
Kd9/D89RfJEoWzVxsatTc4OFs4h4mFPOGfiDm2WBRxU=
`protect END_PROTECTED
