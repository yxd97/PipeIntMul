`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JvddP7rhPfvaAWBNOWdn94ns/nRC+rHb/H++iYvJQptNQIT608Nny/xGrB7JuVbU
vp+9t4rw91eOyMxZRXlO21KB5DOr8L/Y4R+ExUlWZcC215lQKFGCbdG+2l8J25pY
5hj8Syh7BkbDCHUih3H1p03uj1CmI4uxXhnsv0cPgJyAUsppsJVnHVqRf7fljTTm
JOG0p7JC9lqwVVxC1aL4k1mL3PtIoGURfzYwHaTV/2JMBhkxNFvW8Q74gwWiAnT1
eJDciga8O3zfkQioH2bYjnGIXMrclnVm1cEEFb8h9+bVifq6ekqfslprzFrNwGKW
iSdHnOzko7I0pviMDeUNbk2N/oTY91f2F2GhdmXzh23xO5v5ntFaFKE0buTq9UPE
b3eEJIYFgPPIQwiGZ98DKyv6XkQdugICr1YymRITLITTH+94lDv18trmEURPdOmp
CTRuV66nOmKkZ/pl0i3GibJM9qL0xSUhye+t0D0lPduAWXUNlwBQIvpPCy7ylnF/
52/24Ys24ZflR2P0TMffKXAV6YNHEvhkFTvveGOJPREHZkbgH3z3/F+RSXw9Q1Mo
ApeWyYDtsjyxfECBd/JHnY9RK3IRAEYjXBhJMcibcWe3XShl1fIVzQQg7PjhDw7A
+KnWCHIBn+aiWrPCUMVL7d5EYiDHHvIZQofKJIFc9NN8Ks+vzv3olG4yIeJ85iVB
iUZZJSVuk6bf7YQ82wR31T3uyDioWBCI1PFcC+8hV8FmezuR1sEscpyVLGIcVe3a
3PqYO/IUEq+kz7L8WO305SEr0UM4LE+b/wcB/db0Ahz51pgb5gJJ/14v/yrzdMJ+
kmLgBKAm9UbAh7frhM6bmwaLwC6EpO/YEv3fFsimmPyuFadq8COdfC+HXI33M07m
FBIUul97Xk+E301XHguWImMejHWu+LvIXQJnEOMfa29lZrAeO/ApjwwHber3kM3h
`protect END_PROTECTED
