`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaPTqjojYORqJq+jzPId8/cfiUwFdrVh7vT75HlUmvjz1TBmE3J+fur/XaASEZFh
DoDkZBmnxs/JiVufLuKsxlzIATmK5pufWRjFGUR/Tq7pBfk7ud12kjIbfBfs8X/w
KawY9QjADZCEO5DuaUmIBJDURCVZXVichq1ftBSnzr2Trk9tpN1q4+FSPrqiTnkz
Bz/PEg0a1Gc4D5hnOGTaMZmQzgw7lijTUhVdiixz+OZu9mx+utG8z2ZfjmRNEFXw
vnu7NsoXghoqj2dZCHOaDBGeRGoVjojjyhGYM/IYqhzvIFa/jjapp+BSN29QZGZ4
`protect END_PROTECTED
