`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aY5T8RGTeJDsYV8RC6PYnnUDYaVmoToC05gd4KzXJXU2jZZFBUmZGVvvfU3raaai
4T/TuUEYpRWrVJeMSMqc6eiryU3eovI52djsHzGNm1/wD0vbi8+9QFBrj3juO5hL
G/Bwe5mEZ8m9sARckNLR1vyQ2AcE8d3P5NKLqnC0pu3FAVdGhWT0FuA0NMVZG2/N
OMUc7AgNl5nJwvPWGLS4iqo0MJiINGoH6b28mlZtj3HuwzmBfVGGXh5zeBm91upA
uVgUua7feteJwMRlzx3ZxiEtAMFPJIM8mAQsrSuoweAPMkYQXEIHsHF7wWzbDhW8
SHDOmnndDSr66yNeOBtgYTNYsxo9Ou5TjsUU0ZRTwJjZvOnqMg2JYrDQ/zErXLtW
`protect END_PROTECTED
