`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8Tj1+PKOlBuK3fIlhgbhE//5CnsuCYn2tn0IjrixAXXnQl0WtYJAxEvXLDqmEvc
So+HwlsDvWcM6gLDRP5bDb0Ev0EmdP6gMliG9QAHgX+DhR2UcFpGIP9j49a51ZQy
VJAnmgzGG0NNQ5W+uqUIldRhtV7U4lgbrvREkrGS4EZqQiuzhW9mE7tR61J73bl6
dPK4+WXD4vL6Wdo4zOvwkJsKU8NLXuL48YH/SejeSkl+Pi1yWdHvuTgj7/cLgL77
mnGF30gWBXXPvafNmFplDZvO6plJ8ubJBZilVd6ttMLCJSogleCsmrt/Lw0BtvRE
8DLagDswTw5nAjacyPnOekrDD1WAaWQVLyaffUcPkGVFrrWwVaAYABIOdFuX0Blg
4hesGzjCYQSoz15lI4o9PlfzRP0f4nl/4qGgpuYdrMx0FKijQsXoA6Hz53FYgD6o
XyCCCbBMmRFcBwyf+ZL7Ld05sHrQQCFzOI6Z7B8hAqruhjDYDe9hRClYTvfXLI/c
TfYDlFvpC9SiHj5Tt2k7gTcFwGMhyVAEvTyJFjVZuKLk8JdSk7r1VwsVG5JGJb9u
DLokKlG4o3OF0XUA+44DSG5ptC3wRBvVpQYDVo4xUj8FtrRiAci0z7tSxgsG39/X
/X2HZjYWqFh6BR3YQvhTymoQPk1iAZ1wGesrudFfTYQykPNY4Ya1KofU+1cQwoPo
ZdixMbRSmSDuBlaSc11VdyR93jh9ajGjIa3I/7dlsNdag68kBsNwwyvlJ799Is9h
OXWFJ6fHRibKnZ26lrcDuPQZf425pFgAaYwl3P5EBgOTCdsTiCcIwL1X928NLl0w
/oZ3mSR5UWASUEA/29B1An55a3FkRDWglLh/uyo4cj8j4lsLHZT4W2WlfROnuSM0
rVFSV24N+HLrqNS7yWfz2MK+x5spQvY6R/Y2RfdaJzolyXcfTJ/ICde2u5/gptDB
xB0uktkIe2G6Y8Nq4VqmDG7mL4PG7Uq+9rGfjR9+nMmA2mysNWZVLUVQaa+ssecs
X+cwd2hDrVdeaxKrnX33R/yZ2jJl4MVENzLWyr8YhaxJrPjKhq11tw26no0wCccy
/VTMz18bgCaRnJDVTWQhcmwAjwQP7g0MGnbbX7zT4l8xCEzVcPB9wSSdes6GnZ9a
xqEc5mEV58KIFM1sW/X49BlfeOk8l2T5aLt/gd20BIpmf/QlIlMIKX9ubOE9H46C
4kPjKUNs8M4mlPWnZCRdqRFUHzxTnjcJm+nvxrn0R79uUKEuI+E7qx3dlcTGjT6W
hiopIJT4aDlssyl9Albo3O+CCCuDzKahe004XExhKLjXawGBQMNs0zDebXhjgpSF
4K8R6J94OetJ3/O0ICMajEwInYT462uXZa7eopiJkmO85X61PjzpzVo6Am+SAm+M
Zu65w+lnxe6LDMgQQ95rV7bgcahQ+XyQm+xroQbHoSVJqhXdhYIewBs2R221yWf5
FAEAJZQtUGkpYEnq7R7iSy9GJRU49gKpDF3O9NekjpcKKNOLpzrYCAvlcnSmKkCT
rcjkzUvBrLleCWuNQmlEPdB1EaB/5nnxJ2IrlmlgH0Nu10Q82pu3L2CDFoeR3hv4
Tnociq66kLA9F+zJgVA5/PEFVzvTLoKdkY73nv/isctzYyauvwlpwLZimy+T0Vh+
XIJQu/Ve6dZIG86NjivmLsRPTjkfBVdIARdCFPF8ZXTyj/Q6YxKndyx3ivxYrLlh
G2sB2N1S8/d1c+HPRROXaMSyZrTN6oPI39xlGKxonu54XUH1G0kPAcc/8t5AIPoE
kCRjf0fdsrzcAkRoD3EmLIhaWPRPa8gMMughqGpMJ/JSyB9BuUSS2xGaMSI+7h4G
gKHPcfAR8gN3xMV1ewQMClH9soN3JkJnljhrJ3qStug5ZxmcuO+aEgIXs3BkoJFE
0VvBP5Qr/mtB3u0646NeSo15XDFDMM2vW/+eklxepW9fpbL9R9aOgNLyDaDdBEqN
ypCW6m/kpUNLq8tbsXFc9g1uD/G6jrQu+LL7GNKMRDb6cPN4pFJCcs+rm2LzLUWz
DdghfwhELBlZNlxrtn+OpL/HtmrZI4qetaUz2mGRmYiEkDNGtBBk8PMfRuuU6jzd
Biet4ipNozQ/9FXYzxPoZE/3W8kCDT2KGYbZ+e12P8z+N6JdvMk8YlYCQd4W3jFi
UNGfusZK0CkU65AkMbB6fykOJ5oUixGAEnox+/9dl8YrheLcww6kyuoOpj71EAhR
wxtcS6Q7eVCkBCCvEN7Qrk2pMIR/xdo+lpQy6PqAr7e1x0Xccq5kqe/pJvvV8IDQ
gm1xSVrxYDN2RHQoCkStAfqNsX1OupXlWWshyuvm8YTGOPlpcZCbi4SpP8j5Hm41
rNH3nBc2/gA0rz8MDiplTWAYji8UaVYahkOEQUC8fWhYXflAytH3SbfUkKvykmBN
wDoN/KRt/M7Hvs0qNFWMzspapPeaZY2uOWo4z7p8LJOskxtdlNMN/1gsXfBEZkIq
lkps6Fupu0OhEUiqtnVvTaZFMhw7NZM6dsKMl3lmwfr8qU5iTwaK6/95yEe9S9i0
p2WhEds8YMvnxDIs55DkRPtX/Km/w7zpcVwaZUC2g+SLR9r/NLfXWr0AaCpmdEDZ
nn2v3tzmtFD+ZM463WCLof7trDdTmHNOqFqMNt/DXpEtfGMMDaS72s8UZB5pdCxz
/4r8WNldSfN4TYEfGjfOrnVepnWfsdXYTJUQDIIA71KPZQ2jwVz2BkENhSuBEI7K
kOss/U5LNalIXFnYXm0ODCUJsB8Mma++UlVCEj4A/qMloYq0cngAsdlYYyN+PiIU
slHUalMn9GMRzmfy5Rfi7W0iupyXc5zGcHzJyw1n+KYl2x9y2IIUzZ8Zky5gs6sw
xv5KbPtIAKbjd3+UGAyRRBI+Hi0/oTIwp+dgHY5tcdOxOLeH1ywwxWMykNO2HKt9
5gKApIlNI68IcImxfbuOb9l3h8X8ux1OwNiMxTp7iE6zOZUiyXmA43k5aL+G5jje
S4B01xcv3OWFDH4si5OJ5GF8j7arkIuxYFp0bc2IZvzreBDLkpYfIFvm7MP89zaL
QJDiPOXIqGIgsSmDHLTu3nCvAJ9Nxz6sx9zN1H6j7S05eyD1XdyzapM9TYfOMsfV
u6yPDu9OPX/s684LEa+BzUDdpCQszou8nXnBKIq55/Y1uHkJ1bfroOp2Ewhxx7lR
DnKrYo0gWdLRqnOkFZLr9ItnjSJoFPkBlSPQg12B2piD2Jd0D6HO7uDlgQBkhlLz
P8GgAe8Gmx2qQZdNkHkDZkkamxW9VWuJA+rhZJIFVadfBdCBInhbH8e/nSPDY41g
fAUNP14Rw6oNxvzKjyJWugT1B6loFiQ2SrU13V+0fzjLM47mNk5NPw9nYumXyb5h
EPwHTn7kMv6fJfgZFG+595lEi4wn5YB3MQJgpFTZEoOkUGmx5wJGQ7QZhmrhrw9N
jIkd3mdSlhui0qZJgCMCsTIhCA7tvuoO8ctFj/5DW3NGDntJ1gXF7Nr9CSC/Hq7T
w+KpmtqWVgkf672YrgLPwp0K5SnG2awuq03/aczNHxpL7QzNNsPElmgz6TEEQJRO
36Yqsa56c7RLrONiCjNNfP8NUdmSUefmnX0zlXr0Nhsufz07z5wkopK2AUxWwcQN
/Eyssom/Bs0tTq3DLp6yZJXxPAhWcRCQ6RtcggdvOEwU/byJIHE+0goEnvGuRBSs
nClq4kLOCxSGSq1nflI/h4pRYpb10mwRlQlpq1HmW57Q/tkFAsj2H9mYD92NaIuR
HgnYwalFhpUf5JRDw64Xu+xB+QVbGeF//WBJqKl9gGvL3CYI48sn6tJBwB51g3AC
bKKc3HWfMHNNwhUm6Tpvu794v3xsLxW5Qed1Y4YbhvhmXyFCS42HzyuZ+W22kbT/
Rv8tJtZCr9tXevo8r/TJiWnAFfj0JvDJNkPzdWH4V6nBpjt0YXBbOLguSRRo7ifi
12++9WkInl0KPfzhCyoI8/Dekyj0JdH88y55N8ilDVuG8jjzGC2BZGlSmfpb2oq1
YSNDBrVtcze55MY9itMf3Q7F8214KXP7EToCNXohkuypFZ+G1No3BbpwG8Z58b3i
ZAU3plNBdcm3ZWdoxu30VIoeAVitwsZkOskGXrOARq/WiXQ7fpnafqacLFArlF5m
G1qJalb9xVFgvbiv6e+sxbgbFWUIj44KYpxIXzBjEfT1Ctoh1Oq55RZ8xpisLx+O
YWbMdXjBNvysej0mo4l7q6GEFQFYg/jaujCmh29IWAcm+G9lvNGXDJZqYD8ubrSv
6y+tAQM+GDQSYfYXJ3rvcKW+6bF+XNa3vNENW1/rqsrYgLtpkWZgkxb+Pd36/CET
xh+r70BOLf/M2s+Hnw7EqqcxZ8ARGzxp5YmrjwwGfCkXvtkVkKyhtoHvWL/i+6ui
nnuFqvy0YbJDQJNRAKrhhNxRC/ya3Oze513OVc+4BgbLllo12PD1ErLOiaoZ6FKW
3ttJ87EF5RdORdOQy4bPHdOHfK5xQg2SC5y9Im8rS5pz2dSGc2oHnYyF0kXGGIdl
Vq/OO/5C1UzF03SWKG2baNOxmo4Ds5yyLlsjJEvDHSIrNgsXJ2eOP7XNim5Q1tJr
WBZVqAlGYfLE9xBWJTMZE/GZIAFBp2NZlryzRZLeAv+rlxxrVw3LvAY4EpBJ4oYw
U0upMIr3jxC360vZFRPFxxEO/GZ3M/kMMKoRFfERftC7y/vAB30Hf0JEtMjzF4FV
8I7C9ZOriJD3V23T+Y+IGnDC8emK9XfxdaX64bFSnq4sVBntQydLShu/rwRADlqc
onwo5JGhNbS4/W2PQALslemUlCL3+ieGVUPx4hbzappxTXfPEn5wScFYSb6BIsKB
VN6uLNC2S0KohCKCp6Bw08PSTuXT64qfKkxZApik73D/jptVchmrx8LWOm6jlseo
qTeElqoJHqGQZ2YX6+Q3LttSBONScD0m8qhw3ikAAHoZbf6T+yHFW34aKjLWt+ft
Xkt3pLS/N73lvZmNL1txkwBg9BRiSlphtbbjOBca2cMDNxNSD50I6hRZip1IYKU4
9gms0337FKjmZ8JErD4fTg==
`protect END_PROTECTED
