`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CNkA3zJfypDjjdCQIyds3QhGlNNgUTi8waZzkuzzIQoAwroohKFu0TSzhO1+8HOU
iXzQC/Z/KrGMogbfqo+ntPzkwHUxHg/NibDXQZb7QoUnOoeqxJgD2tJnaDDab7bM
lJY0agn/nmDdD9JO6BeG4S5Bh1LFPMkrH2hG7QX/o8fzB3D/7xr/Ks3IXxWbyBTW
05SNgsXsWoJ/wuD/lT5Mc8+DQ4IsO72XJ8zsKLqdekmxQhZU9bShLsuwDYWWmH4w
4iSVQPVcbiyYL6CNLzjwrk4vjmlyhhO24QqYZUe+5LwB3VqMIlhebOoii2lEfs+2
06TpmiAhg/HdNZMNByGFdJnok8CM1bltleI1OE60p785QRhZ95IlZRSaEYJmj3wO
RV2BSrDVTJ4fqEzJ5ROv4KT50DyynrEwyhK+i7P+ZgXu2MUocx3xM4PCyg8oSbJa
8WExQ4eaTEbV260k8EU0Fd/0c0n7qNbvqgwxKb+4D0l0LZJjNWf7LCITRJBWlRL+
rfrK54vCFRfzZhJ3MhGdsHv+ISMI8fF62vCa6sE0kto97Tr+K/EvD1p03axv42MK
HF0wefrqE3cCSOo+xBuFQAKuIF7UEmEy0CEcpOEp7ts=
`protect END_PROTECTED
