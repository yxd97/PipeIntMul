`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9vXZ+M5D3F7Q9K5LT+Vn4ZHe2ltD5jvQGqKTRQQB6s1Fasdqu+MT764PSbLxqhzk
Y2MwsSkTrA+J35fGUKPEZ6Iw07Vz8/YLe7VCMb5N84YpE1rvyVB9SIO9+TyroIon
NPUMxvF3WyhMbov394yr4hxGPybpfBbbK79lXLTazuQ6ZWgT1k1Z7v4WojKZ+GMp
EgQSEOmzbiEiAL4bRgx+BidupRrP6LKG/9xFWf987a4k4LY4UN7LBbZzSUXZ0lhW
yUbsIDgWHHELHbFaN8bq88C/uBTqF2840oUyUke0mcuYEivySJSldtEso6awu2f6
730y7vHPXtn4f9SRkceoRnyMmyidiA+GQPK4iI+oBGOtOu9WW+NHDW1XrBTK++H+
LilujDuArjQfojjnuvxtK5R3PdrC1/lLplCIyo/AgoLmESk/u/mJLo9et7dNGdVu
ZLI+jD1t+G5d7fI7HpT7RA==
`protect END_PROTECTED
