`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JrdaRt53Om/xAFGKSdSGxwdywcAgsTa3ApvKPGcZWig/jME9NI4tN7dZchikHGac
/JG9bS9SSvHke+2vnWreRb3HIFN2R/PoCOHQMdIgonKgJkOKg50A7uQviQZegEke
buQfvet6Lv2bTaSRmrY2vuOKdIsMPQGmIyJ3MxgGOvr81HdBTisTdYO/0hqVCMq1
nNEqo76+GcTSZiCzidIagUg+S7vRdKUafyRQEcoS06fJsgXcL9Sqx1nbkQBW1o7S
WXcPXqhZdNvT+BerIDrxinJpbiYXxYmnYcnnWPzQVgOOtunxVs3KOiYOnIV/KMtf
qAyvy36BDeaKZXLK+aF0UBIrJdjZA1k84YfJjW9YnoQYgL0jqymXQPpk1S/u1Trb
THydws7IkvXC5oyow/W8CGVGPzzhp930gbwgLaZ7cT3zdLtgj/NMQNdePvVAXFkE
YrscbbSY9Unozzf1gVv1w1GQmoBq5gmcE5lQ+HFnSuDcqGJZLQWS3o5VbubY46EL
cFKSARrlzAYFPex14BLWiSAk79Y5jdtOI4LvHTZlj64bWt7i1SxVZEzgpCeTq07I
MJcPG3/5DfxOv9MhXIbbyT+LqRfFSXe+EqnoEHHnAqlmJk6fPiBF26EfTMV+aIXZ
ermqKa9bFcRLjqwDnBTc40qB0xuq0g9BQ/6Kw+REfl5dWLLWgisP8Xq+pHBcpTpU
0hDTXZ8oZYoHQAsVDMQH22bsoPzYnhi1asNYuDPUWp1VuQGAQREjhLIYR9nEidOE
VXulIxBZ7UlntLt1L8w+Z9GcTSgsfZXxcSPym4640+VBLi2qqu0jVXXMnYkRt5Jt
ShaeH/hWWxkiuUO8BVccrQ==
`protect END_PROTECTED
