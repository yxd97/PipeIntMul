`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+coyF+Ufl1RS91wT50tDeX3WLn1PrYuhbmtdF8DALasjMiS0wTXLn0vqU+aXkPi
i4vM5taWQL00f3lfhUsnDUlRzomHwH/4fsriltA0s82w4zH+yUX5LgLvnSVFURoG
KCSLJUgmlxK2LaZDEFIXOWwrDOcbuKA1QSRSOsH8yAtuBTontsV34WApMdVoMfgT
0K7wcQVTGz6QD53zJofZlg19+fXP4h5PDGzF/8iVnPg9Ptqa19m/QIEP4UEVJ6tf
YpeQoLY9LfWwBfupDw8bflhSFcf79i+7CcCUDz0UUv8q5ThPpQ2ZxGO9nbCeCKSV
LtDDoWLRjQcn/B7kBm0wz0/cQAFQQq9aiNau4vwqBbjtGOtn0HeG/zwRxLjuVzkP
hrJgbyxzk5GgHpjxpVCPU225euoOXBudJPqfBUJxNsGDM1WMRQDtg1XyMDcgZab7
++ThcBFFV1A1OLbwf57dxkP8Oz10ghzZOQ6eH9QjYoJuVMMHdfQXyyG8GK11iNLW
TILILSyBA/SKFjecELfg0jBp+bItTSjDq7GAAcFJzJuKEu7CNEcjoDjswXMPolTK
7uq51uvXs3GmCFH/m2139Or0yAwkQro9zz0UPxPMlX5KOlncsqh9XKuhdFxgNh4W
wLqmkmJvZZR1yJsXJUejwNQXHC8x2jCnxt3IfwiFyh8a+xLNPSnyNcEsGazurr1z
zwDBPnJzvYeDoQrkv7NcF5uC0LMma4vUbvGwf9BVz4sSsyCD2PpJUn8D22aPvUMD
jTyuJWkAiETxxMxOAaANtm6zY4PaiDvaMY1F7c8iPAp7HXUEaFo81j3JOnQXWoat
SXLFf+aINnvZ1MHvoT3XZrVX/HVEt2MSQz84DS8T36PDfTWbrqLpYMK9j5lLrYCg
ivuXDhGRrhIYtREfjuVoeM1knFosPnCZv+zG8cOQbGlfnrEAR+ia/gz7vyAepPG9
`protect END_PROTECTED
