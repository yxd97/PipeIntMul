`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2gwnq7WyMEXH7B1mWF6P/dFmXz57d/Chm/2066QK869XEeiGZTfce/ZLPMkR6KP
1OlH6VbzFLSmCs76aufeVhnRQlmbhIX536SZbci3RrXhT1D7iglKez2zNtDLFJwM
Ju5+QMm9AslNpz1SV6EXk4Qd4FFY/Y/W9+FtZMKd7yUdITV+VEK6stD9KU7tZpRj
NmMoyRlkbEERJUbJo7Jz/mK+5xiBWxe5RdDmkX86OuaUgewlpHHyPeRigXF1IeNZ
xhz2FWalhb44KbX+27j55A7P4lWDxaE2RlhGq9uKcxyWCsDA6Z2N2rWh0HYWUR7D
cZkBjAPXRxI2OcT6r8kAxRZLa/mocR2IJPnPKBktOpZKSvC+G7F9oEnjHRneulcp
MAsAiQn2DwgsuknCxt5nJt63/rpHePLX/cf2evmRAPn7sl8HIwX/Bgqp3gIb9+6l
`protect END_PROTECTED
