`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkchclBitYy/w7CECzsOkMynzhnJnIVDhFPTsTMCX2a/Zm9bHLu17RE9BMtPFxvB
G3MJpr7mrQq+m85p7mP1T1CI0plvCIryyj9CIMHNT45fN1yJsravZ+Ffj022tBo1
yUB8W0ZYfMJgZ041CdfPHJOJ5O23k0v0PrcgJu/jYfoBtvTmj60z8kIYFr9PuLMv
kELOf9h/zC2rqhDp99PI7KaZBlguybewHqpbAwtNT69Er5OoSSALazo+Q4WDmv8O
LPeN5drjHMN8AG+75I45gZC8vTt91GDZifT2jfowPaVA42zLCIBD2bZ2HustunCH
Wr6omfdgQNxCaMzk3SLnzGxqVWIo52bUeZwBlTzPDaxKlHrfgvw+HOx0wlvH42sF
pANH4VXrXvdNCi5apY6qB+Vqbs81okee5y/1OX/7U8oWNMtleoUER5HJSvW/XtGF
frKEbn8h+qMtSKc8MIBbC/B8YTpFGmHZBSUtwoB0H26ra564RrFGg4G87YGzhKgu
catQp/U6V+Ib8u61K6u9tFYuyv8CvS0kiZimggkLqCh6vEIH430LIMOsNYiUY3Jx
7Cob8qdlU3fS2L0+3huilxmCXynYV9ttOtIgWsLdC66+0ylY3+qM7oxJbQ1ROD/w
U4PJGNCBpD36O/JwO+rjOkCqmqZY9/eAM1ae0KHszz0t5/MHvftubjNXd4GGjnm6
BZkEDe2LDCwlSYF8G3cHwRcTtlnbnTH9fAOVyS8ZZIpyOCN+EZrWB6M9jzw29bZz
DVf51wiE+bw1DEOWEkIzvyjdbjz41tiiliKt4nRnaaPjzPHKB2hTyQRBpdPs/nI/
zsRqcKbZD2yRdd6WtusjCN/YKqr/IQ4Ozqkg4rjT7JI3f8MPYnk3NM3TQCCbGo1M
QGj/rrASeD37WabkIiS9Y9J+aVs9dCRUsmkvDXteAzL42vKA82NS+uNWMLiochts
ncsjuxHD78XZuc/hNo76KIUiQjyU1leivBv98jFT2jegl345FTD9K4863K0X3Yos
0jd2c3eAdJdQB0d4LvMglBWLK6VD6P76K8/4QbAp4F2sPtE9p8MEhnAb+b/iQBP3
Ibez8LH/HhPZh4auaNmF60PDAmn1LyupVA11vsUE6WUy5LIY64DxarYw6Zxabdm7
UKZub3O/TtODLbxca1ewVMU/q/rOWWg1s+ZUYP2lOcUSI/soIpfqK0DyJJaGsFEv
9Lqc7EVgdajzYsyiL3CB9+S3bLCGPs62yDsnsFr4vC5ETQoc7JuMggZkRi2HC85y
D7gpea1RgLfN7fDRz96nkfpJvxYcQB9lVriQaimBLbwdHBO6VoLs9eNqmZeJU9Q1
WhkogqnriLZ6Q/ar6Uj9JslYVSMrphpPffcvOqi0qMM4xb5NkUv097+L2doEi3JD
zCQQ/5Ov+4C8z/rcaVz40wD17tI1TmB79WgSxJikicPKS6lPi615MMQpldCRf0du
9JCeU1KnBKkAF524fikLXHhEO1ciAAXdrHUHTPd63jyObE43e0Pek2B2vycAVjDN
A7c1XogpSp2m7qvFxsdtZ90XutgxfSImjF7kzQtCEscLhmU1UDrP3ZPjdKGq4PCa
Wy6KBaGqH3e4cf4qyaivg1P7mehnbHfaPpxdDwakt42KhtpYuqmPP/LIGG9Vbnpa
85S/UBnB8SfUBPH2Z7+D/wy40EuVRDLZGc2iItLoA5oocPrwy+bThGG7aYnXU9fN
MJHIjBwtCqAwMPPF16ztSA==
`protect END_PROTECTED
