`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6TDvQLOEi8g+9bzp5k8NbbNdF6wG1z+TjyIuJE7Z3ik6In/jGUengRTt/8U553f
V8rkwE5sROp+1a4lHTMHnaNnS6rrBpjHO6YzngXYtsvVkn+OHWalVxtRZAGbFtjI
WORyipdXrf4rF0ngv/kIufkBRFwfkoG9iyAg3HmOII4DDIjzwtcRmDU7SDtzGISF
b2ITnbjaQ4+4+Goz0sAd2znVpSa/DnyqTxaLR+DLZqa9hk1ql3l3dF5dt/q9SMDd
H9R/pgpPdzNgYBZbZH5AP0rswckFL7f0T+0jcJSdjsQgbZlVhO+NgVC42TeHGSPq
`protect END_PROTECTED
