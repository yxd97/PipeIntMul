`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYBv72rHWP78iZ8kW6HU6BQYATpMYN/DLWFT+RJdbX7NrITcU+5IrMIPVEX1eByF
wK6tNDTIbjo4X1LBP9YNM1frXHHOD6XxIB3RV65Z/NW5cZ8TmfhL4jcXUF6f/YH+
uzYe4jNqeAdra1oBsE9+bJ5dUDKlXzoYUhr36jejCqK/vPryK7QV2wkBSElR09bY
ykg3CYPs9Wghc8Aji3eTFuC7AWN+Q8Thj1kyN42IfBbigK78NvNxBblPTVaK8JeK
trg+SEQf9OIJwZqdlZxfA0EQVbOuuRqwRloAraXqQbYBP8HB6dnE1y45dQJ1/CAo
HMloCjY+yHQfN3DtKqX0pr+AnH8Pju2I0M6FMPQ9N6GEQlBeZyqdJ+nA+gT44JyU
aN3gjLG3rVcAegpy3H42zK2MjPANBVBkmB5gvtmFFs/2MIfYd/ESa0RevEUgysKr
VIs5JcN/akYZb2d7QZTw7MeSTOUlT6gYJ4eJJSWw0IBWnkjDLOGSwywtRqYvcKN+
w4g4QwP/wdmbw6PtksLcCtyteNONzGRNxk44awq8Fp1qzaJju1lrkWYrhX6iQPI9
aCEd6b6yXVJHWQH//m5wmJ1riPzFhPKqiKhaGG2WSrhXy0wDRR4nXFCIzJnrMLN6
te+85GF0jSxSKo4eICRW3LxBeRgw35uX4g72Ut+/oaWgk/hK3kY5lmUqfycU+N6X
FXQQKPHrfaQuJZL0WKWi77nkNFzBFjFan5x8pA1CK5NJWOdkEdGDCvFbaq+vjp7D
W/V6+XzaCGwWDBkaTCXh1h5f1Q/z10PwmIWeVYVfSl6t6BW/62DZxrUmszQ9gPIL
6o/O4F3BXM8AkJoYc9kDV1MHTjSES7MJLRdF+bb4JCxI1II0zm2rusmzVrlE+KqX
b8FVUvoKgoa9E107fhlmSAvn2UHE9XRA466LDT1c9e7hK6aIILxCLL781OCngO33
FenrP3wbvTMNQPfFhOnzZaSa9j3yUVXCKoKVF3lZUlZXm7P1eTyJoLy9PS845X67
Hwor/nAUqIauhi3HPkzSf5gzFQ+wfQR532vdy1II3LphEzLmmTusW/g53GJAf1d9
NjyVfJWJne/R9DBj9xbfcW2JgtI/FwVzQecMwtoYKo4VXMik2WT0l5fCzf9iaTnm
YF6d6Wzg2sfMIUwrr0MqszXTpq3X0TyOy5ykBKfWzTXFCsfNbrVfkITwC4AWymF7
pvdgGlzHoceuzAu82vxll8+/1NQXpNV+7WAtCAmncURal0KyCguWzSHCsCTfDFUG
`protect END_PROTECTED
