`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SmItng/gxIDCGdYtdgm5k41IsFEe+AhSNj2kipYlKX14y4QqdbVrpI8d5pFxc/tA
8imgiMV/BC+AiKcG9RFwe7An+EM+oLrRBTCEZMyN1VofokKgfXXcf4JUzFHudARY
yNja0juI3cAEtqgPfnyqu+yVQYGuPvgFVVwln9YX9i3EmmqSHDeVAp0nUCph5mqQ
/Xa7ic0AMiquRSfDicNQvsUJ70vTbFqxl+paWceS0JoiTP4kpqp8p30YChahNiZH
RAjdmg4lkINAD7DKytrQAjYID9G4/AXuRt7yDZxVhPcTp7O4An1b5L81cG6hjRKo
0UZr4WM4u0FloIHf+y+UzB/Ik+G4ZpsCvahR1BSNmponWb7zRtoLKGZsgZPALNnc
30yXlUnkoBJhxgu9E7j5A5gscJcoLLgFPbWTC+p7UNMlOi7sD6f4aS6c/MUBOW14
e/lvD0T624kONZtFqrO/JFugtJ677aSLiNrG5WT1Ga7x68YdKHXiImCGIXirEi4b
3bhA/sImiAkQqWIzMGHuB2QANnVOwJOQUNV3ThiJ06J5Z67rHyMDTuMsC4/vVX/A
xA1PpnSMOJt0aId2yARwQYiXcxt3Hmijw5SuL8pQO1EdR5rz04U6+ARhFvDKjPX0
TSfdrB+F90frtHv4o88W25NVKEqii6kIW28ZgyxCcw+BZxusEZ0k6UPBuNgwL2uN
QS0ws1hmM81gjO6aKj6g56FXl5sqFJN0MMhNoJn1bs5FunLCcICDHGAI6eW7DswF
GAefJlPJl9JlxhmLMfBcvnZKj/J9oHz9PsXDSPIMbMv2XgEju9HProOCmlVDbHV0
Z9FNx5J+KqoIvJUzhODmle7x4AuxnYdRj1rFgeV/Lo435kmxPERPtszVp8bUS/vQ
AdLG+Xl6eKsAw5jFBSniNfSi77g2/u/3e62RPIYXncQqhnHWbQKrOC0mNObIYyFW
WQAPw1n9+hfc1DYW8GbqqWfiRDuwsq7kvE5l/u2v7uRBa+00q0sz2e7egH036zNc
ZBZzWCaqgN3Yi2VRfR7qErvgcAFj7rYDbQ33TYjsMX97liY9hMCUGDMwsIy5Cav2
MyA86lPtn02Jf4U+kVQ7uhG5o3zJ1evEPtOwAOy00HpOpVCJJO6BQWpPfLDxVbBJ
`protect END_PROTECTED
