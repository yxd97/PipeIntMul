`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lbQdJtoPGFQkLpBKbIjTggqiwAr+asiEdOpRTLLNp+UJR8K6UNPfolUp0xxRgOE9
PCUJzFLQTz+ObvnyE6ipTCQ6QLhp+p+9nAdK0C07e3wZWsxjskr37p8NtvXsjPCC
dh219f+tr6yG6FuKFI8TM5keisdYha2xTwdSVPKVFnDtzBjYmMuM7SogQ5LYIbey
1l591Gy88nncwPEWtm4opHfz2R2bdzvFW9KTpQ3yvsHTbmqeerZzzKkw5COsu1ba
gxV5id/G2hbtMGIDaSURc9cSIKfy5lqhXw1clF2SWTBzt0dlIBWhZJJkahxBtXhE
aagPKfcOiO8xRZ/PTMjUGyD7GvBT5U94HE2R71IBiMVCvMtQ7Jg3tSjc6gWiqePt
Z9+dwGpJkHIUfU/ZziXt9A41MziFTb2Dgb2YHuiuegeJXztvYODxdnNGlYo96PwQ
eYiNeq1NGLezQRtbpDhSgWYks9bOSOPFz1rq72f1xk3Nxqn/1lw2zKI9h1heEqTZ
VUFyFZgOwwnxTuHSorujpFTHn1K4YZH+POFG+fyIy0gqh2D/mPauKgQR6U66Boxv
gftKBZjCRghpx84LqWsn8XEyBBXibtHf3q4pvcchm9B8qsMWiZW4gAgeSuB9Ksza
YgEuXfHhjSrANrqapR6+kKL92kVQDWedFGRAfgG6xNsDML96p0dkwuhkG0fYlxvL
T9t7nB+m2sd6XtUP1D/EahaW/+gXvdj9YikoyrSWi6PEiLNXQglnEopCpuvRtJIF
nrOa/GEbHbWY5M2szozs7FC8F/MhaLcZhzxkgK3bTEc38KIi6xSon3dyW1v80eZJ
9sMGIThlxcqrMrZ4XISUWEIz67awnSCNYeB/yvwg0A8wxPukarE9pI3cYIqGY4YQ
QPUBpAISz/gGN9H2hNDFyRBv2Nj0l/1FReR0a9qcgHe8qCf4i51wkDt3a45GIyJr
/C4nUG9oxST4qc0E7EwBKQu++XZNbALhnLoCc4mYtRjegM1mUlJoX00yHhwmNdO5
KmZZAtU4C6P6asRQNd9qQlulYlqro99kajgjWlhQ7R36MWbp5Ce6TiSVZr3C8s3s
hyS4qbrG0WDUA3GwczE17pDo5IIfF9Fz7A4Jc8/0J0eovnSaJWuUc+6gboPbM75a
E4Nijv6QUWfcSaal086vsSZIhIc/BZdoYu5VxI/iTrZ7tAjmv3WQrrf983eAVCO2
uvItJuC4q/LpyrJZ+i3gtPpCSkrI/6zRJOHMpVZT7zu5FvjAvSZvK0IB3xmKbHe3
`protect END_PROTECTED
