`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfXd6Aiu0DkOMYeMDwtuFApgKRYdtB26SY0zJlppKJeUWEsWdUrVRF+ZWk8DxgoY
l5w3Sk6WueZZyawG1t5wGtZ3goCjxMLdKf+z6QtOZgXsN1fI/ERIRn4uqLeIbeU4
AllXJvyU3GEN5fo7YHu3SOe96v/9SJ53r8RbMwEO4rZSdIpO7xwSHHAvJkHLBD6E
0aXkuLLJhGYET6G+QBXAuvrTgQYx4FS6y3wpX8DRSO1uy78T5LfcC0BFdNnDdd3v
lAIFYYtMjCfcOneBaV1RCyMHZaUB6eOweMB6xysMJwmlb+O9SMmjF4GPlmpm+v/0
Jc1saJV3X2FOpT6npt7OBW1ubvwwON6sCz5y5mAJpqR0bEIhOlnkONRzKheouGCN
jh673RnY8T6vp+c2r1f/eczJpPkjBY4EDzOz1HWY2KSzGn1MRvtRspNv44pPN7x5
Oco7d18ZQkanM/6bSnQnal20VjI/Jrl1M/TmjPLEV07YpRoRe/3cWN/uBhTHoVjh
UyQIvmOdFrCR0bzy/0tx425XFGyEhj7fJMuN0CsvcQVpo88NfQs6X3X8tXUsTZH3
ZNxzaa7PhSOGYXUFWUwC1+hAhG0WAnyv8+OBTl27f5hkIUkaB1QfasFywcv7g3cH
fdqreCZZ0CZ/qbwaq+c/Odz/F/UmtUZEz0k0zXH1OVlbxTG1KPHEldzjScQcVWX5
/rtg6LW67KY3k0JAM/DvI50VA2gQLU4nuVnbhATYx0+MVSwRY9I2uki8Pjqh2pM+
rAcRTPDLkU4MUpAWS87KhdTvWXDWs8hW3yNKPt7KeU9DAU9diP9z6qtAsCXwV/Bp
YDHM22QnHRbsIxg8P91FVSnAdWeZCgn/arZImQl/ntbVrjg7jhWmrJL8zb3N6D+0
rukTI0plKmvyOz1yZT+j1/AvUriWHfG8eL+mScRZ33YeEvmN7xrYywGnAi3nljqT
Me947kU9nqkXeZSmviF+UV4LnnYqSCOBqhmETEdZN6DXRTRDnqpG5UbJKte+cf22
YcSezOWBxt05o+24BDfyqWXtbHvRzXYI1L2pCQyS7fqUxmkwLpG05vRH9mRXj4og
/I8I5u+RKjSxfHrH2YSlofwAvwgDB3aY2cztQOputT5L22KfqFsB6ycs6Vgskutp
iS5yanYyZ+ftTnIKs9JHb4yENnrB9j0QfeDzjmy8a6gl5iXWQ19n2H2TZ2jDx351
IC7/cSJGwDpGUm+FpNDGKjH7lJo9FuP47+vKRBudnIp6mWMM99VNNOx5fwLwx6Ng
BQPQWsiCFRywVrDLp8VFxJylcqlqHB6tnlVfuxUt1SNNDP42SuY0aOyv59052LSj
cCTX0fkB5EaKya4fpyTVpLaVtZ2lUG0YOU+qMfPoP7MN3FSirn64q0zzmShcGiIr
LLB9kX7Zugc9eZTu4VJTYbk8P7Q00uAa9SziPxuBNwq43Pr0WP2r+m6tp+tBMyLL
sSH1iamUgoZSvj1+hrHexINsHltCRnVkPtwHyEYqi8gMYowyRuMrFuDvkaZq5OKI
PY0UqrHZ0P3n7/vFPCgeEBeCS8kp/DvbZz6lTA6EfxC77Sa/Pz6g2vFGU8SDQloJ
D6jjTEpAnv+5gLDWw87GmmLylQGishcXevlySIZipT6F5Z2W5w/OCzztqMIPGmT/
Apyy4ihtPwVIn/Nw0BzBjrPC3hqwFuVWi4mdzEi9LIQNy3a3afRHDGi4OoKqelAC
yvYNzyr3ML+XIQ3gh6cakN/5nWTMABYY6CuOEwkfHW0FAyNGAWwQ4+Km6CQu0AzW
VF0/Xy/P20lXJn1Sh5SXbMLZOyYANNwulxjO2Nf8QgKwB69TYhyqOFYIC6qTmZYY
f6KehKp7kXyQcI/A0UdC7wr2dp50ZpVvJfXGzTe4rWsnu3l/1i3/bscZPPweyczY
5Vw6nUzNnuodmzXep54ujIIQslinF4F7Gm8ws9PZsUN9+oZBNB9P9AYzZBPCjfPn
zVpLp7Kjrvq1+6r5jrg0S9ee/IxD1V0a8gkstRpDe6hJMIh0l0nvyRLH00oZDHp1
tbKddo3WR7C3/v/N/bebMLmwKMKzaUfVjlotRLEOtoMgPfwbbEbVD66G6a6y2TwW
7v9y4tFzyIWkOD+0E2/wn1tAb+18PU/M+zzRo1miAqSwT+v76EzAI9dk8vVyPDz3
`protect END_PROTECTED
