`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XutE0a97NBrzWunkxD5v7QXVbECGF0UuEX9QmHma1mvcpM0rcht0qfLwiNx2iHpR
HT7iMjQXnZwe+AdF48wslNLKoJlicseSSPX1Or2OqzBT//IucqIhWKOSH5ewEWx3
oiBRuVDoWfFoXQQalKS0ITKcQ5RWbxzsOA/3t+dSnRRXeVi/6G0lg8gZ7WxxV42S
NmwVMAj+XXTQt/sdw5rmtweni4g9GCzxSPPGezC7imAqtD76eZH9CfJGsfyMGgFZ
YzbHNPS97QY0eInA75T9Mg3lmGSxTy6Wu+bFytC5jC/MDa5TSDHK7THQ4rNw9DuY
TM30hoZ5a1fpLRYC5dXCjTdYZIz1ewZRCE4oDdfLRFKlriulmXjT15kTe39GspFj
yxPRslKQ3JXzLmXWQVmBHoS3GF/MYZKCMGfZ/qXJAzOXfqGVIhJSU8th7JGyc0NJ
WvubgtwKjeUgPNQYCL/TTyb5+Hqk4hodZmqB33qCpPQTcp9W6Uj4tBmyvD8Sy9FH
8BohBMvdftl/44AX/txc2We7ERUWeVeCP/rINs4pALZmv3QHdR62+kFMJXTM9NMV
W15ykUY7yooPGxnrtqTh9A+3e5FMFjYfekUEh09wH9L2Z+FWT78BMS3B0hW2RN9B
0aqRU6SxGN9t82ZNPpnfMSEt6px8xjPcBHZ/nHCMX0BoJ2Ack4Oa+e6H732OVJIT
PZ6+ev/HJALaZPoYORtcgJv1y0DIqCsOaVZstMRsfo3ctILKmx7TsR1owPSQktfN
My48n51HObyhK+ABwQMu3aNH/g3vEOZIlzOdsTABRPTC8ns8N4vQ4ff4Y9leLqbO
CQGuMunU/tRnf6TpAjEhuAa8rpgc6G5rpnw9IFS+PXNbUjbp51Ua1N1103eWO8vJ
xhtBgq9tChzeavJvWd/6YnVufGgmBaOtuTiBWTrT0QZC4326ZHDTE7IPczWkcUCz
D8+F4O+wUACZLZ8m0f138I/nrdiN2r7OW5trmwoa18l0SZQzulJgulFEQG+H/IBl
SrTUyKpODIJUwaM30V482EZPDmFkihlPcwb/RuwgOZOdXf+girTbcdZ/UHq93leQ
jUn4xZmx3iNCB5agxpLQ0WNn13sd9vGU83iLkTJzNR6oid+nLBJ7kcfSo3XvTeE8
`protect END_PROTECTED
