`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NaCZ77ce8YBI4XALaevugDcBgu34PO/Kob0Ryk1TVrjsAyjCyqidzw5T/YYeHr6I
njPFX+94xnrEftW7jJXTVLmXfnsWUnxrHET1wSkvbArOFa2aIBAvNr/QSQduTMKs
vNjqs1rSmMPdGva1zpkFN1fUpdXqhbIOqcnVXm7rLDqaBNtUfDFrw6DmehMoCl+r
hdhiaw8Meu/l4+KOXlPcHT5mXXyfL2OUlYkmRrUG6Mx9RGQ9VEa/9T+TaR+J3kbE
UIIj3skvL2C7SVXO1vmbV0qqQlJJT7U6gtxrXi/RNGlBNQwXdN4QzDIwF1pmDOXV
KmvDRnUUc9Nb4dp3XvQ0DGG3GD+sg4fVeJGB/ZYauA8StA+xescn7m90nzojDI0P
rlCVrau3zDAI12N2FMsg2m75KuVwY/VQ6tSgEKdBSoQPLY5pa6YCSlavMF6KGhlf
T5Ij8ndsdLLD4pRIqiKTfw==
`protect END_PROTECTED
