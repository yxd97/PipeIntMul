`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29PByuEXiRpdFlo9s7MlvMwd/JbQFr2ozJbYvl91v6yKbq3qBlzuwQ/AagLh4eoO
L+YSYLcJmhPA7/uYpnjeQVKyWpBQBg/UcpQ5bzgJZa3o6FxBHOaxWigwhPKHzXah
o2fa6Suk+IpGil0re9wSa9tw/dCupJZ6vKJarln4EnWDqD3a4Ps9+m4UbCdo2JYd
ViNC16i8U56jkfEWmPJH3lpeRso4xjpxAWT1G8xCh1qS9LEsFpqP/DXNMURPPK0U
WWq/tGKFQ4E74peDlt3EeVhGFPQ+R/UmwEIkTAxQqhPjsuo6wsNI1IUpKVDfDl9N
BQGHxEsgjp5cisu2qhegThfkN16yrrd0sS6mZ5LmDkB7oN5mus9Tq7tC0M0kHtjm
i+F4qcN+rsutq8nXreNLBb9fViD9ediRQCUy2kUTfq6BgDqSm2/QrdZiy7jDIsC5
5wEhuo00N73JhAp9aydNKdsAQeWjPtWa0End4/3GZ/gRkPZxRdAWO1Y3lW66G0GW
5X7g+1Q6CYrLPZb0q6DKRuI8dXzd6q9ff3CtASXRZIpgVCi0K88TYIetFTs6DHfF
8YjiriXEyv8WM3nzIAv+k6l9aT+t6/7WHWpA2gU98iVKZm4O2DOEHQHKKaiVwa3m
`protect END_PROTECTED
