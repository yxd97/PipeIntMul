`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99ornGciDEaFYOmGCowOJgeGOl/S4pIXhTYigsbJ1JD+PuZbBjYn/eqB0NNJzvHG
H2BFOyDtv1oFNr3Oa7QTrDpZPm4ik6mXgAagL30T5Mg99PQA2my2WJ4HxmM6yAoQ
yTqlb1Bl4J2Jik6Xp6XeiwfwZn/1WW14kcIqgz/d3GG/m5uKXmoClB6EgG7MTjFv
LG6jx52w1re7iZdcG0Av8F1hDg2xkcraXDA3cWjeUwkNXGSbmt3cPuzRvotfnOCP
QiRo3KDnmTot+QNBUMy0Ise9o+B1Joyyg08CI9vdUY7GpJmVFaUWWu4lq3EIQQzM
DquozROb+52ctN//vYN+m8fmpAY43v7Zcj/l5Ac30mlbRpcBvBmR7544rjQgzJFg
`protect END_PROTECTED
