`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XSQsLSYDlOBObOagvNDNp8zzBjTrhHFiZOe5i2QcZ8RBEWgUyjGiOOJX/LJn+of8
83QS+4t2OtKzgOraw71Q/SqE49aQfg42F4Ny+tePFMhmlQjff8VHO7Gbdlm+lz09
EudeQzZq4liyMH2ff0M49Bny69AE6U4EeqUg5HOmrjTdRpiOytscEgOdSyxlua4U
s15FtpaZzFpLAPMYnw/s5krZFSBTBc7cIPtsBYKwc4UhfpsWrPo0eakWqmGhFvVX
1IzfHoNRCKYOQdnbat9WL9gq16nnPSwUB2+8ea5Hga8=
`protect END_PROTECTED
