`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09vpVg5esrpT43tqNJhI/ZZv31yBxALNpk7k2gNrZzje0Nj99au1yyEMLszgVqPP
BqfjV8izDC+IP/rZu9GVTd8JJbTsWW5sYff7Ik2dau+MED9blOpKlynaWIUPnrnE
WAIb9KFkoUJpSOR7eULIMDXlrv3yw5uLUqZb/ZC3x45OjVQXUktfHzWUmRSSh8k+
hEeQIsCL1dI049XXpzsW4wOvygzcEw9KvZ5zHzAZKQecYUpKWC3QwZhRosJx0hly
gQwkeDQxg6xl7w0gcxAwGqdgYhau6jRmuV1VUp36mVCj+u2iauFmfA/32bTsEIgT
moSNTxuPTLZ7fBL2SStn/1FXCkzUTZ26cZ265eljlNZkwafS2uVkHOkwVsuhf1hU
tiZjlU2wMxPq1MTM6XzM/b9DDoNinHe8d271YfmN07yB5NzribkdLwnrtM79PDl8
wnnG8pjI7AbP5jcG1e69OCaHStQ6IWx1dwerEm8t6cRUKbIm/XYvHCgANw+Avt2S
qG7dB1flomoaB0eqGX7Oe6TEot/XSiZqQ/3wT6fucQ4xNthm7ApCKeqn+rQZkmN/
Pl4kpuvlpQP+YLcYXoJRlJnfG+DtSsxcvTMjJy2nYppoNHwrBAC+t9r9iHoIsvst
oT+p3ILdWP1WPbdTBJcHIfOTRSBuEa8hiJ+4phzoUrCm/CLjJOimpzkmJcRxcjRv
eCzNNzrKLdKtuiQ1vi3KyuGLEmsJLbpa7ILWwz8/wIpkfis523Fu1ujdIUHQ0vIL
gZvAG73EZKyEOff71nh5DIiW6eoly4xxmUBKH4/YrkseECYWqnCkJY1XPmYBQ4DC
erXpGGZyzqABF3CIhbLs9RrCAtMWdW851jtk0Y5Y9PYja8HJoPghWxQp9KtnqbWh
coSoVuSyTGkli+muUmjaMZ7bJDRZuHvpohQFIPFBl/kAAiXSrLbKUEXcaWHJi6K+
6kssnwzlpHzaOUFJF6ERUmB3dAe4xpoSDu4d5A4lN29ZfO+nyth6h1zGZSzL2EVT
TeyWpkeczOZSlRhcnTZch9mpOVwcyIBpswXkGSkcfX3VPNehyW2ZgkKZ60OGO7fU
0v/btjdTLeOS4SUUcWXlmKzS9vtyEH63+lXegurzhvpfwFX0B2u5elXWfrEVa4dN
2spKhnct86pJq8iJyfmskzc9f/eNc3Th+qW/XgU31H508Shi6Jd9Tw39oxro4OWL
CXZy4mXg5rb7hJNAlefYgHIeS/ttOuN0BRcLtWtGmOl1zFmx80LL2R78+AUK6Shb
wJmeEaWR+kdKGpGe0CaNEjG6WVScmaW1kOxNVaOmbYIXxMtWShyhVCamb9ldpVeX
n7uub13Yhjps1KxjJDt56LdCfF7kRyaYpM/mLOBp0WvLPnsMzQoqVXIo7xvoMBC6
cAR9BOzVFqRrzMPy5+1ROsG/9X84MW94o0b3/E4SzITQz674J5QVS9PQWckO7TBp
g/rLzELzXlI1Eo3bLn+gAgrkU0x3Wq49sre2Bz7k0OQaDqMRgJ4Ufy7NNmCeXHnv
BRqwyx63tUZ/qoTy+Wh8QtAWfe5bW8i/9CrtYu+iRNczm3txB/89jcztTGE5dsww
g6vc//QOrEDUlfCD+H1G4F5ssXy86Q8AQU46ClOYgiY1BHd0qo0wiRYv3yUV+Oxo
`protect END_PROTECTED
