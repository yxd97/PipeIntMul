`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NDIXrs7y0Oty5/4lVcdDdpKgrZ29maL6S7ydEsTz6FYAn5o4SAwDstr+pDY2phYC
v6E7nFxYwRPwqAudMohsTEBNEbIe5xRrmOOQKtaEC6uXtIqB6/vpNiQP3Pwa0CIs
7/yiMsvmg1MBjHxg5t+TVoN1bSeN0zYBliIDKlnM1HLTmaZUZUWinKhFeEUKEUO4
In4YcPHDYS3x9/tJzdmRLVbUM8vPyKe9EPqZgchEgHqedioojR+Bua5iK+M8MxzH
hOptoYprCNW3IXTl4N2DD9z3oBaGb69LTOPIxxM5ipo=
`protect END_PROTECTED
