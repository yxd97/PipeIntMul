`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RTJ2igQznCYCup1cwPJDs+zWyQS7KNznOM2BBjwK1hgzTHpx0e9hFf9QTX3kSysA
kxwqN92vvvGarBBCxbP6WPpPMf0839xDgCAr6ZLUC0LOy4CFUeuldkVxKsc3k8nx
ik69YXuI0zlasqimSm3G/KzBFVxkEqn8Nzpdm4q+uUMcamE16+OOWkdwALgSymn4
mfGl3dN7Okorx7u2aquThCnld9zF3TqifPIzSzEH20LupbWwzexbd8BBiA4Pjg/8
04WNOoHIlszQsu5ZKGZCR8mjN6YwD/b/q43otZObOEJm8bU4IIgPfKqOHKHnZVpV
t1VIuLCUk0wSNgl2ckaN3F1YLpdvR/BjheOC/4aukE/u81pgKoAdprLHP65+wRE8
JU7lT/qVZwEflSl9pn7vdXShIaC3gi/q4MRuQXLPta02CsB0iaTjnEX28ead57Al
uI063kwihB1IVLfMqgd82j1Nz7e9LtxoNK72LBOPuBlPboAhD42whIDwLW3OxV3k
IkL5/rGdHKo5lgaB2dA2DZPny7bXg5EoAWSUVarxGDdgyNvwbrY9nvRQv8IKmSvf
gORYr3qC5Bs0fJEEGX62k5ry85SdTTMFekKoaOG5sDt0Oe20r67a9ekTWo9lfrBL
8SpQC4JCI70eZvHG/MDoln8uO638VkmBVJa9fLFWoZ7+sBRKxDg73jt5f22H7ho+
qLFaX6rmK1XFs+WPH5dq70kqO2T1MJG8LFZF5NB9ESNIAgSyUV31eMrIR6jMGsZX
nhJjoPD/A5AOOCgncdI4nNcZekAg3WD61wTJEk05Dtg41osKI0JTZearwKLGJgur
h6Pq5CKihgd74RnKSK61wakQRWAO4EavYRUSyT/CcmGaQjyEgLi3R2eS9m979ek8
wObhhSiwDiWh/x+A24+lU1w0CgPa6V6DRUx+4UbwkVjDKMB6EcnAacBJJpOppxMm
kNPZryBl+gbu/TTO4UL1cGB6ZyMt/q3CcgnSVQj+rwOvpMpcOqxZyjw0ar5JmtpH
CX0DpVaxmmM8EwIuqXDRq3SMljuhfTOfKVdPvnH7ZcdLXNBTDev3fPmPIMyRjlui
LqcQtZ++5dyaFDC/zeC7e8H7O0zJTMbMf+B7BX4VpJphOjigvF6v1Xzi3SN4O3Xt
qnpAHm2QjPKu/SE7l33d+gR87s+3sQcOOLIihVeqfJe4RN6VlkyBDi/JNQS3jNYj
Ggc+XBaMLkEd0Uz18/bCl1J6YLKQqh7kkGH7DgrZjIiCa3lMIH7vZ5WH9N7bCH/w
`protect END_PROTECTED
