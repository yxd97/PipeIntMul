`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLULNpgmpbU/hydu7bIGSAjyPyxs/iXgcByeClYQMUbIsyqtq6uzfkPzclCVu2qT
m9KdF+0QXpntx2ENll+1AbBamKoXDvKvD+MKDssAWA1h8AqDeHUiVwEp8HGR7vEo
xWpujvh6CJNZFvwATA6j9jVJV1OffIel/fhRsUHGyRkXVo5sJ0TBXgr0cv0AG99I
oDm47VnxNExv+cLgouBcLCCU+8fr90At9y/44JzHABdgKRz0LO3PlVcG2l+SeRBu
AjHQG+2nKhDILfK+UDJBLE7mHdq0znEljrp8dJpWA30ZpHa1sO+rI/PDRocsxVxW
dq9eUmzvEXXQHo9kn/6GqAeO4WmStuUSvkLa5MFn+bArbt6nbWsrJsMzm8rmcp0q
AW7+VFE1fWpt5abawbMAh0vgBNT4lKuiv9TQYB+VgcYnkQkmYr8ZXewcli5wNdQk
9xWeehyefgDWvp3N0X16iN5wgbxsFyT5zchJEuozTpiu2uYZ6o64LKHFqRFAzdvS
gPkAdd0IChGYAF50Q59bQsi0LkWFK0Cym1NFMVahKOLdpTjbIzVw6n89zp6rr5o0
ATzKJSloT7xnngxBK+qzGXYas3fNx62wD3e5VSHu49wkj6bEErKua2qr/oPRenU/
BQ0ByY58QRL81DhkDevE0d9LSS/smTf0jRmgDuxnFTw=
`protect END_PROTECTED
