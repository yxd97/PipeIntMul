`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYLHUApf9ZuyEvI9+fkiaEcwJ/BS+/ju3M4o034Z7+sfCotEyr41UvYnAiy1Tmqj
mnFrmMqJM4p05S+AH8zVKMkd9oDA7jtSYsZpTmVeQJJV+uyw0fuTpx8C4FvFjItG
cv33SfFIV6XY3FXE+skTRbGdVOABcItL9h/W5wnqXsI/bQtfnVRRW6aVlo+ublR4
KjELfpnyJa3TNrRBW8lXHHiaXF2BjXUvvwXfF/CKmMmosGgCMlg0Ht374zCCzQYt
YElems9oVa+J1jZcxUGlhWnGUMdmV0KIVqHOLusK6KJRU30jweiICmdIJwG4mruF
U6bDySFgROvJJCiC/pYV06nU5Pshgd17TI5OkkyGaEQ0JvVCdEqhzCI2XOJLzQve
Daur41Xb75GqT/OHtBSdNNJNRcSpnw3EY7KQ9KGs/OI=
`protect END_PROTECTED
