`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1lAsmuRpVHaBQRHN5M3w4HJHkfSgtmayTmTR7bliorO8rGy3TjVAmzoLidwPvrU
xB0pQXXpdHnE4p1M9yzdsXu+EeN9pLaxFfcCVIo8u+O0yL3YCeWA28dNMRugbiDf
NfAFi7HljMfI0mlw4Vok0elk/ph6b3Kpuhq9idU4eQNTy9sC+JxMwJu4Jf387SBT
qD3cGKrL6rpptMbycvWjtZ4nvzFJn8S3Ss/3PFRfjS9kTNqdcpxh8bkk0hNnSSp6
/kL4vVixLsJnQqGolpNK/iGs1C5EVA5eSXmaeuHgaGTHhIx9ephWE98Sr1ehCvZE
89ZUuCB52fraNafzex+FeACiUgiK8Icbf9aDzcELcMSX44Q9wr2r4zTpGCFTILri
`protect END_PROTECTED
