`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5p2SXjZ/xbzQbRe0w9lX1sCxezLktSkNxDT+tCws3kQYeUXzZdeacJLBbyW/bzz7
EHpK6PYu3g6eDQNwjpQrx191Yx+Zhn+eFbbfXtVcsBxBbUcf2Bo0j7LKOj2qgv+b
tKoVcFkHY2tU3gqf0PRXqE+2GnAugZTo0ViwcsiURWglyHvdQSLsoBpuc7jR+hH/
kueMeV2/JxuMqCMlpyt0M7b2E2UeC1RI+p3dTNfRrI3CIdkUs34eK+1Yh6R6QuqA
5sRtiExNvm3lCDt3T92tPLRdVtWMcxw3oj1sVxK/1m6gxObNFPRDQ2ilhpmj/blS
/X44drMiapHmlx5ub3cRj0zmstyLW+hjPeMK8MEbeGgxFFAELmWWKzf5N2FVlRft
OyPue7ehx0rauQMveBejjh8749nCjIiwPXUjs9hiw70=
`protect END_PROTECTED
