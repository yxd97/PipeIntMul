`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MAQo5id9v/25h2ol8xQ2YpQ6x9D4o9EFhbsqBM50A/bphcW0h4BBPuymJCGVyP78
aXZtXnl5ivvEYOPRc0IRgPf+7A7YpqpKDxb5mIHDSgiGiPL07GP1eQgr8R1rbSry
M4vRmemAuyhdhq8Ak4rcRKI7YigxCpoKWom6GLQn0gS+oGX+e8r8BDDYX2CJ7RFR
rR7ANLzX2quFLO5DRWDvVj7b0DoDHCDIrNMHWLp/RUt/E7BnPXZJ9Gvb977OoqL2
i9+1RO11h0QSjxZfRk1GtYEh9rT5s8/ryWSnTBl3/jg=
`protect END_PROTECTED
