`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXjAfH//f/ihPrDKT9wR0WxDbhAFDKeTxVj/EnQhQ29z8YmrIqDysZZLaYRAxyuY
iPDK/1jFiRv5jUvJdWiwFk/bDiklvxPsLTPTIZFvKattfO9sly4+2HH9LE0ne03a
uYF1ZWxv+xeOcx0G1lrBa2YDRtQAkkzdCucwYv2RyZy64STFQxje0V+p2pW08C8a
hXkUKYC+WVdvCUMQgC8MU/3zJPIZNNGJlrvaITU3TNShxr1mP5Yqcs9EysyNkcqR
9JVkLXwPId4j10PcNNz2hG38rPyo65O1c5WQLx6Be9Ij2vAgbZbxMI0iAgl0V7dk
BBqpHh8EQlufh/KcUsywnpJj1eYJdlvaJTl5ymjQUjD8H12Sdr0GOd9FJUTXLZG8
c3TI2upkNb8QD5xWlWu7XaJAOLH61wOeBZ4uSjg6XOicg0101JF2WtW4uUjaPl0+
g2zPKEkEu40Lr1vSKtiArHl323JqeAAPNH1eUjMgZtCGHquYDzRRH6hDZVZDxQhp
hy5Qzas5W2yX3YNwVRe4J61wiI2w6FT7+ayRfutGm1hE0bAaEjVnZ9XbAGiQ56eC
iRGJTR0aoh1uhEJHOsLXHRC076Hw+fmEzqy3U8TpXn7LtHztYtW3UGvSzQXmPwgf
f7bkaUHOcUV03YDPoPh8osreCKYjGJ1GNdX8+MAU0tAqOjCT9JiRXIZhpxZ+R2j6
DxL/n3etpzm+uryfaYUWyFhB17FuB0VrGBiIFkLhiz/pMOvqP9mMOAyVB7FnnmxP
hPYeS8x9t5JgEff7S2YGjnqGpekQ7zC94OLDj4yzaO8zFSXCL43hLSuvihWxVbNI
fJRdKP/r/uACN4AFl4EbJ+zl7rz7XKN74DreklwJcgSKo8hra5rqGkEAPkTdsmeZ
YkBawoVoImutC+oAoibJTFQioYdDESCriFEbe+ZDOZmh4R5ay3vFWkRFYX8yWxEw
f5Pr1ijDFKvMUGK6TowHErVuMHYHxyluyjSw/UZ+wErsSP670Osi0NPtaU6T7fYH
zk7SEtKICiFfKuK2YYWRc1l3NqMGu+kliwfZ3F0d5WCCjx1fwrVUf1I1r41F5P37
eeg2n41VS37QnIUyqQ+rNsLXmby/cGkJqQqvuYkE1lZzi6pTKSuI01DX167/IIPY
z3FR/TsLqhQSHxoGj+aR019Z16oXKPmC9FYOhSosjkAZpsvGMTZYTsUy1RV0nkiN
kMfaMOBqPfr7xWUZJhwo4NLmTYR/wlzWVkHwoxRlSbeZziZ++nMCTIkliHYQIK4A
RR1a+kEkC+c9Ri8b9i/GhhPlIYndj/DAYzzQiDz/jhrRpDaZAyOv/Sfo/KQgVv0q
a7PseVgWv8Vrm0ULuS26R4iJSwaDnUeIPf8Y0omo2tslEkhx7vEUIYHvy7ICxTpx
uf7xwsynQnLXJdG+cMr9WU2yJTqwkuSa6+MlYGMayuB4qNHCsJpj9jIFzV5tNiqo
NqZiw6htzD6Md7UabuvcNaphdxz+CwXT9ejgJiGP09STbYRhnYETTNWu+oxFvQWT
Yl8INtbLmuqhVmhjpVD8m5+rp3fqayVUS0gyJCIJgBB9jSqjIhmfrCB7EEVhCncq
PVA8MmxMSKMrPMBE+dHkgPCBMvfik9JPY8gwXjUhrCanaTITszkIGlFzxYx10LeK
lKFgoPx4rQtD4xz5LriHSUliTCCHXwOczaUcv+d6KzdgAWpxWzAahu3E4r4W1Zks
xG2Cs73G4CXZkh/IaSCkM31WJWEVf8J70Yv0xIF+oCC/zqXcRjGujkITuMBKrCFB
/ctZRD6j6eqYwVfV3GNUJrpaxhYIJxLi7ctcOzAra0o=
`protect END_PROTECTED
