`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVs3cetQUCzne42dLravieUsReQvDrerA25ZNYRnwJSAdhcf3AqhE4f/0+mEH46O
r3/aLIQgCiF/HBdQ4c8+W3G6yOx09HUwh+/gFB+eAV6aEvwZQwMGIh3zwhDK+3SG
HpBFwDn22EDoy+RBYpvC+SmJjcqlZ/BHihdpYEuWSJLzmHK0EG3BhKecC+VF9s1e
GeNOT0mgpMDERG0sUk8IEaht1t/eDoQwYbUdpjjZDtxYdvxExCsTlToG07XJWuwz
/LHc/CV8y1yFN1pIQ52km9gNjRr8+7AmnFpbkO6A1hY8+AH7ifbr4BL6MtOD+xgO
Q7e3DgOddAWUBBUUzy4UkvhiUtmOo/1A+vlBnK6XPszu7KuJiIv8CRtoUhBHESBG
4tfNGzPczpADXE53HJeiZDgT8dfhdoX0vb2Dzq4LgvXLyjC4bpVc7LMob/BCY5bT
Pt7V53GFHLvpIfDqgiQmnNX+W6FfFciP1IiqspIMQQt9foIhnNsYDaMsfWjpfZaK
twfcggZkKI/WWrD2QAqZPPcRJ7trScvvTUnVDVBoFm4e8CXfDm+inYBCR/WrjJfj
r24PEReJWcqNrDAyiuTrc0aptI7AwXAxu6yWs5+n8SBbp5x7AL9Cx+JwdwdaMyFQ
Aj/WpVt76SG1LbNln9lhO/HTaogxK/C7k2CfEp9vwQ/1vnMcRa3aMsVWAsc27O4P
ewTtOJOiIsY/GDhdRa0wypP3dLW4WZtFEXqHLdIECofoWevStBEfvwyIIzH5abpi
Dkk4e6qg3lFQYhOeZiXbUPal4Be1QLf/dwB1tov79iR9KJXe+cSQ3dJ95vNC/Ud0
B9dJeiMdO0PT7Gx4M/kI0oXGJrc5vYCPEhzUNIJ0ZgamIGaXbBxPo5gKxKG6+n7C
g+fl0Sz7zISGOoN1n/TrFZp1UsYSZmB4fmEo/rnnShJAY3AF9TgF5vYHIKoyGHdP
kK6odntfteZkrEwTHL/QfZFkuCUkNOQv4MkUDAavvhqHXrAWHceO5bQ2Na66AtKQ
ngm/VYJrUTo9Gols2OVOTQAA+glr66tuA6/RNjoan+nojC39F5wqShsMD4lT2L3Q
ISv1/C3DGPMYW2ps0rFE9tdsAcgXo6ANcBcjD7XRart2h3PLcp30eo951bTq6G8r
`protect END_PROTECTED
