`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocYlqTflHMieIQ9lDy+4LsWqaZ6UY6jjxRudGXvjz/+XpzdDB49yuIGsiOKLsu94
si+MKTk7TSzS0quJVnrSqM2pD1il3/R3tAtrHSG65fxDj/SA/stbVWYsEfyH7jeT
L9JrEayNpnd8SM1jLojD1I4D6uM42Vk3+s2zErF12QdoNyVGYEiZAj/tNKmC9Z6Z
TSpzqGhZFgWq9kYleeODmm24dtNy1OAWFD3VvepYOcFIILNW0QEsszfA7x4+i+QU
x9vYxCGQSiESmu+E8gdfOyNFovBnGYVMQKVrOuZfKbnr2AhBAzbzvp/pipJCOl6E
BTl+SqQK6KkRXUnmH0H8Rib8G0SCnlIXpfL2lOY8Kt8=
`protect END_PROTECTED
