`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDB6Vd7optUCojy70jPT4qc4XK2tqgbpL4G+95/MgQl+EeNlYezCjxqcdtZ9uFc7
xrOUyJPWp39mnU+16SlL1ajvK9HIK6FRkzPSUoArPBbJQYQGLLH9vMLmzbPWgVH7
GoIjBSQBZMDV419+kjKPzqsgorcOeSLBs1eUMhZDpQPT0B1XZ0tiv7ROR7UXnVPM
PqqioUlp62p2ORgmWfdDN6h+q40bR+walWTll0A0oeNViyS79lkXLPccU4ghhZCl
ekpJIjkX+VTzq7Xs3J8vUSgL76Sy9YalGaVzoOhjLhl876UVIngjHWUzxr8Uo3Kr
EFrKC3pIqQ0YzLbN/STE6f0YoLSXVkVFAxJqANLGKkGbNyLWE7OCvUJazPOv1ieH
`protect END_PROTECTED
