`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXkGR5ht5ZfVTq8mtoXUrUkKHdKU2/cOOa+7KlN/OqTjGzfyM0xSL1P9gzOF6/Fk
5wEOoERXMXqj6EIxeS0UBk2bpRt350/9584BtEszwJ1N5ID+AnRhkTctm9RYevL3
xTvvMNydj8v793/NSknMfoHG/K2FqTgaxT3gH/q9sFV7pD8TBJ/q4LnzK0IWTfhe
+VPPcy/z4WQP9LgWCt6fe+2ZmYXiSLbkuxSUCQGxJ0CMgcwIkmSzamWFfJqad53V
inco9oYKkol0+ED97OjAsaYIR2usV7BTyfDN8J4AyxpGZXbEKxRxeq2cn+0z4Mmi
ecjoXnUvitheRs2Y9R7KDKP7OysNstmRg7Qar0v0TlZsCDOEKvQPF/ho3WKB8Qb9
RC747MXaMQvLQcvCUcmuXhGW+ohuXSmh27MMCUKHBgfa2nZV8UFmyLBMFQlw9tD4
OcQU4nmVTK14tiq18aR8hw==
`protect END_PROTECTED
