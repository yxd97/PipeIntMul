`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLtF1Cy7YGlq8KDrBZ+7ky9aRUAYaeIUPyEDUe2qgim4Qdf0eW3FwIW0YyD6LT8L
FRCo/Wc6yC5u6FoA03wTyJO6r8TxlXFFwWMJH3M+olc8nit8/3vTBrQgMIidkXEZ
kpdQho7Jh9vcUPEh6I0YgSNUvmyO9Em9t0LUVupqpjcO4zDrUqETx87EN7ITyfyE
MnHz97C7Qrk1gIUW3PoGpWLCzYKn0poRzTXkYEyMEizofvNlMWH1MldkNrgNVFA6
DLGZ/Lw6lDYUFry+gY1o20iknRWCwXmMKiG5XkmmFT6rbivV7u7vbWPK8U8CDb/M
aUIgnmrJYScbWo8pCKS8oInwwVKlZr3DSxtVIS6hxjme8G2rU60sDRCUpZVAbWJy
8agd+H9iXyC+ChFfUJv9t/KK/xZ5geVV8VxPSTVC5mXxpPkdeQiYotcH+ajlDVt5
wnwr13P0F38Wx9wuwSEaewScUqM1CXrO1AGaBz02NNC4jINzNyGOkGk0efyBUlWR
5dgkWR49ZK1VbDgwLKzjaQiAdrNaF7/vRdZ4+VeR36OxtRcR2HjzIaJBpaN5h5Wr
93wNrUMeOYSjSOcVZagob5gsS7qAvFjN+x5S+VlU3BpUbQIpdaKV5nxfLt1lkG70
ngsDE1PORWq9dbqpKMpVcdgkLZcYgA9xufrCK3cmUM/+Fazs5+LRpj/v0zZylV3b
NPb38roD4od6Dpg6ncFLAorQpCROYziwIVfEU36DdXYWhshYf+1JOzYxRZHmw4+l
TAn0ngwsCsGZZHd39sb0q6rtI40IVlejyw2Oi/+PdUFbpPdpSQHzeN9qjABGY3BI
JhyhURCHFbffH/ftg2XC7sEk4Cbg1qqgLD+E3EriMGrzCDVjXY/7Z3t9KE0MgB+x
W600S/iosLPQOwOtztPwCg==
`protect END_PROTECTED
