`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P04S3n7x3Rq9j90pXZGffPAGK3mYCtbp9R/JAh9r7VhyjdA4zCWeaSHQga9GljLt
ypBCgnGi2fHqbl3QglGOd68JcDj11kogwmVf6K8+ofG7kTZFTyAnTsNdFOvK4I1L
8Xe/a68aMxsDlO8zbZH8L6NzqRkGhT5WQuH9PNPd6xu+ytrRxBoJLItOcWjp2N9T
pcLXol9VMFQEXx1Fy9+uc/XqR0tgUyNKHrX0BtMwdsaVydahso87JgBiJlXhvtgt
TlBnwQy9PiPiv7C34WJlX5gF4HsfBVlXweGYFO9xnI9ffIoe9sXDt7gOkAQ6oN5E
93enok4nGOmAtYVjNXmtqpTmNL623qf4mXf2h9usn4H4X//Uh7hqhxiCXY4HCWwL
nqLboKIWG0BS/1M1EzI9xcc3SOBIVzojH54JKcMyqJlXd6VTDRCh7CuRsjQdhbCC
pcBtFytrtFA5UhfoaQF7wY/2d9G7RflAfUckaMf3W2xUa3WH2NKoNy0HBouA78tK
89koD3vSc2AybKT6mqvAYAiwi1DCxScWluH/rm35+p8TqrJ6GA+HRxEdcHYFxMDm
5t9307YbnqOBMv+E6+GU7AuGUgbk4xxu9mUGm8pB/4Mq/wQ9lpp/AT9q0CKvUUyj
WtqmG2uXcHD4QLhVpKHrwMJnMajNoskz03s73nLIedyjybV9mxOq29LcYGkSLbGC
IYK1viwmX0/2b9vH6ravROnFt8JSlj1pS7VwdDrWLAQ0jqFxuggzVguiaFqZnyFE
Nh77rFSnpdo/PxLW1YEJcjR7tUqc6ZSOZYDJBhV6UyXcX5m9PM+isD2X8/jrj20i
/EYTbRXsJOOjjWFlQsqZs+PmcBQ4vhDjQZw8dFose+4c1B3wm/eESexD6DQ0tmLN
EufVxlfBF4td9pKpiaJdr1Ef4cPVK6qNI75EeXqE+JsNYslRo6pbSxXxkQVCJeYf
`protect END_PROTECTED
