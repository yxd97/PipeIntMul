`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2WpxV5q5iPtaVN8EK7qYV++tfjmpIeBqY1iYIn963Me3F2y/5MVH6BZY8RF59A+1
Jd9hoquLN66OWMDImSp1oN3LmIt7EueAESZVoX+0Ys2LQdgPaXxkyndjMagI4n1H
V/zNQOA32YUxPc6unbujiQdT+0gF14RrjEYP7PRa8qejeqi92XUUGsfHjA+YNpat
9IxKOt0cNM495x95Fe+NAS36MUMGQIFfFOQ5vnYuuCUNdrHubiTDA8SqrwEvAUoy
nB2QlsIciElTJolxzhj3rtlaZqNfMnrE5shNHjGuvwa/Y15T8cefc8HUbd7+wEHD
O0T6oKKsH0FQoSq2tAwBIg7QRdE/OTowlIwk9axTYB5a1tc4Y4yi1Xkf8ENCM4I/
kQTo42YuBhuhDCFuaT/qoZ4ZdQEqJOFAa+IPMVn4eq/Yl2QUeMJP9WgFtEvq4wfs
fyD1Rfpk3GL4GXtK89OZJsH3LvaNVxlwQ+8cneuOVGbEY4upSJwtu4C5kQHwE2jS
lmikpQLZLEAaQBvB1FHRMCkU5OEv0bHTLIv12QDrVb6fTXlIiQDtB1YhyLKOS0Mj
2Bm60+w1j8UMoWRtrSHOE/uYeBHZfBAXjB4117i50Nq/41YIvtcIvNgGxn+W0vJG
e5fDS2I6ztZr6yODDDKa2wFrgEsNXOO3cworiSWNzlI38vOKxRLpYNYcHl3znjik
7Hc797cEm2bcT9OHcPGOWH6GiarSJ5dMQHZ5rYY5ubH7CUBs7UZDuPH+W9AgJi1w
Q0K2O7ZwgZGQQlvV9fUUibn+kT9JPMHg31XDHJLF2632TjbUY3VM+yBFa8mDDpPj
cpUcwRBU2Z22d1YP/SwVEMz10neIUuViYpPpIIsUbAI6yZfkJ37pt8WMeEObMZym
Ueb/6HBO1LNRSGUD+w6fQT0COvza40kDRl003QeTb2VD/gzDPTs59yaeu5dntNGq
YStY3xZVOabDs3gI/T1zsafKhza6EL8zGY31rscJOXl5VVwSdfuj1Pk4cHL3KlN4
NAJITD+EVl4lopPe29OdF6Lmt5NftseOB98YrTrUNvHXrHdGDmhUI08F4pXEM8+b
+K0FJEIbfSfDjttHDHCHfPbK65IIkSub8N9FXf2aEUZw5G5mB9wCuPClzLozh/vU
8qAoSEcYC1QTPd0OpgggzybpsU9/NnI5a6NqMQRHzWExuiRsfcuwsYrQ2GUXaPS7
1r2Om6s/eu2YCD4NT0wtGtaqaIgSlv8Qt0LheHSVtANExjA61qiu4qn+s1UKtBfK
BjcUfa8NIBSJzw3xiQVWVX+wGb69aU7XCn+hDGNAjImVrVsYjl1vm7lmkNtb5rVM
efFU8FyxE3TVQqIU/TGeWB9JlWqxn2E/6dp4qk2n2eDpGgKuBMQl9FpSHOaWCxby
Mjelde9YbIgL0kSvZo+jhUsVhfTWkeBQk6mhs3o49/6PgmhL6k42s9WWKN3JNeu7
CyuiEN8J5IFO+G1XNNgOGOk3mRtHEMCahLSiuB/TATajOq3v0zrH6Crk4Fa1wp5+
IIKFl7+3KtQW5JfQtxW6stuTZWlAeJrsMr3GNuW80on86uluU38pHEEBPiNiZBuT
V1MJQfQjR1nlobAlz3Nz6fRpluGqC3ntqK/nAvkiCZtrNn86ObAMgkrIHNiD4H42
pkQQYK3IQIUXF+DM0uuFx1NlYBwZJZ9dIQ+5v2YM+6mGUGPZQLqGEdVeTZj+aev0
JZIAY36/cSucNrYkDdLXx12C5YEogMbe3YPShVK8BJBcP8xWhChj7gZPx4GROEK4
mQyaKnD0zDJ6v/QTKLIOnTSLkwI3A0TuZl+HXdvJZe0YADYlvsFbLI1huQpYkdAP
JGOE/Rr32l9A1AoBs9MSVteELvNKg9hThD9J8yNW805Cl0OQUv8SJ6zRVPV2ysZe
sZ0k8tEDUxokYDReEGbQoCyiOLeOOdP1rqzvgG2FmtfpxTozLTxwhQIjWKvEYRU6
GfQwMO7MWWFtpTLhuP0O6Cdnx/YT8I4rSuqXIiUtaxNOGULNMjvWra9oUOj51p6y
Zy0WxV6Yxs38IvUUY8DcS8UfFgvBLY4b1Xtypobj1xrOQ/6lI3FZBVqdJ8Xi9Zkv
EKlevcvQQxaqmDSEXXPsrLh5K/YdZ1MIHjVfkLiUqfyNJzBsUgwaadrB0IdT/XfR
jfv861/d6GdWt7VJ0MI6OjUsEYC8K4t3bR4xB3X+j29E3QK4tHlGVF0qzoU1EBZ9
8Yan+cFzGzATP1c+CaA7LMcjQux5KrXLsAsLwBj3qeC0dUBvL9wy0ZpFv3NsS8mH
SUS+/0wGxgntvYA9vEmKujdv2/p5c/JCoeNpaRFICpquxZBAsNrLWC8yKH5eeLbn
eGz+jUm2082H+LYE1TVbbq1jzAbNPCVs4CUvW1PgmL+dFsbYQ469kc8ZknhLHDG3
QTVI5gX+AuOpmtqLFv6MWip2JNcPgzpBYCC57qECIoidsAdVsQHyEXt7KvIKNRnv
fAH24iaqOMDhWRwmlYgJNpI0GcPFsU7yHuYXnwm7+mUCw4TtGVO25VW6SeDpG8VA
O+wMjEniqcUvAEkhktOp/dGJFy9l0IMJLGLT8o5FMufMEwaP4HoBvEfmX+pV6ALh
AZzNNorFeJVMBt9X2mI9IZA8ggc0AVRpznrBKktLDcuLsYOXwJdmfTHUmxJDVP1E
sCCzYoS5KgCN+8Xe7GWjBzSB+XbcRhWgnZdnFmgR4G6WHKtMI8VoxODdK//45Buf
dWb6UGPbxQWKKwFlSH5qlN2/aL3jKaBc/3utGLmcdCKqUPgE4TPhdycg8z9AMIAC
lankWjKXR3d5kp2rlbUKJFdEvpdRb3zeHqv3J4G0/1CJZXuG+5g9dWpfzMquB/nG
bzesVLZxEEzQd2Q9sqpfTLB4qGizT8QGURLYFYv9S6pb2gwdhHxTRSgfLTMoUJ0h
trp7IHOoWVYirCCysBayeCIE6v5xZN148OP80oQw5Gnmal+b0DTMeKmYeAolK/ZR
NUvZDHpbvM75rmgnKyIPBv8+96ELCXFWItDs/gEl+Si1hPhR7TKBFl0j8vB0qXUF
1Rd67lEkZmzFIJayC7SM08epBEAy4rF+NAK490KJlAlyO9RSVqo54TeLSf63VRBU
2KsHKj4qdZLk0RSwV0fiQ8qCHSetVuSlrN48EWBLZ/HTmOqpy+kM7t8OtasS12QC
4dv+2d5woKP/29XaLQyPKrUMU/oz32Js8X/I6lg3HYW6GQ9G4PFEErDXVaz9OzOH
SPkNQEs5Cw2voQh0xperPc9pK5jxoWckfdBhrFScoglHFnR5iJSiPzqnWk4c4I71
jG3Gy1691U7QiHNITs9atlC/HnFEUmKqgr8g+YFJ05Gf1LV/2MCNIDSP+KyIqSAs
lSiDUf4K29eeV+/wTyCnmPn8+uY/W0hn/jII1DG221mL+0ZlmPE4Z5NaoO2J7e9x
7IOrcsvrweuKqEZjrbozyn7WoaBBAkTpJJ5OkwDn80Em1wGznXeWR6FaFXyT70x+
pbS05jTrT+DZsYyzjhTzjIJGm9gUv7bOoH7pPKPWp//fq/8jo6Pufg3fxrNHkpT+
h/O98P3rXK3Mh3FrRT966MraK9r9G5fZZHeAYrFNEV3o3gJ1Xp6JWrApNn9VSmaw
H5nySvP+mxfv4/YsnOR0cCpF9rF1Rv48n930n/YFquzcmpu0VhcMYnb6nFJJGHJg
3ZAhW1dMoADNK29ThHsoE5QSJhrMR3ujhB5ZM72SDN1CSBSdf5LaW1E8ORCHYFgo
Cm36udJopWjkq4CfBHfCjaF46iM6gQNE+PN/TeI/36G/jkQKDxnjyYCfkIOKbETb
OER3++7w8axt6HHL8S/aX4EVQ5GP4cSBp3UxxFfxVW2LTJ7Im1CsP9S/vOtIy2Pj
VVw2hexvxn1hL8/dzCepHSIBPGNn3qWjONDG09Oo5Kznkzjn/dDj25ostwER9x6G
uwjvBjksG+EJ0Xl+S376eNR7udDb+bt+iu8Ghj02do2LnajWSdTH6xgIE0b8PtqL
4yd8o4tP/mFs5ymX4LLAsG4mtEJ+m3aAf5O26DetI7onzCPsmYSVgsIQM8SiswyQ
8uxlgyoS3spiWpifwmst9G+qJS9eZknmSx7zRyftQcXkFJ++M1qQJPfJ3uh9IIRF
vWeCEbtfEoOW+1ptL3P4vXcAuPyJ5hKTRSzQkJW1LdNFrg5FoB+4BNKLbb+zZHcq
lOLNE2nh7VsWucIgMx/CWQnExAw7EeO+jM4m+OQROKn/0OK7tQJsbEPPoWxm44sy
n0pZKzjpfvbq0Tp0jQoYL+wJZ29k0FWDrfFBXs8N2NfU6vhdhkvoqZP1byUfurzU
9V1RSZwkR8zpGMuP+GnyDGf6210k881Tn4Wx0nVN0bzK4kF6ZxgTFHaKg2krOWgg
8occVHjCPqhMUbzt0WI4BtWE1luOZ5bvYD21iYEN/t1T1clx5fPKbJ0zcFnOJgPb
fNYWcJp/gczOkToStOvHt8eJjrIElai6aSEEaJ8H8JWSUF/P92h+m4cuJ3MT/wNl
YQneAsamLVfdqxCxupcN09Tv/18I6vt5OFwFaNdQOmrF2Oi4ghHbmcq+VQZu9dXq
jpE0nWT0x1ay07MbLB9s+tTIi2iplj6wBCG0IGUFm3EBAArGWhdMX4CsvfpARgs3
GLCjzaMwBnJbbzKpVydkawDU+4j/sQ2h79mcMLqRkkvfkzMFFzjag1ZoCxBpGelJ
qYaL44BAvQZXykE0rAHQ49LrP9nI6GsyMX/1+VmISFSVgnDzSOFD2jjdjOzxlP4P
bgg4oh0gCELACjIoOflB8HkP7HRBLyC3k2if7/VNNQdJUFFiXRnrjgC4fZXEQQPh
COZkoKXsc5fZJcap3mX+33O3BSjmvhbllQSxpYqWTSGgYHe0n+odYKLTWI4pR+FJ
zt/BUZ43nxrZZsik339glHb9dpMhfVsYqcJTLPoF/BHnpMGNUcS0YB+IlxLzZmiK
lxR0TZqNMBaJJPKAhsV0BPA1ifE3VYZJCc52+F4wJOs+pcNra0uqyE7pGpTJ+C4T
Baih5JXwwaMc+GbnnGZAohN+Lk7VtDWx0ZshdJFCJY/KEYHpEe+ayqQCC4/cenxi
cKltg3dUc0vLntRWy+U1RyhIFHp4n8UqWvk1BCzdezqvMeeeWl4SQKi+aQLKhs1i
cdLySUlIG9c5QM87+oCQTEzBZnqzUdgjKtvcwPnKN4nK2Ck1KQFnS0LNujU9V4eK
4eDkLA3mqrJ2OQF6akkb0bOpelrV/fRXlTk7kRkBJ15PyTU12x4rr7zEEFDc9FIu
C0B/Vb5wIFZZVbPaiD7eoHq1YHmiT1G2sNBANpE1+YtamuquWBZqL5y47ctvMupp
v7kTK07wTEAWiKFBsRhuElRG42tTq2fEfITcRcmLpvXLW/PqjLBwBC2sjJTutyPi
mTxqYkb9fk+Ba18MiiCYc8amEGjpn0ZmzOY//Buc8MROm7QBrNHLRq62xhPuz+/E
Jy6Gb/DhoquHROcvIs4p+RGrjPdAltV6jfGfWJvIKDs7OfgrJwtrX1yAmSag7x2w
UeOeLCJjfUYNmsRD47QucCakBAevCeHZvMf97f4kn3yHnNGIR8+qIwmtgCFoBfrR
jOvLZKIkbURc4FHycri5MDni5Pb60TWAMRTli2SkvSrC235+XJzgtRNLA3jrMudo
bOV7vSb6ZhbTpDj+/6ldLoheH6jA2updcTLwhQ2hKUNmmMnK81SlPCFcNbHwjRbK
cGmcjXnlMDRqqT30zdR0ebclCqbiOisV+wkUP8WbN5u8CCd/luH+yB2kqPd9S68/
nwe+DOfh5OrDZK3rrXZL2hSzZ2OxLtzm9E405eMnbMd4z/NkC31g4xRlxBmYXvVZ
Xz+xxZEVoyRQQiahMFHWjh/9zAkO7L/ifYybX5g9nexKSB/fMkmIJl1T8yLUEJJk
6myvu1MTUW0EiyPl71hN0C9bNhmsNTtXp5hnGAUich5TtR6SoO2yPAK6il92xoFf
ZjuBXd/PGulQoCvPvi0Sax/MK4/cxQ+0sdwk1ShWZUjPb3yd13yg3C+x0Xldx8pv
wi3x0pL6mY2CMYKg1rtmyMNCKArbXebdE3h7WASYPeZrBhELhdJ2gJUDFeXLVfTr
M+lYzfa32fQUO1qJ9NzrviJaKYHR/yeQq3HRWdwXcZygFA7lGi1Td/ZtRIEDVsu2
po3C6AUxdzFLgVYMuoNzE2UoVIaS1d+mga5ZzH0RRIjETlMTEq7sTnIShTRSjxT9
ucz5RUyvcS8/UsLuZQ5OBS22JZNCHK8UxhCnWuRz/D6akDHIkweh9Jg8xTDgrucg
RE8ee2liLwjtyhKk0ijUckLMopFTgr4fHyICLidE164xbcGZr85QD7QOtl6mfxSf
nRgiQtwuuXw/gLJckuEhldzVNs0EsRLWqnpDsngG1gj5+KHMrB62NdNxc9FYm+Cp
gyPyqRq9TY2lVTzUXZ/OM9cIsxzBU/UuLJfHWPQmMDzzUpe39VA3pC4/NfoMcaJc
Iw7JXEtx9FMH5M6IYOnj9lwV7yOTuIS/dCCsoi9csOyeEVGxyGo/KyujtgPhH3Z8
aVzIaqomD1/eZRKDKU3/32n8BColElKzft8lDy2YoAxY/BS13wzit25S7MdSB4Jh
91gRgZ1pTlG1T0jsmqRrvgp6HdE/L0b/mckSjSE8GoXjr5rnr4/CgCwHavOq28oa
cuyV3EoUcVsI/AtYUfAgQIITvAkho0HGx+/bNsDwjvWavmhoL45SRMwgTuYSkalw
xDb+C4W8v0fcDY2m/41chAle851mVHTErokdD2zmFwAyH+jf1qcM2Ywp6ctju9gp
Ug4RxVFM8X3uSaO7NQu7ePA67uBo5EgTZSdsAqKNg6Lug9yFmwV/XczT0xG+Baah
ESUhxpMWd3JKKNQkV2pTeYccwKPEAHmAd+YI3bmaZj2SFMvYBOxXJIQSO0xtHnHw
NEaRoW/A+qOswqjhnzVTeoRQcRDIjzcDnFShN2QH/TTSP8+sq+stk5x3Nw9NC68s
JhwHL6T5tXd9PY2u3NPU2QtacfSZsYrPUIjN8EsNEZ7jWRdhVhpInAQEZSJTw95a
4vOgvsZn/0weZcrkW0CODe0HS62yVAXJrkZ+JVldYEumvrBRGv20u5+R8CM2MPef
1dsyU5OODTuMH8TY0efOg/4PQFOFNNYtQL/lVJCc0/SFjOIR4sz69uxM4KZE3KJg
eASO5eAZPrq0qBSNlMBIfl9Zvo2ODdHS73eoAeFHhP5BqntXysYDFa742i6yJ5wL
cRkBRenzMHWREGeMbJOD0pfd/KFoz+OVh8TLYR8Nn7rDki33e2VFqiQ4GCLQnsQR
kuCMG5VDzcPr2xgeioUZFZWcopHNC1xENhetHCfVREix1+8g9I8553EOlyL+Urai
DhlawB61QZjSKjQPuOkOavhMadlDGGuMlDrRO5E23FLOLn/Fik1Q6lKw6ZvxOm74
6m/pmcB+72GqBMQHV8E5XPSahLo/petloqbYGNjZRVAgNtZwiXtsN7dS4aDJXbsx
yEOkdM1brk7DBTfmaqqmi8s90ydOlQxQUMKoqvqSztgFl2C2xr+jCHq6XD1oQGO0
0LicKRfamL/8XFABlSyq/WX5wtlBusbswX9BpNh/iLq9XHLKW7nJ8myEDxTTs39c
yNOHa4RSrvimibvrWdV6JBRjzTs4mOUV/yAPjShRPOjV0deL5YdD1UionwmIqtOl
M5gMfP9GacsLFRNCIfA5DHDXOM7ybz3c1yAkUzmY0KfwL9YHxSN3V/RLR0Y83IPe
3Q+CHlDApxdqurAFa6mXbOiqYyiXgUsF2qvroxoYDnFSm3qyp1Qj/wbo6T1WF1Il
cJdbKmXoUtNBq5Qn+AoJiMvW5KpqpKwmmwyLm6K24gbbcFnGlnopRy9Y+EVPeZNW
7Ef4FVJe+KXDkDUb7rtOXuC8Bu7bCwsuq34gix2B23FJdBqSIfzRxiR8xm//XseI
YjnWiZQthhhVdjqwmgKTAFVh2pfLzzyQhEWSFdFgBSdxkwMUmG48n8Og0oJ/NEi/
p/bLS/i7X7KRQOfhTe630fgHe90m2GIqZbAVAnBw7VQJf1RpOYAELvXaLYznFc74
/g25XEH3BtUFGSJ0UQF+n3ti6CbfHVxzHA7YU5uB/5kjc86LvBwhJu3mAR2DiX6A
uohPJMHIO/xsiLD3e4fYOOhLK8J5CLMOlQSc4U1G5woHn8KingROlRDsmbFuBTCQ
Vck4KSRjdiv1xnMXu+MoT8avK5Vdh3PhPSSayy2seWVd6vC32RTVXOe0toq2R7Q2
PhnMjmqjc750c+9IT1sDe/3PNP457eg41NZEM25RHKJ/fmsimP9YZcG0k+aetmKe
+ghqcZn+hyJ8thrdaSxwaJsL2TgeVQWEwGiKGdYPu6C2AWPI5IhcE72VBkWQwq28
5Ql52ux6XngWUE+ZBAmKBWSx7n83/S1R915Mics2ZG7V5OCr7LCr0AdwKaHq+qfq
4TAsP7dLH9rJhuPEmCZ5N4P03T8u2xAGwrdEDun85+HHXSdPQiv1GrFuf4mhL3Oa
7hEOO8QQ9GXyklWqyQ/SqYTkuYBLnHVarVDKo+xNfGVcIcpvU4y1qZBnE9y1Auyo
QBfXp4uYJnEHESn2Jo93HtTIiIrGVXYwtfGlyOmUq2tCeHFusaG44T48m25AIhfL
a+yTLTzv2Ly0Nf+g+xEy9QEwkNS4ZbTfRrcBGgmvwa2ztXDoMlZ7Ibb2I3LL1D6F
SxSSmkxlzb0dl6pPN3I2xCoSPaE5yBlHmO/EHFg8ibnTQ/PUSrRB76r6xz3S21FP
ly9yLH5P5dRqcKutG+Pt9D95k3u0NvNmnCkEHDadQXYF2vw/bbZaJG0BwzK/ScWy
IWoKmpjDAcvCGwPUO1rQTnsj4KQ8ax10yxTuAHYk2Usfi4NWupBy/wOIaRC2imMk
CwTSeLtuwD0+TPtNZDOGA9RyfntKqJijScMu2DORgHrcerrJCvDvYbpkN75U6rlM
Xpr40asn1n2yO6/OKVfYTxcXFzAEGBrAywRg8gpmCct57jbMMAUkcQOl353hkU5w
6Z41IrZKK0PETP2b0mFsPoR3xvrcenCMYMN6auB8SSUPIkNdqxXLc2KI90VLMTRu
SA2pvsRFpR5WVFcRNPvKnLP/sMXiibZ16hFi3SwCYEgHdJ/IROL6Z/I1hUooyUDR
CFUfO+cTn7iRgtUkl9YOv5jfAjx8t8sALtgIA6CkZka8ADTmjeppcSC+wwBYutDN
Xc4YVPa7fJVCtWaQ9sD6Zv6lfxDPcUeHOc3ZcLYprCdjjto0X2BURtPmhO/mENtq
/grrRffMims7MqSxTi0WPdM9oEUpHNTPGWdEQz3WH1pyfOZ/N4LyS8puvPWnmNgw
aK7g02Jeezm4Jeyvlf27rp9q57yy5Gz02WwwQnaFG7usXnM414JN+CNtIDsY8fvL
LAcuyRiR/fccMyCcQt+tXXpOdHCfyAI/fSen3di1qiF/g8DfmaS8IOZMJ/hUsdkB
nca66S3EO9gopB3UFOo4T/Q/lms948oH2wmQNRJL0cNKaXONqXTiEQAxG6Ae9PhY
kcxmyasHhRYjNHUaMq4MaasJEa1okB1aDxXjnXWrlhxFPIHKTXufxpLrbIYlJVB7
OLP55wTInfi9GI+OyJHpKPhZbcqfBwtuZwE+UnZxFDLEktpw7MmNw1R4b0XEcdU3
929MHKPEABGLF1RSirzOJxcnBE3c3MY8ppexFqu2EyJhF4e43TVQltsyZF6QGKof
zL+JbTA9qaVM9tGQ5wh7L+d29UmsXNP30O9/11w/l7OpbT3qh1jqGiVSf0WWtpzm
nLTI7bse7EJOkWwOujL+dobO7nFMo50HO/bBqo+M22CNNVbMuvrTAmWFAjfJ+74/
IAnO+f26EqFjpfOGd638+iQlB3YelfUSHeWLpkwdViFdi9eXCiyJvmDHWmnAmcmW
7T43engRN111JICHLWvM2nJFE7HqX5yF0anV8ybZDpB4To1S56QrjJqCDkSm8cx5
vgaC28pTE+Had3bjmdWT870DPTk5nQTNGMfZ3fVHJHAQTMQ2XQf2CG2ybh+YOXAe
5lq7xW44NZaenD2PPE39EGbSpSDoZ1gmT4Xj/fba/pvDO7QVfXXZXzRXa4vE8iYR
+/STIj8sWxtNWLfWrbmY7khs4tGFu0kXhBCbZ37BvIGKydHUHywUytSBfs+6aM0/
OuoMnmP74LfMivEg1SOhE9s8XwoBwiPQsAOEMMXWQF5bgxVSqymdwvt7SM7Wpg9Z
l3W9x+/GZWN+GpSWIRH46IUe502QXbCkJX5DgDidvpGUxbCiTtSe7EUp6++Q42zl
A8Jmj2MEpMd0LU8G+Ul7Hq/vHmj8UPvIvlMuwY4CrrZ/Zeof8+ouRnsifAHHkYli
FmaKBljkuyqNZBmSW41HEmUAaUWk8pFzIAZZg60X+P5oGH3SHsPFIRrm6F8vhmiY
L2EDxlle8szPniCUFdgkEByVeSUQHKfOiOjezYNWDWdjZwdjzkm12s1W61u3TUuh
LSGjggUTyLFOqDaUzXrB1v893uU56YKcv8483tIeG4vEgyXf9DLa8sVa/DH7awxV
zXXNnaMXYHl/abqUYuAEjhXeB20QqM9oWZoCN4bfVpmaJFN0j3Mrd+t5jILwMbir
GuN0tIxb9WwkqN9mjZAZzbDLNSHP6qcRDGUktrfFa+0X9dCF6Tu1AgR2hmzM4WEo
zYPcDEv12mDNexOypZIp/VbTanU3Gi03q8P+Ef+eBqtsmHjsujSoExer9lD6JEHt
YPVY6bLT+FFq5zrvRKrhh2xcgRRqNWFmo2ezG4lt9SD6n4Y4N6VZcxRR2LWfSCwB
tFqeVA4Gve+p+C6X0/3eTFEkYhjE/k51eNcpC1BfYv62o+0W6OGiFbYfxeSndKve
3IO8Lw1IQ5PHrIX6gC9g3biH8w1TSSoLlmHnRpCSOO47OrMvxP+6KI/kMbB3s1yJ
EHafBFAIOdEg+LWL7Uddf02oHzOPzr1EobM0xj4owM0l6ReFv7ps/3yKV4zLJqeD
q4z/b39gE6teGuwWww50V4Ga+LskKCvS7TQ8L5Ob/EzTQif2jzZ/Hpk8NR3osBvV
UxJ+Dvtpa/au7lzOVpaSMsVgbsZaas6U9yX8sRQk65I9ED2cTX3bRJ5k58CtRsd/
2jUBk69bj9WVgpjDdYnBhO3DrTjue6tJbcD8WmEkhBCd/24Cxp+VK2EnizSIMjUY
+B8hAchD7w6KQ+7ZQB1dmrAFmm0Tla+66ogHmTT/vcJ+oL/J5CMO2soXiO6ppgWX
ISMTMHX+VywyB0/b4gc+NEIspfMHkxNCaz0rfP9byNHronb5RJHoiVo/ZdRUbmiI
uS1pZYORE11UjbwWtLpwUVa91pzUzCsYXb1wOqtB10nMcQ9D11beMnL/BDywigwU
FOdk6LfBRLZwXBfTb4aZlu8kTpYid6hinTaa81Prhpwt0kK2WPsWVGu2k9FaL3pD
crKxurkkUa6+Xwf5pA9kpdSRQ8Ss/Ayi8r6S/1c8ArpncVbChYPbntJtmroVgcq4
EUF9fCfqd2yuElsFrJzR5tZzt4OQ2ezyfzJawhEU95UQqQcbrh0P3N4g15KmL5sc
EJa3xwPqtx3Igx/H0orWCmOymSE742TOFLN7EsGk1HeqSC7XGPyJNZoYNAnWh4lJ
Z4weZYDefXMTs12HYPvPRqPoyQOrRGQSnTVV9nya0PUAOJTfESTXvo1Dcrc73hp1
HnPJdlle9sslWRVrhwNbUAQ0m8t8SGt7Gs6gecwauAhO7guPl9U79euyfRev9XK4
YV76QQiSFVB7kDF+p4ZV/Y6Jbev5QZyNe1U/aU8kGgzs6SH1Pjoj1HVNzp0igOSx
bUax3wvY9mhZLlnvpvV3VH6uy1w2qsq86sLnTfoK5JL52cAWBDvjzgijoSTWjqI4
BtNfE4vfcEyiGE06Zfukher2rGu7ay7lg9pe1BU6wXyy7kFoZfg0xmXgjQ+PK0ED
iz7WBLY+xkTc0y/ENZX0dn99sXjboweU9CweORVFmkUjzCt12HpR9aYwbQFXQ90G
SmuMimWfUXcOYCW9qAroJP2sfb3rSWlPGbC4F5bSu7D1pnoRmSe98TfbfWPVbsuS
GPbrsq8J/8pEWqyL4yFlpre5xE0A2nUYEwK5oekppmXabJ8Ny5yFtLPkGEZaDAGH
hXtSrEF9LLadjkLJu7+2dcACQ59NhH3EzpDDx4JnS2LAbhvEHoaickuTpWiQj5WU
TPcnhIk2OnWJfcLTsEFaJYvSF1iQVORXy/zvuIo/Ysf3NMUhirNRBvLgjnkgzICJ
HZqmnsjCzgWAJWnxMQabGSyyMVncRFg9M8nYJ7kcEzd6zU+o4tnY3zrlWznisd2a
dZAWDhQsGESvdsoFp4HLPLX4GL9Ew1iX01iNdTpcqhQgc5tkHre+Y/66+BpYMwLd
2P1QV8U8yR0wrNuDiHgr/4+AfnO7AZbEMyVZq52jpGFazupwnBPAsyIVNPYBSmlg
Qdu4TwW4qEmWlx3eUpQmoXLIURGwijeFYg7a9/ppZbJtD0l94gQxhOhOj24lj/z5
YfHauoTG2xrc/L943G6Djirb1L3zNXIO6udJHBQIJz4=
`protect END_PROTECTED
