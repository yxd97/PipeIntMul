`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scyNlkw2C19lDeKsVvM1Sm0HnT2vi+bkL0r57fDh+giq4/lZ6pc19qZcXjnmNC1a
hIM6qX3OlQFbpYnRyBo58Abb7yM2e5mOQPKV5xeBMDEnjiblAj2jKdrl18raW6V/
OVblN6fp7YuI8G3QQaNX+hktT1Tw9Uncol4NjdvzGZH2rySIIVhB3l95avt2GbVv
1c5t9JVNQyY11kCAP7vuJ6NF/GBMJLQHfGqv1SFG9a3Y5ceDhFSBuxMtNwFg1K5s
nPF6iRqj2xCNMBENCoio6vmjloStUQoNLHa7WJAacjtl83Ft6KWsSKejariZUafE
f6Vivh7invR3DU6YixdRnqQ4zL3eDYGFv1WMa6ukkYtEq3Ct3OH1XmBT5ff6JSVk
VNvVB/Ujz9Q/iUcMTxvgLg==
`protect END_PROTECTED
