`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/S0gjntVrB3TlxLw247ueKJJSyc1IXhPHp0t684XSsGxM2ZXHqRbKX/8/q++N+HI
1wdAG7kH6P1VZA+6MmIe3fw7Kbwq4dctKO1gLAIDQ2qiItCywcX8YPWc/eY3BiHy
25VW0c/ZlZv9i8BVg0DJ1syYeOjWvmMMkcy/4Xz31j6EnqPf9qgAP6pzLHv6XLZd
Y9prz/wOl80NJjEcexSlkSyWiJPhaFnfpofVPagucK+lY2cLg88JSOqEd9TidxqE
V6/B2tIFUZZwVI6TN5uAkF3RN7sW9NV4lu2EeGzqlsJAyeeZlMCKL09kp1sLPIVn
ymmSTDdnVUEpaeA+qKQHt84ijQsD+47w0yaPIN3mc72zfWaEk0UkBCIMvrpVFLm8
/VMLUjmSiwizQFSTOcat7y/+cNPx8D3R6iobYcOee+s=
`protect END_PROTECTED
