`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tab+bL/SQJ66ECs24UcVV6RsQeTikPzJfEz+SMqpicbOWT3CMl8KozP4lAGHhuPB
GGIlOfIB2N7mLHIW2teQLG/eL+09qXGYNmZWFmXO3s7lci2kvZe6GA0xElpooMuN
0VgwPubnHKxh1Nthq7Bg75dD/J5hB6mhX47ZTOTb7uOvhEv91ZBwXy88MKHuB6ae
VjUEh3iVijboONEp5ga/SnOeR3cMYfDAhxokxuSiQJN08rgnIQKOB6B7vL+IJkMs
7B1Um7btn5tLoYH/almaghPBl26ICPFXourPyOA4dUo=
`protect END_PROTECTED
