`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgOVgv4bCjwBi96rqekypMvpFkwO90uzf4iL4KZh5zg00Fsvsva3/Bmt+jH3vofg
kBxEmHl+e8oabC5h7N7E+m59i2fLVr3i8jgckbwGwKpqbUzxKeC/wKMbPg4oKdpo
vWtsn7W9NKiQ6Un48ELvsKHXoZ+q+J2XtU13CZ0y7OOjZl5zZhvD/S5eM6Bq5nu5
FxP27lPiXMfRM5gpzQYYzX3olbaj8Iek549h2gB1wG7e7c7fOxvbhAgtZY0EQeia
8qZXVQy3TfyxbleXDQKCOvtl66Nv1qUMLaqiHHaGpbo8S8RnjZ7rz7ws7S69DRDu
5I6M/EOrHU+b7MhVranHKR39h6YoL2M14pm02CJyKZKxwbuauNdAjd4K1U6pjweQ
Pqscz14qqZs6zwPgwFSjbouUi4Ya4fZYnNVY2Xlry4vgmIbw0C71+RvXgvAhguW9
QcIu0gPOW0mV7iXYXBgm4q6p8KqdXaWc2CDJGCpe0ns=
`protect END_PROTECTED
