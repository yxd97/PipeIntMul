`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmChzfuZF6LfSSLYI3RgCDMWUrfxIWAhlYtd7D5tpIdBKAyL2Vcj9zhrPVA5j+VG
C2nLKVhsNiObQy64D5VhdltN/2EormZcNmpK/CGalua/Mx8yB7JgyuMMn7tFUD+y
RhI7vlG8gG/49xEHaAnlfd3W1DXYEP1+xdGSeQG/v3V4vn55MIhEq4Zt8b47ucHr
FkxH2VUhgM4NMYVWoJIeuudJEi14AnnMkNkANxddd3qjno5FByAA0nsw7ULfwq6M
fZxaWzq7osAv2n/MlVZP1/sZ+zKMc2UwAu9ZUHTUNBV9KaJJAZO8AaZiuoljejPS
sKlQJJyg3VDqu0RoIgu51A==
`protect END_PROTECTED
