`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4OoXwD43PYhxyc9ucAI3yftO9OHnuxLekCuXRDcqAJbAixju+6xx5rsn6vcM/6Rm
x5daHqdRVSfMIke80rx5EBjfBziiYcHQ+3EbdVz5JexldmfWJKslmJoWwycPXNWS
wIH+rsPzdBuQBZlewy8M7F2Kbgy6Ty+t5GM0pL8Ly9KeywRplFV9HFzqwGjUhlTh
f5dDpVXRBbTmijbTjGn6+cb8jh8ObmvIVhyarxByk7K1CpFWB7FtdzzYgFe2jHsX
bI0yjkM43ofp9iVj8bBhkO2kVJ55vfKqdkjWO/aaA2/8q7gEeVV0rV30ym9So26q
nt/s1zNBlPybWfj+IMeGTV16nd2f+6vmlrQamhR5FU2b5Rxvhz1/18orL1rSXws6
sBW85juaklJu6iH7iZO0WK2X6SghuVAxKrK1fAjEu5w=
`protect END_PROTECTED
