`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/yKAfDV0oBqzmWdiWzgYidJMxLvluBmSVbsvtK5U3GqXylc8bMoNoAYDx3FFm8Pj
uE75ckObsnJZSwmF/6WgSxu3722tbbvv41VzINras3hOhpQ8UP3zsb++SFVYzoat
KaW0y1vJouK3L4+t6z9lsopFJ5PUv1j2Gyh1KD/3QRzNq5Hiqa2pcjwq8ez/L4vr
/VCai/hqbxSBQBBKYxLWyCbp7jly59Y+TUQkJk/xKgBu4BCZMIvngHNL2YDZn3Qa
c0WAwz9TbjTk4P23E76rhpwoJf8AHuGR73yWmkeSSiX6+z57fIwB2HULmGvaGCmq
VYM+eI6dAASTjeW70ve0VCZO4B/vkndmWOOZZPBcgLjGRx6jpFR36J/8BONxzN7R
SSNbh3HtME6Cx1RSWjDGLPr1+qGpjL5x1bdyodgcbRVjyN2Yqnb2DD8Kzl+o0tv8
a+fHKEJpZ8guYSCCIQaIuA==
`protect END_PROTECTED
