`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2fNe2r0g525yPd9k+BmV1ezFcpeRl5NqOgbH0wXAZ4/iZcXJHf7izdbdgqLV+ZnF
IS01iwWGIv+CsUfmyTfm4g9MFgN6ORjG5AMnKwiOhaRtTSLhGt+tbnML8hPYKx5D
rBm5B6OIf4K7+DuZXzdgxUJ3moF65m3uMDUB6lFxby1anfPqSjI3gLq7qoCsotSV
tovjI0Z4f8uzuu0j8bM+xtvBNLcGfD5LKXBf9oyTMMz1LsL3L2N7/entjaFim1bG
BRaQuJECiFsMEZ0kQV4kybjZ09edBR0PRSUJAeCaAUtTFm9/QZFv7jhRzPyUKJwi
bcCkwMh8oljx8C/De6hNMKTtGgbIDqPqYzIyBowMTqXPdlgQjm8GfWGbyXLGM2wU
JU06ycJBFTfFOG58AydSPCLjAvwkMKCuZ71XGvUCRfhDGVLka7wUeL7Xf4vB1eKN
TZhus0Qhicwr6Xn3qKt062bcLrXzLo6l69RNGPWLzMnf7DYbnbSkvtq9ZlD0Ij21
`protect END_PROTECTED
