`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olApQ6KqdC8aeQ6WxXWo01gW2OeB4pRb7IvmDCb3SEJ3+Y8u3vDzLm8o/kwXZzrC
sDtylTOfPNPVbI90SkX0m7a82LJICdJ5drlfyI6BKegEeOCw0YevPZNFns662fiT
CkXJd7G77MyeI1iBlip6d6GrwlNfcHH4/xWeiQU5A2ZjxgLZK/Zqg33+RcY02KPN
xbDBrW61Eu1nN+lW298u15jP1W9Olp+ZxM4m4CUFm5j2vVNpF3MP+mFosVf0hPHi
8Pe+SpGVWpFyl2BXVlCCmPSBzHmExWWnUmbGjqiBU/r0KNBTU3I0iQ07CDZqclGw
mWkrlKS6CrPnD6PZ8qJfV4TyT4k3EnV2iBLx2ffy3spS6SQeIP6O4L3RN0RiDLyf
e7jn6PLRwYG0lMeg85l0LMA5puJ5bwxCnOqayypfFk7aBCSaPXrHmRwBdLF+lsv2
N82wMj+PkLQfg+zOfYw58TkeC/WbK+a4AbLdUGXciCNC2nv27WZdLqOSKjilEWtB
7qDBhXY4W5nXWthePSKWmALDNLlUT8YsFbZJR8NugqCW11bUhJ6znerSbyoBeMtQ
fL4R5QF2JDUJIuxPizaumLaATrsAuTFsNsLoSmLT4iOLCovrVokpG8jXJqBiixcR
jM5xfGN+z2UrkoqgT5QGBvoU/HHAJkLEfDkDst7dHzLEFwF1gFVAAeR1Q8k4uo/U
jJy3l7k+/TcploUx/trbr5zZdUN0k2HW484wTloGe3Y5YeV0FuESWmL2CfwuMl9A
mIxBJi2kRpaNlVQ/ECme0CNcZUy7rxeD4g3iKxwSlUsj39vUJFqrt6pTXGpiAw0S
esDr8417jTOPDqdLCHS3UhvVeFfQl4B9w0Pch+XgtPSx6f9pzxCf0bavXQhbhMdL
rsTT6+GpLgGsFQgjPdY1nRSuD3Sos7V6rVrBcfAQABV2HYr2uK1oFSRvonppm0W8
/bbKtXO7vkQ7dbIEKkMV9YZh6EEdIU//Tn9DYxOJ8+iSDPpVdCyofB5g8oHgeLw8
7Yu9Cbw36I73L+bdd+sePKPQ4D146zaaPJt6J71iIvnvuUtm+WvGG7VEplc3H3Rn
GdPdmj9qU24g4qC4o44HP0hQjmwXRPlFpwsw5qZhdPUgrOIOSuIKI5YPd1LccbPH
nXiKQsvxUq7o5VhWrHy3e1iJhhGuTG0q8aAzF76+ywEyI4Mv6r9rEc7orn4IP1P8
G6mWFYufVUYjDwtRB1yAaKkbeA+2RF1KpiH1ZSl7EF2Yw8eW0TJkM4dQPK3H1eVs
MS7TDbl1UjQzykCOtYSR3dp7mnKH0AzIaF5ejFtzVVVv2MW8zn6ZXJ9sUuEfPekt
w5r8ArZq3UeEY5X3uqmtjYZJLKs7XjW2qCfqaHaHX25jEvmQtFwYP7x4225vI/+N
/UJDwWUA/zUMyscEDRhzoRD2N9KmU6YidP0jr/Tad0+QjeyCn75TTUpiImxoAAh8
WdhzL8M5FK/0mGT853MgNInkXZZdGBS43GeQ6pntSSoxhhIU8V5Ow7HdmxxE4xVy
kNRKZi1Ue9LOEyCwgjdsheHw6ILgv/a7nEt+D44CR5swaszjkwWvhbtSDp2MhdMV
XKaZ1BUZb/S0RsQYD5uKbes0y8osZlOSROWQLop4077PAk4+woosHrcLxurG10M6
a/WhVdFXTWssA+5ISTigH6P0QQVOFJh+emELW4s/+LFdKVleGlbJmzFwyXpARMBT
pn+LiLU/LF4ingAUWMU8nvPMW9l6mx4vTN4WbnCZapFFtiZp6PAhtzvRxH0PH/wb
/lzvTWtzTgDWdFE3eVv3l/O8WAAgdmXCAiuspdizfFKM86rzerx4Pg9lcfztMPuq
zByJZXuwxCe8hk6riQLfmLj8TgRWGuVFu95Bi2OIygezHby0hq7oDUPuHK4+MzeS
o4UnKbIz7DxiAs4vZrtpRO+ypI6ftcF1QCGpVxJMzHvNjGjXa00vU53NFMYlus7d
ADvqZUZ1undcr0cPtbGi5ktlh+SMfNAdlAMsuMJyNVnt5wuHfgmxVsHBoODdbg0W
zVH6zqmcgmoJqF7ofDlOBvZk4qsHKySJig4257mOBw/wCEBGmVjkcA8PRO9TkTfl
YVrpfHjNPtG/kj8fWZfOM8mGcVSN6GYD8cIBXAAwrHV5I8HzbYFlyVM6CYfP/cQo
hCb5qx3R4UZ7mrk00gc0UjC06ccBpgr7RQEWIuyhdz/42buKaNgUdEigFH6681M4
rGRPOFMiTVPEeAQbqm/8O+fv+XEyW5o4I/mI9lWbBzIBRSQi/23bYG8Nf0gk7+YO
8PRfSWb6803SU/+mFg6naZrR6VVrjHp3IjzwZsI/kn2muQsM09pDD5mh0W9DzgS9
t/BHhbq0mOthXWYUD36myefMoXZMTFiki8saG+kPi4h19IapJ/IxeJqNDRK6TpQS
cPEES7VIperCIBlK7LsulXcXAGb4rG5B6js+QNNPEx8bmhlCrbcg/R/ilCoztahh
z4HNrGKuWLjRQ7y7vRbbGbRu3oM8UQioOLC8NTCcK3LrWtF6KElyjwAZJu0+oEbl
9/OjQ9foHT02V2HR92zW8koh8TchsZM1M9eKRm1DuUlyTv1wOIvDXmAUp4/GeUHB
XGvqmAc9PDqrIkC96lEfLe4FKZK5+/sdXC0ZyNBgFtbm9EmMb8mqSbit8/q+b9Tc
cd5pa4MJipYlKcCOqyEGyTkEzvqUQ9r/8UvEi86V1zYemYQymM+bZzHk5EgjSbH+
jJnOB1ZvbbaQEwG6tu9YLeR8hmbGMFq+IMQDktn2s2dSDU49705wRNIiGqhBAAIC
XY+ewSvl+P5BOhwiusqrNUkVOvZkDE7j/xvBlRRzX82lm1JUoyzjneb7QKliXy8H
0l8KZiVwX8Ibxi1l/oqV5qZ9UkWNMLUcXXwZ8/dBW+cTET7ufgK/Fv4h6u5i1Dlq
yi8XxE1fPjJFLGRbG6vQPI/Waa6MM5ysDKBrBt5Qc5GdtegGw+mNbCeU1PCIHDif
xeIeS7yt5CCTojYROrohE0uxLDJgF/64ohs/9T1gLOZpA6qNp5N0caOtC+27Xd3D
58Tzdj4hnMgw5dqOuAs6RkHQWO/AvOeGxy3EmKicehaaEjTzFU3u3Zwm5FpmQxN5
XfU3wLCS1Oq7RSCB1FgSr1ebWsax3ZMapDeMmFNN5FEvATBZ93imNeaz5jykCxol
TGXS5PghnqBWKO6FuNzwEe6fWwhq9JAXxxW/Smf7xa3XKqEA4Ou8RtomKZlyxGhD
Mx8A0iC+p1TGgBMykNWQcWZ+Mik8AJidASPD8Oq7+jvQbvyYffEr/A8gf1vwdKa3
+Z7cci5g3gbf0c5sQJ08qkSmIz5txfT/YmUyfphtAzIckmJdMlFYdOwdMaiYmPm9
f3PQjxME3hfPHQI16ork8RxnjOyjaat1H0IZ4Pqhi+G3+d13aR9gQX+ej25++Okf
pvDgmeEuoM5Mm3bXe1e3agxUFOjtZj/Ft82nrzELsszWQB6EieQJq6d07gcGkl2Z
Wn4jMI+pZ0d9apF6gcc+XJSP0FZGX5LSUjhIytBmQTX4knbWOeUWkgCvcJ49O4qC
SRfLQVpSWS6Io4krmaA4EdGLT5zwRIgXywhmOtirw7GXH3zmi/R0hg6ORmXZQ/3D
x7dR4zw61yK6j2kOMYDoTKRfCneXjbYwF14lbBWkZL5/t3v7PFxLpMXjY6M13cRG
gT4cTwFGgK5bJ+QbVnMxwVI8qBXlL+uqfa7CaXdF28QohmE1OBl+yJnFMgePh7o7
cEib55YlYNUM2ZqKahUZT3Ya49Wjj9NXYR22vTqgKQ3o3HYRK2Oc8j3oBWv8Kea4
byKa8O5ZJJAwRTYMXlAT7AGzhEaAxo6zxMFyvS0NEZld/uPfuuQmq/C/RgwlHwOm
UqqNBp1fLS50BWux/MZCI8f0Iau/MMRAMdr2JM3CAt1x1CRXfUxnnYAk70kVtkjJ
C2TPzhWHwrdHajFBMDl7NhCCIvyQ1WyFj8XVawaNqdS+W3PSD8hrwNMgp9vMNTCl
K3lneI+fOhVj5WxMo9srXIKRN1E0JITWjSkGD2dzeiQ6PCZtpNxxcdIql9+i3MJm
x/XThwgT8eF4a3GGcrI+B3G/QrujcIFUtDc67CKNvXYfnEhzsxlQewxG8poOiaXy
FxZeKwvygAaLiKTeZIjeKnGS8O0sdaAqrzYYqg7/z2AHDlXBfYNGtUte0ThO+55f
AwKZY5yqViUBs4sXNujHg/kf00aGoOOTwaBDzLDiJCkhK4rx5tONGXr1gZfCjlTY
rmoyq3CIbtGu1m/skhnUgId2Q8JOqmPVFDGKTXlL1OlYV5IwQmgE1UyG1NPICB6R
MqGe7LkEbaiUISvVfSBjbGRrbD0ow0nF0nlbdT9ghIR806qHQpP+aQolGf2ej6Mo
GJJAHc3AK2Ub92HAkz0LpS0fmn3laVOQn9Jjli4lS0DrWlnZA6EXoaj89ZEBpbpA
d0YyR2ZI4n0p7RNmRLGTgdZ5oyGL09qPkzGokbV/QvFSanElBmKu5xWlnP6q6lvX
uJP8gxuy20ooHvA/p1DidMmA0W4PvxUYih4URNDo9ECjO8mdoabkpuWd3Jv05Gea
+0f5PjuKvtbnRN2iW/QArcgNkfpgc5UsXLEmWpBNOMWTBtAJg909vOQGn43mTjMs
RqujPCLF9izGfxF2G6KhEAVS/laNFRiPJ+5vspJ3kj0JQWwYw6C0f8hMw7HhHyrM
93CL/RZZPkTmMdGAU79y8Vn8d4lXT9en+9vddNnbPanRmd4R8UC07XhvI5Uxd8bK
R5tLf7pNc7+ZQjt/7hVY8P1992rV4GMuyiaW1bBPmSObie5pqLsiajS1rxXqnDj/
4eOiqj6c0h7KvQnRBZTJ+cQq971cdtCBR1VQXIteZieAqFsh9nzpwbKIsykzRKoE
dkGzAmBIlqVQ5jL66KBdMebuxVsyDqOSzzwvUk1kDpHetmNy/ypH0POSSudrDbgX
FdfoIMq7RNXD1nGFPm1c/VsRXmnwk9SjESUpo8p56cc7hS19VYeTmul7wsgNZOt2
/3YeXf8exVaxWA6fjNkDmNt6EbiQoBRBAmpI+D/i52ExocfNzbckBRxDik65oG7I
W0p6IrVWD9UGU59R7dAjCLXPho1uJcQJYQZLICoMhU6yEm8hEJrfxrsHrghpvShA
R2g5Ti8h5DRy1fshW71EHaZufwqfj9cd755/KiE1on/fyBpb1kWKtvIJnvId3Iap
WfvEFb6+UyM2fr1rwauo1HFaruiHhqmbfEA43KJN3NHjfKYYsaXFVMWB7O6BVHBl
8zmKZ6W5ve3EZH7yIURGSIU5nCph67WB1d8xQ3PJJTy4pmQjKSbPZIicuXELpjM2
d62RSCNLuG/xipZHhGAp0KFxG+nGzKn+fmV3EiunIO/sTmkjKiWQCsuumf/eAeF+
VUQh6NiCNYSkjXjzJW8vom+CCQMBS663ioIOcvjtkXJvnMFb74BYV5cNUAvZtQgO
0Zv8trwlC5r1S11WiSXSgQ3ZAz8Dqk5i31dAueXvkU3zTGPajlTVntgDvjb9QMey
agkNPy6dGiXmXGmWWSZTGE4FfPze5kHZBUknvVojBn4jTf3tbq+vsesa4/UX+2XM
orW2f+LD/acDc1GEcTWOQQ0OodVm9yNkn5GWNKrhR9373a9Pj3FN4NVgz5PHcqmw
1TTljmCOUB8+FEyi1p2oI/+aR3+Vq9oyP7lPr8qErV0K4FHTE3KTDf1YpJ6/RidQ
Aitua2/RkykEHOj3v5mv3zx8+C+rbnI3c8qGJSRdCirITKrY1lU1xc8GaYm7jDkU
ZbjN13q0bo0Pkbza8nCcd/tfd4cMzNO+0hehgkB6xPYSGzM0iFHFNJT/t4KsSO28
SRIbAxHa2rynG40tJIiaA/SdGo47CHYSOurK1eIx7E6kbJJwqBnGIE8Q1PjZ5LxA
hcQnc9fmDY4TCYJHMkVVSVWOgXtNj1XIloVSFkwBWY5dNbgkuNHXvCQGNXPikYNO
4FaII2+R/orVvEOygvWjBH3nGjAW4+iFOLX0lY0/amntrLEsuNGMv8/6VwTJ5SuC
vTtCH2oPegBkdaDvwn9Kjg8MV6TqCzRGM4WoJrMUQsfT8Igab2xjB/NajTmGaAbY
0BGXMnOgROSN5lvfU8h/943QMWE4qkryyFUMS5nVyGvEBnVG60R+mRvzMtx5RPe1
5r5dOfmthG20UHTkL2h3HZ/nKUDApbaTOOlLqfUoqvrvIVDebjHeo1S7aR7gc4Ii
pKUzYXhYnxzlO70QZZzsz4W7r8bhPx+IYq3aB+CtazbqVD+Dbf6Ee8g13aNhPBRl
TToqTFBQH7TikrAbHYCT/wY0OswcLnmeyDGwBc7y4ag6FKCmer6jBMR6nu8dtt3R
sflBNptjp+TlqUpasOWV1GyCSIiXQbHKJgfllS387N7oGyg6Lo6SZfOH2xjStFpp
sVPUw+YlXeJLfL4Chnghbdm1+34iohB6DysnW2N3FBPUL+g26AMbX62sPea1ntiN
fZkWBkECmtRguKab8QE/Yy4eIVYJZegou8//ClB3Yz6RAdU8m/Y2K844Iv3TQOrr
wRk5Bc9rGiqUP3Td5PwPWxE85aM7Xy1RkBT/jBsC4Hn7yx5qOj4pLOuYaxGA6rv8
yQExCT0tqeeM4FkbU+2EaSi0cEDpOhntq6ekFU6aWiVT074b1TO60BAPzxCiRvWM
apqbFW4CaWsa9Z8zQi0xNay4+AH66xl6hdJKJQO88mVeUJF7RqaGz4jA1ApvV3s8
LrwQVud951GGQe4wVQNkfj44YTCqqH9mnYur26sClgEn5fOz19uDbMXe8/bVIouu
ayH3LdGqNmpyNw5khHEdY4VEbIit/XUV83DDNBrWs5U4fyf5hRkEgVg6LMp8RXQz
96qY86io99iMl1jKre7DA4Dt23rQvt6yGkOAXm2ZaqtfEGnzH3hBtkbo27l5dy/g
W2dSDkdClhfc2/Zq0t4wxOAlW9ohrnrK0HP3bFPzpqJ4ck2lFWiomjit0gomjnm6
4YCmhAwq2HWA2D2mmuUDahvX5/XEvEnZyaVVt2/tpBiSi0UEDUpC9tp2FcmQr448
4kfJk1WOpj/4X6sDT02qymaHOUqEg/s16SHG0RgN/KjuRgBQ2dUq6+92+g6eAYoj
EJXTxOIqdLgc/GtpfvCXUq6JIJsGGiX6VkLc8K86KgIrONc1KDCZOl9PeLJQuxRn
Aah4DDopGoU7lwTnyYX/nyfQSfFoJohxTldYfMrO0HesVhoQutVuTcVZqRbp5J7S
7vSOuCaTtoIExsEO+6+bNVYbv+Hy7fX54vTp09+Hpvv/qp4TlUen6E5grva3qgIL
u0GCy/Nv6R+20mA88e7MQ166bFvCJ47a0qOnlyeY3SOKNjxCVzv7g9ttlK9FkiX6
yGhnUCnkd25CaML9AcavasgyXWSI0hKHlmuevB8kDj6Bq5v38TWZ8S04o0rOix58
lZ576JJ/r97D+PnOf7PsyCXsc6BfjcSYV/gE3x5QEt/71yzwVFTOBTDvLl4MtIY4
wWP5ZjuRmeXCLqiK3Q4Dbq+Kbq6XCdNklvFN5g5gChxMOgxrTUoYYgcJ4ui4dAi4
6huuKpGyHEhZJIn5A94pgK6wmK5krSPT2BF2eZLYJuiab6a8sEiauvIgDFwkWIcQ
Aeniu5jS1EqB48zKWHpu4CSo/XvZh34l4ptQPopAu0wdvfznQ7n7yTwhtUCGvVq6
e6HjDXCgFhRV3rW/r4mkyHY7IK2cRYIFO+JAioJk08FzHTVQR5WRPNkcdP2nS8tV
7jqPoi0A5c+Jxfk5tzBYC97S0E2LJZkZ/7d2D0dfNj1rR5bPmlz1xwu5QjewhXRF
z+CgsS2Xi3qo30S+lVcA7z12YLYpow8QxM2YAk/FpEBYVAews4dmoHXq89WkionJ
2a+3x+t9DgX/Yb/o1gNwuBiZFUdqG1FnZsemXktACjWFJvQ/rgJ8Qquc7HolKWVK
8qf7NzSE3HJ98CYK/FwWnEIzItTrnjU/+/Vo2/jKGDauo5vRKtEknajPQpuuImNF
OutHUGrpzZSgHlI0Eu6B4XXgHuGQTEJuUO/D5Xo/cB3dXhPGL1SnsmJ5QDwidku2
Yhl0GBaKnd3zogqCM49NkExHoWe/akPj1Kew5MiI047Eoitpqpa5S4wykDmottHC
aOdaja2IgytKsvdJuQtEq4H3XevY9HmfNNoH6VFkeCMdE53vzHb/o7yP6SZevusr
fskra/Po564D2si/FqoEZfhwD0r4qLFN/Qk0lfsTBUNrNeaM6emsIXnbnmAR/fsj
lMNGJrkEvlC9ZQvHuKU76zoWSDIO68glrbcSnU80SEU3YbkE9hw6XqENPuvgFak0
pLBv7/wn15cDJyB0GXS1SGc2gWc6CC03NmxnPhlQdS/2u338SoHufXoOzE7V5LDn
tgZjVJOF2kkv+XMAS0JOCxVIh9Qdmqr4vwBWVDKBvcIK+Int/d8dkYZnqskRyae6
bpjAqo98AfoYq/EHy+2OFo5GU7NM4lxL9Z7fl+1KM67upFHITTCFI/OZ0t8dEJxx
9QQ2td8cT1yC74n9hG5gwMXn/GzK5kwG4JRPDX/In9+1In1sg7zshTGolu40lvOT
pSixj0/95hFsG+Zb0Z7jFTuKA7S/SkbK8dS6NEq5shVSj9i0ud5t0AFYXyEUBRpe
2GOEnrmgCzVsji6f68/5KjKy+wiqYRVnPa08Qiie8xnOu3/fL3oCL//kQLz1+abN
Xojved1vz/vW2J9qpBiCehY3c2BwODdvVD8OcIOEF9uFWsv6NPYj6Y3y5M4k2ZgU
uE5QM4JEzjTbMZ/ES8x9fbWxhahVPEkeyFdyin472WajyAqf6cP3Rt0Fmtm0ODj7
pGeQ/O2fe0wA9mSqlhRGIeHfyFdc1VTbna7Hqqwkqo6jHsemb3Kf+nZn0E1U/RkZ
N9wE8HXD9/b7e6uMa/9Z/3D0c+POMj3SjdG1roa0+ZU2FmD6yzWHkmwbEMEpf2w7
Pq3ZVWzpLT5uaJ4f5zU2ackQlDZw0scPUbQl2HIyd0KyYX0OeCEFkVT+7tm1jiCN
nECB5xSy/RVPLtJRDDVak+6x7v1zor/nlAk4bP9WfFunSe+NYrKzgnOPxpJkgETo
HcmmEBuiYECn63EsGZnD+iIWYOssPxPMp6e4TrMpaqK+H14ShltOF0Ef5oM8ASWA
eNT2QeTplzaKT6wP6OTl4B0hMcrlrTmFmTx2TweSdS8mDMQtZkZsvz9JZrbS0+Kt
Qop4U6UVY5sdKihiymhCm5uzeknDtNlOKPlFc9XDLXNcvu7M9TN9wKxLcPyvfG++
sGWbqs1j8gMU9Zn2YybCTQMFkE2Iv/ijLSNXGzjTVP4DLJoMM2AVjKsie7ZGKcdW
x1LVqv0Y2ySQ1cWTC4HEqrz8gCUahS8yAZsu10b0LhwAAT6LkKgao7Xzt13HnHOx
XLZ+Yet+7n5Q3FS1NJWCMdIIICBDohlQS8Kq1xuHjtdTSllTBVvVRAzT8u9hOXU2
bPOKq5vM3FU8ltHxw+oBqGJsPMyJllY2vUrrJkzR4rME8Tij6D5HQdnDeQCk16FD
omW2f6sTjxiGKJH8mw8TYfZGIVmStvM3u33wH8feDuHrPJx1ltwNCMj3t1CS9wkO
x8pmadZyNTog3wmUIf8gnppiKIadunHVJI6zcemyIZ65aTOO3m6e5MBwCoM71Wcd
ewk4nmYzaE11GwQZiHweghXzKNmtfmXOOYKzY9ZLwEa/KvbpF68kLQNtJ++mIMZq
xmBImg5gPcTynxU+KL0qD/Bf18FFgpZHxYJfbT6gsi8GO/Vhe2QAZcTvwokS7J+T
iN91fdXdEfdmobpwHgdb4VzgLAjkD9GB+PCd0PUOMQ0/FmJtWjpnuJxw7LHK4lhS
yhn9j+68CT0zmMd7V4Aapexv+Gp22PyO+R9iBpiYixWHxpmMzupyc77Qel/ZPuQl
c/eNKONyjlT/khNCZYUtiqRReGazTuayrIp4zkClFeGmTM9m/ZOC3fA9hRfnKGA2
c7kXDcoWxNki2MZS03032jZQDZhnzDRyGRBYaLpBzlLvfhKZET2Y4OXFBoml19dA
WLbFdv3g8jIaTzukV/154SE4imtaYiGhi1uODbDtrTyefLv3bq+YDm6es6roVsne
faNnPZnkgrwHVJbOCRdr4dOyNhoWbS5CJTHszcTn8Y5ApzvgOsU8vkkAqz+LuRof
YpxtQXy/yb9bEKAKxCs5zNwt0pkEewEIlbFsxpENMIktRo7XNPccza+RvQCtDRBX
I2117TkHrRYqRa7uCUiy1nVj4BKLU1V5vtmvdkzulV0=
`protect END_PROTECTED
