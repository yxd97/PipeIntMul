`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OvwlF51t4P7qRHaB8+KeiBAcoEXgKvSFfq+gEZjisal7bfclSFfbCUenWCIBe8Hu
MNv5usq4/yw4idsOQsDoXhX+7QT4TN/+kBasDa9INntP4SJgYxtVfoAr5G8hvwtz
3+klklXQhslf1etmZE2bWrdOY/ue0R4+BVKevxhvHow2AACoDZDxto3hmedxgbjF
H29lhRCBCZy0S46gdfZbxUx2Ke4RW/xEBTMknbaKnqVlyNToAqF6orR6eFyovw1g
ui+H5Igv2/yPlS02xX85FsPQVQ57x8kjNMNIABkJTkFGIMuietNuPB8L4qwS2atB
UbMUq9kVxF7XWFGTE3Zbb2K9acmmZRZfDhPwS5b4XqTNL1QUBNpRqbyyc00XzxXb
EQZm8EOwMcBdsciBgQovl4OS7BSWuYzCWOjMDIpHBshMgS4xEfQtN5vo1y0TvCFS
3AHxRN1710v/xWndSihRjO38YmeZZuPnh++PKcSAe1CbrYGYWPp/R4k7wA2wC26H
0Tm6C0Au1VVfpozXY8Mc9zELU0zPXeCe/4FoiBUUWje5J4UTBCbXD5Ax2pkSzIpZ
Jso66Pfs98HJPDca1ts1emH8+v8CttrEJmLhcc8ubjlCDCTMWvAyMFKRxMsO6Wrg
zKyBHRmhOTfX+5iD0gnITFjmh2Ea6G5rlJRi+l/oTKNXNNhfmCy2Tnt0QAYi6aBg
Be7irFZAKOFSbN8+V7kMVMWWJzMvWi+V8lx2svwln+9+bn2Ibd2fDekgZGh+k8f2
ygTXbbe8KuCdIZ+Izjt3Aq/Zpj3RGE7i8ImugJsOnrKczQCnOUJj2jsgDf0BsIpe
8d2eNYny0I4awMVjDpqM9+J7nzDG0B7FTFrkOa8yqQq0WS+BIdGSS1MCbrA4rkvg
qvbkB9uD7y4uaqfBMS+sskjWKyCevOHULmtmxZUPDpjuxstujJFSU9WXPzkZctjC
r17buVSEJ+JzqZz8oVFnMKlWk8qt4K40j3CXSYPthu7USTkZ9sa3nNtsbPAfSHQ9
C3vp4t+Uc0aEifjujBai1lU3Q4b861aS7D+HZjMQa3TeWJaU5fQqfsDRjcjnFZXU
0UkhoTHQ0Voj+sASgfWi/wvzyW7QI94PZVcMf4KsVCU=
`protect END_PROTECTED
