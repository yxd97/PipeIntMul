`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJtA7gVtNBByLiLWKiwiij6lXugVDbSsubj7vuEj3cP/Rf/ZI/AkO3+RGXAa7lKw
L3lRpGHp04F7TBoUr/WPf2Xf54gAh/xgiXda/Mjdj/v6t94h/nv4fG46bP0Oyzz5
V6AfTL2BhbHor9DC6STqelKH/reHFt2VTQuv63pkj2Q+rRqRA3NIOzBDsVxxPFcN
DMWReV0CYENY9oGcxLJ1rdhf+h3wkYvRf44HLbzWBv1q/JPohuPw0rDbxrzSaDh/
RZddvn8aeiund/+eW3Zc2KYSRKsIVg30XMSkqwwRRWTkYwRzL2l5UFhKTNiE/7d2
unBOAJruH80PucI7HLilWdtePW4nxcgXhcnoz9DqhndYfSEBRUdGwcPOL1qOO5H0
X3d7cZQi2M7K9ftGdRqyyo9mKb/Vhxt2g9Vc5EfMkEkJj/7cHF1UR2jA8ClZ9Olg
VtEwbVV+XbOy5Hy0LCo/VYCaZifV34aHw2PixdgZa7/AYsGabhAfZhVy72bU7Ywg
PiktO7ax8yUC9uKRZ5h6eX/Uqn5p/0CFO0W+rOhGh0xYFBMgy2hTYB/3dGXUC/BO
EnR3oRek5lgEbMxz+zjXaHB8mXbSKqrApapGXABDGSJFdwnXtnVrjZapxyum8G//
3psosczLa6uCZApIm+Tw4qnPaku4sDXWzmYH7YSfRIRWfL9US2MvVnVrKQV2C2R+
FOfHZfBh+dHxEw/rGgy9HkrZU6pzrZjiaqPhiBdLFVc=
`protect END_PROTECTED
