`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I5SdwBXHpE8Fpy975a4FuHc2wGue02MjidYIV8GUEuh2WY1Wa06TdMAsdHpaOVAM
T2gJCD3IC4ASqmSDr/T086Ys8op3/e16LihU6Pgmmaydo7Qap6oVQ3e4b7fu7zVp
Yt6GGxgRsRqZoP3E6jsAnhBlE5vD2IPj6G9kuc7DXTiAFw5QHPH9UMRk4r4zBrf6
F1a2SGWZqNIXUJXt3Te94hjF3QW05vEeiONpG76UccWngB4V85G0uRL/c7p/Devv
HWm/7eWruWF/A1YfLG1HG1z8vnAp3mESk+37VzwWjOCdGF2mNAjEDG6x//JSySY2
ZDRSQl4UhLhUg0cDUTlfHua8Y+nTcJXFOIOTOJhvXmxIcCDY965m5T+cpgPAMNu0
NhmCIQAAJpF4uYxXv00invpRZD61NtareLeRKSZkzim3a7zav+16bH1zUkKkO73y
a/JUU1eF4xuy/Y575EOSGdvL+vghJBpeVlbMLkDkw1pFzw8tpT2QF4FH+jWHtnYi
+mwNbaJEi5sNw4ltnPeGYjhuh3eNT+wDlVi9Vw/TiG6ZNj6jSQe5AmpXjI2oThW8
4lqSZwTQhtlDqa0y2vPHejGCzD31JF03O8IoVhdbj2DXTQxZvIMgOkhOSNrbE/Uh
2LCMdBOZlUzRGPWDhNQwruKR+Ad+S8D8Qi58zSwsGFZ6cbDEaeIs2vSeeGJPVjf5
lZ1rPDxgoYxLOvvajQzaoF2HbIkKWo2PvzS3MgYE2QpOrYPDGhj804AtDPPuL/Fw
SNPzFxTCDuuSWodGjaZSOaUKA1pa012Kdg4G2SdmDxSb1oRRhct91DaMdFvyE5ob
ABeSpHEruXWvNnWZRJ7wcfzwm5G+9hqHKJcgEAzPlMowYx1itccFwy3wrDcwvf1h
qQhydT77VO+4l9zborMsYj6I5kceXCk5f7puKK/b0shMA8AA29r19tiIv6AK2O2c
I737gpR/IzFT9tPwO6mFxxnp+Ngbs2WNhPTa0s4I/cf9S0DVB1Xo4TLks3ePRVfM
lBERCiW6ncbfECrBsHiWQtWMde1xkUtRIrFz90tXf85X7UKIV1l9e3lBeWWmZeJo
FZfd/VPYs8+7oIEX5qD/5HXjBZeSq3HEo1Rf8WEU5iTlu2pa+5AtxKcDuK1+orQh
Bw9kfALbdjfkUIU3V1XMJ1Mla14J0c+0wB4PGMBtMB7twULKemSzfEhgtmzvEd6Y
iWb5sllqQH+RDN5W0CSneKW1G69FecODxQ68pE58d8C9Srk0xqD9DqISgk8VNDUM
noNlHome1vCtRVYusu8jA6wbU76RvhFtIDDVQGtVXADfZ1LSGIO4MJFdgI47lAnw
siDXZLNKAMuSBpCRu5dnTPgookqXkm5Zm3bZtA2FkPmy+OXPUkCJy3OSf9EZTabT
AbtQIYwBT3cDjNWJ11kXUQ9ZPT587Mo+Mrlb6Gxws03M40x7s/Qn4va5PN9hDEyp
VEXU/qap9EztJ0vr8IIIB9nA4hUrBaqqwnUbjliDLnrk5wx543sSMlqUF8qeH3po
NoL7S+GR61T9wwQ4sSugnd1AC5rKXsZorz9maEUCPOpJR9jNEF12tUa5PzGcA51u
mWZ4K7/JFHfgnOdztPyvuMKPr/czljAoImqdQZE/Y6I8gTYaJQtYQfd7oLnADj3n
pCYvjfJJK2oZGJHOm1B+NEgnMKxISacPX2iaKAruK5pbmUWpHH7xzFx9OCvm4PFL
TwqGHHKjMMXLD/UpB7RIzqKmk9DptulvA/U2yv3xma76nIUTH4zNP9eRyNyEIvbP
3HO9udMHW3Hf9dygwAgTPdRD1ArKyuqaXjJ/o5GRxgYxH//cw/vNf0ygwmkzIxrQ
HFW6ztJGyMdFQjWQP/Wy3ecajdTpxfSp2pJMSJwOLC5dCtqjHQOjTSSfdRdLRQnX
ZTi7JtcksYBflNbsyUqrwmCU/FGMla/JAIJlSsZDpCoN3gt3UUW7TLSJad6Jgx+h
SaPzt2sDlUuYKtfDCCx5TaOrNa3Z7Vioz7AZCsIfxiFcS52E+UnuV6VnQqyzEeHS
Z1mcgVN1lvXL9T7sCuFFSz5sjQH6NChT+cpL+lF/ItJDxSuy3B/zMOxfOcNvNZBF
lz/0bnMsCBn7onnDPjbloYP9G5dVUEC3MbHabPeuBTaZCfreN3b7Iw2dyYhWYom/
w+zvoqkXtCfZwH9fxMTv35Q+JUTKBEQ6A29snblcokQBy7VYEHlLsiXT1amForXi
lcw8pgnuTxKPHPBqwBDxmlB5kUpYX1FGiinzmCJJsX53jzEIh99MPU23eV+EeqjQ
PuRc7ow1vu8NlvD4FgEXBkQrQP1IG03E+syEX9dHrJ50pH1WyxEA9/vC7J0OzvPT
by2Mvk6V/PSS2vADMvujyLzpqHZM2zVrVAmtRkYiE9FF9BMaIs0dUScNN7a1ZMRW
1SIB4mC41JJq3WPf/xCkwfQ9Ud31oVFR1XlHKXz8FZ3ivpZd5UICpu6msZCugfdc
Xg4NT9s1JIN3U8jPd78HS/Vd/nugOIYTpo8ADPkalARfcvkf3d9ywDRySHm1DZDk
IS5iTFKZryh93wSeWwTprUoWS0iK7WJjxZiY20qG8gWeiXNuNmv60nZvL3FhXg04
8QP8pSuJF8LhjzYakSmqUP9Tdl0Tobcdk8tNhWDc46SATW4ReXYoajTAZQvNwcnr
UIYGXJRHK+80fshnqi3mVpO47OnPNEs3IgvnW9+w2rulEwt1d1dk+NeDLt3zwn1N
5i6nyeysEZo7oUa1bAGQFg+nrinFtqbiYQzBcfeCPtXAXes5/n6YiytFyHJrGbzQ
IEeG6zja3pxcxh5myuugGZqHGgi7kVONOv1o7D3F8tJV5H6J7APKNUbSDsIIRlY9
hX5JnLEfljvRRwju6OUwOfLdEi0QnrjlCLr3OHYXtX/AFQDbqvxoK+UHP8u5mbDX
GqOOLfLgK2ewdgp+947AvzNrtyKs/B4QIIfm3pDWJ0SX5S/qjnCCN50UmbCnv21g
rU14mNjnjsEBx0y6DRZgwcm9+c2KPUcusN0q35MdcytHs9lCsWYLxbQd3aElHHAk
/eXIWNWWNbqYNnOAd3uInlYzUCueRWrQuy67dhoVjNLhh4f0jADDazT1R3KjCHVx
wzOk/Sm1e5ApBqiPf9+Giwg1aTZAqHEjr+ApyYIQM1huxHwAUnKCiV3RpOaNKxXY
iq6rkJp3Tdw8pqQVhSsuw5ZXDjYy4ge0RAX/RYCLwSb5cpL2EUjFWo0mtEV3Vhge
sI5cHcF5M63yxH9J9qPZ9OQc42UOFA7G52JGgMbPI3rh0575Ug60JF6reZ330riQ
qeHBWpKHpyrIVEqbLaQoEpTFI5ubpYrnzPz1P4AlIFRBjxAjPcWYSRciPEOyKqww
iOBE4NJsf4WQkqGdWG8wTMXZ6Ml7jczDXvZWFY7PcsBCkRV9ez9alFxeU2r0k3ou
9iYEbVSw47+4/DRrrHLORcwHdWNFrPjfR8Z6A+/vriW/ftCKcFXl0dT00ZktKQjj
ZHbpNxo5PDl+dwSHId8xkZ0p0Y3E2f50LoS11ebfre+HqFv/4BzU4ut7wP1d0khw
LaAvYo2tRGcymL1PwWxakxCuex7lMwK0rNSTBCL4yUzNl3rRGIO8sMnGTmZcIOMF
+2B0Cw4kzHYYoxeho/n8e85UeLOK9BOIvOPQb9ZkhHUgYMl34hjdXXGeTkQf56/j
bglKa4PNiuSCKjM0mjFub7VpvYXoJ86n4jcGYU2Kqy3+uRaU2UqKd55uHKlRXU7/
oitOqvUQp0poPG3xD6rgVee8UttY8gIxKoxuybmxrhFIxo75XWE/yjKh5/oDTD04
1jWs1B2u0CJZbCNPEzsNPlaSRBPo7+tUCpTfQgZdEpkws0d1Y5JMe1k5UG+S/zLT
iO4G56M0y9hQwqc3+wdHNiu6Efa9ffaFDayWr/39RoVDduzLuxTa1XUfqXSDLX9i
yiO6nh//ADHRPdVJ21H2mttsDrjYlfloWIyY2qF5W0tW9Q/0riIZYPu5LhB1xPm4
UKmaxjXungqdRosTJ+mati0F4i4lrid9G8CxcJ96lu5Ewkx9xsXhbXF4rhCM5J+N
nE9higItFtS447wqZTPjJD5lhGdOl7ZDO5hh+TsEvuKWXypr8bwEFphHVwc4NXi0
z8uZiwi59FVtufyXTXxJ4ixaMLREvQZ+OAT9XGGvzmpQa+txmRObzMZdl/oL31/k
hfmLYJRWWtMD65CvKQ4Lr2hzbagqiUUJM3xUd+8+gvyJmy5k8y1uAjJxCvWgn24u
M0BBgwIzwMaWAfxPRIGFTGL3c3IBr3Ft9mNi79ohcDK4ny7khG2ya9Qvc+x3P1r1
j0+Kd6YTQVbi/v09WJDOJKHONtmQhc7a4GjluUIdfTLdWzwVqb6NgXdKv3fe1H2v
9TJl/n5lHBJw22s0VcF2NJvEZtbzWI8q21yuhxgbp+bdmVF0w4oz2PjLkzn61EBT
hizPw74aY/ETpYclnMZondVcLrT4wer1/J7orIG4SRdeuudqu4oeaCCG06JxHWRv
nVToyH5aaZZgtwzy41XXi2XtJ3oqB1xM98ZcGQNxfTLqIplUjdYQEgLWlUf463AK
qH28/ODbieREBhkUZuMa0lX4crBPvYtit4YgKn4el2MfFd2fF75OPthqjIcCnChF
d3KJCvJdYkkE3q1aBbCFI3lG0HYrWu3DM3u/SPR4InIPzbLvS358P6v9xQFjYLtv
8FdQdoH/fqexyW4jEckVSMp0eEWxZrvjNggXmIt9pSPaNZ1Lg+mSvuIOv9bxSGml
BRLfa3LgdAOWGahrfd13taYB6IwJ66wGJ3nulmlCt2bF0lYMglauKLaJx8N0Z+rx
zZIbEXKdBTn33+OCjUvAIQJRWY0704Mgl+4axdoIpuGMaYdHg9+GC2GoNJBUbVA1
3p7HqWCpDhHylCOgnH3fi8zzSh9DYVxum5ohdONg6NEGpaQzvSep91gN9fxv2Chb
cifi0nFPEUtNXlfpoKxkmLsfpllKaDDQ8wxFW109chpYdSvEiLnyMlbUEaLWLjhx
j/WxQX9RBr+m1RXNkOupdwlxwh2eN9uFwwgtkrfisBsCxMNWOy+kIZKAcl1cJ+dy
jRLjQ/R4Xjd0jFjOp0bdevEp8jC5vD5gjc9Udl9dy4QgeQXohgvkTxrWXfBzmsMY
LAWsIRex/HCUhvaACx+QQQy92VI8XFKKboxjXhfr2YdRcWurTJGBRb24N5t9MYnj
VmYjoDmB7bLYYG/xokYgzieWuXyiV2ve53UbqvEmdLTOK3eectxkl/XrbCZo4Kso
fVlIDQS/WQi1d7Eanyw7a25FweA1YXm0ifFkofj60DG3+Rlu1esOhDcW0hED0UYC
mouHawoA3Jyf0m2tUxmzNLZNa+i7aprvjHhX34iZ7nceRcrvtszoF/agXADPRuW9
YoyPB6w8uLL/FtGfWkk4vGp4Z7siSHHJTo2PNoinRU8c6y2pOmpyXpUi5CMMCf5l
DvnKk58iWZO4KVLiwkm9p19yFrFdkQ18H0ynSwBKb4njOXEJ159bjxYMOW1ufbJO
AOBGyrdtIA/5rajhTXJdKCUqtNyD5NU+Oi9cwUcnEQg=
`protect END_PROTECTED
