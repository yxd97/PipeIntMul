`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VUbbxU5KDLymIpBFanOznTGCY9DOWofSxToI0RFMK4b8CpZGBGyBU8ij9fDOIgOR
h6AT1ne2EL65km5DyRWOfzFYbnrw10KwZ7ebncgHlgbQSk/05CqbbPZMjJnyfwj8
6B44fTmzeoj81LZJWkESk/XigSCCcx0V2Hf0sTLN1UxbwRKaXaBIVN+AU6bdUXXp
FAQ7oiLlF61DdMVqnrX0dpG3sp3vJKR6tVxHEf5Q+xzNzx7gpfWES9voriCboIMd
KmgCOy1ORnB6wLsBtGextFErQcP3AhalEmlYay8gYauOLQjbOoCZF2NdZohx0pGx
0EewhRo/nmsAGT5b65C/IOkLmNrVr2PFuXg8oJzgnp8lZSliXdjiROVEjarIXEka
CBXVEhCcpqHYaoxL+ZMrXpUFcPNS+ZoiYc3n0KLbxE3TZUhQg0qOagvtA/ve43oi
`protect END_PROTECTED
