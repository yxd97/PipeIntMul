`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMSWDC7qPpg5QyydPPHSQi+x1ydITvuOwpYOS7OhBq31UwS2OigD+b6WK89XBz4s
N3EfuRscIkvksMtUJIdGfdftXX20DeWpIBgwV6RPxjB3a8Ukqw4uuguhZh03V22R
zjksahNZpnvU+MQJnHz0iADzzWvtXiainATqY+YCryKOi64ReT+uecscD9/ojig7
rDgxo0EEsSwhxtUPrBx/J/CHYhvz7BYvDNdWQyEr4L9EK8x5620374UViJs64GRk
ip0YxtR5gCnEJLc8KG7shAGrhPOAB/5xEeFajO2qB99nGewml3N4gowvvz0rmt9z
lX2fwlItd8nbw+xkqg1MCJpajYcdylTynH5CXJEltjCsIMGgTKMtexIGkX8uk66E
cykPEPSddYTlNmvwz4DzAf8UQRd0DdfRsnS8gAnHFVjWwY9lkhVqdMAV+RCIOndj
`protect END_PROTECTED
