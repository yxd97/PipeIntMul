`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2eNYUpUBMKKVVqtaqBON+GzxqE90xGTS971THi3SANKzt9hi2UX8ufI0CBXnfI+4
pm/rpGRjkMHs4Gg8ozW/3QnbRP35VGMz/ycrWvAlT3Z1t6oZo/EAMUzTi8Cx3vbY
YPWK/y1is3vbo3UaQL5Olm+CbkMBg/E42AhW9P9l+hqI5/EQwYQilJ0sTcrzRgTQ
utUjUYR7gmBytNmR6cduzFA3k3DEIr+R7yA1eyMrshbRYQtZBQTElqSIG4k50JoR
Tbnl4jhWi6J+JzjT0C/Hd2YanNemrIuG+IdsiISZWMw=
`protect END_PROTECTED
