`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
31j25ppfcdeZJEc9clh9mNeUfzYUSALlb5iY+SNQAYU+koSREKV3YglT4b2fqSgk
3uCB4NxCFC212W6JOoQlu5qQYXpkpfHd/Rfoei00d7/QtxOwJJjG4eLEGXYDxqz1
wT07W0jMNgxbhEZ3kYswh5UoQI/G3WfoNZ5hKApzei4m2XFjYCAPLgjXJWmqtwCo
Dsq5bcHhyjY9R/FQBvpOLfF8XQ+ahWbLTaUp6/cMjHQgLxEvmG/+ZxcKKO0iNtGz
9O8dVmWofKtInItyXbP3CziAu61jDkRFuHeN82YWakUlv8TaT3GHlL4a8elEsKQp
fTGH51N74Ir5Wb0CcIJ7k0Pw4FG3Y/1fbpP9As3XT8/WJO6wL7wzCyR4kcLS0ii+
xn+vVCoYUmgpUFlMA6uBjqtRfuPSwImYSHe0Cwnk5jNDF770CAW1hFNN4v6bYT6U
`protect END_PROTECTED
