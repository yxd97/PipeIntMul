`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HzWUgcvoY1hQLfd33vGF4C8qQ1EhxRR2olbz3oLxuQ765T3zb2QrHFPnn+FamZOg
qFpxfsIH1ZSOzO1wEryVFxncZHFxOFdKtHvmFb+Ght0R/8owNJWLAZDc6To6+j0W
0Awn+ldIcA5qB09Zamg14fL6mwP/JoLcb98F9lNFMjoQ9YmXaulhoNE/BWTm0xjC
uV90fYVCiCabU587wbFcdXPhaHWq6BR/mXuHYn+boIBqHFm6oQG2n1s6y+WUu+qs
RjdBe0Q/VruK/sAqDtDTBRTaEEIkvfmjlP8AHd3k1zbs4xUTM3NR5nVQnXEu/95k
WTZaL7oTDTSmkE0IrDgMAM+GXhFeg1OngJH88EcYKAU4JfnleunJFKoPiQVkIdkV
tF+m0qJLjx6CeULXC9FavrMSxoAAmWdby+YKR6ubj9Ad0h4zkaHFGM6lycgrAQMf
SZztp1zY6uAmR3ENUcgYVlq/qUbH2uUiRPeTafDv04Zc87O6Yaowb7Nb81rBbsLv
/2U3xHpcDDhIo1NO7r78ZdVyEzHT4Oj2plM6q9Eg8NNlZ4oaPH+c6ST0GSppxXtG
/TCwMu66D54rUuBdjGE0mfctn3Qsip4hI3iu3laJmKePzHmT9cS2eXK/eT3ZPXKg
pJ1pyyP8jDZICPdbwu8/C6IRsXsEUqE403/LtDFTEihAVxU+6tW4TEvsfrZTN0Ez
l/djf1dOZkfz6nQtePIRHLktyAqad+W93EavySxp/6b9BT6I2oS0ogA+EJxDKquY
bHbIInxnnsnIcA97u5qs3yWe27JJS6FWlHKV4J2TG/0K70VqxdocEMR6I4rFdSbY
dN8WpBPh60wcuuPL5A7Wxdqg4mO/FH0aBgcIdJcCjWaFsv3JgxzSXk1c1Fiqxou0
LxdzmDEiG/KQAwEO6wNpZRCAp+Zhxr0a76yqT0Wjrctt4gbZcFVpYKrdjz4sr0sQ
E8UQYdDmNTY5PZqcsM6gzRzrDgVKaD4ykQXQKXH47kOxFEqaEatXwa4w2Sda45YQ
vJvGsc1Iu9zKaOAYSbwBdcc0Gvl5GmZ99ENrJFJfeeuHhScmUWQYKl904/lmNC5I
4dnaAMKUMbLUUinXKsYv+oXx/PJR8zkI48mK0rh0cWgQml1P4ecsvbenwGBCexcx
yUZag2+VuJF29IOQXmqEd1/C1P43U9ZWDoXT0iUN/6n3C0FYprdPezoK8AJ7Vya/
Rpo/x8t8sddTnXdOAN5HdFX23F6RJSiBMrU+us0xKTaklLO3adVKlLXKp4OV4RVF
ghn672DN1WdUh9KyQE0Zjckpg4mWbtsloljvrb/4gA4ZoZDCy5sQuB8rSjmPqqyv
bntcGIA5FvNBWdrNQtT1YMkDR2PvGF9DkcX/TjtEb2w6gVZbzBeHfyUgHW8iG1l3
LsLe1drBupwTHeUASjqDaE+NPFLzFzC+lhT9LWRtjs8sRPgtwHu27PEcqsrH1CNO
Wo+Mzx/9JfcpD3DSlUlmuQGsulGMAplcQnptihj0Vq57Lak1VWBg/zK4yCpnlOJ/
rwqbPdgp+5PNN49g9+kxzrrxTbCAlmzcV5iUGgNu7XVJV9zBV1SnndKadZUl2y7z
eVx1OlMFi46SUQ66z1F+6B6wBylK9Ko8w9kUAR4zgGR0wqYZBcX8wjAj2W+19fii
imIEUZE0+uStIzznsp5iKQL1i9uetZUxWf4vbwdOXLpJ9nMvegykqFa2xbLaP2mh
YHTDSfIyf3Wq0GX7BGsZhQiDoNOOPg4iy0MjEZI4mNzInvIk2O1N+L+326a8ROv2
3ctKqTMDKM3XhKoWi86wsWlbxzaWge8pHGpdPG6edELIhDwGdaRl8+lcdEQUxBXz
TFRu368ODTHQlb15b5e6V/2c/tJ+SP07aiXV+hgWkMH98KDdaTxMC+HaJSndHEEO
ZQbNbdpu/SOUbJyIRjmTW3FnxSv2OqAhG/8LpQgP3H93YEhm5o9mYnWjFyFEPH/h
6bWmljwxcxZdtYvRBwKMcrWU4YsVJDn1iA20FfAMsQeOifAbWzwHDN5y5wrwZKBK
Symy49VfC7DQvpiTQwIAdKqAgq9M5sHyo9ByDJ8rXEsI0c1QxpwFPyxt30ormMT+
uoNNUB45/SckD9JHODuwtWew63/Pf528kZ0OdyvHxDxQ7omouS4EQc2FdvLYrq6s
0E9nskWe1DVKR78q+g4HpY6X5RaFT5A6J553cLIdCGTqXciKwhaPKXgnvd+O8dp1
d+muSmuZD/vgaBvABFO/oHgu2lbJ0HgsKgJLbyAfWr3bJ7OlXMIk8EAb4FEve2oG
LoZLNPzPvUT+HV5ZAbO1CchoO1vATqZSzKFgGO53WIknNRg3oXjf7M64qJRvYny3
e+tWrai2rTiq9DjXAWjodh+dT9hquTQcJK+ISKkY86DH+/Tfd5QzUeXJ1S1bj0SL
XbzO2ZxiMdpJVlZXzWdMQbITdEZnlQsrKdGPQ2iE/Tar4BE9mgoXHcsYfjUKIQV3
W1dVg5VCkJ2Nz+XHTWmhMQ==
`protect END_PROTECTED
