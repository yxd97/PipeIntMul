`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nSno4N2F8W4pAKWIgTF4QQijBmSfTdM+Y2PPa9g+zbjVL8qA1XaECM2buP99MNql
2VwXvwPqNRcjvbdp4O0tGjXTsrdI+oHxR0p6dmgp5KswTaoUeP+kEXQt31EUapRs
NLcbBQOEaWiZRhW7e1L0jpji5/EbKQQI2W0oEN8XPj7xAHy7AuyWLYQC3NPchjz9
6TW/5FYH5OlkJZkzqSAbxJ8hTrvAO348Wqmct2qw/BfdM2bsVqvWLK3sOJjLi9at
UBUmK2l6lgQaM8JXgbVsvRef+jL0cqgf9Mma3lVBXxgS2E8nzqhoqMNILuqH9oI2
VmgGgIcGKW5ZUrWfNyE9oWJ8KP1NfzARWZ4kExuS9AiJOB3mSnSPa1AYNGt3Kx20
Hm5ijyJpuhQJl37vE5mViHxVlIlowTXoXDXAoJeYJuRMCOcFgS1t8Rab6Vf/3fCN
lb7YcZy8y2XKRissyToKyKFCDhqtFTq8yajTb475Tk+ZgTHsQrVXM6+HuC9JnX/k
uNyUdjI9EA2zj7iGOJiarwz4MUCrr14BolMWqztVxxyfTlpnyzfHpX8B5JgUunHD
shtxJM7NXmeMwsQz9QLLoupY2BDMfMbg7AP2zu+4c11GxKT9nVjSGVmdrIkEngfj
lMholMk3ApkU1QzdsqzRkMkQlhgkpAuMk/tYO/FXwKbN35d+xaZc+M5uHgD2bF7D
I8MmbsQ8AwYl1ubnofLlNMnx3xZ/fqu2AnSFlNxGrlQ2s0PwUmFzbpDiujR6nmoO
dOWBI6bG5aSsNdNkyCCX+ICfWxHy87NQo11lw600GDzbTyxtB5xhdLtLSutiteCO
7FbPbPIz+eySDU58MzfuIYMpAshaSyK5WpFfCu49AorBS7UYBFiwrPpo9RHvIr3/
cB+2U7l1vuzs2zqmdmL0RAFEd4QHcuh6Ke0wJPeAcjhHzJRQyEEZKbmAeSW/RPCT
iHOQ03P59m0ruIUwlKASFFkrvEeCZBdnK2ZCwk+kQCczL0oFI5L/gI7n0R5wsNtK
WihKchtzMdSRxf7vi/2StBBDP2yk5ov84zV9lUoqmmyOUjucYSUvRWjduO7HvzrU
z9ravzEiS5U5khnbueRmW+qvqJQ74tGNR9240phrjI0rl/sPBwHjJ0lfVi2FNGWw
HEYMMxkWLbcrM0EZ4EYaH5HrYrPYdahReSsIn+izl6OIX6aOqKoZKV93/Kjh21wZ
BRVjQnTy11Q/TFgghHgfz/tJUCyWaSSy0sEZ2i+cKhXJm0ysnn0vDA0nR63bYnQP
cbGHeHstkiNJvfCQ94YuefrnYky9fPXWOJ5m1jbML6otVVOgt2PaV3pMha1r2/Oq
+RNkLZt6n+ClsCp5khQ8l/3W9nBoerJYP2oC+KYpXmtvoYvF1iurdT0JxD9I3iN9
gfCTyZGMYqwtwP5JDG4nEJyO4elGqAkgQ4ZelpGo9yxv2oizN4fl651h2bqx9O4c
v0kLAHHjAORPcCklX0zf4QvAsrJX6/vGWl8zXkMNN84jhtbHoINBtgBOEFgkWFAb
JHnNLw1eOcB1T8nNb5DriUJ7CVH9hr+MzKqKlkwDSSk+eyAqn6L8lSY3SfIGPH2r
FMjlcrJ/jqJGq3CkSQ9uK3bQd7ZZmLX9iYXy7kNJxooWLxqXcpPwbh8zDGwPbnUb
W6q1jEKktPf9MpwRo0odXnURMVwVqQMKHi2RFuiTOKaHSv/iL01kdSDeOsKZhTwp
`protect END_PROTECTED
