`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GLi+No6TqEyoaf/nlWjRdzQHKBcipZW2ngk2rf7SGpimA1qxkCOrZz+iuEYa9/Lx
wBHa2jHKC7/lN3m64Nc81+aPrRhY2bliZD1kfT6OVBvxIU7DQfeuYCjHgb1zdYNQ
kbE8Eq6YVRe29xujNfXQFGussBdjsI4zInBMQg5hwdU0wU0puIy0+VPgvkGuCxnB
UyU0ZdjMRfRAboTpXjmK7hsIDaVEPqrfX6i/vNMRdcKClacH2mJZROA/nJrW/c6R
VnwI+bAT0gdYeYusprmP58PZkQcTRHZh06dhZxiOHyrpyfxDFTdYj51I0hHFuAen
`protect END_PROTECTED
