`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
akc3hCZx5/KztfdVIStYRzaJPpEFt90gwpQNQNWsZmAJoUiLL0VLZeFh5S0H9Rx9
jf47KRRrKk8bm5diJLoq8B9Cov8b3A3gyeNjIXEDNsHgzZqmII/deJ9CLDfFJ+fi
FjSxeT5UiCr7+NV1Abr2bPaxAm6BXV2ZvnNUBVfOzoZWMIwYQRF10xONWVdZIxRZ
dWj0oCKZ7vIzjNIYUw8EmzRAnkLi61q/mTkjAjOOH5axEPWwaUMYqYeyBSn3BGjF
2oh2iBimTJ6DJ/1iClZE9KSqyyUZ4WUrhBBDMeZRdkl+yRL/3HWryLi/5ObwXUg1
xmaMZ6Ttt02JTfaQg235Bvnc34lmESRmuea6OaDIVmHxwEZUfLg1SjjZEFnvgji1
hlysDDRSy9Tb+dPEVMt+mA6LTuZ7E5MeaZ7hFUg1sOTHjXCvc2pAF8e19QipIjfi
2vfP9EeUPpjrZ19yYdGQRB7PFyc1SkRQOA31Y3LR7BwRw8E6FVjtXEN3ffCTMH8Z
zuFsyiQTtEq8jqX+zzcjAfkZ3ogwvut9zBokWbZ+qwR2G4uI0F9pHDFqJOqmCOl9
5mc20vDxMg3E7tB2jBywgn9edNwYe9bZLJId4PS+3HZXlnKCsQSjvMgrE1cUHZxd
939DG2Ula6pa/HlKTojYSQfny0YdzG1AsQC+spOwOvQ9QcrHqJXnnOx5XQA8gJkQ
h1TnAO4YNN31aj8wY6PVdLVCXXj5+9O1T+h3/Le7tuZldcoteSjusgFU7anqq7sX
wTWCTtv0Lggk/Rm4SBPHmfQXXBOk5MMa7eH8xN9n63G7OhMTRBm/SDxLXYidmONy
QzxJZz4INNyXON5AEdlzIdSworDBSIy7+wCta1RcAffgN4Pk1jfndh66Zez5BM1f
ActFvDxjjeFHnzt3lFBsHQ==
`protect END_PROTECTED
