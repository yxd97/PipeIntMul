`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1A+yLWbUbrTErBe662zQqDW59Vk5AvgsQqwCGpc40b85Z4ggvRi3nscJWmSea0Jr
/Dhkm97suEK1rWb11nLe1ORKJYWk4wK5BSnfu5Aqz/NWqWLD7/jdqMcdeb7U6ZUp
kjUqV119uYH2UKX2h8ErN9XysOZHz9TYWZuFsb+q56FS5zO/OEcS+RPyS4dZbbWN
7YVbZtiqlWF3Tndevyg2kdNccWS4LP77StuORWqVasJqUozdRtLegWA9DeOnqfMB
lpB1O5EBJblvhQwVUBfCqAQVPoSivakUxpquoQEdvQKWgUKFbNH08jOohzhljhFp
SORpgO+cit/hyD16bah/ZpQoQ0IVVaoW1w9HXF9+pOFv61tKfw0LwMUsraiXQoLc
9Nw3g2k2Z6S7A08NyXqYGkj46ZDogradJ5e2/fY7NxCoagVuLSbtptwpl++AU3JZ
BdWVM20DAOQp5mRkBCU2p8WSpZQURjJjCIlpdFmJy+Z9VYsJRqp86jcaAmPa2Q3x
q5MJOomXLipxcDDPo8EWKyRWI264fDHhZBRDcEen0gHMuP0kD/QPqtAj7Wi5S7P+
Fw2hwJ8/Ev7AMfxVABvipg9GTFs4zxe9rmnyXzoX+FVVwvBxpo9SnCfuvKkZS/5a
Pti8zIANQc4sKhT7JJAILNq8hlwdb6ZTN3/sKVh4m4MShcKyAhAA2PbA4phcKsX3
+LOWkjCRkGGT0hZiO41b3lMVQTtpJJivIvb+o7as1+YZ0yKB6dnytGLPzMAAgWT+
U2j/W0s6yepgs52EFQkx8jc6ZW7dHL4Rw0KdjmqTl0z0FZ/+sM+TUfsEt84Fttzj
eVRNRD99xmWSiOPzcUwYyKBMdyG+1jZfVBropTjBQPYYJmUy2UcPdYCWnMA4FXKA
d+ykWPoWJEvjCOoBtyy782QSyKvvx1o4xJoef0tujn+OjrtNvElQrCJgiG3cLChl
eP9X+dq40ZFoQ3jqSWKX11k8FVQGVeUeizscow4MClZYtnSXO94DuEgyHbxxS04z
ZKz9MqH2ULjnvx9gsjEkxtfJl0gOE2S5ITR+XWiQYQXYgkueOvLPYVdPgFWCl/Wt
ryJ+pki577es44EEOuAyewMeQsQfQ6ChLK4sf2FnMtC7Vti8GPYkGkxrfFmjhxSk
QgryVl/ER0ZJhLcAM+A1ujcSvwXWZjy0nrHRgkM3ISvng+yrv1LtNejPEtbD5a0g
OqQrfVQLrmPN1ZTPNoEEAAHVa7g3UgDzENUaa2XKZZq2eifsbVZj6MVPI/9fw1UM
4a+dvq940n+aVXLSmc0AuTVT8rO5Z3kPlXqKV9uvUY19kg3HmZd63gkb5uNCro/W
EJCYJzQLFN87k3kZDGCF41FoBXvCLH5xjndHbj37ekHiJFgCM6DNC0ehX67jbUzN
iKzn95xHGKIr/O1HTjfa52u6VKY/knqp1tknzA+3cnLbiPkj5Jx1gwhyEXCPlP+/
u9DwKvvwZE+lFDemr1u/s9wzB39yt18YHGE+0xqnekzmCcj3N5JZxoQPUBm5LJp/
yf+yIR3j8UUM3bDePH4PU0DLpB9a0yAoNvfPYR+/k5EIvoJeyfXmtvSH9L22jnyR
JymsvkY+RdLrMCiusf8soBrDgfx2GnORjwNvbDHnhzl4+1IqaUVHdaGIYkVp+xg0
53SRGyVfxn0gG+U0weroEwVBKkE6kgc8fh+SyRXeHf8pjJoaVXMYwoIciJp0MT6C
CRXg6FEDa1/iEqG52OaH4MWhi4Tv1SNR5zITfTpU111T7stJOSmMrNSp8kQtkV47
YiOJykyQL6NOLPn0HYxNEO0eJXt/17BFeNeBx0PT4HSt6xulKGpgHWfq8S25TZME
WojgpLmvQoEEiQZWAgz+L2zhL7CJ+pUFtT2fJySEk4nEWiu4F7uBZk2ixRHszHRQ
zdkytpRlRfTkMgW8XCni47oMP53uLBDD3eiRxjFwjci73KBbdHkifY9/XecD8J++
TdIql+HmGhJeFw5zXXelK03KaVVdB6b8VZdE4QLiHDPjj/TaYBU5V6xxEwjotfoK
xFxa5I+PfhjycG3kiZvi2OQ+lec51SxpyeuuBxRpo8e6L7s8567cuWEJ9MgUOllj
0jxx2Wdls0bh2+2BPIwVvY+NRyukVR69G4P1P4ZKCFMdE9xrjH5twC7VBNNIl/Jo
wDWXSb6fb0A1zYKXTkPYBQ/NjqtK/3nKIvko27IvOBMR1SoivovlI5AVgkxZqBmW
xPdELwaqFDzHphPYNzzfADsQ7D74GmSykLWRN9SapPNKhv3uISOez3aeXKENJDC3
UkyoxwFsae8s410Vl3ugDt09IxRZ7rf/ce8ftyp8yq6sJUOJXBBuV8+I8v5rZzY/
47o5kpI/R2OHH+vlIn6pfVTJys9NjNp0hQHLrSgq1uLHMVVJOhk/d7XdFJBMt5c0
Yq0v+FLbqs7f/aBkbylvv+aDtOrYaM2WIuB1y18w9SZFhIT1BqPs4USvsOVphNSj
HLaw7zschSfv/9D1lphufxtYovNhpkn4N9mm9LwQp+DjXqddNbEVHnmY2k5fcSTB
dahx5zg0TTq/lSujqNV4qbrJUGJ3va7ti8Te5t5CUhfIC2zK8gSSWargTb+QhB62
noOlrC127RyOErcqMOM3d8Y4mliCXa28qwT1OMBO6m0ZJl4wcoRzqCnq+8JBAzS8
6P9LwcpMlAj7JMaIubwE8/Bs5OrYw7u9P7ez4zALNIyNldO4ZL7yzxvsDWSTN4lU
rm3Q/dzsZIOc9AKTJ4Ni/0TJisg+734ui9O3+0+K01LebGyODu3LMB51xknWIDJv
Fz87WyA3ow26PPhE806wDiXOQRitur5S5sL/OvHuk60=
`protect END_PROTECTED
