`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDsKVygm5OVUZuAOsM4o7OS8+lz4+DnZO+bRuBnF9bWzrq/aLlgcJKLQYxLvAmL8
QTsDC9/5IWAxtsXUlhDcJDKLlrppJqraJM41msM1h3xGu1SKFpkJCSd5ckWdaZDs
XHiSd0D0ObSYtN2hdovSd08WcyiZebdOmfFzVtNfxTGgxybfXxmk8X+K71h1dOak
d9omvta3aUyu3ij4cmkVLqvaTvWOh1/a4DHoPPGtidkKO0JRoAqXAGUGEWSFik9F
qhP1/MwEuesGz+Hi/hihTfh/uidwGlf2Iyy/WQTbb6E=
`protect END_PROTECTED
