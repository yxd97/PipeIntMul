`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7kHxS15+rCliaOdUz1VpGLP0iCMAYqAyFsL5BB7UGiDBfvjmUXTXE8c/WRbMJGM
tcHoto3ATS2v2zS9q+FvYpHhDiFa6oVZzefEnjEPixDA3Igh9vkVpgjdBi09TdVT
QovsKe6qoLDg2gjS9kqivBVhFlhe5PGDtmk/UZZSyC+6zRF4YotWQfUKHoipOxSm
OYfjC9QfbLIwhiUhWzerJJamOri8lYLYmagy1oYXX32/K5StpZmMV8wIorLDwfBV
fFuvFgpf/IhyJN3yzctpNNlhxb/0KuzwoZKg6IsyRUEnzRp+NnY8DwXEWYyWrh5p
7pL4D/hnh/eJSSaiiEVQlK8jXsfOGByefo44G181vmq9i9BrVEjCD7cJDe/aJrTp
MYZxCijm8thMlzj8kE/gSZaYsC7TnO1QF1fSTgNcM+I=
`protect END_PROTECTED
