`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TWhU+T46oHtqyDokwJDIhXc1Ov58zY+U82+4am/0kl1Ov97s63QLJBtfwkRqgl7N
7Nf9eo0Md9KCt8wHLAY3n/Mblel1Xx8sOJKMS0gZtY6ZmpY+C0dcj4tZZ5KZu7Ga
CQD7xj4GsJ5hUwzmt4ZLjqcupKVXb/4RAqMeDCVk/WbShlpnp/qHdBO5cFi7PdRX
ljWq9RKZkT7fRaj0WidVSGPDjEppdV9VxlHQGHAXNN8OdTXgMlM4DtCqpcaHAe3p
YJZMll/0L1AksPqQ6y4UZ9Dk+hWcox6m9XP0735t4xHRGpWjufKQsVbAjRbXD7F1
j/stdWhZqP0gyqxFMsE4wXyCW3rzZmHu3zNH7TH4OmreexPILaixT6GbUnTat9QE
xRpGcMBNBDNFWfiHMF8hDKV7d8YnoBJ9eKgb4LunYDS1I5YyAKXyJt6dEgrLAFil
fa01AuFdKUVZh1yMy9DM7390QGGcsRVqkc6o4x3wqBPM0uQ+dk2L6KglSeIlIsO8
F3KYCyBjDSqZcBvM3McvmpX5dx3KNXKTSmgyE+IkU1HOLpOYoT2hytXIq8rvTJUP
jmWAIr8khfWRQNr71jfmeu6nO0LdyD1PXfwmXhLcGKAj06UDdTb+ED347ETD0CLB
7Eh1MvP7RA25MBVZSghrHn/xxka2MGxN8pBC1uTLnXWiI1W6NyPo7ZrWUjsGzq6o
C+0qRNyd4r/nivZZV038JQlrJkEe7e7r5DvtbGlmeMYilpnH+yYo1CaERcDqNI8Q
4VEuQ3dyCySTGLT/XL4zkFIidu+naNtXKzgKAJdn79Cl0ith6ZVL66VGcQY/RcAX
HSBsUuvYx7+drQN/hJex8kx3eSGh5C7L40ZLgyJOBcL6MH6lCHCkxzg4A13MGgJr
BUvFhGE9SHsC5N1MbGmlzK2+RRM5N7c4iXQ8BmUjlyEjP58J5KL2iNiUoAhHtHNr
GfU2e4sg3hPpKUAouVzs+nUMkJf3SSmaDriV1TT2pUI0guSkVbmhSjvq9e16I5P9
9NuQchuWZdf5qnknp+zWV8d1YNFGaoNvftqQO7J42m0iF9gURdQfXnW1NGFtXiUu
lpbuCeQQm7owwKS9pZ4+HJ1q5p2ptGXQFYWR4gOnR2LNTFdZWEpe5Wet43qhWN/V
D+2GVeNS+VehjjvvxIImA8UaoCTIwpaj6T4KmTOBxPvs1aY/tDHp52Y+Ueeu25RC
9LMfR+Nz6oLkLdOl9F0ywJIX4Ulfq2KC72jEf8M3m/qDkPQRY10Y4pFQLusKZszk
uQInp/iMYV44t1ykJWRh1/hJ6AN1pmAdlejaMo624AcZK/6eZwyGIoH+NR7bMHxM
rzHjVgxwVwxG1q6tHcxkDm9lU/IY+Bv9ZcO18tPIDQY0wp2u4BYHbcXNtlraufsf
zqrL8Jo/txz9Pk6r3EO1Sl+rj/BDx0JlXWWvUfpEuHnDVwfxoWAup4sEj/tt5iwC
fld22uzszWrD/E3hLiZkvDxNook2/tBmNz1GMWCLTncHtFZBcQHWn/QB1fHFBCHu
C8h//LKyIMJ9BU0tuquopIiN9sKLQNCuhY6bFHxkHzoAyV8iyADJSuN1XMYa9xZr
d6U897OLBVmf3SDm6SD8xVeBkJwcoLu4GT2fKAaxmoHXdpofgKqVb1CzG/7ml+I7
XdqVseWJ4lEAh+HQK/e+2GlMBu4yibyv7NW7E8ECWnbVo/u0QVSdd0dntmAed6zJ
NAw1GAffIAWutI/KmuARCk9/iiUysB3oXeMN7j2TcIzn5DtlWVpzGSICGcAOubai
M2NjsAONsLz7rV+FCZzFg+abP7nWzd3Cd3jdrDrxG6rh/vC4SoWny4WwzD2DD9TG
w/GsRNQ8c+xbuG1JVeQO+H7qaIZGVynEBAOpc/G96l7qUh/uKGv2zKXKKHHw80r5
NQ0u5QgahXKNK2LBwWIdanOuOsqRgpIEP6LQqKHez3Ti5ZTaA5ZVTWj0/7quXpdV
7183Q9ODsV4Wgp8RWCCvinTM00slQt3m+HEusYml4WJIepoTn3G/UH4DI6P82Gd6
M8hCRh739E/bQJjvqV3bl4WLlbsttXuzhUgBI0ax7lCncgiNy4H3905r5koS/4uN
VsfZE9xw6yW/+vJK1viFNOQSORoiTZ5wLupsXScp+CBrTUA04OKxjEC61bTB1RO1
YIvLGFukERe5u5lqshcJs5YCWor5ggWZgjBgzcYIQ12o9/axjyLQ/DKF6IVi/Ghj
9KwM04hwydNXNA9kDXqkGgShNKCuSd2RpvfShMq9jvtUzPEa78H46FW2tqQAQ3Ur
NoygBs64gDgNYyjLP83iTbK0UbckkrQ43pJpq4CY4Dy9eOOeJlWTPNfOkzyn2Uxs
xG7cmXAGQzsVRBjkIzRYBw==
`protect END_PROTECTED
