`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBZgrsRLNPuMkN1qhLACn+/RELMC37MYGEREub8IPh96H72+pymZ5fRHNhWBcSlW
iqac+IOydlEJ68ZbuoDFKnaI+rRHyHD6qNZ7XAMqAn/JglqhjWahEEqO55zBEotI
v9agPDtwpY7a0R/oyUcKMk3kgYvOTM37l/PMBhGMqJE89kI9k0C6kkcr6e6tPk4D
dc67k1khgXe19fQjkEeawxjDZ0sKkPwavxLFrJPwRKJePGF+cfHyypf3YsT8eTly
na5W7ccXW+64KjYSJrzk54fnPPvoDeQhX0K1v5/rL657vu3p3etE7X3WDYq9V5Yx
YsOkhcZ4gWx8duwtpk1YaIRE2O0MjgwRUPU1psKAtwofQ0su/EevqPnCuXAdm2w2
Q7MaE1tW/AKXF5aOiq6H82mZU32sqBHN8QQunnvVw+GDsS+Gd5n+U4EMBxVwGB0K
`protect END_PROTECTED
