`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p/8RgCh/cawo1Kaa72In+boLif3sGtG/FRZbl6/b/YJIxKZJMt5dnCEpZ7shNNUO
anWv/XQr+gkXmaNCb5zUaZ5qmXRBlUr1we8pIW8EIddOK9eZS89/g4W3CsukHOnH
rgTqezbEUTpfCgJDoRtMXowQS7x1zeJBJQq1F+B/IWmDP+rzfNHj+UslbY9hhme5
mZJ91uByRW/g1tn64cUsiE+gRBB5fEUQbVZPFHYr38A4kOSESJO2f5jergkucup9
8SCUVI+HJ38AYB1r+Y5wbkJR/2kYAenGExJESHlibg/pZ6WY/AMY8jiXlFBfDDDH
gHdU6rlC7Mx6D6IShSTp3WRHpT00BAGCFlzmFxHD65K2oZR5T5CxV+PnNeQsAZ/b
a1+uVSqcCCdnsjb2QYu14+kkL3iD8Nlky865H7pkwiMWHAQ2dorS/sqQ7wIE64Wi
ilOT0kPWSCKNWOUiLRy7oKUGohRNNgy0gErbUzecGk4m4Dpz527DDHSbsRyEdSfZ
V7TcIlqiUNLHNBhPP1/bPh8m7RD3UGRIwRGx08VpE4CmzqzzMsrmNzmM2/BHmpHM
/fVKsFb2Sbox+7A2UKTy1yK4T6/SsZ9DFZnyLA9TEkL3RdpdBR9IE8ssKgGw0fPh
77fj6a2TCSI/tNSbDrmQoPuh67ShpzIBUKrBnBy9zRaaaReuC7F++WUkbJTNLhai
VKScsEKDLDEUZkWZ9oPsid87HxqbfngeJvxf30v5kCoYPqXYLlmNePL6VEUV0wyJ
4CJ6FMM0Vw3FWOJCXVRrxqS3M7puFlrR+lREQx+hNAR2BzszxrvsdGtJeM5PX8z1
1iWgkcS+ivlPzru91UxkPrpmGWGxmUvtxGt5DBbp9EE=
`protect END_PROTECTED
