`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fO7/wxWscBid7kW/3N8nKM+zAGRqn/G7WAp3vVHL8Wdg6gsuZhBespU6XLypfn8C
plG6ljRPfE+MhVG0CFmcNavRylLKiMVF+M5yi98GNDwQSf5FOdstOpXndyL7tUPO
eGd5AW+j1EeD0WbJUcyqW5UKFfHNLX+Ix+rjaF9OhcNX8xvPWrnsksGhV+uz35zl
ayD4s9u7KIeUSkbTVrRpLgl8AmcYvRO/bc2KbMvGP+k3mTzIFTp7xS5ldv9BI0hP
B3O0Jl/vD2ft5jB2OCJRXob16MqfQ/aJRHws5tYObn+WT0JCPvppR9J179PzlXHC
bj9YLBEHLF7EEGWxnVzoyJ4O7Fd8hD2kR0k8lvl0HY1FNXbQBVBEqesHtLPk2v2Y
RJw9I0M/lcGQBLctXHE02lEi+bay6yRGlBuwlf9cFQ5g9se7U7cZI0MzSH5eg/DT
ONY8Fn9N3Edy6Lnno8oF4aqjSZiYS204o6P3KK/LHrEUSLJkb/FhDSyejUi40g9a
bncXvgyu3lkyNk34IooUhKxhviRZ0YRG/efRgfgR3LxJ6eGGRc413layomxTzdxu
UrCJrRU2zdr4cW0ucVOMdwA3/h4EqTYyWqllg/1NlI2cFME/C0JS1gq3Gnvvdfqx
sojpZJ9Oi7DY3M2Mx529zv3DaoTPXb/U2SGD+M5+mokhdbJybGIg3xBlxie4R7Hi
jSleQyzCiZm5bBAilgDkjaEf/LDyGkC1zwC4SffC7TcdLuOOamqQ4Yb+NSdLq7K0
TsSjcTZvxGpr8wr2tIcO1pb2NasklTyQcwpoxHjyUpj6crTlrmHd5rlu7uOpS5fO
szHD9WHHo5ArcSpi2tdxc3E0Py6hKxPRZsYnnM2C/1at0OUkjWzthGvOq6FcTngZ
isa8MZFWLR22n5CkYl51GGZkAL05ptcuH1nJ5brn20x2bdZ9dCZFW9da2hFGlOUx
coWma34YV5NUB+g4JU2y6w0LQBANUChGiZxulv+wItyNslyc4HZ/TKV5gqJzwozy
yi/0BdvBAMSJqC3uatXVGFgqkcCV8JBNzlK5T/MdYh13duvHECtIxol+ZZ265jie
zmq4ugAKLRlOWYTzuWAtWUpeLBQrnl4w8US7ZkMark2tgFFCQ7KAdDq8CrY7Urdd
HKdxtZZMcFLHtvu+xyhJUm+px8WmpxFIaU8PFoEGZsCUvZ1xm4SR0ukTlJEejegT
bejMhg+FeIjlhAfFnx1lgGZc7V/aY+kUQwuQcCjIlkIxVp5w1StDRjrTdQq4ITM+
g46kZyteKGqOO+5jQ2y1hAPEjo7XTqQPyaC77D0i8CzLx6VnkrcuhcGdnr0FH+lT
MqmJ/Y/0yx46OB4eUHvo+qmuGtzHSlfwch4FrZYbiZYzG0k62FT2OLHlcBo7WEYx
V9g3Uh6rRVdBu8gN4fzmHPcIIHFYyzu3duSDHx49ZMovccoy8ceVOzKg+4w/mn3K
N11z0GIOM7nq6qBwJ55aqCEemzR0C4EgDFI889e45cpM90QSH40cfoOu/nl8C/1y
2FtP/DTrMGGOPr6UFtboHVtnoOiQ7sSd617dJoPmpZM1uHxlI6s/R7OvBw4UOraT
fHN4e3hCaOMWrI3/e8AzC3owaDDYnE9wOwdC/5ixHssNRHmiM/0SYqtyale1Kb8v
kEg1nd4NtM59joE2cSZ22zV0KdQOqvapgEDG83WudSZGkFzj2iVH2eDr7smV35LU
qymRxKrPEdk0nFsSzmLoUjfBfcLMR0BBLIV8q8ZrOrXY9tjCqe0IQdOSjW1YlXKj
EaAy+ybh6XdXBUBDICoyltTOK1rRwPsG7P5eS4zoP+YlUAPtvON5ppXCgQaDw0MP
+fbsF+e8LSZIqLvOIkYaW62+tAhsqC1LMvRBY5LqeLD6KAYBh0SlrlbsbbC0SXkQ
qwHtIzKCh2FWuG+/t7UvPZYAhrWcRolt9YD5UvhxS7F/dde6aISpHkFL0Ex9iDEu
LnENCGWxd/ffXPeMSUaad0YylLjDuQVyCS9rFRThX80CQwjwx3wK0JhnQ+ZISt4d
JW+sxiu4v0RnLOFTt11GCwkUO7vMfjMiQe6l+QHfYEOIzaVTG+C7sMV1tgPtICnS
35Bms2kquIkxBbp//SOBX6UQuJ0TelHwNpa2bvxiqXo6LNUMfDzhY5uXt8dzWCsd
R96cpcOUux77mGAXhtVR1C0BTsa1FUnMEwudID7AoaCkRhCX4Ms2jdNMcjftPvSU
nm2hAQmHFHEu6Zu+bZhzHLarNf6sM0z2T/5YH+UQCfRvoRQFhFoR7Um4bC2ufx6q
zvNNG76BrTbv+ZJw78wy5hRMYXaoKETPXCbN1xUJRzHVeVwjoSwnZby9bRvlmyF3
lkJ9EWATycPt/LEX/df5CfDCgW8iqlagW78f97PVrEAi/r1ZJ24udHi/OIVqD74v
rnbXihMPTJwUPjvk9Q8xYWcl8BnojQ7F6BUs5XdxWmFzAikEAqb54G3MKBJHsjmb
YNPIdjFrXD76XFl7qT/K9u3fnbLLr+Lm9qZdudGnFSrZ//CHWT4MYRvyxEMPwTgv
CMpdvTmBLeJcSFQqRXaEbopNQSqi+SSMaY7Mw+08jhgbnEBwu426iuEbdK7Lswei
n7k/+61ruJE9jYqTqXmESenHBYuh0JX4ywwvdjJh9NRB90UHZ0WNjbyFovaE4jeD
UEM3czOdHr1Ln7gmOXucukhClr0Ohi828HdEz3Y32YF5O0VzUPbJp84p9n9nZIJY
/vKPoZrcNEA4eybrN05WIbNfsWPihiEe3ArMoQqicIh80aqgzbZN0q4gb7RrbYbR
9v4BUpHPbw6QY4TeqaYx946qoGEdvDNqIvIlVKWnwdOqAi7SP/t8klWX313k7Pl3
uGaN68RY60QHUcZbPkjF1GRiihOPTCENJnXbVZbLhBBzK4UOfaFyRrrenBrIyHgd
HI1Gj0QrSaw9WuWSppmnsmTm0pXvr4FtwZYALtjq+aLEqjRsRZ7j337ILfnk4+oL
63z1gvAPlvj8OH5dNRnyKfI/LSm7NAlUxh0MdtGNfXGEn7ZuUqsjwc12oyY8xbHX
PcLSfCWWnXrxeclKY+dh02VSg4oiAJTb0X0cZPr0hyzvVXOJ8EEP//jQpkdUt5L9
oBxybLlUEo1cF11bL31bIx4+so1rLdMvmYQWCFXLJbb/fsDQmX0tcx/XzDoLapFR
1PGJm6DeZeuve5UmZ1lLhwCtZE8MRNMPzLSV1B6P5Bq555NR0T61ZfLVJ7Zt0xH1
bqdlYNVV3Dw5H+zIdUMBPPF1hAtg3QdP/0Lw8WEGs6Gz7fi0hI63ObxQolX5GW7r
i/BRu8LtcyOdEnf9uBtrNEhK6oxuMHe7RPmbsNi9INqmzXzw0c+RTQM58ED0lhzs
koXF9VGZ7bsMM46EA19SQrVIUGbZ9VYI1PqHcXorm/lxET0KEMsBuz2HFr8NCRMI
P3Q6YxFMqV1Po2IM/ozIXEd/0nbNXalPN5SVlq/OyHQlyy6WDhGS1HS3l05orHOf
KA+FbZvcSSXSV/bmcBdFO8MwynKnzxz9q8tYPjmrC7FfiYrBQuCAn+pqYIxxGZt8
7OTOIvGCqXaaCOr1vYWlA1iubf5/g4UztK1SD0hSrv6AsRsAkxmQ6vrYPfv/mto/
8hXCAW3biyUkqAh8fluz6YrkhrJvxrz2RNJrtGa6t1F0i1H05usvttcPL707w+0k
1x1yLsvi3fAURd3tJj31bA2XH5vxrEPiG3tHROnOSshBRnpDEtEA5vqscAkNV4Vp
Rv7CotlytWtP43yX4Y028w3kKHsucRs56LvA7AaQsZ7h/xwL/Dz+tO9N2bGtUOn8
PVc5tY2qnvv3riqEWPdOzIbjNQGnO4OJJBIfhkNoXye1FJ59U74hW/sVtPYSnjc/
D31W5pyTlKVkKRMDXunIJKDGcciTnQYCAIyANfUcHl2H3VeSsX99Tly+hoDZ4r/+
fA+FhSHk5dkHL3nj2YStCsRp6a3cE6oN0Hf87EopS4sU5jq+3m6lTtzxQ1+7+Ch1
c3iId07ADglPLAlMxftNQrW7YTdbDoG21eWZolsUxgRQ4gs3wP+TqWxoRXfs4iSU
trUXOiIT/BT2ZwR/jPMvXWh5C0giKEmpxteikXbGHej1eNYjfRKUyXC7uvFvpS4j
P9yxtlrcysjPMxnmZDjarP1EFd+yzEOa747daQ1pSdIIWRWErtfCM7Kwpy6TCkDt
3evACl4qvLe9Vi6KPKnyxQqCJy0u5nDOLn95c0hPoewzNFp32/yaRD29PwJwbHtH
1+6PKHuvFk78eTiZrUEhxA9jmjUmBochfQOrFW0Ks4fajNoG5Fmxt6XtnkKHcM1v
9f8XvHLpku6XRIx6Z/kW7WmaZ6iow/1b9xuQhnAex9kibSXGg5mcqctIqHNl1y/L
ee5x9jwbzFJfKLoJsqAtlSiHjypYa7+1aT2//dNRoi+ynIw7Cz5vpPDMs8zo7WIZ
SvoyLEgOJSGehlLOxiL4/D68d28pkjvKwF27fzLD+X87seda61vJPdTBPO89l3/E
2dfnNfQcN38T/WNjHE4wC6hgD647VvK5Lr8Wb7J2KLawwsnNeBy9K7y5lwYOBFUc
wS9WmLh2gpbIjAhwd5jc+SwcERZir+0RKoL+p3ZRYUxzYn8uSkTvx4mc/GzmVmgW
9D3b6SeK30Kk++Z7lBg2/nE7sg+q+F61zSM2FQ0EHpu140pVCCpjqXv46/qOoih7
eFNqtPxxcQXFU3BxyosYUaEG6mMEHN+ahr+J9pHmiOTFhkyJzJtzgZ7BtnBZ3OFx
IKNzImhMUk6MxDVn0qdET1MNvOJ7mcA+U+CEI3Ck5FvtcrFYsnLEcBNlesnInqgN
twXMyLy51FisZ1+Nt++oMtf6iayhg7QJH4N7bCCTsz/P0rFv9IYn+7NRmj1BcTDr
CHXAOwZ9vCLuX715s6A7ria5dyivlk2r1sX3S9anIy/HRafMo4vgdmU1pzoPTISW
J/Jj/zGp+pYkTwYByRout7Ad8mcsdytojNczbmqrZ27LEHsym8xYQnYP0FUNp16M
BcJSX2DqxIHb8IZ2FkKLsk3a7m5OOR8kFIvJz7W2KAaXsimZQsw1YxAb2qnOJMVr
YX343pw+8QPNBM+ZqnHFoW4c7l52YR1+5YVu5G5pUVbPWAVr1BkduK3bxlSODoE0
DizJnd/3IZ9G+jwJ9DY1UStJodzFWAdb8UUbHAD0RBBzxhh5p6OoC87C0xGXMUbT
nH414HiVVjO209TOC5cE34pfWnnAfG7bLJo1uJskclVKNsRZlNPZ5ceoylUfpP8q
aXGi7FOiBYiFrBHA9pit2AJokfNUE52IlAyToAjJAm92lEoxUDurSrGYx95M5+X1
/cdRQLznpvtpHI7wpjK40e1iikX+34k6Jsr6OxspgM2MA9v3Gu/+8Ki2cTd3MFxe
pEWk/uzaaTDhwo0LSqEFtGBZ82FFeBJaRRuQkxiawXeKY1ox1FhxQ1oBio23kwcf
d6KNd4HUBgeri7M7D7Ykb2MQs4MgVF2P+jR47zU79Qu5ly3656+ixTy/o8oDitH+
OyQVYZgdgtYmQQkAzv59PzcNrbJGqzNi1fOpwGyyFgUCByXxnak6sVXpIy3odJjf
3a9kioFYtFQn0NE2Q8EQpelVcFAHQLq7FCP/yNCh3gXff2Rg9I5s+rlT/WDUBmm2
GH5lWL/w/AWAMVsX2deJsRIkOuqCT++dR4hvQY8TWR89TW7eM9Wp1WJ1eNhCno1B
4h5U1ykGKE3q+pNKR7u5Xse2dFFliw1ly6cTxA+wAE/FJlWWJ1Mfpkyx5lsQdlp5
5+ca5OgfEX2hcDR7Wo2hiwjJy9S0A5C9IwJ08w6ZrZkKvHr335rJ3bZZLKUBSWGK
XIGSUp4QcsGZpUYUdMELJ9tJr7IGZIGcYUDViz//NaWa+pFS3Ku6osS9aECR4SWr
URV0gB50sNpXGSEIUniFKhgqapBrU4abOQWj0roavkRKgbQ8L6Rj6N5sZ+cAV+su
iLesm9N9SDe9S+ASma5hYQl+XLB5P+booBnFccw5UbZXBvu+aUYGUVgSAb6lNuOA
qcKvXiibbYkfYvzv7WbEC1Dh50+eIIr1mMuFKVLIUxcPQ9DHRzlW8xYZD50Gcswy
IJzLaMwoTXq60VvroYYBJ8rZwX3sn+3gbq35v91S8yC6wWSIolKA24/NlFu8hxTe
75I9lpjM0j8KqbZUFUg1z1NJcO0+g9gNgtDhSm63maanYVnFOupl57jXF0MId/gd
0UhFJNEPnzQa3JoCv2NfcHi6TCW5Gv8J1EjIFWLvpIMNDhbcT3+TSiRCwoT+rJUv
e3AmiP23rd9utYMw1DTCQHtH+GAWbcPTwkRkb4xhnZtqHAe8JT/o24n04fAkVML0
Gki1NEoEz0fD3GYPtmLq7C51xzehdgAm5wCSBEgYecKTw1htwFKdl7S0CUNEAvTi
m6ceo4Iox6X99XuuFrISa0+W9mZSu6UaAX+dRzsH1iMu0XH8Xzse20Qs1APAFms8
qOmmrJBKp0Vt6vMvfocSC5H0ZpB6LYKzHoQD5h1sV+/T1OA3IpHgd2isubaQKBar
6sdXR2T8h22OHgZ+RvJ+rkmf84yhAe9jWaxCArR2kPH/MkgfytWc63GQKmgFM/Kq
JThkGX0hwziByh/n/5tK0PYJw2d04FL6UMXVHHDPnBASSCXCUyD5nN/vWKRCdmOr
G3joeen77thVmcPh8cCHWHJKgXHpxXbD6zNIv6NHdT1nnWtIswnNjLuSSxSJj24Z
xeRRUHSlgC+muwyAqxXiVJyJEKlXZeV51mpvlcE/IqhM5ZpsZKoQKxWkqK0Kc39S
wxbaoxBM96YbXDqo83+NuAzeGLHpB8dQmmkhrfg+l2tWMhpHx5fwAbt8Mqp8ZesM
6HKlIGEekZStAQ0K0rPeFAolu3KtS97KPpI+OjBv+Ppg3JelAYR4zH8uI7qCgotO
FeiDlwjeR8PP3V5vT7HlEKld2rzqmfyca3vOJ2eLG/tTKYESoIgbCYNV/v4q6Hoy
L1hEoXTX6W3wqdxfzaXBbi93mjGLx8nPugQFtMCnG4bGjDXCFqc+PJE6gaHn5mzM
567n/0xX5pe2pXn82GpNFkiKz3FOXP0W/U8zgYkaQIo5rDxy6fj64myEAZmZ2GW1
1/A7QJ8h4qSXUhvC//VN1hwyTG6qLu0tXTiqcbb1KROaMVh+RH4f6rFBfKk8JHGA
mnPUujNgkxQuVGu3vJzfemt2ftNIZV7t8QvpJg3MjDR4f6tNMNRGf0jZyxWGcytw
ouJot1ZYMXcAXphxGHN4ix3Yv3IlCTJU6hGiZSn3/lrPGkkHOEy5EWj+TkBIX0p2
gnXpw8pM/+VaasVypUJ6Na1hWSLS39czPSrYYDokLe1WJvjzr1dghZ1RLHLBxYm0
eFmZF8cgxAKepFzr9hcVDF+1+BUeDJeIENvlYD/vmf97Iqlk+QAAFIq7AzvV8of0
6bN6ONyUnagphcmSwLlscyh0aUN+AJCV3QbbaD+rRPddkAS9xSlzZU2Lr5QPw4Jc
kln4UDKoMmpvleOj8NAzdZToYivwTd0HILZU6VjOfkt5KiJzyFXeuKly8DUYY5F9
XfrvSm2vhVYy+CzslfqvoJMUaivkJxpYDerCOXPngi7boidiR/QUesVHfpKIykLk
3jYQ+kp0ooUYMuRRIRckTDSVGUQhuKZfzLS+URrUFdOxPqyPIQjduVQN4Puv0hCf
L3rIwj/uLzDInglmhXjYvwHirIRC7Yg7W4qjKeljEHeD2x/Mr3dJ/S226SVcrZUq
bmY3UFIWOUXnwM1+jp+orTvWLXw80tj/VXps7XNYJkd0bvwwCNka8xsrGx5yK0Ie
MpBv/tpQbBBhyBxfQivo/qzd91lZS1oNhSoNAZBmq2lWqbyu/vkVkdiosfmW+KUY
kDvYgskS7gDMvZQqCpmKaTazTMIiQfxYdl0ue4zOGQ457JfihGXoxh+OKQOciJk6
sbri2SLUxpqsrRLwHJQ1+F+qd5CpA1969YG0f8umtYZNZLmZn7BjMEbYzGP+aSGj
R/rvgb8Atj06Iwi0JYFUAKEiPn3xE7/g41BahW8uyl/MLNmkzScL9WTJgNuW+qep
18Pk9VGNtN5esJPU/5yn/w6I8a1nKxGfEYm+vqWXf8g0iANzThr8lPFdi0xI39qU
CQ31ob1mR6CU94+GEosvTfBlwOXUZS9KA83O6D3xqr/ec+d5ok7o/168ypuKWU49
CMx8mMTUvKNKjEAtCjXLa4swb8Od7B2/+MuQkFPBgY2Q6TCHfNNVRjHjASoMYCWY
QZ/YIFKoqKdx/axRxen/fDYS/QCq9SNYNy1keIsynmfLelkiCLD3NxprV9XURWum
XBTYyjhNI3K/dm/3DgcK7i2da33hUw6b6IciYChUdwnohf9VADAPpdArqS6QO288
5yPjbfT3CXpWWlM2mztK4g7LlfO5yC9i4XnXdz8ZsKHZ8Z2+kn9wVCnlrbmqaBwL
oZFuBgxJcIwzckRlbUMvAUrePICvd/PL4K1XRJwor1PBDNUQ+ZlVm32IljsfXLh8
2AEsD/xSV5oeN1aUqKceXQ1N3d9apUr/ZXJlocOt60dvk+nIvSJv61o0exVHBMRg
z6EmDrDmJzHUpUC7bBnDZ5Kny4RObnTxy4c2arxEx8m4VTMuxBdua5ZTedWnaWkG
IRblU6Rx0/4DdY+43hyUz9ip29yYeBxMsoI5OKcMPwpzw+r6O9IY/PaDSuBPUGyz
IRoZNY5z+DE6tyfYycEqalzmkCKI4fm3mpF3A3wSfwJiOWltSZEFxXN5GBek4Nxx
Q0DrinZz8KkKtnTYiP2cXFZmETdAqMYfZC8HSd/aVOiYgjCJDcDXriTnLrT0QLVA
Q1meVkK6uz2F6UORwhoslMAyxmQPPHIbDR7j4BijOxiZJViTcAB3iHQfhsK3DGEJ
uzKZ63TG09C8GeuvwFO0GXx1vmgDOm0m/QYSI/swvyphJ5RRESkfOMDJLIW1Os60
rIeJMG0/LlAA7fGo6zxil5uc4i+Ywg6QVDatm1hwcDjO1YbYxS6mJtA9kKna5yqa
e+VLmhFTLzj35tL93uVU5x+9/9nnJYGfMhEPrV8f+oR2fRN4Cj6GgMel0G/c48cH
d+dDZNwF9qPg7mvC+1NNuHq+7d6P8M12KfqW8Whh0wO0CAbYgvHeccqG96UoeF9Z
/4gEbo9IiflkvE0Xh8Ob2Q/F1sdS7hxs0DgDr88+VfOR4ta1ltfxvq3v61yVnGbH
zSSZjkfAWXYsrkhEGJfW6OXToFIIcDr4TeA3Yxyaem/fCFhGAiVpJp9+H5DgO6nP
jQFS37m8WhgxWLqvD7XG5PS8nekop0gEDNF5ucU66UY7GIs1Zp5O7UxeMATAPHdy
W4OSTeWf3mq+ZivBOVmhLs88B1inri6nPJYTMh1NxxWulEAT8W5dEDlPdi/yp5P+
bRUUFSz2+uxtf3U27j0KGVROfzcwQPl/UAI3N85Y1VAw1mP+nWIlbf91TAN1+Ril
sgU8qTPEFh2h4ewBS+g4yeTBTPGCHU8XMNQU4QHldtwKHJsuYh9Qej03Jyrvfwus
CwCIixcwmN3D4sfw+FWKPFJSzeZylFkRZavXodxbPf48eNjo6EY9DY1kFAh/j/uP
iZgw/LQAkelQB6fEV5MzYoLNR7vUvyNi9C/BzBe1sQ1NsOpeKLhJ2JyMTGlCaoay
aJfKlvQS+2cEX2bPb0Z494QoVvcI3YiPtl3WeA/cClKiRlP0wrMVr0L9L5cvFxz/
bePVF9tsepcOnvS2miOIY39wAV4l6LQlapxvkVJQIZmvxm2rg6UdBUkMEkmzlH3C
ZrVgxdyoHebIwWeR+zGrVJOdoWDWifnXmMUdb+kTo2IaBfq90t0HGPrAgwVVTJe3
Fg3L4nP+XFUncEzwcN2AU797ACz574OUIpQXPQrpLj/rKkEFCUzjTRiRSfh8bgNx
MEylF6yxi/v4jUSw9G/hnrhK//j9bt4sdtr9zr0zKK3RWYhhVSN2VE3erXkPleeH
9MrTTlkRfCiwSMzYmoeXQjtYqmXd+WIFI61IOP+6KXncW+mktIxESbPQs41K/Sui
7BW2j1wacxKdQZeDI58oDaJcaaeRD6a+IcxuEFRfJ/baqTsm/zgXmgpLZQ6Nenij
M4GdW++hEcpqmdWbqzpom/evZg70YC+MYZpB5nLrKvRdpWq5srC/WLlRCz0cmq7o
af4FbhTeCwiraO5hgqAAuakCD85+pV9eblsc4LkrPa9yh9u+Wj2Dfh/ZT0ipzKoq
9cleG7uXdhuEzPwsPtr7Hz383PGOCO1rOd2EIH9tkQTArFEQC3qItOxyKvnjQawX
p+tDXPCU9FPBuKaqOz/CV9ZFvCDCFqW3gvfCKj7HCw5tviXAwLCMBJLctap0374w
6qU2ah+pdvL7i3FJt7FOQxoHGi+gnEI7w9W5C+8gAuuRPX1n6ipXy4Zpozs2GN6j
5gj8wUosc7oOuCVdu74D5U3Pzig4wQmaCgDaJOT3VSRSgpTD+1RlFYQnttNSH3Db
Qr+y/D20NkCd1/48aV0N5OgWVKzD4h/IE96Gj3Yf+NFyhRiThHlLLF0mac4UMcPO
JMajlhUURADIKTGkkre79Gkg5B/kOjs9EiqNN1VZVHiwf5/HatdzXabSmPHVZXgi
DSZ0hcEqgHhsmdyQJbcbaGKjq3jHdMfb88RAjuz347Vo2b7M784eWIzubwPlqVgU
MEpwmv5f/ldueE9MQpMi2ktZVufjSBQsVn3diPJdzyvbG9dY/P8HcJhiOkV5PjWD
h7xfBvv7kgN76D9GEv/p0VC4P45pM7cBOZqdRXp+8dXKEHPza5NXBoAIYVmRZOlz
5bnPmKg95zY/L9QxplmUafiOP/4g2riNv4geIsZZxLQ3XAwoh/cb5Lxyg6t6ghyB
xs93LJvaH4PxUjea1CBlsT5h430txLiQP18D7Ojf01r7s9YbEKkKqfSJYKy3OmFf
EyV4GXqLkwhW81UG+tyMEuLJ4Zw+8PAHMg2PluycfQw9czfXBYqLwlygPfXv5A2M
8uqHnmZ8MJDRZNV/hnaXoWzReXsy3TwmMPYv4r/8/wngvAjhUa6/tMdDCZBe/5uU
3HhjBynf5atZiVQCovri65/QprAN/BxFWUJJNPIwhTz8QqzuCGq9VyHgTmGpv+N2
xU203Q76NiJ7c5/jUWcuyGwEdRYcFy/NCPFbWqp03gGkhn0w3goosh6VBIcYJL1h
n7UqsLgAE9WBfd4OWdw28whtAaKEdk9/+bfSZn43a8UhbS9q8g9OHIAQdEAfXnbM
TrlGdBKjBOSzKqOOuQpchISDTNy+eqYWQPMHfgIGeZE+EaJ6g1UiNrXqWbrnRJxD
+sBN1pTwPQaKMpv5myazCvtXFv2WQxoMNvMD23i4IY9AZIjH1nMVpVvog1s3PkB0
KA0aNuqEPGYwmnS37EKcZdZoYTrxOlvUOp/e+Qmvh8Nr1GGl55Xn858xcuS60FXr
v2aqJxUtBr7IJPhoEfoZzHsMmiq6LulgV9X97OnMXyEX6MdVa23CsnTIP7prLRUh
57MUw+973SwfFV488ryGmKrfD9rMYqDPgiV9OyDsCnpY3LkrREqp0qX+pK+qKZAQ
U9CdDq/srrFpKzYwxHREV9YHp9u00wZzS8PD+zs+Db8NHq+KhJsonQjqZTZIH5+S
6w408Yu1w+tF+Eg/XPLUyqTQryCJPFhh+ILWIa1TX+2KYlXKKHcHzVU7BFcs0CDk
762mZsji57O6zd6SufWAtOMohaxL9c6A1Jt8/Yh51R6/L/hU8oyroaQFJxT2CGk/
msqPHFq3ytdUBd2hsQtHwuOXJtsj4qR2tg3ekRR6zNizWGsfppsFdOmEpX6IgyJJ
WYAtk4dH6kD6j6DNMKutiWPkxg6Ws8li44MiUNz9W/B7EJQlFXMRIm4CYqvoOG91
/rQaaBidnoCyRXRpwRzKTE7Mkq2Ohtm15lW3AF+MATYhwJ/pjuDxD0wawVubOBLl
jBtQEeiac3NwNb2T5Kavc/pcJGLnOMoWzbewuYHRS3RRlJai374k8AmxAWtnhGOh
/FBAzKhJreMFD7Td4k/PMMuTA6JcR+dmC33B5CG8kOtrjdTvE4TFqHzv4lLD3Dja
ohfCmckN9dm235vnR++M7TMYjKt2ycvQAYJYB78bxfGd2vPnVWcdQUC9/qzvFTn2
b1XKE0i7XXqk5p6gtwJMUHGUHTbv4Ek9+5WvCFt/zX3jrB40HQyR/4i8lV7OOiRK
CrUf7u3YHeqiOZLDHYcVOBZUnRsEN8S2BxhVrid1yvJcaR66TnAVrunrhKDv/6NG
Ukw7p/EctTmfNR82PAmXtTvSPk1Z8+O1T4Fo8fG0Q2e0JV4ty9ognKoRag9kKref
18oy4rFU0IUHalcfbATmSZ62lNZzADdwzSIQE7akpid2ip3hMWGJPAWxZPlIR0rD
HO8cHr6a8fw29c92RfrgXupejJoj1yYLxZwWjV1z1tZzWFU+xAnN7wNQpTB2US3D
2Gk7KKegQlCp63w35vOmtMh5iIWejctn0BVaSpXzhE12bVtsFzS/gVT2wGeQR+OA
cNM4xOT4AFYA6BY9IHTWQ58jQArVALQnpEJI0+Cvj2CMnqg2JRD+gsz7mu/CL/jE
NGZuPezoHNjR1a5zQUTbKcfOGmUJSHkLWrTLzWSUIe7sl7/M+jZF47BqAA0jpr/d
59pdRAWYhbWLxqKypd1/aDNVWPtVqUs6oLW+4B5nYZaKmEICTx7G5e6CquRW5PfS
5jPSRw3eofVhC8CfIILxM2dVAK0Jn1WDRADbbkhBmhpjgTn9DpM5hH9lmyHnkA3O
kDIC/ZImI+zfRScwGo4Szg5b0aZYgtjj2mQ8XXLlFxIQIeKtS6bzCbzxqHXfTjNX
X2+Gd0sMa63bcCqoKQSb4235a9M5cz+my7xsi5yU2OubSg3WfNJUwcNjWTUyXwXp
GkkprYHD+HSUo16oW58cRvQvLBUFpnChkYZS1GLXX5+Vu7Szoxrq5NWpT5oW6Pn6
DmkgCK0WxsJOTlMotphRuMZ5pJFuJU5QHh2RJHD/bhMp9CQY8rPKEdk3laAv0kw6
PAxCJZnzga/Y3sVdnQxr1jNo6rXYe6nEMtCgcFeqWxopG/IJsT2RvER/0VykEr/h
h4ZmuoswQLDSvUhe7mfbRDSHymfcAkwgKG+5kwZ1gvIay2/EFByzR/HZdLsI3jWg
nMK7fv5+FluPQgQorNZ2IBUw2ByEnwJgSeaXup4/mUog3G7LA99mfqm8bYy5FfqW
oaFhhGuBHzR/QU7mBr2u8nsTlnOIVlptPnXTqYP1uSitgC6H4fwbIs84xkR+FS1f
5O1XO7bP9hssQjMaHU2wvUow7Oa+OanvV1DOVQeMIHFfelauRQZXXHJzZKPNE9Jj
wBxrEpt9sSu8JQdQ2EU5NehwNRL+GD/blGEEI0EIqhlHzgyep0pUqwMzC5N3ddGZ
d0EK1lXF6JEvyxRc2S1g7D7/BaKodSv6gJl3+GINMVuLW9BoyNh4IF+8pp4AQzRF
rzwjeFor9IUJxYiH44LeBrU0x0OnBHYuB/+efdV81lqmniYK+09hQ4HaPoU7SZDx
DFl3junu9/dSih7l7CpwSBDmuCePrCw/LGL/q/j09cTHo18gyDqXMN70VZkI3XYt
IYHNJ+gF5LJkdtN5Uqsmfrxmnu0HZci6Bdnu2vs1KIHPCnUKFVlrAbptckXphEGO
qmQh6ZYfOXEC+Qs5v8xuAG1J6MzwYS3VpSUJ4rZ8fxQWukRktl4hMwGPMUNcNXAS
jNv3/ExA/mozWmPZ/eysUpuWmo13WcmHCpHUKIV7FZzUi6HlO/1xItkTB6Css+mI
JKl6LPzL62lQdx9eLvQdkTqOmoEMuPn4X+VeRSLsFWnMR8h5DCjOTmCBa8kJ9FSh
zxeAsR3F/bsN6FZAU2vpNOjvz1ApYnqSjBCBGBPq1FgzMjAY3V6FqKGy1T83RYUw
HjPnwZqPT4qHeCWIJ8pjjzu8sPxktyH5D7KoSNBf4gzK3nhuednfxf9u9by0XcIa
qLvHxG/SUAsEFByUz10MrfauViV7JngPXKpziQwCtMXJC6gGzWoREKPPsnoHNszy
HlHqmbVvqew5boRptg+/3zwt8raVhJ65JtA1ODABrFuYnssvVfTf4KfjvG/CUWcH
Ae83gd4+gj++3wNhZfbNuP/PNtKrAgcQk7Liql5q8360M9kcs6a0PUYlTgYoQoEZ
1hSGWi51eTjmQ3yv/G+nkuLLE09jX8jMwkrd0jq02SmfkRfeqTrzUuqTGBWCN2Ks
iufBad/+OsjNYyY2K3QAka9qJcMK31P0R/8IWs3SSiBFfwghliiQViB0IAfqOctB
aEiLSVmrzymWUFx60h22GInaeUdbZ8XbEIO1HkhfObhbAzXik27r5uAtlCss+fL0
rQ3VxMjWL/hIsCq9A9soNCGcLMfsf/Vbkh5kkiEXJU9R5Y+fr02t1q87I29YlgPy
XvpAMMcNPDVracJSQkoIxPtDHLe+Ti0o59En834M5OSqIT105rP45+u19Z++Lxyw
OhxmPw7OAx9rnyCquuD4EH3AMkAVPKyi7s2BKjHlYcHryiOACkOU3gCMNI1CB47z
6kSbuX1NZHm8wNo6Y+/kOXHl3morSFj/2VALzArV9V3hcv9wuOAv77/EYSP91HhC
YKI8Es10ikKWQ57vAUtgKH8CBZwQp/zacuOlrymhK6Y/FhP39rErJreRbSdNpvj2
QklsTHpDp9ubnpCuRqXOuYb1d42me7nHrRnWbZQdbhWLamomA88N1lmP/BzcP02J
1q/z95H8+7tSeKy94+eiIiOL4QSSH16wGHkAqlJdTqmg1o8TG6LYAapYH8pmZVcj
AaFHfGQFKBJbNY4NdAodSaxorbMQTWe5o55erGMol7jHVhZM0jIScqvM1yVTacB8
advoIq8H2zomWeCzxEpRKhrHKIEwclA3VdTeeEA+Cd2DFoqRcFCOKWCfeaz5MuA4
2YFAGNXGRQc0zrXFu63/CLGAhR9BvhdCt7iaLrSB4SU64UV3ncTYKx0SXHNbCYEU
WpngYjLNiIW46HtjqNmJS5PBoY7kZmgNbOfei2UhcrDhdybEXpdHI0y8GHFpHLHS
LJZDPRUkdAgeisIa1dSY7NvKp4eXdY50a9d5g2JDe5m0AY5TflnsAEDTVXnc2jcK
Klk5aDklLei+mQBaT3sPqazM/XCSWTT4r9cEvENBkIaAW+0IugS8KlRSzA64H/o+
/qyA0yYZjzP3EI8R6nBnoOew40stvQkvrOekupYOTmvwPfhcnWQ9O/PpV7sA7fdb
uJNebx79IXYOfMenrB4c8sCtQZH3Gaj+ZQxvjAsCPnQyv+1xDPZ7mSanrNSVQRf0
5/bKGZrSMeYg5jvJgUm4kPO3Ubv0PrFjGzGeiVEyL3yPUSRf+AkJydxeoLFtLKHb
B+yDqvru130XyAAAoGzLPAAp/UIn3x1LAWscRxynVu5DGjGCz3mwfItrm5i5PFAc
aR3gOtktyeVv07TIpLCJwpezTTk5GGX7pwSPPKvWv8Spbqijx0GpPZl1/gn36w1i
U5u3jR4juLqwiu6AK5rhoPQ/fgj2AkEd0ao98fUsIke064JhmeUh72o1JwWnqqrd
IqpnM0BpRf9s/7zSKB7TgY/gp1hcn1XlFRWBb/uboaWRwjQdD0ucZQGtTw/pAEgT
GxbcXVIACJZx03toIL3t+Tjxp5VCrTyNuuaVR8TS58+iT36ejLzwAT3exmtLuIma
/FCZdYKvzc5wgk+QyhLMfxU7GJNN8Abfm//ov23zg7PqiwTI2meJREDGvJgh/XRN
PQZure1LqEu55qfP30qjGmlD7Or1VynCGg9Qx3VBSqTCmAZKlf7ORNNAPrMS6FOz
RkCXpGnd/asP79Oy65/vq+ziURkMjWZ5eOeU1+3+ZN1R+8dLiaZAqZCtkmT6Fdxb
goDfNk91LM3CT+C9bo88Vk/XoVJNETWUGxj6Lwimyv0TneAryW2uETVCCGIHNwrB
JnFq0kOH27RXYc/ugT6WTyXi+ecYolBUlF0qEaoZ0rvgoUWrrwZOFufJzBxVZXBJ
iFRnlrF6BxX+nxEzh8jGWbw11BOAEBazEU0oBFqUeeW3GdNh9UPDwqHE5//7fKdT
RfEBZLndzsZ/fjglAqSAquGcVOy+mNfUOPCXe3oPNTYQvh7nwUscYyTuY0BCOSG8
I7L2viTl8GugdJyqgLU5LKbbrdNVLX6SZ7+E6vvPjEMFcYAJtokgb67FtRqPdKyU
DgSvxBVqjj31so7QqoPp/QVAj3hCACn36imL3/6MOums4EpLzPtb0gL4thziobT6
3SZN8lrcZGbkzh34qPLih2xtvK31eNKOU2ZKgS8mDw3tZN3c4nGhfOJrwyr8jQNZ
02l+VuVGeeYZmcuStu9HMzYukEkYUaEZb7XrBS5Sv4eXDcwmkx9mKYtGY6stg+7A
gJlMwAZochs+c+fTUBhZLSI0NCZFG8Fovd2afCY7KgCbBBpatm23ZC66YmWE4jOA
abKf2WsCTTG3kwzl4uX3gzz+HRL5NnFhHk/LFVbzOTkv930FePDuehvT3hXIYr1s
fN9GpeZ7+i4nzrZb6Dr+koEE02yWtphuD/RbYIvATgeJe4dawMxQleuuCXwQ6b9J
jEHVpG2QU2TcJNFUHDIXAQwl7/BNSG6HgQMZd08XVt/ueI7DbShQNKWSM454AVV0
IXlsOETKi3JVWcVqc2f+s7S4UdYWzceirR/NDvSC2k7BUmrqO6CuiXyV1IkANySB
3CKh7ZCZmELCz/wzWjuHodorLbGZlJhmCyzOgRimFTOzvjUFzKwDfZT250wSO7O1
vdcScWlc22mP9GCn02vY+nZqdLQfJ9M9MoMk0CLUigY4QXHoR5o+hNcYBZ6ARotD
mLSDEtdxt3W96iVKg5kIo+NujKngMOXTNqXVYNiAs3m6h3fc4SRbXZhdINXLvjCh
6NKnlswQs/kFL1kWz6Q+UOe2M8GO5SODcnITfmJoy8HHMDrelsv1PUevzobg/Wfu
3Q+/GKe8oDNzhSxaOcfnakCKcDxBd8MwdG0rFR3Bk0ftgWueK5gPVfePhtRaNlqx
MyZX6RIv7BDMx0UjgEryJj+m+LmBUwX45Wmcd5pIZ3lm2aTxSCDSSdB+oSTWEqHb
mX04zR/sSfjkicGownrMFYKfDTzSz+Ioa3KE8vn22101creXZwNGS0+tMNyIMSgD
HhCLZODc8/F6Pd4GlxkjnGkcIJABbGVdxLOIiEXOdKdIKsY69MtoM4QdQSJkEnXu
EDzRzObm2XTCDXlaQxWwzNDJKP3h5hv9YxVZJ0jfTCXfIY6RfRY/OnDePegEw7P4
eCfSuuFdCAqFp7DXN42wiJgBgmbRsXYDUkOXNwcFbCUqKHMvZzM0Sshy1QWHHbFm
1IAKTwqf4bnxu9SINhbvj56q01lPysOBtQyQu1xEQ3QH4h6Nayfsm0vbYFRJjScw
01yRh/kyh2RSys7bpVqPyDfzLLFCQZDSRWbNbqTF1dMzdz9gGa06Lxxh893wFG0e
489FSije6oetDH7stt5O0XYEMvnneTACmzWxJG0pVP84e4yKJl6xhh/0eVnBkHVQ
iPOK06rWdhs8YgNx508Zh5Abhcga3SQc8RA2AvQ8oxlcucTMDDwF00jgv43gaZst
BkMx69c6oVC1iKi1Jabj0R4A9RqcbOILbsOVVajkX2YNZd0SeGQVU3RXr574cQ+5
wmMa4rH+RJ/qwPsEMjXIsCwEiJPdzyuPdXMj+plx/QYNURVQg8Et6ZqvPXXBLJ28
R5cxuIf1NB3T+L7xoq1ROEhqS/4/31eZsPe55sA/tlmN40GhWMLVA3V3ZD9NCtwr
L3rI/JafpyCHmAVHljlIj+2DLnBIwwaoeIPtIjHfjsDWkWtd0P/4eFKEtjUYkejv
CO+254qapmCHkLmZ7PpQ5XwgD6+yuq7SMUo8MTOgG9gq1E8V7/obkxfSh2CF/MMp
47UMqnyBxcR20F8Hx1hMI7V4Vu65GhTvnIXNJzHECfgNoy9pBauqGVmhMe+ixrV0
E3lfd1pmX3k5ZnKUc/kkGmC9xkz0yfnNhQE8SEKHvXWeT7u9dTwNgypj9+hjBzib
Q9uIiUlqhS8DhSJzywNe6/xdYMCfeDfB7Uwn3L1dc7NfdyeyxaclxlfWBoCIgjtU
IP6oCZ3dA4p5qqS6tbH9yde3Ha3SimnmtsW8lYsGuIppG6eu8tfsjxnn0GOTBul6
AOy+grN5PIvLGbC9FlUvDKyzw4KW1OTJrO7KU0T2vOscwQIS9NCCLaMGSbVIrJNn
fNwYdbY7JtvPWigqikZkqVWp+ba/votHFAwQRVhzXC1/qOpRkzmdQyTEmSEX7NMu
7D15mLcJw5G7RUTt2okR2lYD4fe+HF6zx5UGfDV+eLnbTRm59KYVqHKcd+4LTvU3
xuS+kKKIljpqyf749yaSCA6FMkasamZRpZk+gMkHyAmubsry9yedGckIrGDRGC0j
/9ruZjFdK3SX6PYUyO9pzOuFa3jMSQE6R9TUtSmQmKZMDCb7wDihSKYAMocDxsZQ
OVvQnBFA7BkS0fmajd6urkjlJ8hMhpV/2q5EhsYtZ0/nsSB5372Fus/k4WV0/VJ/
0k5DAFOfOivu+djHNXAdNPKMzIOdnRslepm1L7yKhWfjLf2fDmNT4rTug4IPw6sc
XxDnV5r6Ith+tr9NA/Sy41Go9/Rgxp8aJmMX4ATfO+w9K915LiSag/So4rqIe4UD
UxSQcyVKrTzVrFM3osWVIC52e8LXjGkbF5JXzqZ7YH7XQPFU2cikjL1jA4K0HCIH
3VTy47iCMHzIlmjDx1PZbljCqCbkXioNsS5ebVcSzEaIOHa2E5Dpr6chcGgv0pgC
cGXF2QSlMYoyV8+JC9fz2r+XjxL4yhsn5DgI2buS0kG+ffStsgys5rTPji+wJwlE
65+S6Jf2A0XZpLs+f42YXsLELlbizmVQQa/lLd2WzuL7eLRjSpjyhzbh58ULXXlM
sm4hLks15cDwTnaFlj1j6yKBtnAt6dL/7isc+fADJtQF6lf5/wmX0qOelfUr/766
WSlrezWK82ouiRo5yzbfWIihiNRfKWUy3S59JE1vEyUYQEGlI3y+Uu6hwxcbERiz
9l+49CmA9P6CZb7QfyfvTS0S78DurAZc03VhNGtuTNLxf2sj88hGXIk6ytppU4kE
29uevjr2rDnvgaQ1kzzfOUvVRmG4mDp/NOnma47Y+H7nnorM5mTwkqaatwScV++l
hVX0zgm2vMG3UCATNe+9d0/OE/ymcBQTyRxTjmbf0Hbsw+niKbUUp5rAcxPd0ymj
QN8wMWf2fH1OiUuA3pSDp7KCWoyPqpN96QqCiGanF3HZ/2KjPtsvwcT87nm/4MNU
zq3sUx5eTfjm0z1iW22zBMkBu5IJHoy+b5BCABdI2/JDtoSlSeXMUL9Do+cA4SN1
+ly+3dq9sY1RnbVsvcjn0HfwyueXhHSFwbbweztLbyoZ5bExog6/OM+wds07x9ky
z44Trs0EDbFPhNiLWsxrKyT2KIk0z0kZR8xEgIsDACHxEI5nVF6lKiZ5lxSAvsgM
wIAkrIFXA2a1mbtnLaOWXPDVGPRkncY4LAns7nnuBcLeo9ijnZA8vLglLZ6yo0QH
/T4Nw4vDgWk1aVoTRux3K7tNP3LMh3CUE5OOkL2O6QgTSYkAnjRrYdEnxOdCsqbr
HTNC6B5QU5ASDBzaQpBOsUEVWkVHcwjJf89jo9KKtBfrK+LkUgZAHMN5jyLgrDbG
c52B0vLCs/P2bMW4CnKvKG59qDaUliNr3DsaE//tNWNz2wIrcoC420NF4li+TkqT
Gme78slMpbN+SYfK+q1oExCBqnEgdYyZ3GiIYAAaGBY7rlqEavQQBn4uhdz9XWtN
s8oP+WwfgbEWXtaQIX/SHtmrAeYe/VtSgFYdEu2H+1rF6RsqNAL0yrFUmKgPolb5
nkYIc2BJzuOgOdfymWxG0qmLjzIT9n7ecqjhE9PgDbdENcxP6G1nr3RiN8s0PoCo
DES+U+51E4aHFy3Zy+lqXBqQH7r71ZIltkeOKlBUDK0X6bP0xBLeZRW1CE9uw4VY
xKjygZOsUwpxxYEnPtXAzz2NSuiuKuNZRBuJEFg1sFf8wYFOYSksL52IMIxTxE0c
n554t272dBBbhCA4WaI2e8hLJkP3S9fVjQuq5RFqSNYvirLwKHAdPNNIPA9wFet9
SOn1RlJVdkOfyJWZB6Nnpl9rL2iRx6mvXxRb4MS6RsBug7QHgOfWCSeqMQKZEs5V
7VvcT3vtd8V1YU9UZt50F1gA6s4Ky1AGlqKLXu76U10MmMHQq1fOL0cJ2B3BN7jc
+5h3bN5WVrhu4Ibnzlm/b8NXfbhs3JOQKyjAHVGoGc/tvM62VogvwfnM6BVIzEIk
PiH/2BuV171qENhfkN1NxEv1TTDDjTSrXCq5as8k/M/Xel5VKnAPnDqT7/LkQV+l
9olyCMvQ5jZbNK53GqnoFlTveb6qweiNLQvwSfTmUAyCkolFfLXQ4brYUTtjDnlM
uQYgN22l8I8cul+hCq/RF4XnXFaKmaFXVUmrmQ7mZY5b4xNsUZMSwXkXD1w/Puh+
Wb3BD8FuiEwE4OEzGnRNu5Wy1VF+k25/ob07TaZxrqxB9VtOesVuMMujVu4QQI8y
IcQJHso0bdXF+yz5lyt1QKVXFEPIkbvvnH+3JzCjDn5WAfcfDmzcCUbi9Hx3yOjh
xPNAzSTZtiC55Hzoo9yYeRJ5Bq8HzObIBT+qeN1sL09XIgL9RtpUQ5v5o7ya9CmX
VV+H1Mj/ATmYdRWEVN530ejaIodp7+AM/u6HOuVfl8EN3xiRNSKC2gYbS43CPgz1
UPxEckv0cfu4COPjSiXcG9OBokncqPYIvcB01wHSUccj5XJHw/XlBMphalgX+RZK
6HeBr1bfDdBepQ/DTE/oAMNrUGRDfrx7Y/Wn3TfuPSFKttWSEpUC7N+GWrbmidlx
t1pRQRrfxfpj2VlMHX7aQimiRFDIgFUXn+5dv2y1F/ll6kvxs5gfRxzB/1CGdQA/
oGBxFEbYP4sWyoR9Cl44dHKVq2LFPt160MLluuUHVylcL+EH0JaCX8XR/kTYsnbD
stqGwKXVFTiNagHNWIheT4ARRM1i1t8dxFroyGYYLGera9eeWOdLH93Snu9UkMiE
WHZqfksylyPaTaUKA5rjz7a4Z2KztF2ZMYsYnU/V7B4K5fqN2FMZ1jy/64Zmr1+Q
szaWVeDJoDF2L37/0395ttW/MqT6s9Dsoi78+u3rdl0r8tohoqiEPqdwNNfiKExj
3g35G3KQ1wUofpNMhLEq38xVjN97zDeTmr7fJ4ROtFlS9w3ZakJB9GQsnP2+fcR2
fwVKeH0wwMT9LJAfyUlqwPhk+HuI/BUZtg+YaD+RlCIfZVjBECu8zDc7r6/Aw/iV
VA8Bb1+1bHnz2nJWfjUBx3Iw9hzQsp9SNMc4FrJfbom1X3VjQBE7P7T3kRZX4tti
udfLOlV1a/YTe71tsVvWd7PnejeFBxmxTM7Ft5Zs8NF65bRat4p2wdDPtdPckDFz
Mi6U2lyHarjVXctta09yfTaPPYQ9eZosZVy5tZ4zKwhztqb0EIZLqMadbrNggL4M
DqvktTJJDbh5HsXBEI54Rpv9/jgTpgPaw6K6BJpRMJnRTJOWI/Go6FnHXiEmwjNB
n2KJ9HiSX1GATe9qQ1Ns2ti8FtvhWDIx1W2bTv2MNk33hznGpiCDrHpKNpFRk6L7
3n3Vd2kCXoL8xzr5RcgOAAFJh3JJrQ3w9XTbhuj2fQmCRGohF7CMU4b+vPWO5S5j
dE63S64zdOhCj6ae4suZIymv2/IwAgi6DaRvo+kxcfL51Y/460nuDTRRkEO9iaK/
LsZyu/2tlb5uLsPs0zshHE7s7xjs5nFXM/ZnIo+JrVC2mKns/AFwoqtQPVu9zEDL
kxGhaTLFjmQ/oWxE3IvXHQG/lIcOh0ZZH4Y4Im+jU4jh17bphSBImxNWdW9plyKP
wLr6iN5NRSKA9mUc9OIVLODfLrOalCcyzUajDzgto8XPv3BlynECcccDnWoH3920
finfvT9nu975+GS7hVWrIe87CSJpKge3xQ+qDxmLEE4Ej0mxzLG8ZOLkc4+VyuZH
RHIk8QxEQik4GKAZxz+6/71yHFdoWKg4XLhyKL/3lt4WecJ/HFUoX5vRlbUVoWsi
m+aa8UFRaWvDV2vxeOuS4vygn8uNCjR6PB25tR7R+CbrBHP+LxgTv57VC1NrG3oi
oNKGicMt8DvPhDtrMU/p3VUKW1qGPNlNSnALfpEqi1ya8jZRE8UEbKRUwbaE14fq
aNA7XUPQPAkxTfOIiR4Y9DXwYw9+rqtJcfPwravAZ9yMTSV5G9OgO5nigBE2uFh9
89EzwdT9AiGtZ/staWPD+5k9+0jMls34ajZHU3Mk0VjXpWqYQA9+VBBOPz1FaHaB
/1DGe0tXAsAVhbcUDUuQBEZ67gLobyM8tUneb3OYuCWxfLYYvjZU+TN7bjvhBE/j
sF/KMBoj7yunAI/60NIo5HaQlrasvNB0ua6Rj76W4GqoYWI8CZ6ygBkWOBXDcGLu
Y38rm+7lNOyDxL4DLc7SGx5L6/9ot2+HorzHzcuv2lCLl86h1LjcT4VDYlvOd3SC
MGU+vRj0Z5quFNzcTJnpz/XGePwRXpeVy505ujKfvlwqQd1V1E4NMPQV52tOzvSW
sGk09WFM4wNkzZ0qlKVbGn3JlYiUShymO6+D6BefH6+VWD3K4IK/7n6qHhh4ZJ6+
pNpQbjkkKjOkaq4UwssjqQMvhZRK+2RsBh0MqBX3YH/hsGnxNRwL/nfg3lvuyTSt
jG9HVPLD+AX4WCZwbxmKcSwzJB326Us5qXJnPphvrmtnfPW3y3Y7UFPGKxw73P81
wNVHqzJeN+zl7iZp+xdErx+y/Ttq+ZxImWRFJT+XCy20qy51peATgiIZgfGXniuR
trJ/98BUKgNoFBR5BjA3uqGybzIaJ7weKPCD2yGZJMeQWanYrxLJX6QvY+Elb1gQ
fv8CtAxGBvmOM1/zCPGvSUtimYDSstmEHC8IImqoiNFAohhnMZNg1sNRLhsr+6Dl
BqHJIennhxoIdsL3esjsHrsgpxGVPHPno/a9PH8zJE4X9+vBKpa289EMOwbr3CBR
79KJqIxybejU2MB8Y0kDL8A4xQA6ZFLKSR6MMnrCWHw03kgfzW2iokDwAKJ5K4Nv
dD9TlqQ5AiF6E8lMtT46TsYpZGnMwbcQb9hV+aiGWkbOHRA3Z8pZcWtez4WVmrec
/8MEHbCgCMiJdCJ71l/TcS8pcGCmoh+AHS3/I9/DhN2hMgZMQS1PF9YDA0026jc9
fJUft5IxVp0tjXOnd2qR9r5rcPAiAijtuq4Sz/N3Dk+810K5doflxPSc06NzrlJo
wFzcsgBgGTaaqGt95Rp1DVv3Xi+8txOjNRaSHIxlU4YEvOhMWaEADq5aJtnuHZ1X
d/U8t2WSm/Yap/MGhsn4nB2s0nl5coDUAyne6g2TrGG4E7Oq0zCO0DyMdZ6OVg5I
ElN+sSw+wWM0c6lIO754CmOJGq+8HW/SXqZ+981c0SfgNghPV3Bp7fgRr1elsw2w
y4NS74GmO3gTqyeoWVOwwK5GLRUBkQLWunRKWhL20TrjLOBdBH2a+QjxyUMIRt+d
TsF9qIVBous749SVw6uLEahfUWmz0M8hjf6n4W6HK3TzkpsEEd84NPAXBA5/G05E
tAEZsI8xbPPxxuoS4FxLmVwGpb+Qnx9PWQXRwN6fGcSn0PtRWlz6TPZZ/cmVRWqi
5+nur3fwoM6WpEod8T04FUpp2L+h1++ydFRBYUk0qxIH3viRHmVHZKuQ2XjJ7zqS
UXtHRi2o7GoFf+hW5sXGPax3en4g5wa4duwyBDWtIhiKPIr7sQ59yhfILpu+mCOn
vU3c2CzFaxl9pEcUrXBlpRJ52c6CS2CnbPvAeN0NhmRGYafOQn42CJ6/BPKmJFBj
jLReJ9UuvK4LgyXGtBHbZuzIW7UkjoKT/VT4cVDQ2SxirTGQ8NYgQXimuHMTFpj3
Ti/qECcFaolkqtoDQ+65eK6dSuRsT/4cllKjus4/y9UubIkiEzx1oiebbCshMUy7
L9w63MuFo1XTsnj4dwzUhiK4MSSvjWUyTxNtUEQi7HCC3eReDzNgt++L6bID3lOO
K5c9xKME7zlzc92p7fHVn+BP8AGZrMiilLWRSVk8I0FY2szYjGygB3m2SF8Ptyt6
T9iAQgKxcINJpXuSLzoDPClYuKfQUFD3Z7JoK03zrWvgD2dhNfkFoKUffbGH62DI
aOpFoYdgTPABVjEnFR8upCwdEpDrpGmOW0NjCQYlI3EuQNgxwPTzidLwfIo4wQgS
4UFeEgs9s8VfWH9r2dxrkEhnzUp1pEONrf9e04B1/t7uXb8HhuiGbrGJuvy2d8bo
fGe7hxMPnWC6egRCCZzOsoaQShM4W4rAABJEO+1/evYvgH88VSAJ/YIzMluYaC7n
eU9x7uR8CQEBfSp71FF/rV40FmWCz2G2nOL0U+EVNGjbdDmpbVvsc8kgFn+b9D5+
bkfmKvtNJz4KldKxG3RE2IRzY1viykjlPAwac0Myn/kxR5SzPm/1Ks/cJZitlPyJ
lZ/3QOQJIhJy+VSfhxolmUdgRm9EDlZKKTlbOw/D6w0Yo3eOX2ejRo2Ut0b92jbs
QjxCdnowp3rUYWsGEJlyVUndJGJxR9pQh6ASeCdPZeKMoOEwqTLe5zoJowJQ2kb9
10BOfdSMLCh9fkbH0ZWTHiopwJPmEsFr8pjBn/xgR/c7uRnL4+NME5go2Y9GIGGv
oHDwvJhhX0Z3YkLzdypXIXPpvBb5PdRCDqgo4EE8a9P4vk/BwcPLdnwGZT4yjamR
iVbW1JM8BRX86nj1un1i6tg5tjdJPN6rKN2/mAQZBXX95mEL/+iTwxO24wjav1dM
avKPU7GsKJ5dG/jJRH+W326QZ3NwcUfJxSWwRxus6t+H4Y/Z7hGgH8pbXz8z47L4
LwpHgzdyXNbyBodQ8ke77/2USqBpPmc0tnwBsaScG0qyRttwNXTG/+PPVm5SsnZ0
Ir47JsPtPsCpdVYNnh3gKxtv0gbqpseZd5RmSZP2xW32zosjGUZHx3d9vSn4ZdjR
P55r05XCCvrJ2tjspprokpJJmdRwLHJ4UYEVwiZfpm4FAcZEq55L2Lp3g5AzU/ig
w8gbl0nXef2UjJrswFX13Wuu4vGCb1zeQ6g/7HBF3fqSNIT5oUB9UKf0WYecShxD
fPZuXog+A0KRFW5uH4RziRA29RzHHggzPaTWHUa45dxbR8hHAA+TH1/Zz3Rf6q7k
GtJ6O1nLy+7YQjMRzrA/8z2Ns2GDpqRgNfpVutBvyHoS6pddrnfbc6Z5/3iNiLDy
dFcUBk5JgsfcLwRIvnECyd/MhWNfPhhFOwJBkD3z4tX0Oo/4ewuPqg9pZMXhHkR4
pi5bzJMLCFHv6FMjB7kBcXM38TABA2tfgCqQjeUm1veOTrZ65VrI89K2tSDQ93wB
1zR5KfBIopAzS4GMRFOi1FCH0IbYbFykTj8cZLZ6yltFlX2QN+/AjfRwWZ8ZIXaZ
VPZ/fTkaDHPed9V+CjxglNbvwY8BTfeLkxOPCp/hgYyFPVKZ0c8iqqGmVlP/wSdG
+kGmZ1vgJkVNY4hnnz6rhKVwNLry6ohDMGWH5pYIhUGGwMGopApL/u0W1PXm9PNb
XHkB3p+Rz53c1hSogvwYOS2tIxgEfdHeP6wxQmUaxruDxl7F4aJ+8frb22TMw9Ln
VIcb+Ala+xvRlqKA79mpCynBBUxhGEtykCYi8tJmynu3MCvHzmZDgvT3DzAjOcky
DVi0EQL40foOLppf+YgND05dDd1eSp453LlWj97BEX1nFMbtWPwdol3mTkiJIasI
sJqwfrCnqMOKnNvuMOIJV9DnDREOXRPB8dbEC39cSwJOgu0gdr2BAyLkcucKjohR
fMhgRmd0+ssQKd/FZzsgNBQjIqFwL/lhRaKqSa4CPUzIIEV4aAVHMLE+64ZaJLIu
oG6PvFRd6bNFerWYwdkTc8Ixx8EerUV3njjFPWSXa0yaCCRlVt48atinXLUZOa27
cJulaLoE6ikUckq4o8uIlVDdeQWl+RZauH9zK9KtPYp9tHvMcwKNCX7Ab1e+h48q
ZwMTXbwxsx0WvWa9zG3novssmWTasv9CllREaIsbuh+dcv8h4fkuA/bqoh9cAm36
5mpJCh6btQzENszBnwYL9Qc8WU/MNVmscP1SkFHyfJuIOAmfOfscarWo/Wmz94pf
7Xz779Js2fAFjcZzQZezG4If9waRRaI1mUBzhDWM+gB8syvMwu83QRqhWODqYtlm
/oE+d0vDtQQCWNMPPJk1Z0DgREuHc/GdiCsatq19gTNxihMM6umu87sL28d9smJv
+A22gDPPprPMjd+JmcIpVoLmjWlx+hMkEbQw1NkpI96Tp/VSpp0Rg950rVYiQeGv
z3E8QistpQ+xdsH4CNN8wgFtlgSZhFL/MA/DWNHOEq4GZ85fLfN5TZg5Psdt28Kf
V8GGj/33qH5rvvTa0ySaZQJ89aTE1Djqu+ZRuXCvZcMQEyxWyyCNV9uc5b89A81O
SDFcv327iwN4D1Hifx4//u7+6rZF40GXGdjZu54BNGdaAq0qEJSnaaEjP9EjZzes
tMvyQmyrF5k+dVpmAn+Wx7TmypwMCXAAAftEMvtaPQuVI3f8DJd3TGXrtfaGM6s5
qRv8I/bSX5eOK4JbpAJCpZQuDdVuwA4zScLnoD7GOmAdAmXTZ9ppPl/HtuwLZJJx
qhUDlB5aHdsQutkl1sYXmFFj8Ye86cI4B3uRw34yDgMXXmLtaCqpradTZYoi2QQw
g3NjhGmdv4DARt5EZ4BngkVo8h+rHOOgdVYwmtcgatBNLOp86kpydoQg8Asp77CF
x/U917SdyWuvJi0Bvzu8dTEHMlxsSOJCtEY3gSvl+c38UbPzt4VEyQXjaOjAu/LD
qrBWiOctOpB+XNUYwhNqU8r1VAt/OexraRjoWioxXyvT9h5cX+4O0NhhP+wGKeSj
0oqS8NurxeMiKERhS/u25jRl+/XoO+3wSR2QRpRCNCnEt1EJfPTYPmuN2cK014+P
b/Tj2oko7yiW966gF1JdQ6/2DPrPJ31pTYgSyD4pFbYP+vxLcncYLFPPI3G0QMut
mwvM8vjp4BgO9g+h8KpPmaPwO+WY0gmC7xWHsaxM1BYf+zRKEv3pS/UgZKzUOvy8
0mGf4JLa2hpA/UlQFhKzxtJwHZ7HKCYR2GnYI7rYei6ElH8MtfKCl3KQr8BE6+Lo
iirK0sy4AXQdha3YMCtu+1AXCslDmOQrj+CXT0FWsCOXmUOQ6i8bOwgPSpffU3F4
TxEMIyuU3VD/Hb9ECo1Un+jP4xTa/XoQlJQu/ti/clMNbsacpL1LpAXkzAWuL6Yz
yob2tbeBy/G+bIZVGEimx3XklxdbHRin1ODkBCeCCDf6L4dPrggNL0B+fPdSeoy5
GK1+U7AUqptsE06Q5SCdDZBJh0e7G5nJMJu2qyqEO7WqeBc9xP87ywLnPsqyUdBF
57hSHgrh2Oiimj21x4k35Dvin1fT2X3OMpE0N8htrKvT1VfRxgoHJFq8oUYwOz4m
iFwk7NYXUSWf2kwBjCGZvFQhf1MiKClcUy53eImieZcap45k71dHKgYX60flUbOR
ImNxNXcvVVSNO4ZvGjwZZtUX0RY2lxgKT1ELQz8XLDALyRrWiE3u7/+sIrXZqckU
9C24Nu5CTJ7MVT16n6PH+bhEISPo7M+TiUEoaFQ7HFBxs1qF1ACzFB1LxTiSSE4U
n48G2iieZxXJAyWA7F3gg2VIXKGY4dIccCdV9WnCJBgLN4DSBeJZqbtfaOmf7QFn
c3qYUO8IdtoaQ72nfsZmxHRFE2HCgdWVyaTOp+3HfIfwMQN6JgGcLWAtC+gMeow3
z/8mjrGBLuxhE4iHOPEMrLIq7dkGfiP4pcNHohhmV7lXlHrtypSZSAnpzJaJyv1+
WIt/KOYxS49hmDLtMZibucDfdHragff3GaWlWb79M9AEk3Suo4t6nZY3z0cXOu/Y
NwKT+EYAt1SxbVzakp9g80KCEcSQVVbOXpsdC6pzvwSQv/M6qTSC3HE5sw17vAWU
PzHI6ASXfloQGI8WP0wSV/QXNZskxvO9jJOl1eoEhftBVvQtmYzgUyrIne4/VyGp
WlSs3MCMEQYoXqYpQZ1BMO1C+PGQNi12zyKalloPX8+u2SVZXGVcqlxJNYLdo2eb
SVN/mMoiLVIBDUvI2SFGPShun4GR/0BLqcanLEuviilwN6V6ENA11AyFwrWVyY3A
2on8lE08sEjrwUpVovRBHJcP1YVnIIb3dm+Ika8HIrpnijYsiXsIHowmUe34ZLo2
5+GkFrkLhciZW2+3YC38Jp7AjyPGC4/b0VUQU+ou8OfmTZtM1/sB7Io0tdLrFJFS
aXhZqNYJlkYvhN6Ud0/R1BZ22VTdNXXrAfF0Mjev302SGEcaOiZvezjGBBQJa8c+
+DQxneHfo3omuaexUcJ+L+/lCL8dLagymc0tv/SRzBJCBVTVTBF3kCpwyJEInkwu
IgIEmtGZd2EEINdv945XH65If8wOo36FohvWZicYo6w2sg59FTwb/Y+4yzQpU0rg
dT4d9vDQsXUCwBgb2fHyKPd+PX71nxeBgL2eMDO5FBWZhv4tmywTcFEYHJ4zFpoV
T2lNreFwi/EZ7t+UBy4J8k5eoFHQW4diktudNRuAT2pBIcgQfJHRPWNDAe83XAcE
8dOSw9dWpxszhy8mKQQrH6j7y8wnULC4XmWHLFYFI9QYr8mOyrslxOhw733n3k4l
b7FDgHulYfiBoETbuRRV0l33JhEr4NceUohBbg3jIiFZSPbMwf547IoBLjcA7vqP
rhDEVndg3a3nsoS59f2IY5fEKdKf/Bhnj/i5CjI8LMhEJDNsN0WyvEmLhDlPqGBi
2udlcFUT0yCrhtKph/KmALkcpsXq1u3428Ya3U31DzXKQXTwjaOAxV5pehtEowQJ
R/QehCc+Gi5wcOiczJO6ZKHPkpcBpRLd+S/XdE37mKOhdQgrPk95B5tF0xL8udND
M7XryQi3LYMXsiSh8uD0cgoJMuad/B6cVqE/+s6f6W1Nd2jH7sXVZCiOQl4NnRaw
p2Jo6WJc+ZfDIBu1Z+E9aXQC/EYbrWiK3RlP0ejbREhg3Qfit5OjEdmnxN+zFrDs
pKKioMVhMe+OATFtLfH90lQ7uFHY56Fzgx1WBc8+mGzdodCq9Lct6n+bnp1eTUq9
ET95/piLKtfaUBW8M27hNObUzfKg75Fg+6VtxU9HAM6gJSXMbeIq4EEmRWIgw0Zj
yNhSaObD55mCbGt/QtTLUqW7tU6QczQHLVxgVZ3AiBWPn7ugGKhc3/inAzEWLE82
z+OSKTK85FzyuFZNg0TsoL6FSy/v84fIHPA4PTSFt8Zv9jlE63L+fzzyiyKu5CZ8
rVvZ3WpEyIbRUfBzsDi0DUy8Wl8m+TlE1w9ykBqtcipVG5I9nLMJ2hf0Hx4U9SjU
WGfPoFQmuhR/nvdZt+9/GD+0q/mqTaUmEjlkcZtivc5l4pBEKw5ZQp5hmj9XLehL
Dzju6uHxgUqs1H3DgUoHNrGQjdvS2v04sDXEjwdwIyqjZxmq7RYe5BciuKYyf/PC
c1Rdwy8qdWcvmkjnQ/TSVwcQvxcWpScod+zSsrSy/aynBNchRs9FHsLXXdicvied
qinpxImwhTBt+OgTt8o3pZoka6uLHEvWwvX+PsDfqhpjOECYB3yKFqz7DLRpXdB5
dSAP4QV0jyiAkieWIzJQxv6c3WG1vAU95M8Inieyo43eP1+d22hkMkig2Jko3wlx
xIg8TJqJetWEQLTvYAfqe6bhSiXs0dvIZrlEQddmgSA4zNsXeqXGLKyUsyQkdtsX
heELsDdZSvkYbOIP9X8Ag+lTCnYJ9PJJZUEYMaBDwfye8ApvNSU7aSvmIb3S5z9+
BdgfLuKlEr7/2Rv8QgWE/DjUQbXLqF0ZmCpEpMz3n4lF9ABIju0Pb9PlkwPTVX+W
tiEwEcrHALFZTzLSnw2dc1gNxNEuU6QbPH3W9T3+HFQ8gJeetS8+OtgttmG/qKap
4nAI+EJXfAgYc0iuf2yQdBRDtD90zUrHB58JYHoUM1mP7ZdUkhqLmSyAbHlsOYUX
Jr4CQ9h2u6d8C3lj6SJpYziOkphvhoH47uHde3XpDqz+BtVrc/h6awDWG/IyCcTg
YuJo8kx6k23htE/lN2Sq91CYcYgTDSl1hRaKySAmktgex07oU+Li7smVAs3FEZJy
KOtWzgUC28oEj3FNKklbkshCywUyXZaD4NV2K98e7aRARLuvhy7Hc7X3USas33CF
NgfoSLHzaVyFpdMTZa2wDln+7wYDnYlg/kEE08e5bLHJx3gHhAB5QuxgWY2uNTPC
VaNNKqMZ1z3ANgOCogjHYAd/ps6YkXECWmyMhyJ5D2evi8DOxpivOF5NVG4NGlxH
8Q7fWRPXi+rKxoTDrHtmwsO9aavKgD466ae/qzzvrn212NyOd1ifGmiZG864dqMi
a51zWWfAVfymlF/53N6d/vsPmhX1XpfW3YlCQuQLTceDgu3k0JoW7+ZtRIwuowvv
XW0tURX6DkBJXSjDDKq4L0TibdCk6fkjfjLtXrEtlSaPDxNANCMuNDXqzIqJCWuI
yEgYgQ8gb6kX7EJci2/MBdUS4twmrkQgG/aQGKar1wNdehdr8Y0jwxhTVGWnrndY
B4Aw5Ofd4VvGHCdI5Aip4Gi9Gwc/jf5euvOZy0dUDO0Ad0RhKw9B6ydwAGE+Xlh1
18XKfUqSfC7NSXz+KjwaJKTUfW3Bpu9aLOrHXOY8gZ9kqGlFKsp4HXfMnuysYGEs
fXY7BbfFwxS7PDKE9ozLzPmhXqqq53sbTvMYtap3Q7fQpSYOfjRJ+gfBW781gjoA
wTfFs1SaXR0Y0yCWDzW/3Z9yXFCKMNsK+BAS2jb5+c+bWd3KZmhrkxA7D6LnSRmH
c2yPEbd+WyHwxTuDsQBgqOPWQ+xyxAcg3y8VHto9qKbPWqQCbAeomWPWwZiwYeGf
XcuaC9+UwkHUmEBcObNHxdkTHCAqp3IVecFeNCr2yyEjY/7sMJCVETE0EJDuCP7W
+rermtSG8jFltqVg2Sj+QGVNOMLhz4nF9iMwPOajDPnUhJ8mInB6oIoh9Yo81TfH
ujuNZx6mMLWY4KAOF0GauuZY17zegvA2b2g4uAP/hbgwFelJYEKPWQIz5FZLDVZX
rwlOcYyse6OQ3oIYYtZnEgXDFFBVTZ3eCYiMU/hQnIN6Xnn1dtdX41z6g0ING0kz
Az748vAZKhd6DrcFg1bkrDVkcARfbBR6ehP9shkkd/tJ6hArz0rJud84KI5F9Afj
qtlgEaG1mJscC6+WH3q2eHI5KphZSARgVnrhZN6nP8svJXIfHP/mjKkRsEAvKJli
NhdzgPeH7e4YiA/CnwxtVpnrr5R28QMh6VxpIrnVptkuEWxU9ra+K+4IXP0HHhM+
Zln12hdACHnmhS4zm4cGIolG581J6EhYgirZarvE9HxZhwR4hp0nFQoXxQFJNJjz
h1uzfCwwHjI+x+tDDoIXwxUfHry/R+bdce1i1PJVR1K5a5hzJdWhoiQF9Jz/7oY4
QbUb+XOCDZc2xjmyGr4x+YF9x5B3dG2kank6g+weTI9DqwLtOeFIOhTUnpYdhqmo
aycmMVRwMgvaKlauyNFNk5YtLD/ria8KlEMeL8A8zzCHqhiXy4AES1IzZqeUjb6Q
bKmTXBm5Qc2wJH/wTAfDowA/r2XpBkS15CTFMhvxU29ECtAk9TDPYziCOhWVNU3t
JKN18tBx0ljtr/J/eLOlDRXbFHn6XP+ZT2hiNYWyPRSmwz1AApXFj0LKqkRiF1Se
WcvDOg0k4cG38/eRZW1HXy6l898+PYA8QyD8b2IYI/wIfvVpBmj2CMBiLE3zo82X
bgGdaPpenNlAcwJSNuUyMq9X9+XtdEaoqJyydfgLBtq5acAozgLmt2wYdhwS7vfy
h0hy9wkw0gZMMSSTHP8Fm3dKBaTe3bv+pZZb3HkgpiHqUKBGwP5yNpmeSjGzqOca
fMe+2Zp1xVBKh1KYQHtpJVuGoGEP8cHl17QpnpRS/iGP2LbLDnbKfxBgqyIf74jN
5ypvZxWXkAJV3LiLCW3IGp5r0WEJPHyuh3oulZiY+eFWB0jcJT8A5n1HI2sKYaFy
W74IPPdcwUvTy/u522/o/bqhBE8d5wtGpvjKqPoHFlwMJel45EZskK9a5DK3BzGM
Ov8Za9OlZQXS8dXV+nxJj5Ac/9QsytlJc1CxMj9cZ0wbDeCQdWVbEC9nnNNQD5DX
L2/beXh5XuYX03thVw5xOsRhAl9DURkSiRq5I223LlCNEGHDXMT3CAVkuPjxjMTK
vqqcz6COKmZUtipzOFL6Gu/SlpuCxmif9jv8Bjg05I3eLuzvPbdF/Mdf1oUYKufi
aqMnxUO6RJCpSBx/qv+kKm0xJ4hEt4j1EY8rNaop+ke9jaC0dm+K1CZwEHofljLy
X/6uHfG0LYKr25eayn247r76pJgH8GMeHbe03NK415VjA6m8XcMGK4xUZHi6Ia4L
k5Mqj9rq+Hw6AgGXrBXmXzWwscPn9p5P3GiTFhRw+H5yzcZG1QufppME2VNMS6f4
4nGnHaKTw+7kSdZBHnINnEnNdakwpPsz/9S+lZjwp1QnhOFyHl2/1BW8VW67jbtt
smzGhOYpEJ/5b6VurGDhWENb9ygUQ2i3e+v7a8B4lJQgAufOmUQp4QRvYxWITmKz
mGii+wOjfJN9/ozwQUev2w+8i5px93CTaz3HvWbuYhtRFqPiicDKmZ3UIbdHZj0m
SpMSud4nGi8p852v817MYrV8c8ROrAu9trb1hm7lbHYkg+bWXAGfUc5H5tGsgpWY
R4BCNPm8vkMEFAFdZ56aBUTbD8THNSxfo7zi2F0jhu5ue+MZHZhgpi4FZgwuBScH
0WvtIufThxZ4WxVfsRGhoUYFYyZj3uiTVP/utkeBFA9SCQa6zzJ3BonM5zxKl5kk
TQ1SE/7gFnNwA2u7hVM+j2AT5KlR07KZPZC2Rq1gv2ZZGH6ZsxSKGauxVNkZzyhU
fdJ0kbn1N6RpKtZcShJS65zdpxLeKvQLTTslYuEFB40Ln9eN/PelilkYhm32Tl0Y
YM9K6JWW2ZtOr2NYbJJz6EJfut03WhF2cACkczSh3P38OSOhKVnfS++OCBMbVkRX
17NvgOysFv6Y3VTaS13w25PHqaN4ULT6hDb5bcl3gM1K4CySmuC6jpJ37H/b2mwZ
MAnKu/iXCIGQQYtsRDjT0VSr7HdcXJNEKamWgQHvNig5thL7G3CqbSFL1WVPYw4H
j1/5RvDhQv+WAs43VWoZ4Vb0h/qApvhhxcBdCUcADVzd5RszQUIwLATnuKjTEk+v
WFAykLkpLWOgbN9bFJStyAaAIucDkE+EQr6HVEX8nZGVBLuq8HhzP9AlkGouBfGz
t7XngQ0gmMRKUwjRkqRZj2wt0ugCXBj6ZSsKvyCpZBTKzzkORlz8UnsON3kS3LST
NRm/RG3Ow2xM4Vl38YjEWQmMTNsuJ1GkiK0QTU5pQqgrdmf/f/Z6naFOBhffkqkL
q9vlLDITw34arOcDqkx3Zul8cwI+TtPiry0YGE5eQ7/2OJXcW8pwgH0SiCDJWkAd
UR6fj+ejxnzjEX7BcdWf1z1dD6k4umi6/oUdemgfAcPkAYq8UYOdPM8Dc/3Fopzb
5r7sPOS+8+fZAmOk2dAdWamTu3AecMa+Frd52hBaIQL05I4UjdGBJmEOotSLAaMC
OCq3wTFvXPr1+rOMrYldjzVPQOV0Kj5o3jn69To8f2V0Nv7tfo5MJYyBU7fDNeC0
DMNzxcK+SWo62YskAscqNMN7lMeURk6R0bHmy0pChw99g7+KiNBIz5ua5/L/QkWm
vO+tH2/sDo+1XdmEd4CjScI44dOidUgFQkgCteeEH6iSiWwyNDPnIcuAX7kgv27i
PLxjaOef5v2iIqOuTREkdnYdfv7S+kOI5FyP4N6uPNSap4v5qDIPEoUtNxHKtGAw
oWAx/KxVxz03svxX1POY5Dt6lThfT+wgdU1/VJxiPndBJ55pdSRcNNS0lttdo6B/
fq9ffVeB5YY+nwTM/A1sULrrVUhyDTOL0vJpMhfaufGMVBuEFPowP7vLj1dt0Mo/
Z5enfZmT50w5NKTCSvtFQNsHy4/vKmWinpdvdZQRKzXo4/XmaPXrWY8NS5AO2Nu5
whuoUEDuGJeF7Eb6z5PXEOJ6agJ9rUrJFuU0SlrhRuqziEu3Ux9qVJqLIsBHhtxn
trFJPxYmg2c4cVhntQCGWdQrCupENFJbZ+uV//bUZyf+m1wJvdJkpeDy+o67u7v+
mLzaHFzbJVsEARHuMJMXi4hUzzF9euLTbnZiAYvx3VOx3bA7kHw9Eejarki/7e7I
OxMSQHqYd0QDGN/rEKC4L+w2ylc+d8LynT7oPiwptr9n0SNWyoWxqxBZsZuEKv/u
ScZfrvH68IOVLoiHNXLpt0kYqcCpsX3SPfIPlOSPsXlgtDiCTxbffmpSzCWUqqKo
2E7qAr9AyQnbGl9mSxIa2BleYJoni0J8sX/g0b7X6oGfaAlBkHaQHgPoV04ctypS
o+IxIfTCAuI/fi+DnnHCfrnkGnVtsZ/zAtuUfUHfSw3qZUKYEgdXMmH0olBqVNud
eDd/efduA191Sd43j4F3opSIFGaid0+w6wI43Ot+W4VHVgpQG7qGvQA0wyazoIRW
tlK2jBFw17ps5NxZ/AH+0cO38K7AyMiDvSb9O6SahLibQsqa6SCc2hsCNFKpha+t
TaXPeBLokH/KEnivtv3qHxPq7+AaY0BKFaKt+QtwhiODVl0Homq602SoLZfAouS+
Xz6qnu0BmWpSv1ialPkcG0/QLCuNTMRW88eDolvPP5BsmLMQsLrBAE+HphNL3zfr
bxe54/6Gix4J6ndSyia6VwYO2l5aIm9vsL4jFqte/NmqH4T5M+rkhZpaLwQmJ4OU
1BjYl4enOZKdM8vNEnzqZ0+0Y/njYDvWhmhUbfkoFGPoB5+B6DoA4OKO7+dTu0Di
MLHaL5rdxeWdrtnUc6sQcuClCpzrLF4ua8nF8bGdU09cQVf7loOFOta6dgsXR5p+
wu2I7s/p1iSYWVaSAFsRYQ+CHOVEysE/DCpVDGSCFI/2cuOcIzqg/h8wlWhIH4VT
4rmnZt90xHmUJpIIcsPxJ5c4vHRWtYDgipRZWroUUczGkDSKFuydJLl+9rrfr6gn
e2PzmqejVuqouJKcE7Z/K9dXRetqk118B6zolHttdD0UsK51KdIUw21aAWYO74TI
xttj6ZhebBrOUF+usuq1QiWIaXeEmdmrTgzrsdvTbPWs8MSb0fqN5aWZjpeiU8W6
D/bOdeyf53zt2SPakFLiz4pJbyibXCJ7R9KLyGK6Yzz4PFtIxk6A6ZYS3F9toyK+
j5hFdHc5Iwd2aSiatHR0AoCiWkO/WSJTd2eBdYkkBlezuiu8Zy27m58nZHyGmeuq
idjgoj+yTX58xMmtSySLZnvCi/pyw+qhw4kRQQjK1lG7TgA6Q9teM812x/0fh+qw
hs3+RNYGbA8bEXlmx/nrr+E7Yl88PyaPTKY6pr9qvnIlnOJ29SlAQAc6NW4SJ/2Q
yRmE2YvSr+ZlaLOIeQsJs7/x15WMKLRR0caJ3gx3Dhkn59uQ8a8sFhrBNj6dwXi2
0GDmww1ReqVN57rsq2Y2dSsR8J2irzffE4XQqeiQEOAswBxzVmuMLkxiDy/I++KB
P3DHNlMKV//ghjHnLZp+3uE0Aea1jHlfUAY5ot7r0b8YYCanINC4U6zTNp8a+nuU
PQ5yXTnkBZGgHGSMF8x15xrpAgWXvi3nkTrmhbd/zCGry2Fp3OVJcc04qMG7UJZG
nPRXHQD0Na1PsOtKWMu2d93KKlK/iH3XA+K8/85+tZHlYHtdEAdyju3O/ODbquHu
iPLQRZIwt5lQF86FBFqzDePQruZtV+8ZaK7cSdwM+IHx9njYTap90mno5xorAeG/
MGir7siNL1n4N8zcZLVytzoFJb03fdsUyJgY5eCeuD87Tt9V9A7hiSRIRytpKj4G
PIKTVJHDpqRaeaDwbOQ77UkT6HDRvRyuoEW4jGdUM8GSElpvszSY4w3DxH2Ijhqt
X8kyCexhTlzx+Fm8NYBmYDMy+ji7vyw4mFKGqcrKKe2s/qruHuiC76KYVdhHExJ9
qmbiFTHRkUhhlrHUyFhzhS3mhp1QGRhPsWE77cpP3/BleBPQcx7aZV0Hlnao9Fzy
hfmhp6/6AJyt+KnwS5Vqt1Z9ghN0AM8ibw9YMQHhndJB4QX8WHnZoVf8WqbNASTT
OgSkC+9Qj/505gtqxe7L4m0JzLE/P4tW1xC+UX04q/6tXrDq8ihds1wh9m/F7RFz
uGolrjPvFAOpHRfhR6CDZsjK2Jet8ZtBJcREeu9RzZRDwG24/34KbticIJnxqUUD
jSUUOlKQzkzs1vCLTO0tPlN7qxEY6xBDsQ81GN7V9ZKzEVR/qBJ02mwcX6YC8uSD
6FH1QNpNDVi41I+pL/LNmoXL0uxOpZjeXR21H008Ot1JOtn5+kAGUbV3tb9MCuLJ
KmNKRcMfMo9Yu5ATbz3e/hkHaQsVvxL4rfWtMr7VBABXmoMLrWLyza7uvg3PTU8e
4YrX978nGnQC57Cx5lYbP65V7HXxAjhwSYHYcr5bTiEY5wy4/mwZTn54ypJo/hyQ
Q+9t7gTU5Bw2Z80EamshGIBvnBvkQmh81GH7TBpM8S/YmLqdlTUsj5uG8yGcsW76
e+ts9HcGrFNscC+xwE5RIRpYLtF21+H6dqwaAhd4Dulv+GROZvPkavuusa9OLbrK
f+6QHPQRcVbIFO/Y+wS1p1F36dvS27AUPQYHbU2eUY0ivjJcvArQat71ONAL9q8t
jAwwGFhOyFGvU/XpXye933e8WhM9UgxiNFWYcEJt2JLyh/Aviohe9+9zka4tmf3T
UtX8tkBva4+4aKV6DyIjdCpSYiDx7nYx+2I1eYSH3VYljDhZ0AJUuO2vGF9gHXim
alsz9AWBeREbZVfR114IVmRG4V8+eBO9AfzIwJRyDPwSZ46ZWCRg98OiwoegR4By
xn52CQ+v36WnQMnw+8y3AawROaYg7zhLI6TOa5D4ItNhCgi3Vq0yDPXlXknEglFa
u1xANjMWOcUf+F6vTI80j7/i29C94oCdJ0RD+v0WKS1IYtNJLvChcabxYAghFc3V
O0Jly+bCwl2B92k3wFG8E/hAv6wkFSlGdcxUF9wCgM01qqGiBxACXdy58/r97brw
TYPxE37WotC56jmMmdGdAJS4z9QX1j4EClIeTm+Q/gTc/8hrouJAZH9l7K/SWF96
AlYSbw3N8/cRfPprm79XWtTaLuYMD7+Qw7y+xPKiTUo7TzIkRat6czrdlHFqas/e
riO53ff58bFhU94IHE/MllPKdmnaFicESuOBS9UP+yi5T41n6AcXf85RW8XuOV3l
AkM2bKi4lN2M4m1qcYv9teSqL4KuytFVyLd6eg7+YK9GFABLBfLq5CuzilKQ6qq5
3CzfHisrj/TIKvmVDCg0Qk/S+j3JNzjAQ4pcNegpV2oncmwbNDb3OU0kJe0mo7Iz
nk578LtI86F+lRV5GY1+rWMaxEnfBeEM/F8w/YrmvJe4wklWXqB7quC8x3ti1MXr
tHEBGVGXKCzX5Uo9QNuvo+CjRFmbxW1eb/pOtSryDoi4TY6vYgA8lmnaK3lrAtk8
zXSMgIt/nqTuy6BVkq+O4IspZvu7CQUp9iLKzG26SWDwyu4GK7GUrBG+5Z3kp4uA
RQSdlIvOqMOaRZQKqbetBrIAaFckvJ1vh+13minlxcR3AGC1zJFrGvob8qhjqZyq
H89aJ/xLJMwHxpHD2MjZRdvsAJWmZELrbzr4vtDOQ2FvDaFNH32OdOP5ooPAXsDB
oEMwaQoWJap19z7iGC+vPgTzrbytzIWrf+keiWFk/SHYLl56FQNMDeoNBaWgLiXJ
NlRZ5PM/1bTWavVOj+CAwo3QhGS8Wm1yvv9xheQry6pQp5JSq9td1B2Ay3rxeLft
AcFxuya6qa130oGJktfup4KgVFE0I+r61EkDKVqHgDnQag6eH61DXHfLP4Feuq1j
IuEsp9LuchlhqqocsxJ6wIcHvuCylVdeR3uSL+981ew1dSM535Sw+quLTFx/fRp8
8TAK1QSPeAfPayZUiXUCOk91f782SR4RwscoivhTMKJ3WxeexfGN4xjXjrIQgfQ+
IACwkV5A0vHLWqSS/O2oLnGJXOwG8g3V2GD1d6alvgQqNZ6lyWLB/Th/eBrOm76j
FEVx5DvtvI33rPa+meT0AOPJrwROkcDIVcsqxtNi0UVjnamVwabpqTqz9YQrAoyJ
8CFtjqMt4yv749zPZ5uB0eJrZx2cFuGeeBifWtUl7iWAExnQ4QIqr+8lDRUQDCiQ
0GkGr93Slb4JY0SfmRbe0dU2eQCgEckBCTzcQhiAIgsaiDakkB79SNKAKMbNg2vY
+hdIMGpRcWKd3CxIsRwl4QAYuqyy8s6SOgem1m0TyoT39hcrkApRFlAson0yOTez
aszNay6rjt1YGG/LHnt/CHISBmfKQzGu6xzUnGDELXwjtPN/PeEg4R2OCYM3VfNe
WUd/gR7UoTUnaLGVLz3xoi2jBg8jaKRcz2T4E8IKx4vcebk+nkRnILOe9DA3/ubC
Q8pKIzrPGLg5b8jW/KN31JbwOA1ghRkCDUYF4/+CJPqAi3g8Gq18euA7yJq+/6cU
4wXNSk6EtNwtWCL//+d4/K47fkijotA5hHLcZpedzr2KCmu8JoSf/sVAjlqg57y8
SyjGBLRQXLO4C6SKix370NoWDvvYBIaEwHXzFPrlGvoBxoutQUsYvOnWCS26OpTT
Y5ZSRBkSUL888q6y5FrHlZ4H9VJM/1eH0uNfrJECuizaYAkmMw9LSUhuPlnHEJT5
hKkYaxJAtbEnbstmTlhGP24SmUMAQyfwVGB3KS5juyeLiweAa7LfaSm59eO+Gdyw
/2ka6LUTIZ5JCHw3xfl/IGSKVd60L8cY8ONmBs0G0RL5T1nm5pQ12EiaqobmKsNV
R7PKq+7E8bN5kqBTDKMjgjt3Dpr7et57X6CSybAASFw+UMuvO4QzE5o5Besr0oRs
p1+SPJ+I3fnNs2yYxeufFwcHlIRf0kKWewOwz6kMtkmeRIOm1DLuIU0BJLZQ2/s2
4KJ+IG+WwLz0rCvq7aBCrLUCJp2gC3dncU3wL9Wqe5OL7jMggrC61PdZafWqmld2
3zYq7bEQqU3CgyFrai5vlm0mSuhIcJ9X2S0gNnyAxr/8V7kMx5ugO5WzSeJ7BNKf
wUrlmyZQ5sRoZF59C2O+XnU0dQ3VON22TzKT/fsIUvf4neyLY4e+P7KW4b4iRZ9V
tMlNaMQjMCi7k2zMIR7F5DKMidwfn1nIMA8lxCCLFKWtEM4LtF2aW4+w+8M/6bFm
zXZC44+qLpAy4Orb3ZSdR09mxdKowN5s0tgL1VOPQlfrMq6dcgh4DO4nsRSqEZx/
1qjM/5a/mPV0Xj29WE0RWuorawZXFwEabxh/jDlhUTDKe7LYW1y+hsRleA7eoCNP
8GqoDC/UttH7ZWzVKeU167UFknC4Y8szx/QDI5ji5wCLvLTJi0HBWh2awalLPCF7
BjLP7ZL3cJ/WU8HuAQUpxP+L8q3CHSzEp7KJYsJjLS/vnKG068mkLW9b7TgGDTfO
2kxtbC03vXuNHxx/uZRjlFsZLEYxmIIXsOpAh9XXAEVbD5/GORfy+70I3byMXhiD
FweXgbDEZeaSRStjaAb9Pnowwcbu+iXjNiSe1NHwffGBWUhO12disDN+8Xs0RhKh
+tMOwrnvfCogCQpR+56q6LbC1lyaQESSHiCHUwX45emb7LDe/55BKkGZsBx25QF0
zPuVhzn2EEL0eSiDgzWaLkifVQw+rDl7hkBDv0nPfzpD3A2je4WAa2JNI0ra/NV0
mImEfcG6MUtKcUHRcms2zMtCF6mdJ8K6hdUselSJi4/dMdi3m0GSZtZIOuQApXcq
J0eeeFdsz8E6B/Ph4+Mhp71zynJNCkaFOJeWlXAQjhDrJQDcV48styow2pUWsPUY
QtLJUCzUvrl+eGnEXc+B0cH505GwcxQZXiCL+5z5E/wkBt4LFgu98ZA6uW8iSokU
adfVNGOOFXtJoiNpRF4+n+/VPqVOQfVtx8ZoR1tpCxNXprkaOhkw1Ux6BD2H8l5T
zp6IxC37adu1dzMCt1hc76JWtiaqKPfwqv3iIRWwAn5hC5gD0LZyG8ALZCFdx/vl
j47kiQI3SlwZdblcEPyatYaLZXdTRjkK74r8njqSlXaR+1f9a/iC7TWPdtjJFyXL
GlGQ05ZIIOc1AhZZgtQhWNfVa2Go8k6080jW0rtYDNePFxwjuQCRbzpPMgjZiBSO
oJBbq9yhdVUGYaYiEN3e/kvAj5/2xgFliqN3wDGQXq8gnpzQmaab942IWQZNpXar
/3fa4ZBYVFLLc2H8BOTse6k25dCsxeLh1SOqYRIn35Mjc8AEgzPU+Nji/RpBzTI1
5ihbB4X2wvGoXKvlXTUI4kp4WbD/9EORGZkTO9logM7GPyr8PoWEmYEadpIFyiqO
tOqSnXtLwVsjVXSr5Q9v4gFJylnHtWkOZw7UiR5LIgszl252xm58eoVuZqQZyAk8
EmqnCbJUNhlH1cMliobNzR296x9JkHSQvBCsGqhkY0zBHpeianylOkVcgcNhHLFd
/DyeMOsMOSRdZQieIiSLrWcn/oLYxU+Gsh5bsbbiixEMM+cnwWjal+xajburupxs
w9l8lG0nyqRHuZZyRR1Xkq7PmPPvXTGbX5JZuPMWoxagzHxvQ8V8xo9Fq/qkmVEh
k+/G8nrhmOI8AGxTjXM+GDhx6CUzcZmlDuPINmHhvDVGr1idUbc08unMGghVXpkQ
OT+3Ni2MmcO1l8xqgNGvV+n6QerDKiOAQTQma5guGAt0W4LF+UBgY5pD31SAnsVS
JkGWmNHSwt7o5inBU4uuFtvpa2UhFe/yfPs1ZPiYiFQcs+mV2e3mq7RO2+8u1wAK
uSuFq61k4FQ/YLjdEFBBDF5TrlPddGQgaoDEzkHarCu/9xwu+qkIRsTg70464kVK
KCvUQznetmSxDuqwUodjUEW7GirnnKZFqLlwZbnTwowurXhz1bIza0Z9dwH9pAER
ZvlpQZLKS//b0nfq+DbB7mQf4qu7E7AB6lGE6S2SCoXcDnHQ4dfHsJWO4sHkw/ra
EgJ07fZYVrmvRWMbC+1qVr9gbyBr9bo+Rp/7dv7ULE/npSXLfJ9n0VwR9g6XJhzz
VN1J2sKdxVb4jxgCIYfclE/T31taQYmq3SA/ei+ChY71MuuktAzb2OA4rsRMxELL
3fM09pSUw2fRNEjHzre7GWPikYXfcmFVxE9kDIeEsDt8ZAn3XEVdLxTCC/yavtND
xz2CEqVcTbS8gAe8CvehU68M4nsPDSSec/GJluLeCVs/1dKWWl2wvK1RtynzxjLY
J7r5/pw9guEo1g8VxZKI2dktzgIne8HEThYqeMYYWV9mb0YwortiEYgooAx+vQeV
Bcu62QuNcX43kZ5ERw29+X1AwRsQqAsFfp4og6yUWdUqRWcVOihsqCP/OBMPqG83
/rZuMmEnmdYGv9drhxlSitxpnIOKVU5rdcuw8Ck4+A3YuakxxsNNoQq2dTr/5C1V
aw6PyMEKbpFSMqMCSTdK5SN5XK1yCvrGbZBwFjZmmkCnzsOPcV5NFOSb7q5iNe2Y
lWZ1qgbOm6K7V5rPllOvjZv3VP8UUR+KguJ69jIuiksm++Wokp4DHyZYhaEcNIr6
iIlWxoBqQFzb/QVXdxmPP8d9S73b6mJ1U15bLEn8VGo0iMyFc/bJRtL2xjeuU5AZ
RnK4pPhOEWNpweHjE7D1xTNRewPEphHG3Zch7/XLQrzX1vFGashfa2UZV3lGfpN1
08Saoi4RBtDUvVzUgc4dYilTCLI2LH47QzT5Ftp3w47/tF3du/aOPA4/dILpA0hk
gdzJLtHl8zFQG4oXXisZHsNEyKk21k32dYmiFsGgPpKV5s+YjwIJnokaF8Rv6Ffx
4DDSpJnakC4zmtCjTQPtT9ffXNr7oZXBixx6Juf9WBRFzKRSTtw3MREYI6wyjoyG
AMWAzdSNpGhRYg3BYLq35dIzLANYhdfmUwpyE9yZacw4D06LJfCR2jIfQ7Nqw1Qc
fIPg4nndJ7LthY17yZdO091TFsjdhx/JGRt4WcvGBFfKs4V6UVSmzoC7zJA+PEwL
PrsGvUfhw8NRgu9TJ5zLuMLrYaXgJaI2q2ISvQ7jUt/lvhqv5RXpA7HQ24bAniZ8
JWpbAw+E89RTEFkzggD39xpZlqR2YujJ0zacnJCed0WwAoLStU1ui8I3/29u20tT
l790d9tfOkiTW85O4cH7zi9M5SmoH+o9Y3FfI6/nYO7gwgjgliFmsHopj6gC//xY
JHRAYE/xDozgyiyE48d0cVeH7NY5Hu0UR+I9yaK/43jNAGG7QQDwCF27XBz681nE
GOe3ObQqws5mRk49XFfG9rMhe4p6kZYqUENKDSTVuo28NONme+nK8MjDcTL28EZi
MRtiVDdVnIAlYrovjFxCITUq0OlAn8ENdWf367MEcA6WaWemJ995D9nbBCxH9qAM
RHVSrMtlG+9C91LueJFjAoi7sngvlta1cGipQf/uKe8rhKy9ZnkC9OZ/VRuV+lVc
H1UDfR0wljfZseWZhlOODMJ1OY0BZSuVU1XA/ISD9Nl5eBYFgD/gOigjH0pFWobj
QiRtwwrihGDQKGL/bdnzkTQLHK/GDvS367BZJsSsmNEpasGOJ6s12BFyEWpDqXwF
7AXcwIY2hhnTm79LWOFW8ljgSWxbnVGBcBelPzjmq6rejs0JnmnEGBxIP0F6kfki
7RX64jYc+OEpzrCDZMBm1wK7kscN3f/jmQRFUvjiQiilt0kB+AJaBrzmHIiVQ0t7
UZyYYQKLDfRO9URb/NQhAe7PJ1Wt78O5RU6I3cFREbNCEx1oPur5FpKV1S2iiLAS
StJ7iU4vxaU4JvM4V9qY1rXSF46t3QAJaRxj08q3E6Vx+tLcyy6WLkFi5xfwXw6s
v8m/qRHKV7gugF7qw2xTmo/vOAKjfTk8BaFUr/g5igGQhK8j8TW2Lnnx8S4j9Op1
zj6Pqb2z3Ntu5VY3sZA05hB00Uq3lHTgFh8yoAtf8oC1y2kPuRxi5Lrkg+G9l+/j
nY0zJWezVSOT6oTSdqcxnTsJc185Gbde7uOZQv5OaObsU0CX1mpAqlk5SS84v4Nv
g7rGT8D13zMa3dStE+LOlPPkuR4ZCC1H4gxlYBcexWM2o2ZkKerV3DzaCgQHY20R
7mKZtzKJVmvovI3/wwpry0XaNHixvwDR6W3+xc33++/j4sRNphx2BHZg4SwCO1yp
VHh1l+04tnSY5dw1uhdn8+uhb4RWYtaqRN8y7dGwtPqmiADPU4+03IGrc7ssS2ko
VCW7fGTMW0/6IrDrgvcv167v6bSU4IbjP9bnH0gJ2wvkZw/HZerxRwY0qUpBiOmJ
bvN4U2XjAC3fbMCSz4L1ZyuMS1zWeTNEL9y7o3UzqOVHHAng6mtLfkbRFSJtDoAp
I5ZFFbPx17Di6DKskZPvaGLJSmJ9bwgg+lg8Yzx2gh8klMpc4PENME8Tcd1pjEwa
Wff+8XKMJoz12PEJaZLu1buXOCXZp/iPhUv8VdFmpskl8vkj99Yv+S2EaEe+rSuD
x4W6S08XT0d6lO+dKA/VTyd75u+lhW9rEOhzjEyfEET3h3aP5d0nEoHStAZq1CPv
qUMXpVOLicfsgcsYjC5RS+TaUBPcqP3DRKC+Qk0fD/mn9MieOu3OAXGCd4WSZ/QW
BkKTLtQlgHLa5aa5v8fVVWzsKvXsZ9YQrhvAirNFjh2JyvJY2Ea2DWJwAwVtRe81
otCSmyVGKXY7cWmqvMMnC9p1bdT9W1Ti6RcNx0MpKt9eCc+bd+bbFKxaKy2WIH52
+n04Ws2MxNubuTsRhFgDgj6zEaCjb66E69Qod5oNEOsr8wygCgh95bOOaUa5BiuG
2+0fvpsxaVUueHCeB5fm1y7QcPmwItYl066erydFUWLOMgk+Xbvo8c/Qta5PGqJP
tbrYITJR9vSnGtNW0Mnrp5ogSiPc03W8RjZXVI3VTcoGeL9Tq0dK8miMWyqfD8W5
zOeXFUwJzVYuSNs/i1q9Pcd/QoWSCvvLMGBhh9nHqQ2WsYy2Dm3Uv740HuJYzIol
CMFbxaLUxHx2I86OuLMd09L3mCJlu73mNdf0dli2FpBlbgopS+AJZzl9UZVPYh2r
utTjDOziL/X+j3YR0fLECDoBwjJ18RMJKEzouAPQRw+FOfULQLL5Zm0bfK/GDucd
M7EJ3fNEA2e6Y6OzP5snvyreJL0rr/8Dp7QIpeCvysHsZJZuWUssEHsuUTLWWNq4
mAaWa/yHSfTYH7IG5WFUveH7BdoFNcazrqxQd4e2F23zrBOzurCpobbO9npPx0vF
HuIfYR6Q3ey3W+JoizWcOGFDd4NXfIkOpqj1BsCKpDpu8cfiXzp+ru3dV+CqJkGX
hND2foHHzeGpf9xlESbNYUG03H3WORAHG8Q8/oCvbLcDqw2ifc184pPcDwsFZmI+
GlQ4SbUxEaQ7AIbry/g4erkIJVlKF0lgP4wvKYNavQsV1Z29I5ZRrvMnQDXfN02h
bWh1inhXTQqSUd0NxyffKAXPN71QIlU+Q/gpVIy3ppcFmxKJ1ByOnmSSxxbGPc3V
FSqe/UKne0IcpCfCvG0e2xzz4tUyTtdu6ehM5B9Ff1MP0lxm5hoBC+W8NNB9p+9A
Pv0SBQkf3Ynok4Wmxakone1FQsNGAJK5EevoPpb7Q6tOhP+a5S+cuszCADwAzxoe
K2GC1vk+lGKPyGuafTkIV5oGsmeZHy+W3rnoIBYuilFgzFxTNsn/MoJw7OX/of0F
Fq1661LaXW3xLLMxQ8Qq8EGPQ1WkHsbxv0iwiTeyy5iHBrkrTeRrdnOe/VBT8tmI
nMlRFoGDwIgfIGudulwAZXtcOLqsGRZ8DRCtft7cFxSvs03/DBa8bFuZvQ2B1fTr
NoDMEJCYYudTJ7zcSRYy6K6ItDJkkxiJ6O/19G9uJH2+IkQYORJhPR79YhVQNWHC
tXN2WcuDgmcQ0bKSRnqVeojOeUeFbiABR8vLN37u33hwQTKwO/Nr2be7aZuLAute
szP1y7Dag+rgUIAiPpt5cKvaqFrvPSM2FWTfKOlGiwJgNPy77dGfUuJs3AHLCS2y
OmYwgP80SaaLEHJ+pn791qY9Zc07gUu1U+YBy+0lhDO8gGV7meD5DwMNt3xDoUPb
7SAeZIEgs3h4y+vBoPjUMd24p7rIScp1SYGvSsLuLSw9XDGcRRiuaDkJIUK1bKi6
NPZyEYYHZ21fVpzTcTk2tZM0zzuyqpmQ5+Ddx7MERoHpqY3z8DKIzqy/WMt/zan8
yX2ovz2qGI+9XJDrwY/vVC3rY+V18u3N9spCslMlPLKqcokFEnoLZshAqU0ibQIZ
Vm31/9giKw406F+EgOEYzpedPCO849nTpBNTTbrjlnZ1tTRO4o2Ge9WzBVuYqF0I
LCGbn4yC8anFne9YlKoG5KGTbBImTSjzBpdASPz2R+5vC4p+LzzG2XlUUa77YMQd
LfovLxcw7Yh7yUCpbbSGNIgqxpl0bqJL+vw8P3vXDb0E61NY3qT0DAU0IquT+DH5
dU63UVsUvBwJftRJudCeqdSZ+QdwWQ25skSXDlu0n7Qp9/327De7l/9LxWBD1PaN
+d0A762zaIGnfki0awU8ef3YWy115Pz1jcRsTbDjaUeNnocGcDEzAortlXSweO7/
ekZF96rIn5HiLQ1AuufjsQY6d611RBvFxYk/ylE5mJLpOsEePzPNsn26HjhYS056
d7kpwBXs4Jeszpn61zP3OGN5plPjYeVQEN+nJhMA+ugQwReHflyGLsf4nafRbu8S
VXFBXEV0+EGlDtQeLuw4ToiVLHTex7cYyhka4ZXiCKi9R2kATlDO2bk9dZ4M5mjK
lUx/Xelr7wE8tdZDLHXXCpNEAFKztjPxLNferYjePO4nLNDlWloTGwCkHdHUpLLI
3kK30zfqrUqt4OCK0koq+S5kDa4M26TK0MlWCXz9YPUG/wHxMVvPWRlbJ7Chyvol
uGf5xf3PWxJFHJvl/jPbm1MitEJIriR+PshDhgIH8Ys6LI+FUxTUqi6ndfvgQpWg
UD3/qE6XPvOWulPmBX7Yyd8bexusPYK9JKg+/QFgDq6af2uUvHX/jRgvcRHP4vfd
VMKBBmFTFCH3oQaENPbUFeV9HcAeGVEBcaUSUD1auc2zb/uPrtZuLKmpVnvFU25p
TKvIECOgNaHC/i+2MWTN96jE2wL/UxxX/NMaBW/rHBBOKOG8JXqMjQWRGWvmG4fL
kU8fMy4xBfQvbEZQBZE5q01Sc78vxKc6pW3GlzEqbkwHHXxClmxlS3tHL7+2YWpW
5J7dt3rMdC8+oI0zm86hAm1cSPfOKNsf64BK+dxLiIG8tX/jo8Svgcvdq4FONknJ
E+2Aqdn4h1whixIN9doGGcvjQZlCrDIxAGPtvXEBNwFkK38FqrmRuujX55mHu6Ge
fjolM3Fum6z2ICkpFPqFbVGZNOa5lGXo8kHi60j9ABkv3tX5MpDLJPsGWXAXgK+s
2aEcZxGR5glH9epG4m+PtnZQhLJi2BnLl/umvBw27MKygshNhjqTUfL55DXYVdNK
5d2WB/ZgrQDPcXUi2kkjlnQBa+Q4wTM4lqaRGMyhEuaphtqmmj7eb3OEmb/mhHoy
B7mntUut/qWxZFAOHaW5awT5Y/gJiDeO3SLvRHONiXMFXwcwzu2XPrJmLVb8uAE3
bSnOsH3YnujUwaF2f17CNq2ZjDg2DtGV2d1Iww7gyWLwJb9SqtdGOYUbF8Xua2Mg
e9r1FQpiuWmeCjrghV1uXkbOKFCFDQ4mVuM52SykExa8EUelNL+gSX0E1fdcVDzG
LVn56uYy40vwa3qn1gdbjBXUD0+apbY1Y4o1Dib3ZH45j4KDkorS8lKMRJoBIrm5
3DYOl9l5d/8Hp2x4TvYiAQbvXf9pQQRdjRrYrQSaskls0VaWn4Zdk6/uvGLdVW03
fEj9XYi8KFsG0Qy7NVXzbAwIKuAlL8KnB42jHXlQjnGV+AfXAO6bbZiSZN3sx4YO
l8fNkFwrGahYf4B9xlk9a176A9vpmM/mZOc2zg+JaS4iTWRS0ZRw0vHrZWhZ3UQv
TvyIXicuYSWkWC5bwZvocBt2GhEjoCE+hdKkXJTxOgcJnuft5Nldh5EkjmHGfqW/
F4quvxYlr/N9wzNil+BEojVMsKcxHY8V3dcRwM74HtL6yQto+wFHdOE3sT1oFt3r
e3+tbeswbbWJ/z68DoEgY2ylOpGeerZCRTo1OXf4UsvzV7TjNLdN9y3/Z39jCkzt
U9QRi9nYyRyVO3pK9kG70HMP2BYOB176qR80og4HBDHP9OdDe+1dYYCEzN9sFmwL
XTyVINT+GQ7khBOk/Zou1gc/eWCXFe6/Viz4XniLz6fuVxNoAjxVtVCkE4tpngZm
+M1Hf/PU34o0owE/812McHC6lMlTuZjm4PU7+GxK/V+g15XwzzgpnDH6tsa6mvtd
ccSw3PfSTgEilgaNpEyPvgdS1rfKqlCguOPcI/tinuwQlnBgw9EGO3yqnoVKtfM/
Biba/mrfwtKsF89NdWz2nIFidtvRlzw7K2H1imdaPI+weTakJDnhpD2VGbKUNrFe
McUwAMag2om01o1Az9eGE2EetIWL9rupTGTHDbRVhrj4f9OhrvJlxELxRwVBg0gW
vreBnKXVtDjBUF/+XU/lHOuGqOm+dWdGqejT5THXEmdgRn0qTLTMRuHLLD5brB9V
eoM2TwH5Ksp1TJ+NJdswcGKIkIj4T3u/6kSLgXSargS6053gf5zO5Igcyf9a9MQs
waktabUBXyRZ1Fqi4Bn7fuHcXhyXVcotMVZNTdAGHjLgur1FC/JOJzmljawBDcP2
zcmJANJshzt3uMcgd52wTz8PsRqMtcaxZN2ex5evIuC61BqZrAA/AEZotYaofxvp
V1NgedhNKfUIJeIyTu4bO7psnVRkwEGSCtkFtnGY+U8RJZEuaJ1Ql9ZWL4o2RZUk
apwIyAuCN7q4vLajOXsX9858KM4/OyjZJlkhtQ+k/FUZPFStznAwImsSp3Q35Z4I
Hg7s8Y8r9kn6poIUtSjD+R+ZC1F1UD005C41+3kvvzpg0D1171XB761/lqASEuH2
wYFNcUjAqIDAoCKMY0CZR7E/upRrI74Rr329SastQLFKAvpRgpQbhFIhaBHHgIqC
1j10bsDUIiJ8dxWUXlFIJkwPdMHc/ZFRFiMXPBU7pngBBHX6RyZqZVY3ayTJ3rvB
B+KKSAS1zqt73xLSCF39ovscQWiShQ0Ln9wVflqSDGIvzBNcj7e8O6T0o65wo4JP
fzhW5XTCmdHnDyM4l8tYxn/oYh/crIfwVT4QaicJ/7howokL4/Bfk3gVOS3iYq6n
arnvHxhSZy6P9rWf0nR7zY+W/I61pkymLV/sYSt2Pdh6iGmGTrzeA2LoNhajFhNG
DoVU054O3wbBIixnw2InFuzdwzdXy7OTHL7VxdEZbswxCEPkBGvF4OCedYQaJTzF
WtEGJPa/a78vaW3OxIQUIISBYyPI/S9Jrz4vV+6hQLutpInmxF70IJdD2jJDhG4R
snlMjbTVGBWudSa3FjhXrk3GfNcBGl1O0MXYrEimE+sbr+Dzl0UhLVD7/kIKUUDk
qn9cm2WZELDjm03K9rUPrOVEYbQF2lL/Qip+FpjWbx7SmqJy4V0tZ10bTGrSD3Sr
yup0g2o+cL9ToaWY7u62NhWVdRdrI8EJDJGGyUZJ7U/wsC+9gv3/V8jq1+j0bthg
lJsQvnhwyrtx0IjYOicptZE1Z+F0P6qAmG//+g5r0xbWgxoQfMl6Ug9v1MjHu0Z0
7YOVfDaNVakFqiVhbePixCUUzOKWM2RjTtxA6U0DbEmGgmw1yx3NmC5iIxMXJAqE
vZW3sPxQTHd6SaLZmJUSVADOK22BNUzukURPEODgBD/e600COnmAjXua6nasK5rH
atQnTg0faaFxJHOauHcy9cjmw8egHD6K+chhW1Ml339jPZBTk7GrQADQkXMInXq5
K9eZC2ttDZHY289PD/iA2n6ncpJjvQI4P6kgS6mBSzcjXnjUbwWW/ANtH/Jxwl4W
+5nbsrl/aTD5SAiFThJQxvVNXX/KD/JPime2C/DgvPoEb4pws73ZwZL0CbMyQ10G
wVA5ONrHZbEd37XKiDG7X3MoGSTrqJFgcFYQppAwNh6KYacPSxEi8VO5Lyk04O3s
+mscPbOGN9jNUXKPKJ2exHCSw9ShDR3y3lstpVrZGskFiT/CaX9XJmMy4m2HuKbX
sSmtAcxUKt8/Q+Qf4D5wPAx7o7Ka49s9Rjm7KgQ2Vsmb8zs1jOWtpX9SF9BgIeDJ
mYhCyZ0Q7e+hgM+gaYlOeIUmCYL1J3VFM2VhggA8dxrrfEw0XZ09byZZ6S02Hu7k
8wxy0TlhfUWOYsacCU3dm0Cf3AeLXHsPx5ho8FjPoQMPJEt5S4VARaR50TibhNWZ
kfqGIhNKx0I6qaC5cuY918b6eq57c5rk0i8QbypPu9Z2D6RyecMrLgHaUe9CA0kE
Y4IhBXNliTxDBVI7wNnnHIFTp98E4uf2dB6C+3ckas+V9PeTA8vdJYJ1eN6XEtmA
G3f6EVM2co+jO3BdkVlLmOHIykgP4KT63XMNcZBjObi5tWttxilYqZOZEWMJVzbR
uIecnEHM9GO9nIHAODul7s93gq+qzFSys9srpOTeMYGK03w+czWSRCuZjn1fPLdc
0UZXNUWqG7AOxS3IAoR/uBLIciX+WBRMWpmpw6jyeEF3o9PLy87KyorDJ9FxUaR7
wSDeEhioQT9O4/2OYg25Xwd6Z+fAmU+cWiXMi8Flq41UqtatFk4yj8ccojHtvIyl
nxkSukV4VLG02AkPmIlRNX5b+Ac4MoErYU9x580S/MAva1cmnQaW29Uh8NXdKs4m
4MVXwouY1dpx7U6Tq5wpzkWE8xtqQeYzC9iJENh710cG+dkUlDYBu8zYBT6Cnscn
l3U9eDVvLOc1eTp+uzTrJV4t2jtD6X/eq2A4G5P4LwoCZ+nfSN5rOWda5fhJq1O6
rVSiuvZ7Ln6v5URsFWRS2RsXe9ya/uu35APelSWqp3Tco1ajh4S4jD6Jhq+EpZRv
GDpmwTGYR6vstDG3LzPSRXsj5oRnAlpntlKbTyExz8OrVjyi+4C8/AYR3a1lZg7T
/8kl2fPf6RqZ7NiVI7T2pmPGYLYsdaB6B2F/VFi6hkwsJeeLpaS96rA7DQRMqYD4
KXbNP5klrWv9Ubg0JrSlLZXR+92v4ED29excsMI4pzUY1dZteCQGEZYRI0il4V28
MqKhdRywaRjZmYvGNvQW8itxtZEIDNbS0V9K/nhfA3JQ0NvU1w8euBahES/+cLWi
B+h6TLd6NoLWHiXixe4bfeU7vwK1STs+nGEwdkd9anSwBl2O1Dlh6Xmq24dMTGdY
xLRcaCsFlvmOiuP0R+a/iOlXjxlzQnaljUkIEj1Q7tSd1KNxqPpazsmp8UWInpLj
6JFIcDf5621cf2KAnH7zxOyzrqry1zgdKhWgCE24JnV0CEAorBBAoUuawWSzUbTL
ygUmL3O/+brjYOflZtcxAnfHvXwnegO4gdUAb2azDgPsGGfdoA9pUoJ1HqNvYdwn
AFs1lv2dLHrn7C3O41qKdlQt6VAcmBiKA5EVJ4SnpjG0RRf6BinuPmXppQwOmtzd
uZ+00j8iisi2pVUq9t0Cp3OqmZ1vmWwuf8eDnYWo90tXhn53KQstf51zb6bKQXhy
QtCMIwCHMWVZ9dy8ZS3N8dsFJssy3NNaoBH2z2cWg7D3xbwYSrnYYWexfdc12wfJ
Eoo9F2Q9qvzNHVbWrxIycaUoEo1BckPizYBx0yXHxZGpHJcoTr0HLGRHhbwO1vB7
49zC2BcdqRr92pbSehy71xnWSKQ74nojtfGvegFwuCkcvq/li4JAPxSM6MHeFZiy
JMkCUq07YiI4Rh8k8qlr7oF4B7rfD5Rk+3WeTs05uKgjbiHQLgRP+JesvLrP5Dro
I42ii7EpGOFYw6TYavmlX0HS1o36qWnkdLiASDusd7PuHw3H7ntQ5CzGqa9rCDXx
1I19A8XHyDw4fyQfPpdaeYVk7oChkIkF+cyNVcv37T+1fjAyh2S+4xjEW7hmkz5V
rZMNn+YkApJ2rlRIZSS8ZRRk5CSUJ56AlgmVK1/0rp0ROqFaqYlCYBLar/hLW0OV
96JJHL3fz9rq6ng8kcUSK5gEFRPch4Lu8ciA4qb7/Qr3Cj6yyAkJU6L1kuUSi/ee
I4swwg72aiXdjU2VPjlAl4eTtkwJ0oJ7WgSUi7tYZSUlnlg0idaZfJNv7Mo/d9XP
dt99MEQTtvRflzxRCs6HzPyyeEmNVe8VsBS/YDW928bUSUiTwLQqQBzloZ4rhUWZ
vlcnd3OiBo6PKED7XjTl7x77MUBqGux/gaNQumyNt9r4UHmT1gg/HbaMaAD15oZ0
2Z41TZHA+oQ58iwVaDZ4c4wOxGVGyjgqBy0q5tfATT95TEUkSRX9l/q0l16XDy6r
K1ObTZiWzXKORhXGLsB4tAhNGsS0FMbN69HNWM8PEA8yt9NU2xqOzV+0Damf8FgE
m/XMmZYJCBfARixxGvRXoT/4s3O5J3TlOdjHPf7lFpx0ccCk0GT49rjgDficGcm0
6o79ZgamltZfUJRS7t3HKdHzIkqNfS1JR7gqmajquaa85yjwefiGOsDtqRCACpmU
+eX0TaNM9k3zVTt13V3pru5wMZBTvjrd0kxJbtLO5NZbyNXRbmDHMuwFuaG2KQC4
JSkUBkL5xG4Xphko7GHrkULabJeywAbTbFpjLqyyYM1U0gsJvQiUqZi4CTNWjbn2
UTYsT6KPqdRGX/SS0IPY3q/FukDgG/yUjGDCKM/P9IoAAg33PIQpwxNwJJh4aT0W
4iNqaBjPpgln4sBWwQ3rO7GimULhR9Hez8kV6NdIQTeu8CIR2Cu2I6SI4z62ba1A
1xaP0hq78i8Ptm55Aj7EsoUYRkI+5kvpcCRJgXWLI+lh3n7paHCFvWSK9IehnacK
0dfVO24Zo0MPE4fQq3K4PP2p8Ew2M9PQCfHos69Pic8A+3lnUt3DldTYPJ0PWNCt
9sHhurBRuaNJHDY6B6H+t6A3GMu5PjqfZnLWmriPEMbIOFgkA0+IBOvAYXISCetK
ZeCs8P9DEj0kQOTHxm4ISHKBmheIjfNxso87cZ44mtYSgq3iCxzIJy7nubMpCOcK
YHrANtx4vc0tbAKmrfSlCR05VcrbRcDlluAoTFnMOhULYClp2+mturQezSkvd9m5
Lu7qrJXQV2ZI4xFKj1lHhxkzlqcATfOONyuxgMz+2V6hy6/p5h3A7cGlW99yO7JQ
A9G4QlzUwu80n6n+9nEHSmgj9UV0xn8cHUBXzdpizFwhwZ+2WRFVqpuvkd/S3Ni3
mttzptQqEmGnG1sik8BYA1UFOP3fdXPl8YEeGVzOB9NfAeZ0VQY/Il9TBoEJofhN
HIplb+i07pyXud6sA9adOAxzS0Ew9C4PXhz5istzgSo+N3br1RAQf46DOaSr+mwN
lp5KFY1+EQ7FLxCVcsOS3YqcOsjstiuhQS8kClru318zH5Js06uAcgVBf8mIK/sI
OsJ/5WT+uBBL8h4ktsApfeagaPlYRSAQvYarlepY1qh7JIzI60GhuojZUW4gHAv+
/wZBDfwZt8HAkHkjSui4UTaK3UmklCVz63upX5ZNKfPE7Q8utM+hGY/HPkptkhB4
LZnr8KSpAgDWyAFt6U0bwbZfobw8USScs9iMPLFFeqAsCqyqAPu94kcyNGj25uiy
poF1BxhgyPDO9hvjayAiF/Mc8zkSwM56I6/ZltpghY5ea4owJnTOxZ/zawBmkvOK
lHg8Mmi25BJcEVrTvEL4Gaux3FUIA+/ewxEyRaDlq537J6etJAYVIRl+fkyFA8jr
3Bs2xvHYaRrsl2LleXqoh3VoFNV+Bsh4MjxaSFdHKSb2fKTcaf1DnOU/qcGgkdNu
RQxToWZiEHxqXMdm+nqCJxUYCeSXrVzYzs0KhCdA9wCx8u5CJPGsEloLK6JkE+ee
t2DJoIJyJtMYSMxaYWbeyT/PPijYBlfWq30RWSBjhpFQB9isOy3PJa/Cko/mJtb4
0rTjc8v3AME4lBq/1z6EuLM85AcNIheE8QOMZPTr3I5Vs1MXKq7ZlirrjP2dyOQQ
yVIYjk0HOivGbsaaCEIj3lZLhpQHp8BUd+CCuaxl7kIaOHznFhi9iHOUfngh+05N
e2W1T8eqNVVdTXBkMvrxAXbTKKIdoOnLERhLfIBecwhc1LGLwoIcNLmttuZK/D1N
YY5O7XRjOu53UFyj38GAdICjjlwu+4FpQx+1WNNv7cgdhPQb3sALZ+gqWOrMydbl
rL+cK/jIss+jZu0QfXmOkP29MxXcKqzKevjXM19bvcQQVfHralBDT/I43quhuDgr
WfSrwxBYVhUs/pt6/6URuVOq6MzpqkqyfTxI0PIyK6s6bNUIvQZrLuBHVgcWcH62
vh7lHrD4GtAQBUlYKutBh9aBbcLQV3rRHLDnS3eu39oNHMLGY5RiUyB1zcuKsv69
mF+M/apkZlt3nfanLK12cEipdjg7vM0AICW1OO1qsTjYSRbOBcDWszk5x5UtH8Je
cwNKEbzHJB5FNGcMMJ7FCG/okaVBuoLafCle5GOq0Mb00iR+JI/cA+TWOVzfhewq
hhOYC8rVFgV8vbwXIYfS7GA1SZENqFnkpP0ip3+ppY90Y4ZtFgXjIXgWXsKQCJys
iFn8MLDtSb1uSt/c08nXSLBRSAtEpk8HkqWUJMktVxvVYwLNOi836ox1nOZlAkp3
7EMeupA+d+D61epC4OanxAL6D09skopCSYTBQWAkH23AEUb6NJ37gIA4CnuSh56U
4dA5DD99lxdxykmlEdYCSiBXuxI4kUlgIQl9qB+Wv5TBEu/BO48mGrXCARQi0jT/
EbzmGiqlmSYwT1uG5wcdHr6Akk2Td6aJx3MhVQBPtDvfYOXuwrZNQG5Bx/HdF9QJ
8WDHHIfYmTa1nrma5r6+Hcy/5JPfqj7J59OVrFEXo56928sXVE+Ag9rUbDXUHCPa
6gBi4CL/VSHFfoPRHu44eSlyVCadGeUZYGFJG7kKXzpq46OXanRqeCesc7HdUACt
Knt9T9z1NBAxKr1bfjDpF40fs9LPeUiMIYIY6bKGICN+ED6dwsy2pRI3sKYZCyqk
gXm1U/HcsTnEEUnLiB2N87hzhtEyEQWxPnZbWyN2URzyOxfmTZiLKtLazcrqttqp
Hj1xI63g8q8jJVVQcb+0mpfB06q2HbWQ5TfDxuOqdRRdMA82kHgOrjauI9G7nPli
K4KbKL0+/00tl6+wmuGMGJk16tfDVuM5F8AHk42qQhw097Hv+sTrI1lHv+AXAxFU
JPLF1I/qzBAZedIJB0cuWW9LkRIgWOtJfYgHtiP92TI2a/GSth9gqv34WaDsYmLG
rB5iSUc7tJKZJDfkMKeqvYCqBumv7xxtjEXAkRBTgI1N3poTrd2bswGsGhaDZX9/
kizhfSAGH8aKC7DuX2lJGp03ah72nf8fASYWWXW9rX38u6nI+PQoJ5ffwXTPqrVR
3hLwkRpaQTftnwpAV9I44g8Snzn/hv2NUuYLQt54aa/ztKO4Rk7OWw0HE6AyUrvJ
57K0qGdNjXu9b2iYfW77jofYb5Fg908MkcXcVj4U9YRY5Ml3R+cno9/lPhzDilEx
6KLT7ksucsfTE4ATEeHhTRhJ5C2ER9NvqkfVPNsjmpBUbcevaklzu4skd6s4M3BI
rwaonow0lh/6H5Lz/8y04wubDKgZxP2LgAoK7PrC/dp9eY4UAuH181j4bbm7q+F7
EB4TCJrAvGrtfcno9YZg0DtP+0d1rcvXvG5y6UCbpAo69WPRm2PZxIP5no11tJxR
y4HA5qTzMk0DfNAggEv+s7cWSVy9QwXUgStemAQ0f/gxASaS72djuXSP0UYpmmlG
nYuKqef8M9PM3sdaK7rZ+vijpWEUBYkUYeczcgcc1hAgfh16hT8IIU9Siq03l7o4
mjz31I//Pla3AebIq/tlzWiVNbLelp4SnwTVdO224hFH7j9hMvXPKCjleWtF6mXO
8Rr6S48fLkTI3nIz5EhDxH/gYyfgOxq+UQCTftQAaNKyGqaH7SyL9RizVT/rlvPD
IfrxtMlkQiJkSBOSGZv/nUYAZjf5jU7LHtPM9ME7oe6TwksZyamX1f6J2FRaj0kH
ZlETVJ209Y0ulwZX1Vlgk8bWblE+qQFnrPdxtcFOIxlm81cQrFPvZ/V1Lw8FdAN3
7c/LNjZmZzmEBKHAGDrhqYdvekK5nP6KKZWP3o+u/blpoCrb7p1m6muP3Ck7Syz1
dKsfDVM+C0fuqgvXDS8n8kqrOyi9JIHekXtaRvGStlIHU6uDu0CoLVcgdrTk9pim
SlAOiRPRoL5dKGEwWI22ABYU4sj29zEgW87Uv4vObSixT9G1zdJ1OXMoHqLjZYlD
PNndAu5pRfFRc9bPLB8QgunnBZ8mJwflXt6pgdxtpRTnPjACOy8CUzEL/jwRIk8E
qHc1sjEnQR+VBkrQjvvvba8u8/u93/YSgzJ3AuDSKgeCUZAxWqbZBnoMH2/RvAnh
Q7f2y66QDcQBqzuPYz6rBDI7yQZm1oJXmQ/Inr+vmLox7F0EX0vrSsK9ovy6p+UZ
+jrZayh19w9mQGU+tc9GrYRQZjosKIwc6+0wAZmBb6baHFQ2OyZxqodBb9GlbBWn
SZO9uqExHvn9Gt7kF6w6cGwUMMBIHn+zkszOkLQPzFgBeW6rsnYvMH3HB1BExkW7
SentgWr0i75dQWfHA+LKZcgYIOabkv0jfoJFjcqJN8ghXk3JBJL8/BdM5AMYAGPb
IAUlXZPZ3F3fMxi5JLJqlhCDV2uz2oUrhsjQHsJg4iLtw9CVO30X9nWWxx5O4Lwn
ux65E7JkqgJxaDdN0BW7oRLkjkZOSWF8KURPLdpni0CaPfFLkjd95y81Fv2pt8o6
R4WwewuzKDvpG2Rzuv5wef88JCfuuQKspJokbeHxmI8lMVzuTYP5QzEsDbErmwPk
H2jPTQvMUBEXvA+XtA+dyo0TPrhU/OAIPqobaCFWW+badvDMnkc+vMl58WGSsnxR
/y73t5R4/oQ3E6pPDGRZzSXaS/6UywYg8/dTix+YvmEJEi1yQ9tb/IjMQq5KJ2px
EgC1m11fofsBPCk7g0vGapFBrDvSM43ylqwutG6X4DCr3Zsb0MVUjt3DfgykpsOD
Tv9mZIeakzGts63Zp00EBte1oQwIl4Av4eq8jZFAMo06CD8ABJbsSbE6dYXulg7h
4Xtywu/gaG9LPJTO/4UQLmhXOncleV6LXJrIr0mvmFd/FPSW1rxqXuEkUvyFilpM
rgVlQtMNWXMA4lvZPJN8er42W/rRXcqgVLB/r3LHzkulAME8n/CltMXFQaq48Ljl
NGSEDUnrZrWqfAwfETB2Vor9I4C3vt17o8l3BmIDzvp3fCi++IxPXPtq6fwWjFqH
FAvItZYPKJyo2cL8VaPyhEgnC7pmKGb0eB/b6hMvtuoAhkXo/Bir0u6SiuiPgzSG
5lXkijo8ZJwGnnicuFOXBBGlrw054tfWgJW8g768tU/xEE7Dr1PYt5pcyBwHETe6
Ro+cCOOnXHTS+8oucSm4exw+lMBKBTA6NR3b+ycVqxnl4/dmACthS6hzgpjd2p2Q
Q/rlaNqYwNSHgF2aZCs7Mic/wxRi5VmvOcFplcLd1afvD8sDgeCDxSWGTLGqUlJv
Yp1EL7LET1NLlqxTjVfmVb5N6n9mgwPe4XuXC9D6NLNSYTPKzk6yWAoZAjvKFY7F
cLzeVxBjFSFg9DMzubRZgsFPYpwjN++sqABTwxGq0+8YduJ7q/rjb4goScc+WTIG
26R1OjPqKUAaB0ox75KD1RgVwKJ5nkYMSSKXFBYnnKwF6AgXoYFPiYTcI/LXE4uQ
ttVrbwUTpfTfJZRh8uHvKYX9jPV6/EGhx9e+XgGGT8VC9lCR61daUhAiD49Jzkgg
a6oxqVqY6etPk2kt5hDADRTquq5EXLNupYRajrCx+bzC39V+fdulnxJBbNp85f0c
FyA4el+Qntqwu1UJdy4TQ7vnaf49vmPvu+A+1m5OKUsHzEcbzRdbNuPGi4Hiz3F/
8FkLTCvi1rvc+/P4ftn1IEmVPJmP7gQoT4KOOBtU6LX7ozL7RD5GnMVug+NTalhx
uZjVbtHSzs3Y1k7iF3Z2Wetp7KqvowDOkZ001uWr5ngxhT+5Sf2Dhq1KgHHMIffw
t+lrqnfA2QvS0wLz+2Hgq+zni+6zDMFM+gh0x/zbVtvNXPafqIC791f6BeBI3l3b
ZWdLKZddU3J5Qs+ZHYHKxKByfIBnn3yyzbup6Ohs9Ye/zCwPVQInbINHrnhJMDKY
YATV+5l7ggbVWMkpbEGZ2wVNhb5kLiX9Tb6YMxYUXwSjCgxCH8JPoPQKXaUAjF3p
aGgwNkCj54XzaQoE4V7nfZOhQ/u4PW53z33f/umx6mlx+FDukkm1vR+YjVirCP2U
7vYUOMNK6rNIMplCn36yL/4ivE1ER+ajzF4MUpmigTFpU5j/QhJKBGhZ6KUf1goZ
t861CkqqDlw7YLSSIkjNOjE2/hamfPUmYS7Ne1tii7rVNkY/vGFJXHBv88mnfuJA
GO0yCaYEMz3InSYSCEgsbcstEtovN5RQibmLGbDrtld3zsVR0Q1mLdNgQaUeqv9J
tfUCgsRVj9uFqbbJmHG8Xj/FShMoDhpRJWqOU/DEikK7eGsZ7gBW4UOPR5+Wk2+a
GfgTEna1ifVaJ0mmcDMHAUi94xQKyoKrZ0oSHt9ug37aNqkizg9537/As7nNaUqF
bDuYM8Qa8b9283dd4SBhL3V+82S60eXLcFVBp3FOfv3WzW4DU/5uAuzu3tup7Fmy
N4Kf4ZGyPNZFCASaAGvS99SdnH7xK2RO+8KN/ouMRQgPG3yEbu1iM6i3YI33opw7
9MSS6lF7ItroRrpb9g8bRkAeUD6UFp7KztG59+f8ASV4ZQBJd7foanJjEVhY/9W9
tV+oTV5wK4OCQzg53+3DUOgRF1+jV+LBNS4FtFRYuDv94NkLrYAJjVQAGaAAigTg
2L1f7YkZCNxRfZkjA3YjuLT1ZHkMF9VELvvqGz+uarZ4eP4a8ui9MlBPJ6OqtPL5
2zUcSpLCAMfs8lutTZ4IH6iHVfFrSAOZ4aXQWQG98qjOqq0kYk66v4aGWQ2EMb6I
odnKaHZ4m7hxonup7Zpw1/ElJCwo4ocrd3AefYbK6KvBviPPJ5DiBw1BWmS1J/5K
0wkpX1zpsMiTakeush0OGJ37bdFUANE93DV001JGpnfs9P+Ui53f5pDjEM1j1z1B
4Cmuf/BIXixlnqbDbFvAcy9A8tmvR68WDv4FV+73iDw=
`protect END_PROTECTED
