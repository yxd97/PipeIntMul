`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pjgCzGNfYxJWmEWBnVzUiw2Rp52efeKBo9Vb23A98u4Si8hsj5vi89uobLpMnjbI
Ro/UQJdGw7RQqxIZLmREVQnb+xiHFdjiiLh+toSaFDrkKovWI4Y3UBCtNoUw7KaK
Vamt8Sm1B2r0qmfwY4ofvY3+/ReNkgr1Q1NEF3in4iDi6rjJhBfddDa+Iz8LT5Kz
SmsyHML0ojeg7cMXxot4uirO408ylc3kuNQunxCB9DfOjUP0cGUWtzUA7kZ6GuGb
AQ6SJ2eWtk81LrP1xOuexO5OYvi6+kQRamoEireVefs=
`protect END_PROTECTED
