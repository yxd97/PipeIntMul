`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6fIleVzDCPdx/VkNd5lf+DbJNd6FYmo/YqvmQYGNEBgAWX13UZLoUlJgXsIA/eE
Mqau84km1RThQem4kAYqH2BRYuZxqJn/OGsB1lRxwlIVnNQ+RcZ9rHQBvnnAO8Li
HezKNju5OKJu3gLtq/nbhQVgIhRiXFAf67i+50I615jB5YAlHtbgrvXHKKYlGiL3
bhdwI+v0Qd1FOkz0wVUXeZ+JoIYaRS6FBB2TmYt9B7CbhsuRZ6+ngpbF4OlRgW1/
K2ys0GBAe6zHPZpfi0FBUv63KuBjMbDHGb/Jz/REqil3JVlbuSLysF4VmvWjLpQL
eTkha6eXY8VvV7AXQtiG6Q8ZwPw4cf+HpeBHeF/ou+AHggqD3N0Pc3kmigtAUcCN
C8oL4bYpRMlcNfpBu5QT/qOmmmBoEnFjFd2TtxGohmAfDgYKD94ikEmLIoIHtIVA
e8HB/pOr/f2lAd5CPv14+DcbLLrTsZIv2L4PG1xqNlMWbIyN//BcDBk1WCX6jwS6
Hc4JOQG5DrYHUxB8HZpLo7cWdMmWbAYWYYEOsYOZzfP8SuTDlR9U1h2ZfIXhf/TK
LxuO3YvbI3CHCONAqrOhy9gvQK2DEryyayvJg6BCN2k=
`protect END_PROTECTED
