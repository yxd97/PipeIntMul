`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hxM5r7ftPNP/Gxj71SE0Og8+0WjjgdyGcZqL/ICFqb6WrhtF+i78yj0GdGj4PRja
a+bjy0RuNP053hROMKxddQ2+angtzktAMdgHqLROwCnkHvpKyM8JGZpi/glYua+4
MxOMqz/R/DqJyLgDAOiP5lOQQKT8WQhsuSWW/JMbaCCYw3r3wFeTRyb4fz+kk/tl
OGF4XcsyUN44YT87BQ6AX6us1pvRIh+jWIt81dsBUunm//vBvgkR1c+ADhTvGu6O
9lLPnTp1QThBnpXeP1J4VyZrg/ftWnE6xJdMeVUerHoECMZDVtr/FdCuK87j+9h6
DBkdhZfolBNLZ6FqUmaisQq4F4V7EKAAmCKS11slXFYmuBy5yf6hkIbfOhngQNqU
kxhbZFqp9RuOsrGvctc4GZXHLcXLkMkz4JSrF17y6NB7k3Jt0pjCC9k4BQdxX0U1
5+yoJTK6EpvDqU2gXfYSADbwA7p/UueIDrMyFtT5DE3Zb8DBLs4ogU5hhbjjA4x6
`protect END_PROTECTED
