`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IvpWxC2gjxNUhF71lLjAI8nUOlVQoBVLu9sx8wvlhk6eTTzkE5HyelEik/jtDWqm
SYLxRLXeTFqUxRDNxN7gPZpCwAopeyvPbfz29RJCMWLiVoMi8pCT3/ekUSPD/znp
okaoo8BQMAlp0jv2z5xveR6E4yFF/6JH2r5I114oea3ZK1Vh7gAgdPdM9StvAvLF
pHxZ0xS2i4Sz7jWcewGa2Htpzd0MpPd8Xajs7K6OE/eIoBv4roUo6agVxF/X8B1f
a4BRwGCSY2mSLIdK00sq0dTY3k/hXizpsykU1vp6ZwFe91Wi9VocVCuNklIufDof
l5PgD5SL9eglbWK79WAbL634IBL0Pg6TBJX4m1E2F6b/PO2DmQetB79LD5r1P2Xf
2ZsTIc/FJDCOMrucakoJI8iVM1soB6oPEC0+dFh06dJN74BYIRojocinZAlIAbPH
EXHWG6TNcCxNMdPmC/mM9TGoA9ncxrFfTefT7X26Ysq06/otIXalK60WttSN/ZFb
UUlPbrSbLQmQwxAHQTLP28Tzc5Chcs2U6FKDLJ+yYR8JfQQ5MIGP85g6MAWa9E2R
`protect END_PROTECTED
