`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGkYgum9I+Rpr2waTLYxwJp3/7r62vD/nFjEFoYXaI+CNgxQubmNDYULNB2tTVKe
R4pN/rmXX7vx78OZ2OztZhhaxL0zGE1r9jg4kOC3P2XHdgtGTxaF+ilzOsH1Wibe
wDdQbW0YgxB572zBlhdYdX3ZlpUAn/0fiz/DIyhWBqiwWsHSD23Nk0TEO8KkimMU
WdYzGwk7Kw0OXnj6hmrFJqVlvVKtrkuKMEDSdZp1RlJsokYjrsb1I44miwRBns29
/5cHZ2QtG8EJ1/eRPJVikg==
`protect END_PROTECTED
