`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lXhyEXnmGTWnWNEueb8GtjQb670QgiKfAmang8gPafZqXs6lTGOBgCHRrIYZ6Ze+
IzY9MhhxtnQDW1d2GHThnh/UtG25denPsjfsMAb7bqbjm9yefipmrm27MR6wmVOg
1iAJq3Mh6+zNASVJAJqHvpTy4A/iBvytsxsae4FG/LPD569QMQwwkSyJWQjPtxEp
yUKhFsoxyWhslORte0FGr0VNkl06DWJ7BVzCKSE2Sm3kkgeHu28e9hjLnqfikFYV
MTqgeYzLLpHhcHmPfwVfx3e2LRvO0a8cVxGzNjYRThk2DUhcxgZ+TKQxq2Gg93Fg
DSUknGsfR4c4+NO3oV7+8EhBgPOi9mWPUf90FLwQ9pE9SqPFknJwWmtjGICGo3EB
erkxoIuUlxAFMvpjDsCtOdXWJP0xj5oxBhdDZ/o+BzrwGwf9XL+hryTDZWLMce6C
w7sFmnRwJfcZgoEBIx7UyCyFt6CHU3vhBqk++31YDkmD0hOPaasU+fQpLCawzRM6
jgso/5vljOHLGVlPoNK7SAVrh6JvgicpAV+FqvsyPQbid4L7+cpw325tr9Cj9/7s
kjDSPpPl3ELfPVdWKTc0aU4xO6WDOXy/+5onqZ2dbEWsygnaMIrvNCwaz9c5KrX2
pZnM3eFaIxHwDXoBLI9yiUB+e62YBD9bUgTbnxAd7OaM5pSHdKJ6hHeD5d0FYDkJ
u6hpzs5p34Uc57IUCEQjMz2E2/yOk9CElRxi1bl0o3xfXGiNzMEzbPqte7G/KQHy
a5t0/D0OhOIPa32bAWwvSMMQVod+EIxZuBxiIhC8keDgb1N5WvrHRZowxgVllSuD
9kOL1uvZrNzoFhixVMXTisuoylKonpdlIT8JGdmdH6Iyzs1SS4+Bq1VEBHTIMCwl
hnSXGoDUmBrpBrMQt0qAJuPemXE+SNO4o9mtiXsiOOD1HqhNSdSt3Z9kTkL6C9aL
gh/AplEhm1w5jntO+yPN/CyOJM3lHuN5TI2ufMSI1pOcRZ3pG6/6oJaWo4cNM3Cc
17Z+qYlVz6YxR6zAZV9Lvd56du0yb8TiOMxOL5Huo2j0wVAsATXeaYbRlm593/xB
Yv3wiNNwbH3aAOgtxl+waUoUM5yRVO8eu/Ot2/FDGpyc1G+Xm0rPjtFQk6kK1f7b
qAUuXMEqjZ5gdqU3enVRUCsIpcFIDsLDQCmi/Z74V2WCxMXNnqrznhw4ONSKpdW3
G2QtJ68ucfv5Ucro+b0Z27UBDaONWblPkeic5cxHVZmrfXGg/BwxFOE7ijTLe+XX
oqgNyS5XE4V5y3Ls3Q+xnNYyquEKVi19tcMlIslNUeuACEwjsKClcAZxuMf5M/OO
hCjIjxUR7GFPA1V5AADerli/a+805BkA38JndNwkaFJxSmWHGVwosEiSoDibVgqW
GF4517Td0wAEp5lNscerVA==
`protect END_PROTECTED
