`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tUcQwnkLRNdbK67kao5u+5m1VLxIRQhJ1ZnXEmOEybN8wlcz2gcUZYBci4kJEj/Z
Sghp2lWFAIsHvQ3/fPu9Ow58MWZfJkDbKgciC7epsMPbgU7I+x2SbRumaTmPdGTS
WkeelqqvP0blJ1mYi7GBXxF9Yi49iC7KD5K4AZK7Lo09by1kSdyB/yyZXAy/WItX
FruMqJAlCHofVJGD0jipv1r2FvQzR0vu9MFqMWmEOBTBj+gPKziQ7KqkhRPm2w3y
rB7kX41dLQXeaRYbVy5QWgxKUCXFn06XhoJi9RL6xhwKWRA0RNvsfJpnxPz3zjjx
d1mlxWEASZqSwu4y69sMHzaLNy/6Nxn/UxwFGYDximcBF7degzEFXT+LjVfCBuvH
dFuuhlwHLMiF/NZPytJj2HPs71tZTDWwmqVByX4Nk1l9Q+5DC4YMZNjHRv6Q00pt
ltUdZhhrH1sHLFsehQFH6OkOPaNWAxszAs0/9VnRPDeUIGiaAVSWDksucRq0JCF5
jk2qtSRbGl7ljeTTuyQInyppOej4eZbE/smqKUINoQdLaFkmho0AfIjc7UqHbADs
GsI+JQa8KCM/eh7+4rRWQbkqvkVHr32fTKQA0/2NbWC1DkyJVfK42sCAcAJwxLA6
FyB0xLPoOBWavQ8096GHHH8NhDk8ymrHiZwDm90wxitnpR+xtbxh3qf69YS8wZcB
y39O4FkeesEcvVz7/v1f3NRw3RctyBqDqqIhf3PlFAUxSb8L4a1fsfXWuytu+APw
X9USl+1M68LbF4BwxEmiIgD5S5zixbf42Y6YuNB6CPh/R6mKCx12mMEqN8zwsd4U
Y9pzsdIq8kI+5xVR1RrYo9Qy/dKy/JJ/IHbIdMYCVuY=
`protect END_PROTECTED
