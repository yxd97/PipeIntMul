`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ie5MKp1bpcyju3Tnq/nKrZgEdkzY5xNXNRs7H1cVNHkuBsIFzap9Nb4m1A2klg0W
NLGBwTdKjiTwhEYdUgFDXFvu3HHd0MpXqbT9qFIpIdv2Kh4Eo5OYWXJYYH3DQxW3
Lsy6XG/QF1q5Q5o0+CZmEBRzezQYcHuMQqZv3GL2G2LwpX0H6gBNZ9bZpXlO9xsH
dG1o2TYVCbB1lMaPqJqFVa7Qq40Kst7MFpIFJDJ1BtUjlZ56RKBm7Nk+TuxCjMp5
zmWwSeOdk7/TGBATLmH5CGT+qpgtZWmP37V70sqK4tE=
`protect END_PROTECTED
