`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TpopopNQ0fMsGx8OpLvA3PzZfo5ELE26c4cadmHQpOlb5TMuDzSxOBY0chLncwWp
m+TTNHPAE32Pnt/Gf13jY4TF75bSvJ0qUuqi4HNJEKTBcfJT4Z0e6J2vSZS1He1C
bkRdApmXxkep107m+Urpzj5Ru5308lze6JxIJIibrgshc0mAryintlP5j3wlagis
P0NTquNAjovYb+jSVFc/C/DsaOLwpA6BPQV5bGIawetcOScnuokd/feFYDBJZC5Q
qncU30sl3Qk5WMlAaXKNLJ31L9+sDTZVC1F+y0eFwogC0C/1BjRVDQNQ8hm0FBvP
PbPofMP83/lLLMlDoy6uC5RxvPy6YsESPIDW+BJwEU1gQ6FrXUKWzBgSXNHSuMM8
4a0sIxtwHeP+h2je7vMf0x52DZOIuTjrxhcndgsy5AUVSzZszIMmInIUtefAkYud
W2ffvNzHhcWbYxkkpDQ6u0bghNgvDYT40b/RQNuqUnrm1fqRDKuaxIc/lE+GKMxJ
zeSGviVcN4MsPj3sKYSxySHC8SWhlmxSpoJ0JTPw//NU3FA0+RRBE452idq1JMxc
B28SdQ75gY6Xego5jPIsWRokUjK3EgMh3EAekfZS+DfoTBOe23RvKpGusICOmKLx
XW37MnJpX6L6vsndPSv7AnL0gO66KZXOITErIg1dViq/grPlqUbSNelWQTZ1G/AT
pe6aHBV4SBeVZMZByFBtU8fk5vPOI9UO+cc8DD01yco79QocmvyFYHz6mCQorryy
9HgFteBiC83Gp4s8lJEwt9o3BBYtXOg2NJ9UA4IhpnUKERj39rvf5wpZ0kbISvmp
EBhJzuyxRjIcJQG4tExq27AHeARXwScVy7nOdaCFzzjK3UI25u8QolG4/D5kr5fv
4VA/h58w9Zj1uNA3MJ6kiehCzsekRez4uy6J/WZAWrmPZDZMO9j+oL8JKGR5u42L
i6mEiyIzVxBIblpTq2qUievLMplz5XU7jZc7+87yYSGHWN0w9GosMf+BE9lJtR/r
fJWv7I+wcyc4BBhumnxL1uGe4a0RFsllga9W892blj0r61W5aBkTRSBdRYa0EOg3
bQoxfgwUS0+AeA3n+rcGFmgaPRz5Z4Q/RdUU6nrJWpWRDsdhYiHZ2KF699NXtxx4
G3aLCuSlxt3OTXb+y0S9zTmoW6PaZ0FIonaJAMVSMdwoFfVa8dPWJL2J8zR/UCYk
hSK8Se3ecKvVqS6TK9DDvOcqxZvc9MbnsmCPkO74T/aGovFr32PkeTkiijtuunnj
4UxLVZ7a3FhZ8L/453YmTqrLRwt84OeeHYN4Yn5CbPiWJGNi5OnPoGOR4rzTBgGe
8pyjyfr4FHgWwZ8brRrlib39Karkozo7nhonFB5syNt0BfljoLjtx0OfMrJmix8L
ILfQL9Hi62IVWyGtmD3DnK0r98TJet6rDYKLTouY1vvUm/6P9Y2NaHoUPR6dAnZi
8fayh7VnO5fjKxYs7jLEnwDysdSkNpecWFUm6uY1nDsYYIIBuVjIcDErd5y53r6f
fsCjmswe7Obq3yySz9VoNXH0U0Cl8OiTUaxC1VarmoytFAa7VLYytnuFB/176shl
mtWujviB0w7iHH0t3oig3XiyLHX1ncz5WKENXs1vUhjgVAEr58J32BQbpUJbdO4n
opPc1pyMlzK3SyFSEEZbclmiOPT6QXUJSjGo3WK0P1Nr2H62m+Vv7JpzwYzMxIN1
jJxqxczcZwUswo1nu/VCPxcaITYVizgCdrQfFrGmWbxAA+BLMNkz1N+5Wii+2tba
NzyOK2CwpxJMOsoyoaJPY0Bk4y8A5CfP0Y06oiDhRSpjVJX8j+B6c+L9aTGRlEA5
6XmvczrMfpgvTDUv/GZu62gBgp1G/eN+aXP3Ukt5ODDKFKZe1ch+1gag0sAHBwe/
LPnBcPsyCR2Id/11QU0XwYrk82TAHZoX3+jL4A16+jG/zYyCQsi/3nP9x7Fqn+pD
xkxsOCTGA2jIjIevcgj3w23Q15Xb6nPgqr8Ywihh91zLNroFTBLxBmr0STcQrpQW
b4ffVdg2bNrlV1Xt7iib4lzDd2ec3L9kd6hFYjT7OR7c7lm5kvRwLJ8xaZeU/OmX
jpOj/JGjhXE6U8nbqKBB1tt1HHZG6CTcdrFme+JOwv3hScafAAwrze/yM2whX/MH
ULu3sti4oV/M3hWLEQWdur4qBCdoUDgIei32/xfs3SbMsUtj7zXLGTwxID57RS0o
Eq4dwfjvxDTRsiIZjiCm4rszoAhFRKaEAqdgLC+eD4kHp2zJaDSEZZzmyEf97BRV
zRjfBVxASCU9zEop/djV2AvmSdH0/tvy6C+pRX81a2Be0UrVe3KzRM3N9zE1wsTV
E1HGm00Iryh2tP8GuPAjuFj6fAwo8zSpPSylHfqSKlCFNE8eUw9KW7BJqB935GIe
Xijk2j585vqJY2dD69lClWsnzQujSNU/uuut3SAhn9GWiJzBtQDsf0RYBVfEJIBy
Zl9c17EC3iVFWjcPLsfCPwseFI8EVr5i+w/Igv53oN5qS82zKZjC0AKxVFZTrI+A
lED7AD0QPmauxxlMUDy6g1y2vEKCsHstmhiL6V6TPu5SfbQMMvvAqc/1W7DlYZhC
/gmInQA/GMHWp4lizSORKEei95qKADG0KuxSGk/fLbVQVrkknfLXusOJPhOSSm+4
JJBweRg2TpBUmMPY3O9zegU5T1c4nFSnXdHmaqbASjhvlms4w0n4OM6VSdZ6UZFJ
Op+LNR/ksYI2kDVIVf+RG9F5t30h+DYtCTJ9BIXSWw5iyYZshkuF2aKkQYuADvDh
R+YmKA8XJoVMxJrq0XuX5usiZEibM3ak7qe72CzzQfynMhAz9X3t8pkEpuOUkpVO
vyasM7co/3zn+NTWgmKJAcCzD9bPCCAE5ly4HUZCq+IqQV2a3vhZRrHoK3yTp3M0
IkZeqIrQD8f4qsm+dFuMfZPcHAbqk9P7TgZFzJfgQ8v1KIMVGsUuNsABz4DhmcmB
wfqARGT2JnuyjsC29BN1wq6TvYf+mzgpZWM/XKhoTblTlqcCjYUOlT1avb6Wo+0e
+ViyjG+OfoScZU6x8G+GjI7ZzP12NBg0MtWicwNrdUX2r1LLlaKzAFj9zQH+NBgn
ixOsQvsLYnYWDA03/Dy3E9zKV6DG4/1Z2ZSSEZsID5dcFMVp6tO7uyEVSQUcFR2q
09DVTFpGKJrCN0IW1WSXMg3BZXSrMbRffnPXZ0gDvDguotYZMUuU8ehhryz6muE1
Q0sy84eC1FCEYfqYT6bW9JU+7Y6BSZXBPMZs3H7E3+UZZNy6/IK8TM5nW1/udzI8
vWVtsM9TZyacQtsePYmjOeqeG1aoOSvHoD7RvlQ4ZWFyCqqWw82bPslsk31425qi
rsRfMMv+383zdMrgL1L286lEO+lPoZNdRqM3mgY1O7BI92VrjtM4wcb4oB8d0Rhh
Mefe4dn4WZFCgOpRRoY/uxO3UA9Zvg+LjV/rT38Ec0XeJoCFsrHhXUH97tIcXjqY
TaUtWmVx/o7AMrLmxOlP6i20TdmyRL8ti6Ys/9LgjKxeZVkddhyO4Lju31zr6Wps
PPvI2VoL83bc7XjQO73ORGm8weShgxY6djAtc7vfnGeajL8TAolsVhLCmKsmDu1O
vSfugLGsdlVKSawmHn+qh5P5/A3GPPnlNT6IS3kG8rfaQKkjbQGVc9DjpPBDkGza
wU/dJtXd12AL2+luvdNHgp6egZc8+29jRn0Ovm850KyTFA6h8YPoCyYCC5z6tvKq
eJuiFlAV5scRFbOL2WLoVwQ9hi37v2ZgEJHGXbHSF7HDFlRzaqmiSO/kxa1u2ZV0
nWqSL8nd3qR9B1FJSP0xGvnJ41Y5CtkTY02oujedCJhmNXMT0fTcyWXGNCbF51pQ
hJWpsuCJb1ZVWjzfIn+DuD8hhpe14EPWqKDIHOZHwRR3pfqlW3Rc+P55DK0kEFw3
uSD9YawSyTTlLXljXO9stKAuCOG0nP8KiM1KldQmEk5ZJnjod36biC8HwF0rXFIf
orUm8DCSjCfgrgRD6TfMg5Ft/lmxgFk2WJ/jhvkUL2E5ZHCSbCRq1GaIe3qj//1N
h+aBVxfHKIP6TZ891nY+ocKSCGL2KiBqnr+9dCrG+hjOX0a2eC/LEZGwbKeuStNh
TmlI94nO+2NCwCuocfCQ9pOuRkUbbDOibkRaPKYbj5WUCaWTiyS4Mwh013WwVznA
ZvY7ekXambPdO5SPm84pW1AgrVfv80hDNfRbadTId24oiP5Nri1dzVDXm+z1jyNR
OdqUOn4uRehq2P5gkheKxXGuzbBQ+bU3KqA8iRp+zglYjd4tHVPgOxxvVUWCadms
ALAaO1RmODGnDMfaNncyzJs/kKKTDaQkyW8g8yEWUAugk5IneRRjf6AQLm8niMwv
YQ/apnLRftP72BJ+wOJIilHPzLU3yf83TpG3iZprNB2azobVmCp9Gcem1uo/4lGc
g67M6riUVcOEtcfT/ohfrLtgxmeMnMJSN7Fjv3mQ0SFpGRg54vFy0P8lPMq2vQP+
iznyyWISRfN1rk2T4OxfajYKeBfuFLQZFBTwP3M4kw40DGLawrhwH2PBg/MmUl1a
g4f9UFkhyf4dtWGPp2d/E2VhcPM2E6QSNMYOEUug2WtuvYmDih1ladDIyQ4crCvQ
Ht+EQMR9TxVtaioqA1pfHcOm6s/Tu0fp5dPG3EK0cIrq7tkEuy55GgBu4+CVQmN2
00XDfvXRPaxB5p1LEQoWk+aA87ZmXlwq/wPeG4Glz2FBlIfhjzhXf1oQ0BCva/FC
uoLkFKR6s1txWXsXgI22H+80stVSlSb2HyIPsoZpGlMFN28fQVNVK/36eMEPJbOH
rxkNiCQxDOhxOJ/nLVG8+cAjcibzhDIYVJnITW9IBM+EOCRIg4yrRrwmYrTFTu2g
XZmLvkx2qH0e1MKal50hpW3tK97nz1M3lkJGVJoOmySTl6mecysv6T7fqeKoH/4c
L8CXEQWZZXAaJWLXbaHqrVG5BfH/iNz09sUgQeBJ1Rl7XpHzE8Me7Wg3IIk32I4m
KkXU9McUJG3XBjiuyOiqVsEZ+G+qlEhAsoEtCAG7kTadlmrY7qve5hcTPOHEukYN
SCGf/SXSayq7VZSDdggHSdSiADWBJSTMEVEQw1aITfedSujBSHF3I3j5wQlrKLx2
LnlXkJQNPxVkWRmjw+FkPC6nTjbULgjjfENOaaOi4BtOGE9EdrgCiWKn19kKB7VX
5lvmGBppQy3BlN3bKW9JYSFuLo4M3KGAQuOk9YdYM+RDuNHbP+kKoR5UZTCm2s/M
U4iscIKF7DkzAWjiGhpJLsvjV3Mp5/k1HHlvT6ArrA6YWCQlfyoZliZyNRYvxPoV
OZS2+eLQqVyzPYcWHpS+44xHEh6U9mX4M7CjnmPEox2UcsIxD60vIiCPEYhcd7SF
rZ0LrsqsaiDHs7bBuiFTXGXPBMzJAXq21SFGLB5i41ALzcYcrGIKCUvX7G+rRQ1Y
kcAqTxYDfHChpxEVhHAGzoP3gMDsCucDAdLvUr3X1+kH2SWgghU84RrEMzCj2w60
+W2jREgt6HQ2EwU4ygauxoLm+3NRt81apprdfvaIeDGrNHG1T3lzVhWe4Fo2d6/8
D9JiLts5y6C7W/wifLh7qwZO0eBv4ZJqpir1no3jeJGSyaepn8GfGTrZOXt1k/YI
A3sDVQBoWiFkAXzAcoU+pxnZlVQRRGK/SC2AEdm8bUr76ROFjcSx4RymqmZE0vtd
U9XGAK32Mnbk7karMEF4tCYv/PrhmST4rIy0ML6e7wbOHo4eM2XAvR5gJamLTFem
72kFSj3963Bv1NXB5NkU0auq8RxtTcnvfl97kkQEvosj04n3aD6JqgiuxsWknNjf
dtPSaJeeAI9X7rvCOOoxo1jJjVmlSVsg+aAef/PCMKjN5CnmSR867yNUodFYOwZZ
1YB6I6T9VpOODYgN5uC/jG9GityxO5bVryJISUK1TbiyM8a0qjXkLV3p81Jk1I9W
xa8J7f2EyCGa0V9tKMIPnQYhGilTSiN2i0wuKi8D3Iq+3WicQrAB+fHd//fzI6Uy
nEkayPNIg5EqDTQZjddHj3s02zNTlyfsKsnIMkuDhVfua3uX9MhWHk4tQaYsMbg6
EyPstH2y+9NpEpXknF1aKVRvfDuC+kkNipzqH/9T5jT6+jogyoUJoX/8eH3eZRks
lWJ2l7Rb0rX0fol12Qwmz0v+9Wn1rdyGOQtzmDqnkz+bE3YQ+rMPbNN1ntTRIyr+
lh5m7Xdq3s5Tv+sFSK1zVNzN/gcPAWBWWhy+35RgSYXI/kuDtjcGUvxK5/cifycT
UvoxhrTTixmJpK5T1GaxRDI74YQ6Qrx/IkDpISOPU0sLn4A/4l1mQ537xOKJzYFD
U61iPGq2uf2aoX/FPFG1wdha0FT+bgX2Rj2lD/XsSSXfnJI7Bvb9ERW2aVhWtzWb
U6GUZwlHkEsjytwZoJiAS0VjBxNe/qBoy4in9hRWI1QxxEb9kLzrCzmCM+N58bxt
k4WLS8VU5mhZXSUUBgW89v0uL98hERE3b4LgpA24Nqhw3EKsBIdfl1hUILoU2BH+
ePudOH4SbLmUiv+0/Swz4gMNHlLFBuezxUGbLT1F9uCidYA/iaOBpK7xw57tCHQe
OGu7h5eG8q736QLQ5KUQ1IpurMvQvfXY5yFWCjHLdN+bHfExVjyy/MeA5PTUaUGI
oN3usgyqGzbDTyUmyWIytl4MaPFHzWMe/e774VCIEB+4OtvsMAoc8tEiB5Q1GbNt
Lnd4mIbmxVUUlG/G2w/jg6tAo5tl/6TVH5iKBf61a3Zxb307WeMk2ns1tUBo5PGx
D3UQpk128opCX5DFfaolNE4IiamvIuotaSrkMCdMxIIthV9KfWSpQxUoC4XtJVFN
Oz9GpK1uatmZwc+LyeIoWS1+xgrGsPhWJZAAAg8I66gb7sMuF3jmfhBNdcY0Cl89
VWSBQk5TG8KSWqQaolM8nvK9BZmOILEV2qQEDa9hiLoY9ndM2c19L9IPqXy2U9Hz
becL4ylHwAeGr3ChCoL2MzO09Nh1Lfz0EC88g4utYf6zNM3tyu3GXngeE34fbB2j
jVXPYgEgDpqrpJpFU7dYT1lin9DXpt//yaCWOjIXxEJ/3KhK3ykB3ws46VNkKLwY
zjhdoo16u/dWbGXwPoW32AY4nD/kIlqCxhDoBlwcNi1mi+Iq75mv92VdMA+x3G3f
qSD99oZkJZyqzxNd9GCPT/wefC3gUtdn3AdWL+Txal9bh3iYTP5bT9mJweTJedPD
xAoIO4RGK3J/EKZovr308VYpDi0dWykZXUDGAQud1v3gCgVvA2NX2VQc7oUb4XpK
mPSpy6+OKKloS5OWYJzSwYcZjjn+mB3PuGyKY0wJeX7G7tm/xAPfpnXwD33n6xhR
Op/Jl4ytwahC7GnMYDCkxZDQwZGoDjSmWzgugtNaZPNs2F6EirJSI/kIoociqsWh
ZThnzS7oytI6LZu17C4KvwJwDjfpOpXMud5Z5Uz0SweFOZrYQRZTudZnB/lyWEI5
0KPE+ffm3AGF60cQgO/nXYacbSTe/15N3v9eEVYStYQKx6moEhiG8d6gqxmOomuQ
wILzPs9N+9Kmh7wFQaeEilVocqV+OjBd3e6EPRGdNqyTzSVfI9wdQzLq5mVyg4T+
kAkleqB65HkjF4YZ5gIRaEW5Y4mGv41ff4SwefyVHIA=
`protect END_PROTECTED
