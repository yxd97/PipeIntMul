`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gl2QIdf4p8Ul803ETMg874pipkyZ0K44nJG41XXlHIjlpghePGO7+yA75KwsT25r
kCnClL49p9zM80WjZtkT2DsgS+n7ZtiCDKIX9XZjuKBld0Ijy0QOsH2eqdu2rT8d
4LF70trlJ2JaiApn7Pr938UiS6rck0Ci1B4jCgYhyDhgoVXQDY1INW8GGPYjUtOl
CQkH/pZtnIFZ2LNmS1wpj+tN60eMIUeII9N8qHZ62CXLFuzfICpMcykqmnxo1Jix
zOlXpW4kfvbJxNkQw3cux3hXmO0vZaaEImf3VBO8p0WXjOWBytvHa3CjT0IGPpWq
cnXumcY1HHDFvR00t7txAdeAXRWp6fv0H77mfd2jdkEu/Ew1R7lVs0WE+XyPEXXQ
Jik0JgFGiJHy2C1H3dRfMA==
`protect END_PROTECTED
