`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meAbrP+wCbGIeEaNA+/i0J14JJ+rChe8fDMQePCwMOKjM08Wni1DvQ25+C33HjHq
oojMBDajCBK4yTueIRG+TQcMgSHwWYCJEeWJwWdiEexDK189i4QwTCZu4h/MJ2J2
BXm6eq2QSReqN3HxBBBlBe8Vqd551iF7jH44VqozUcUsji4WAogmm9Aq09aa1A3k
kMmbvKwN4agQbPSlpwLg53rb1b6zaN3X/i840kD79AkgkodlnVMBBAXO8tVg25Wq
5RDJjkkkT9bTfH36CWeAv6Vvn1V4UkiLFzZxyUA3qo+Beq8wl5IYcaDOI1FsJowj
IrF21i5dBVHka6dN8TQOalQlPlk3hf82cWvlZ3TdJm73JufdT9SRnFrK23YeB5WJ
EF1Biq35qw4pngD6O7fu+SQavYTFxsfzPGyMSMw7GhMhVrqHl2uqtoJA+h0TubMQ
gGGel1pn+Xs8Dmb/cHX6Y2LECSTwlzkR04PCt9cS5QhCaAZaDP/Mz0O3tY/7ewXz
DN+49P3pKqRkVUmt1Du+H5yEj/PvkI5/JyUqy8tg8oZJobh06e313n3JeMg7D3Hb
keu2v6zcmMRWE2L36O8o61rDuhN0j+SjGPMaLf92kQipsQjUrqGU89L4IeDX5x9L
KIynankoFzeMRn3efwpt3GWsZSPfatMAaMtF5vGLAgE2dvb6iXUu2iWrbI4vadRn
n5FRexzOy5A6BkAnGQhDa1Y13QHZN6MWoKIom8bp98nrgRWWweTG4WZ17f8WkFe5
L8Ns6kwwMzJ0Fxx9+sefs7qHLMqfE55QFm7TFHQEkAM2JKlAg7fhdye4cHyuIMpw
0eyewMc1A69LZ+Tx+JwUh3y3RAQosKsSEVfhHdMWba3cbUjBPxTOkNAXkhsSTJct
cwbgOZnWh27Tia+RBQMPAYhtjquzociylIRv+omnifmSFnxBZHv7gqliOtMR25Kk
`protect END_PROTECTED
