`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mgq0mATNaxzvr8bgP2PLppcH8xQBGlA6oHOwA4HMJFa44vJ5lwcjbNx/aN8d1pnd
iPX4Y6SVviYYDFYM4d7r/iRWXw/tko0Twh08AdmFG5IjRTvQOzF73PodwbbaLDLU
SH8u2UVFMaa7qyNtAId0Lg0858tiA9ymJOtJC56jYpAIGcnjty2Vk2FI/YeD1PIH
u/RcrGinr7q0zQUGFhbwpbUEf1VJRhstSF82NWmPIcmo6/2m5ittpxJWrv/mUvo2
YWOzhQewBoAZSUKazdzH8C5J6ZTtU9uePeO4Dq16FhhZa2xQGu3aBe089ba4naXe
GYCZWwKYEJYvqVBx5Wq0j5WhEKzRMJjkMu7EKEyUoWOECNSC4elhtLu5y8qtgcEh
pPtc9l3uXPBoHwRLjOYUVW8cPWiY1GawOKeJqDLjgIZMp6mRl3EUAwXANlmlo777
UvmTPQtiEXOWKp9FXsRi8PfzVuqIGzUHS9eS7uC5FMkNGQ9h0QDKs46A15yS8DEy
PTBbUUhncN61ezircGe/1HmtSgbLFInJMWS7+qp7sneag+2Pb34EiNCw4s/YpQnu
dc/NtgVvDrONYf0hvy+vr/3Er9EEkayiti+ssqeaaAwP7cOWMf1He+GHbfPRIiu/
TtoG8BdmE4lZhB6uGI4GdzS7gFy4fr2Qbu+jWSiGF1zFBA5u5aijdBSzr2t5pC7f
WLLbjMQcGEnrCa14z8TVBb04XcWR5UZ1X4guf0b4ID09Kl4bOwq6DrpVXFGkPpOu
Be4l0Qwc7AfsqLTv3DX2SMNcfvDlgFCIqButm1FjJgo0Rwxt35kAHlWoRWKKc5PZ
u0HEgZpHuA0P5niOw1XJSkFhrw/bhvo3bLL/6deg7Fiet3KBTkXA2FiI78o6YgpY
FJRJTKidlc6FPq16VBg9erEgylCCSjbqdepxxxgXrsrVdCchVuM6F58xmYC2CXhe
MYuUH5vg6pM38iQBtGGBA10DLsv1ai123rHXYch5eQdYoLdT6ajlV0ahOtM+y9Tl
6u6gGahGXUkETtwZRB57264Z9rFY0wRNDlR3r4fdyBPxaE/E11EwvYi6suTV/5WY
4XAD3hjIMgt58mvH4oANHiEtwGwZ3xnWw0f0kWcxA4qWrzstWsljFrGT0sjgC/j3
riLBnDsEJN+VBe2uifjAbQluakhStT/OgGF4+UmiFecpR7Ytr98yQ3WI+kJuYncR
BYK4Ll+tNmHPc0V/Zcj22MIC1fzhhFYD8YfKUWrO4gmzXLnYFPWgOj/WTK0AV816
yh1dfQ/YTF/lJh1pnkLUwTQZ43c5utKwRPfQFck6rCpC55wx8s8KhUsjKfDwRX23
C5yDUEfeaoVfqy9ziM9x+4naGEGzqxCJE24+bMDCcwPp0S3tabaiTKek7TLe2j9U
WTWZcRY3pSiQA0AhlxMWewTruhVDOM2Jd5D9KrXsVWc0ma1xPtPNO9yYlzdna5bD
l+VpJ8dOf7QbY/3YkMaX4emN6h7ciAg+4rWIznhx+nxumymsfDht5On+X+77/k4o
9blTg0Wl48EYuombp/3cZL+BOqRU6Nxqx/MYKCN/ogn5ufsxpXMjUTjejW7LhCqB
S+iBFHKfEeJwQ79jrWrwqxe12K9xmF6w0oIIGafpkzb5oQGH0SEfuabX70/pkrfq
LMrGngud/e17UNKJbluKR4jFXrSK1EX4RpJATAV7/zTGQMq6kaIdoqRBN4maYWOU
VlfqXWzte/FzkCyklqbThzPl4KbpW9zktzuayHw1NNJp+F10JGh8CMXhEcv+NtrR
UPuBKZqA9rO4EV1CMz2Xk5vj87PuqUNNmwYU4Fp+zW7GK5gBQv9eygug9/5R0nN9
BXvAznIkB/Fr7w+JB0itizXlmCo4JHM928bIPE8gBQI9lcKgdF/0bHveaVpcm5l8
s3jvFonoQJGgT4cEnGMuWDPZaumnvT7d81f6NRhSmK8TTAmDwlnRK7V5z5Q/J0bo
Ym7BprM3U0MwDJ2q59pSM29dgfLNjQ2/RSb6OAwPsYkKdbNVeGBO2hpLFPmRZVrK
wmFeLPSLYyaP3qrukDMeqCIui94JOPrRYcjodPUJgHcTgWbBLs24GoOxbl0TldaL
bsRiimZdvCyP1rdJJum/05mBIyOgTsuzBAE8/oUHJc1FGRjlzG0rjpJ3m+OxUQ8/
nh5UpoSl8fFTXHQP+Ngp2HcSLG39jepH5jBdEcMQNVOIXaiZwE922NHATCe5RySB
QHuRMcH2bpjsZdXROUaUCc5QCjvbAPv+ZJ8WGfHWesD1mVV9MFjXyoYp58oFN+bH
1KAWngGcfmhkfcf5BFB/kVH4wGGFIBSx96Qy2LiMutHINU6HfBNe/+e0pjRuVsck
3Hl386rJZIiWWWzJ3XtUiU5DXlESW2TCIj+hMPCNBfCmII9sWLAZUshshQMSVJbI
ThwC0f/aCp+8cgazvNq4AnMzBj0ISN7ShOOj7f8huXq9Bfz5MiOP9q+ICLYHxq0t
EbNwwri2B+D5mDkMtFbF7v2kQxKzODZ6xJYhLsE0Z/hVhUN6UinnwV13Cx6KjqW9
Pk6KRtwpePP8A4zL2x8VU/gQDbGeoVPNQWjabfNHZ3v0CpOmbnYI7WpJToQIMM0F
4hBRRFaBQXYZehrt6GOjqN/HgzQhes+BtbqPtzv+gjCA19Guf/lKvV55BNtj1jV2
X0mSUKwqM0RV8SF+hgb9pxgQu4Je4csNe4ga0EcMI9Wzm1nHFmtJXX+y0IQ5oIPb
A3EKnzEjuJxy6AM9cFSKqBDmtydjGJ3waO6XNiZW+k5iOIPiyZy+tjnzs5MsQrfR
6yA/kqNYImYgZrYDi7bqNo8AzNqOiv+ZVRT0DD8TRx2KIgxdo0MSPefytrEJdTyi
w9VNbF+jXFVZVpZtk3h/Wppk8bmy6BvTS0HZBclFw1KfiIwwf3zneQcPIhrB5c0x
J9ftwTFlfT2XwztwtCv5krpTN8gEJZfheSLWmd69dxACwIvM/8wutue1oS6PGI/V
cUpchs8GODCxP1V79ENKYJdquPMcBZ7Wx+npGjBo26iG6CEJI6vgYq0bnWVpDtSn
m6uOefAla9b8hrbR1OUDa+JBW2yaMuLfFIgdBVSInkO1ECmNJSwL6xK/gVyY10yz
QAAcaTprMQ1qlSWcYrCSEeTz4PMUbqsB1bi0lVqUioFk9x03cHoIkU7daD1KIUJ3
zGW7QKLi5RlPjpXf6WQ7kcf39lnDJP0lq6jTDz5SJRpTjl7f495BKVJFV84Uha2z
JgQcdLOJAnZEHQFns7kR+fS9PCzKOnMkxHTcRuX/UuCnv0LNys/AwqTENYLbVQrP
jULidHEslXZzxw0ou6VpfpiWLrDqSAIkr5ZNoJQSFYcFXAow9581ngU15QCo6awE
MIIYHlbFdSk9F7bVAAdJ0N9oxfN0xJjzDXIx9LxDf6Ms8M6CvumMD9p+tT0Z8D+6
UdI7g1KaqLFLc6N4RlsLbPfAwZuhxqySIwJc8MPKKLRsLRdlL3aPtSBwd6mz8fOJ
5sgICwepO3UiWWfIjL5yQVfmn4W8r9noSDK7q2gJrDoEr/CQ7tDYFNyQQ8QeDyiY
14RtLKRRZzH/3OjPvHlB+HIzil28k3tcyIcTBOR30xgVRbIFwfhwpjOcGRJkQn1S
BqX9lYZ9QWvo2w7hiWTIHLVe0wZnZgaMXydwwmt7DLBdwt6WVHIPgvpDZ/R5LeWq
6+m6z7zZBMMJe1gGFVz6rFsVpGeZyWYMt59ZQB1DTnJS6U34SLEzzSE3l+uTbNfM
L98wyslOWtyFnxYX5rFoZO5aiwt7n7SXoCxCTFZS4CAK0166oKypsWpHYqln6KYV
QYMPACv4IiTqzKWUGhG1zK4XRMxz2RvTEqEsRwx3sDKNInKycilm6nCXt1DTOMag
c3QbXJW8axZwY72Wf4uUaExlxoBNcyjiApsCZpgBiHOXDa9yNpKFxbISPYSrMT7F
6d7xo1axZikpvjR5JavfVSI3TVC8Dr5THr4JRMCHhn8f9B4O/zVmFXTMShZWgQrI
VRbFNqkYLWJ1Ow8Q5ks2OVcDOW3Khxe3Q7AwJ1H/3PQxj9MtOPZ6SyKOFWNE3wff
ocxLD7D0gRgdRAr1L/poDBzIzad8PE5JKjyBOXN4XcVgpbhBPdIJI2/p6L1XE0rm
tPYzqfBhqiBT0BeKznUN5FOLf0tGcHu7DXZ548GHtZv9QKsPknxAwHnPgT9TPgty
3pc0rh8/9jP9+qN2ZbMk5fGAa6Js1ISI8BKTUP01zjX1oj2B6Pr8MKUedy/MpvyA
iJZkUEKoYebBQdViFt8dCFXyuJASH251kUhbaNaxO/oUgAiqV2/DcjTj/fmNF+Zq
iFUAp3QXWICzmKmNB8TLIuz7UP3dgmT/ORfTdN+AmzTIc0G/PoK/maZz2JRqEmLA
jlu/uqaX0ajRnsfdj7k8n6B3M2FajHuHsw6tIhcO8IFGRWtfMrnIgr/voW9FIRBP
D2+GOiQZUGG4KOuVUOOqBgX7JgiumaIsqpV0JKSNk1SXo6sH8NMMkF8CwozACfOp
GktGez1MFvbO/U6a9ZAtEFqlIEvYyX0USEveg7qYWHnr3oYiDHYK4wmTq/vVGs3R
b52KZqY2nO3FUdHbyiCNQ1rVPibxgvHjSTG7vq/53HlGJI21lz/CnWgdZGLFemLC
vtLBNDUR4DNT13HtxGYB58e1Yf03WhrlC42B0krCy06Cm+eLfavh9aaRL++I9v16
PYeS6zJ5jY/V/RGacQ+f65F1aHDqqyzU3Jw+qZDRR+GNVCN/Kcq9679zVF8zhnwM
Yym+JeurUTEM0y3t4udHSkdNsbbZLxu6WijONjjwGfWNAaVt44Phthx+h0JymPSC
cjZX09x50x2pMD575eXzeuHiS+m2yHgXvX2pdc+VxXzPhlxnP2fvd+FHb4EB7hPH
LCRbxIlKVBQ0tMJiCNawvw==
`protect END_PROTECTED
