`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hDKmj/Y5tdAOaQkddF0sXePVpVtHwE4gw1t9S5uoAPt6EHt2kIrVwJRA6in5n1FH
S6sJzVWrKDYe/0VyTLdAwxDcAyfFlg9/lhO2Jli2Wgv8uEo3xsthzvbVNMA6myD6
F8Yde4BMYkTUuaHYz2sgNGHKGBjR9uzzDeDsDd0avfmQ8GOWDdwk8nxXuFHGN2j9
gJSgKQBWilQCQzcowz3g4Py1dhzgpyRQLgLB336In6sQ0Vb5oXTQtzv7eH91SRH+
9Oh0r+X3viOsbLABCH8Lh563nOITOUxqismi60mDpRFaMXUv70ooD/BsFgIOKjcB
pl/qpZziqtlGXCHpqndQZXx8gTimf11TJqoPQRpjqfem/dm2OpMttjhBvrafGKzW
LceYpmfZ8AbZAazM+vO7letqWRnYKIiHdvZp04oSF55JUwGi3Y9OI6AudTRaqLIB
28zdKxUGL/upkq36/vPZJixjxGE9tTJMNVu3nVUrp1d/cNd5E6IdsQAOOIP9yoez
ANql8EyGWXyyYhWO/XicDSpcRSXSk/6prubxtoizlllX1vVMwPKJx9PuQP2RUWkW
0mLZ0Tl4n4UaBokXmeof06sAzxJ9UkFzXwgpju1hMM+I5xnQsRB7BuU9Wpd36T38
SsnXJ6nISnw+iCiD6+iJMIPGKiqce5cKaro7FTY41BqXbz1HizEtfOFcqzXehbjT
LYzIB6iPdOGGNg/fsxLtMckPWDuN9zvmC2Ng/4ijaiXE0psOPF9CCz1+k0ZVyOqi
tCDfpqOoV7di1B39lh49iMYbfemKAijijP6nPoti35ogmB9BHwOjEYXbR9ByGk1j
OxsT+tcOkLaYZfbjVK9XLd4IIlKosDgdohh639uhwvPUlc9a1xoE2BVQxnKgqLge
dq9PTlH2U8raQ/70ICXyz5LyFYnkzvsTt4q1aqHB7S8gOF1MsODNmhjfbgDuX+xk
QVO893MNRBc9ZK0OhmTiJN1tW4LzaT5gVmXALMNrpYLItGTk82hP+XtVZ4pZu2W6
8f/LvALQ0SbSTSvhYY21uw==
`protect END_PROTECTED
