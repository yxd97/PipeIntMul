`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+KtgXToJ2f02mWv2i7+pTnIO6NOLdGQETHWS4RJjGLHagGrSQva2lbSwvm7dtlun
9HbvqAr6LjdoN48JJU2xiK/M0kvk9L+DhLdtXMHdiXmkZ24sLLKwTjWUE3+nLtWe
a4b/BZRG0jD0xjs3dCI4zQyJXS3/C/RXBLwhgsD2ESyI4xeLkCPRR6cyIxhKZCAI
xizTqVsAXwW6gG42DggZP1Mu4ccEJI9SbBTadA31qkuVzP2+5242s2OUB56te1YW
9pctgZ+OhE0w8JyKjMc4pCkEPJNAihyimEAGTWsp+ci6IG4GXIcKgHxyBL0c+nQB
HaICrdehV5Om7BxWRk24bxFrSXHfn1o0NjXYROqbpS88/7Q8pFLJT4h+NIU2TSsH
IQ7PpPP7COe80VoW1zBK/7AOZxHOSCnFiu+9Da2vDzwg/OWVxRsL+zoAAN7YsuwL
2PE1opb5UIE0A5FlkUpGurUAlvfciOEnLsGhLI3E5xNwdnyVTfUHoXJ+nt/RDoMa
Ro3mwMa/73Jc6b2iWptjpjLq9nGcDnc2JWzKljfyM2/fCbCahUPgzaFBoGutH+Vx
ZrX2Uvc5P+cMPRpmV7RDjWzV1rD+8X19aoQteTlxC07/BCdjJrHYuJ6DvXyRamPj
siMguonzSe5xLOKAHe9bymlGonCgaZPCBWHOoi2oIQKexddMJ251oUprzCXgkLMe
D24n7dROh9b//NhynRmsYQMPbkH5rft4DOudJXh6v/6xSyy8LoAlUjtoZuo33rAx
RU8zd4dDnpCq7pzWu3kU2pseGLcnTAE4Sb2TJ49+A9QjdqNo0VVyHqQYBkBUymbH
Ob/T0AQKgwlOFTpf0iokR9/LNiYU1OhlgCn6zoGV14yrDhi2oKqf3FrGWcbyA5EN
Iu0a38R0x6+4sBB6uk7j/xXcuIsvFKD9l2rxPYU577tioaTe4W2HKQj/fu5Rkzzr
kz8tQZtheiMTuGClq/mZQNr+qbgR8KXhY41hLRBEQVDCTWPL0LtX9q9p7DtPyuj3
Ho1aFIy/o38nbUrZc+aU34mFNtTf+faesTZ3ehFasOr9Ugk2iIjjcZgxp+rFUIgi
S3TEVKmelEORHYfTdx45swFtpuLAty0zm83lU5e9rvXCUTgB0FLN95wj6ZQieXqq
A7DQLkODNGsewxfHv4v0/Z0qTyaqlttQTw6ta77htIkjEo0+nMZmS6LFDJBb7XhK
6FR7oWZ1vmeqz8sMVR6KeTGhdF38KNjvbHdKjakeI634Q1WkFpFlMfB2KepTvj9J
JLdctAB6P5tIveBteB8c8pC1HfvTbvmghf4Mx0QXZ+PsRrXs1RCJ9btXJeuj3JNs
JHppMX/y70BP9aiTEpX3661FBUjygd7qsb6rSX4Wqi3EibprN7tywzT4meKIDbod
2xrMzR8dGeSFdapHxYJKif7I7RZZq3mDiHowDOTN9ilgJ+ncS6jVsfbvbJukfeUp
JJFJlrUEwKbFSI3YBI0Ks+kpgPOnoxrgnMMSJ+tV7ZzuAWcCFQ0HCAID4b4vx0RD
+MIW/f3cS0FbSLidGXA3SDsQJ8IVHtI4qs1TXvD7BwVuxyUy9suN9GmgbZPIKiZR
CWLbjOxgUqGhHg+a6Sr8TMo5fRs0X+EjxmlA+nI7C1ulEuqeqV53K2Gtvz0rPpYT
0sUhMimgvQLB1E3CyHjcotXsGkV43ygW4IFxfKK3pVv2vAFPMHoucgPghWxManjl
MyYDQx+j8Jxvdzd53EOf/TX8nyO1GUkpo7/9pXhgbon239fVyzy0CaWKz9QK5Y7q
6o9df9fDZnJq83iZriXo6Z7gTKbp0CtGgg+Hxgf5ZVFaXi/3Zh4wn6qyNYA+MlDU
/RSg2e+LDy/tUabkbEPItHMN8uPW7Oo4274OENkoANagZ0lF9ibbFT8TpYYtStyX
Z1LVDZomJS6qQRH6HYkDAhcw3I+jMBGLGteWSf06CZYuFUkyDxRUdaqPT67SiQzr
UpEkUXHrF/M2b6VV18eRtjh9yL9HFxjrCoLnoXHgf7CVdtQ8TTgLFfw7Q6tvAdqz
EDBkGTs5HRWq9xAd9TM2Hswgt5eSnhJjTVF2LGAEAI7JOR3mjZDQoG8he/B7qaQk
8rvMH3IVL/Ns04itNiXd4svDxoXMtZKA18lhirVWenSlXKrYlCMclqjmBU/7h+ff
cWdEaFIoykJH9AnSz1/9cMmWUbOnf6vSpSKoKIIptqtjmeiXHzh5YD4xUQ+ODf4K
16KmI5IFTreZ5h3RO4teehUa++ykdUi5NmKBaBeYyqhY/YauxYAI3spistwxUQgI
zUbu1ynuEDQzQwF7HILx8QF2SKf3qy3AlLJMxYdULmooHkPGuR+UuQJc1D+MXe+Y
+3Uy8JlrBn8Fo0BIf9tzmv0+DtMSb3Xa/36jQDUxXNPv5NYAIiAeJUkmoBq+kbyW
XzIjIpsyktwKmXCSwGoWd6+Z7o+5Zuvr8AD1DopiESY6s9a5r0KUOiFC6IafOVI1
KT9ZykkeyurxRZNSbsF01lq7egm31hnt/m+eGGF8FHbMHCjidOYDxaIxDdw0/Dkl
Qa/96pGGLroPh0jWuk6Nx2N592Jbxx04x1ux9zP2JE8Ody03Zf1tIy6BDgRFg5E3
NFqZCX9bEtIANeC8IyRSiT6yc5HwosrwCNii7jPX6p3oTmk6wEiELTewDVr7nrHo
jQdfMaIhGwWEf9Ud/iXAVTaXVAq/94KOBbCMxi0+ctpkD6HTQSruvD9SccuTvxer
KWxcO7tM1TEykGmGl0XBkh3HpUJIjkDReF8dF+FAB9hb8DOr1K+n6HKBCHv2bjuV
wDtNFd9uSYVxFdReozm8qP0n/sO3oU9tyRRcv6aIZ0ibr4yMbcsZC0/t3Rvfe6KU
+w8R/q99wpY6HjpgyQHq8xA0bkempQ2Ywh3Uz3pssmBFqBYmEGGeHRFCtcr34WYn
LoHJdqARp5sYa5c9Nh9gD1klI3pU7WA+Tnts82OHeG6W+79LyYm/bpPkuVjceAy1
hqyhbSt/EfYKjJY2pZZaX6MEEiHG/lp/7k2WUuS8yULy73sRD2MlD1iwNo4nt/P1
neL6YfLp22Ecf8m0enQGHXUIEvkx/rrWzxUC2/BAcbhNTNffjRXAE48o68QDtlCW
wO++rJIWvHC55N9r1wwbv+Q8/NwwFPOPe9DzRRr7p07QHEZXwICggY1mqVNtqZ9q
tRjPm0qKiE6XpBaDdIfa3lYhQYS/VyJqzsHjq/9G6EQyZ85oP6/XevRZwyV6aemR
vb2ax9H2lZOo8Oxuf+FtEQ==
`protect END_PROTECTED
