`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7DWSp+P0e+kHSGJMuetD+6SK26RYQPCh+KBTMSLb4OOHo7GN2DDMdpnUqdaptt7
cwTn90bBE8jz1hNvtEz59emHcdsiFHTIptE3f2kH6miHk1O5uU+7CsIlIIVObIpO
V1WoslxdjMqZY08Gqp6pFcvlg6fEDUxOBPlmbmnIfRQP/1Qs6VZHvTy7+QPT2CuU
ORPLzdZtWVV7MGhl3F54PvNF8dDSL3aqJ8RQv2zURA5RXXAsljPTqkGLYcRSQlkw
tIFWh+killNA7yaIoXVLCVQ5GmHQptn+bRq9TcONkoNYRvtDB5YOtUNObgjA77AG
pJuuZYF8W7CP36ghmIRejzeczKxVk5ZbHXVB4mZeIx88ZbJuEXtz1r/Jyhvg6DBq
Bc6rR/8hgB0Y1SxbBx5thkCbH9A3QX6TGMe0JNmYpXPS62lk6hRf2IJdwYuvNT7O
TrFX6lKbrDJtOH7PKOVQKcTQ8aBgogYzNhNN4DFrXXXIIbNyoiwZ5kYtCT6SSiQI
ltdKjg65OAyJNjy2ZQRKPU4jVOLplAjxku6HbC3gLbmHGyqhOBP3eGmn8Q83Ce/4
a3Hdl/E4bczX9wiac6xZm0hf6svOeSZmtqmfew2xTwEe/N7PtOSWbtprHyZH42HS
46iezbNkZJFeaLukQld6sAoa4xFf1J08UfCb73GiCrhXyxNs8rjrAxxhnfU1r5pL
rhHy2alzEYtwjqaWUWSvEO1AlbDfwPVT3LXOKkIIbunDV93Gol50o/XfrwC5SIz5
dlLR30+A4Rg+Y8XBbOXJdaaxT0RTZWZt7k7ZyWLPyGzX9rjYeeF2nt7gXork9T/G
+IRC12XJ4x3lISqdYa33h4x2W9/9wmVfuzuESfzcbXFwM4seG2sk7/bN+z/XGN/Q
gMF4UdtU/J/fuXx9cAjOP78rx4t77NdtnZ3dfmHj35c0F4HtI45R4D3nXQQnW4P7
v0g7hwXSsno5qMW/Hh5HXyC/dEhHcbdojvi8ILgPy1wY3Kxni0ZP2+wcb4dpAdgD
ROKcNohGDh/WOSAH9fXL1Bi6QeJ0Ujf6FdOQbBYuMX/wtn4Q0gypyMvWYq7xrDni
wwzlDKD0i1angDLHchDnMbHUrdStihs7p3v5u0cgl8M0rRn00zcIRobOpsfoisl+
3Pmzwv+/3flv35JyWjTV7Ufqlk56neJgiB9p0sptGrBiLvNViwbz/A/N+FLOIH3L
o39Qm3SZZXNS45zSF0s9ekQ1kz1rKNNJPvuxZbcleOPNpE6dehkO/Xsny0PaAfxJ
stBlM2bfMoyl6wScA7nw6iEQdZ+UJwUPaWlhLXUQFik0sPQWZnuhz8IL+oyblYhT
DN37LutVYs/lp4BI58irOlK54Y8xHVeXWZ4QS5JLKJgNnDpc3IhEjqEBbXvx6TK7
NGrp8FmT2Vmpai3awdGLZG1fruWFlyDECeD+f7PEiBduU4vdO45+7icpD2wBHJI9
XI0VyNB45XKCuopqJY4kHh4vLvomrDQw5LVoMfxDIsdDoo6V0OsVMRdXFKgeitFs
vOiZfwRD+p0NXZVQPyAsC7P/z38wdPZVgO2apRYJjacN1FDbr09y01pzCVqRFsOF
snj2HqZ4Y/an4/vhRO8gmigkqJlFfoceGqCiBD5GVg9IKKq3QAAdJ4ymPrRFCV3z
3TdKKgJQ+2J6sMB85U2eB/KhDXcduLIB/8e8jVh/097uCOuaGav/3+BB2pHSx5tI
v37Bunc8w6iFmSuKH1D58oNznXrLNQjUJ7ejx8Lq6pGsH8oDhdFI0+KCi+wOS/lj
KGdwDc6ROTnU4LXPU1ceebflGbuBvsI/ruHgcAKYBVeTj/P5ofL3POcEIL9wX20n
di+E7KXYuJoKTEvRK+71hBgThfKmdmHsdVMLdibwXnw4OpPwqcCvV+QULOtFrV/g
1uTpYbjISaiCpr3BokdCik3SUal49WnjwiG2RgFDnfV72o0uwjOFnuDlOwL4N0c5
B7nAnpKsRwG5GFtFS59yOCKYXWQz5t/K8btN8kXwbIACnDlgZvoGhVNIuqLunW2A
D2HnMi1fFVVgFZjGRftAjbPVoUskrzMXNAzmA+ADXtC8qXR2s3zHS1P1GpyaUbzr
10ZVRVkwCedjGwJwZTlcdhNrpcu1zCjt0dD9bX4wxiyyAZbRdyh2/WZjIGF9nbqz
0/5jGM1K+DHnXRj2A0QcNkuP8N9s8pOSwttAak49aD4xcvKih/jNWRtHhg5bl9nM
Glbgw7q7UJqaLnFOlKGgaJURbXeDMLh16Ca6Ny2LrGafFsc7spkzEQP5N1Kh1uoS
kbPsQdF9+bQQYgIWvBzwXr09x2eEbgqb5kC8eFfSZSt8RoDGngb6aYJAEpw5lmoP
0FDRqa7yKNabef8j9BWk/0oIFVwKOUuUzd5bb4NufzMG/tbrbZXSb2z6T/fpB0W0
n5foOGuglUj3fKoIKXH/CE2/GgsKSCbRPpEU6faeNlWrCU5n5wlzRkDEXmuzSUZ1
wto/drTbdPnN6RSTIsGyXd986hf8B2cnSge+CKSngpQW1w3rRYJHzggJFYNNDAOT
IU8LdMpduTySbPSZ2asH+Fs33JX3l/ckS/XHU37oFZhYm9W4VM4ozfWflImIOklI
IR77YNj903LvwtU2ukqkwOBTK2s/edAQSJrWNcTR69GoEupS1KOId5RtqqlA9iQy
//RV0xfMUTW1GrMABmud2IHM6+Z1oWE4a+LWabG2a7eWqGaNl9mFcMSJVcnnh8df
gUtku542P9/C1O21FpTB9WDYEe1pEdfJI0eljeLOO31dEPat5Tiyz8/lLtbzABJv
dI56pR1p8xMumeQgaMvlw5jLmwAbzb7TNztaL4Q/11wgg+MpvAHtFOcHC+xpNcor
Ia9poUfFZWbjc4jX2fg1sGxtRytjKAaRCVT/5Ga22GfD6xI4aFcRWGm8ZSTByvAs
4d8+L0WdNk+xebw1HDClNo5SVSDL2sAznnzzv1zSkNLgbkufBpHfmm4TypEIyDCx
mQk3WqKluVKxhfVJOYrer/oeFfvnyi1Rs6DR3LGe651kcYpGG42gid4nZ6QR1mB5
uhm+b9h0hb3UBpWtvxBFrcoLAP3KVp3taX5+2v57fZrH/LU3DCBsBuWL04GIxU6t
wBpgyI5KfKJ9+1tzgiB/WoYPh35bVXmTeGm45piejLKEbAEU0BI6e+wsX2A6IRiD
0pmHB0qHE10Bvg8Rz7CFNYrSo6KrQYtI4N8vAPxB+FuPKcxR1Pn7IdaUHzNnanVE
sxuwmnsd4qL1nKXIRKeiSE/fYb7LEmKtU+L1lPC3limc4IqXOiQy0VDzSoYlm8np
8yy0qOTfCKeKBobWobwYCPDNXSkP3BnOZfGOtYtpM5O+5p3eDIet5Tt8vYbB1NCb
W18WxcJHqErLX3fgAUihJExsQ1sngsHk94x5Qj0TBWz2c8G43HA+wC80GSRry7Br
u1j+Iq5IF1xBdofXThpceEoJ8xYxcsINmqKIxEOsPfCHV19XcfIUa1I3mtAY+pMK
O24I6GEMvgPA8n/64jdTTwM1Al67hM1QIjm/5NQdYQdXw6ubZiomcHZXH4gyoQby
JjXu57ZLyeRsFjqNnDZ7bkse3eBDi5vibZUtSe0nAVeXcyscdn85hlX/lKj9D6n0
xCiGmyznHNhozbEtqBtWg5LAaBP1XPswCVwaDuFUE0wxmkqAIyUlDEvqSMck1oZ9
YdJE0CN0+9GP46V12uf+3vzRWDehjmZu017IRXTUkJT/9P7H8ltaUlQWIjLtiBOn
ItFDipBOGYKTGXnraJ7p83PqTi8icNRcBWD9oielTYsSNnaIZ9DKoBEC9IwXh84E
pX20isgekw8KdpdtifWDK5g2UE163GKuLRqR01vyWPZ/T87vrw24D9iLeuvLqudV
bdBBY4jrackEJrcG79Vg11Bfa5ReWdlk9H6W39dW+umHxlZN/Ow6UHY3UA8lG2QX
iB4JTx7M7bt/2R1z/c9fXCwhKCDIFP3frntB/3bkXkjP5uSLuPNJElZPkd55AUvY
LOvrb7a6Nxx3B9r7rK22x6/t/f86wwaPIfYF69cGHKVo2C6Vp0AVodrIOPoX/O8W
/XSEghj7CnZ7MGjUS+SBzVj/lScAEFs+jnXUVGiFiAKT9TuXgkWA2xpNXtQoF4xO
EzUhPJ1uvbRWRoiaNIA5JbB/2kdvU3g2Su2RZBX+LaFtnh+6xbugbwEUxMLDN5MB
OA/fjsVVZCCasEHvh8hRoP9z3r8r06d4i+UEpLimFsyMmCcXOXwqXoZyMlc1WaxZ
C+AgWCgJpqhi1TW0VC+r+P9HNPF5FLFKtO4BemO9Xl2JAS84OiISMwU5x/i5XlhX
qnHidvSDG7vU3xkvMhjpjQvxEPQxG/Etuqr6oxhNyFX3YfdGll555MOLCsJ9UBYZ
RQ5bCN1jfJ/Jh7mO7JvSv74K7ZP3FAM6UQMsw6ASyXRgymqg7+8UZMZ/8PXPzAgq
ZSjhIB0i1BizfPTe6gKgHSdGyMKLwt2rhZASB8FQ4Wyzb21TbCkUlPXZrT79Bxxd
4E1dVorPXTb7lZGrIxk0BAmkW+b3+vv0Yz3R4eEyEG2BtIezifIArFVV8X+QG/x+
9KjfeFC8gNUkM3Z7xXc6GQPKNBQqOISgHGhQoj6m7ayaC6xKH3bZPyDca96+jvAP
bdLe8dELSAhBztyLYoVZtNSpFS8kuTqO2WXkVk+jVkXC2PjYrjWpMV6xjM3zPhrh
jNlP/0PS1b/r2kXwwsyprv8UAljBwGyKrCt/sM0yjIIqzDuWClBAEAZF9L9ALnCi
8o5Nkvf5Rfb4lUjc0KwctSR/+3eoN0GzQ4KcTYBLJ9di9FMjy2IjWew2bKloN8hg
omB0Furg1lF/qBzIRpxftstS/snJ7J/XCxjmNuEV3CTJhFMbOXjVPUoNEyLyfFEk
jtmIigZtnh9oIzo3CksWRN1dEghRXYYf0JdMPh2TRHQOWagB8wECMeIpeRjPG4l3
Tj3ycnsCBcpoEwg13qw7e/ZYimEmG6/oDKW+dyz12sg=
`protect END_PROTECTED
