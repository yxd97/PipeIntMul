`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7xkDSNCA2M9OKR95chCrBZiFxoYewRJze+3ZZVdm2q7p9vXUhv2E0aFYTYjuwW2
N6iPuRjiseXMmWdTpHUrGEoTBeDhxjbmosfE4OfSYspGCFmBkOBnUzJwxe7Mf0aA
48q1WBnp7mSCCkC7uVG5dDzoAoNvgd3MPcti6Rhqb5Ko425A44ZLicygKMl3OrJQ
5FymlU3cNevkR3PH9LYkvQEQbGSnZ9IR0wzYXH0rI7QOMCpKfDu8M8ZtHXuR0zQZ
lxBP0n9+/L6gEJvDX1nY7IOxSrN5khesyAxm0Nr5PzaLVk4Hdjiam1WDZg3UEztL
8oYbWgzvw7AM32yihn0JqXycQs3FeU2akWmHjnpeVtW8KhRe5Suu5Jx+zp3AnqHg
ZUHCmd+FmT1f+aAIf+h10T8kiVX102wkmKM84NCFcLx1VUBe9x0vJzNSjbZuR5r3
`protect END_PROTECTED
