`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNn7OpFxbtH5SBYAA52jWjvgrbALxoBL5E8qHyAjvngOCgvNSuhbNVit4XwHrQPX
H39HKAvSNpf94xHivaUstFupvYshvG4izMKRSQNmysIfYrI9/dKWm8CW1WYoZoKo
TAXU3SYTudlUV07lKJBkuYZFX4U452rfHI7l7+VEqzFYCr3BeA6HI+/YpRS8Opd6
tgcJwgpwCMDkycd5o3khqLKS4Ws5CG2ieru3m+DcsID9Iii8qXMDwg1zEYj14KOD
eIWzuzqohFWaX93CL7CNNIka9Tsz2CV3M74LKs3taOB3RG0aNRTtMWM1C5ZJm0sZ
2jRJ5+dV5w5z8IEKNxqX9q+SLllm/EqOOUFCcbJP0EnSx1FfVrNPH57bah8I8QQd
8pzPsSjr3JEpYnWSNVhs88MlZBn8KvZvMuYpzNoLuRSqzY3kRUcr8A9/zsQfOFoG
xiFDdnQ2sm5TRzIb7+H4Eea8OgN9iQv2/IraeppB90zz6PpVVECfbcFweWhmoFNo
QXWKL3i7IECxY4QIzHrC13A9FVPKKldiBYCvKRevRU7jFlj2rUIXRrYfWai+IVtG
H+8x1ZwTHoIINq4DTt3WwO+hdTNWimZfVl12dVCVQIuo52E8iEhpQM56Pq0fP6Yd
dFWLKEF8sUW0VYOuHqkewnPcACeJWjREvQkq5E3U+YbSXwG+I+tk+TgOBoujwkUi
SWqxOCP5phlJNceYizFqqXTIGe0srFGU8Sw70g30eSVSZjYkvovRONogEcsjLxNt
ZwXtA2EKXI+3YnWjWx3GMqH//ltbSrVB7P9BdgEVssr8V4X2BWOIITTCV7akkHrC
nzq4ZWqxL793p35iNt+1VIRYu3izCt34a9vhWdx+9liOvAK3Rt76ZoqjFWFftfdW
bvaOGl8elt8u2bzB8e6kr5yuDrHXoUw4X8H91vNrAEXHRkTVW21pyNY+j4AUyhQr
WbSCcos075qwDz0X9152ZQ==
`protect END_PROTECTED
