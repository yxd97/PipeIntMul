`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+cxevlE4rqGV8ld4CvO47O/02XILUbN2ZDpsGYHtla2LqVfaY6R0GXl5ZhvlSmtY
lrUuuE5ejFvO27xDBggOiQvOhJ0uON+EjTh1TDB2tcXR1jqDd9Q3Dq7yusCJeDFa
xfwpu6UaeWj/+DmTgYw5IvEgizP7spVh4dRPpFkG5T5L+QM9V7qsQwVcAGxIoybK
c6W2PuwpvkvaxxYnjfryU1jz1VWdxFmSlIgSey1OvcyLxrcF2nlSPzETn8AhkmMV
KZ3QYW1aD566evqMaiKOdCcnmclMdTaPT/U1DTFTGvFjN8YSyqapIlEgivvIiOt9
1G/Kq9DSaiVfwCoPvR723JXz+cpIJvvypsh7sgf5eJ2Lc4Eiihbv3BC3fAlJgEm2
tazNvcHbBNEm5Djj9gekZOvXJZUa/Nbuzx25yzTsra4=
`protect END_PROTECTED
