`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeV21gMME44yzvdAVQjlsM1WspY450n3zO0KIx3toE3qonkxnBSco0eS+RO1ch0t
J5peXrENvjzQFzDxUEpgVnLA9ow/g/EZ3bpnyrly3KwC1wNV7jFUSFv5jDmMzHj6
4P/GNoWLY9XwIm+yfncOTeiszzQaTO3DJqwBTl/rDYA0RAix6kh9enpflwhjfyaW
yf0ptpNxHzkbav7U+UGuXccPVINPewp5hGDzknk49fjsQr4Iq5F8wuhhRr1hNdI4
hGepx3CRERarWo3WJu+baOK/B/b98dWHobcxGK7H8mvkX60oWsBqgKV68Jaki6Hj
hl6NPMvk/Foae23ebOsOD1vWkTX8yOgff28YKM88GhwUknX5I1auyWzKmCWI6kc2
y8K22Iipd+9yJPl+r1CM4j4pJO2V9TeWr27FOfmbtcsqrTt1SC//uNRXq2IgJmJL
gG+DF8sY7xZUDH2CC9rZhIp/FiQSAvlj0Ehcx/SNtTI601ni4B81PceL5U1EeULg
dZUhGCs0Yj1Kb2/NRSCLncWRR1R9SXtyyuan7EOLRB0p4XklwhwyXuMnCiDEMiqc
+G9G4KuJggCZTCt/HKDMc8nXSLFJDGCsqfYfqQyAukqwH3d3XFH7p+PgUAprTkHN
nix1YlxMuRr9qfnaoJYkSNEZfRWzlUncmLAd8PvBdrxP4B8i84lwO6ez8Xd3AJGg
IIvzUDLJsQEg+OKsBSANc+0Zl81u5k/f3BQZJMTkks7eM8D0/lM4eVy/UV/LOLAF
rJDvSv8ZjxAvdd/ZKKubxfyrp51d20iz8GBFXpoyD0xy8Tq57/vunWNHrRM9UaSs
eXAR2fQll9SzybWM9uJAJrn4qq+Gf+TUq73xASGUf4ki9pPMvuSzMS/B506c5OG5
QWKm938pxacLl9NHqru0hy0p3ncGnH0SyWHQ4dmhnibmQ/FpI3qoPTdHVGcHrDH2
p8yGieSUbzGkcOGYFCmRLpQFh3H+hHvplyrYNDQsiJT72yLCwe1uLyLHthHTwbtl
gt1MGppciu+CgAVox6hTHpL8emD5yzZ7UQaJOCJA/ao2mx8gIVn+DfM+ApiEVT4A
j5PHgRSjanwLjIc7nIB+onYR4arW2aHNLPiSpYu+1MwPMebvNpRG0NDkr2esdcqJ
gZzA/vTvMoqwMGFWPJLPL+BYk4rwTSF/N8SOF69XRLTfjjVnGOjZvzCP8+RpzntE
dn73km5QWQkSdRjkAgQZV/2dOGTQ1/Qc+7heWSVBynoqBEfotfW0lxoT07dm63Ip
uaFdqRzCZs1uzWKAJEhe7/AA/BV3P81GoOXDHi0poRMvs+2PnENEiafTY6rcrqsm
rUbff3bl0J7jeCpEb6rozlvwQHBNMUOWaKOIO2UyymQC67aI8rq/+lzRisw+KU5a
xP6sAvMWldpDXWdPlfGXmgfMFJLdXim87vVWjifKtezfMX3kM2YS/H42a7YswPIg
Pk79NOzcOu2YEkt1MjjCb+lxYIaenb64++lqGFOVWBc8VrQ3u0LAU2sS79ZrySlX
BghFH+w1moD62EmvGWDinVtFhKmpXVvba0dusGtV2AW/edwWMjuNiNrUIWE01PU6
xNJQkr4rF/5GIZjC5PPqCadhEa5YH19pHyOTf8oIv125t8VrIIqAaOHy+U+jwDYc
VCFDibW9PIE/DaqrMUKUTeA0j9b2gFSXA2tcfbgVZRojrGQz737U6J4v9MVa9fkH
qj7f79bYZl6VHhjp7uz6Ao3RZt6RzGHwmjZWt+EkzodokruCF0g+5m/6prDgZc45
wkaI7qvyvkOPTufC7/KvyAOlv39u+4jN2+JZLu+8C20Xwt2Vp7GTudaDAMcQnfMw
HsZdP6xEPQ5B8EHOJIqN/6rkfa0QojlLsL6sPcgRb9uoLFT7wr9wZQyQnhGJa+3P
+MJ4wSMJK9eX1d01wMbja7YAab59eNRMAJYBrzameqMhO5yfE8WakzuwEiFWbMGf
BtnkGOWmwpRZ0QBUVYD4WnSC2DDoGFZhQ34XU8g5d0Wq88y3z4itKYQn56bGlAAQ
M+mB9MZq1Pmcy94WsqihiT7QqYUmIB6s0NN5oPEXEEYbdL1n7iFKxzIpJoar/YjT
V+qngoka7+IFsOYZ3SaKZARrs0sj9Ai8yG6INwx3AcZHcwUyzqlbHEyeGOYvBAk8
yx3EwUk9YzAYF12uT3Dde4o4td/U4btGSKMs1DNXDdB9fKOquC9QGEHQuDTSHrLg
6ZDjfgK9PXYCAR/vuToAXyJFQs72Ei41coIm+3u67rgOwy2WTwduG5DSbEky1o5M
aS87bA9nFTWYRt5NmBln7GG5rOijAuraZ5lcaHA8XGrT8LqVk8orjbKGYdHRWMSx
Q1HdDur7Bj+cF4D4TxLLM9zt9PBWqDNgtLy7Ci0sUmsQShKbIXKYYEDnz3rowsVd
HoBi68bUs0qzDMo1iMmzhQCeWJzJfclmf3dkfnBCwdRieIsB0+B6CYWTmFns+IKJ
6g0zQ1RSqUsoAYFOes65AHbt+NTlp6BnZG+y5mB9tjDFT+my9Q7fYyIymS02bRVw
gyJ9h3dmGOYXZXvGv9+vC4knmyO4B+1vQ/2at+XAVtDzR1IZLZlm86gnyHL9rga/
DdoppsVsvwa3vYQRHCOLzYcZRsPpjM6dpMcycKX3vw1bDrxXHLRwYyrqPvuT200O
hqZTdD0TkKLR+T7goqRxaJGJy1w9f93J48WYEkEWqbeiyn5WKQMxdllK6UZNnhC0
65IpRh1/I4Z0ZPo0OigeNfuU6jL+JaCOiXbIB0MQ8Mt1SYqKbwp07KjaG28Oa4qy
af47WXLEBy6zpgvwQC6yzltZWilE1Ws+1FoshEv/Jh6U3v2VIktMXkF4mID7LBGL
J5d9SKrIcYt6tRJgMEsHna1P7/WKTg7Ma5QJHBqPKruxd9JMwRJxN4N+OLA17n0j
PoTye/LJJ/ZUbDZdlGyZpWVbOdKEV+J3X2gw2vsCCdDm+nPoXVF/Wug2YET3D3Ka
wDTRMlk+Og9ClBJNrkOdj1WfBVvKpu+QnZRA8YACbXUDsmhoD6opN0tylyE2PRoW
V4RT97TXNlqIpYj5eoao2b5hGbBtkG5/gK+b1dilMHCA+o2HHbARrvB/ewHjIkJT
1AlarIxK578Rtc5WgQFE+Gv/2cmputrAPB8p95LLma80O/EREuSFB5modtWSwzcx
5wHLVRRDxgKOBP+GOZgcS3+bxX+F/cpkSMUUCkHw36GTf+mV+oYoduAn2a/FfeNi
tdvW8ZV1n3XCqn1juSv2LzgmVHjgPgG7NTTLfa1qZWzjM57ErBnekBSt4WMwQq4m
Xjei65K/o0Bm27VoHUU8Q/ifciKuH1vg4xCev8KkjZm7XEIAWfXd67R5fVDwgtka
Ccn1LJh38OOwVFmdRRsnOxzcF+TGMaOW/iM93SMgus+RwZdzG02Fb3p/tyiAJgep
MfbC+NRVY12xuvvgkRdxvVI8SAaNCBVBnocDQAtwVw3bXn4TIQ5X5tIKgckwWZ7h
JzhgyqhwfM4kE+Y71MJH4OpaDcDlXfc3mPjJMN+q5snYSy1YAbBHLrdveEfXE0wq
UGFelDUZTF6WEh127TjdGuUa8NhQNjEiVH3Su9e0zUhX7eH3R/eom4lq3PmMDmvg
018piO/F76hm4sM50K8nN89GT6yh6RRnZ1bA0x/4RR1j6WzFiqDVBrD0E8W9NYyq
ejH4M+qnFIq1gErA0rYLpfaGjBYahkFB11r1W5GMvcIykIhM6VHsGYuI5Z08+zxq
qPjxlJcQVFdtV1PYf/+5ZXo3pvCGPVKrOjqN+WCakJgv1G/UdCip+3dVXFD4/HGV
deSeYF7LsOCG3pP61ueppHh14fhA5RqylrMwKTHyllJSOqev5dvEAOoLVON4B1EX
QCn99AP3CbK6GZXYYWGCtNwmqzl5QDI9pBtS9d6qHoTKMjztPQS98SJBY1ZKof5E
iGIaixolnh0klnnOHtsrDa5zgsJH/Q2YVnbV/v/BeqA2FVy0DXoe2Sw6adAn58Mb
09v94wXm3TjMeXiCfBgp+z5PrZfHF4EQaTQwKiRyUW1tb3aUT6TJQHWPqcxjq1Ym
m/Xr7Mvl2JqmH8kL41jSy2qd1rM7yGrXosuf+MMMtj0lFWmsqdvvfeZKJvGZI/Xt
CrkNXjXpfZ8jyFpgGm4Ysnr7laJnOa2X11zDC+gUmG+RTKgwdWLg41o4ls8sb29P
v2AaCHNUBw5a5+TFRx0FVB0WX1EdcAlau0gLixNGR9EO1OHpDuZzzAhF8wmmBjJK
VKbBxVEpjSeEHqM+EtDPAPZZOFd877jIfSatRizYm79NpqoswqUhvDOviRmQY53Q
D5BuGN3qdlM3Enfd0zk7NoxvQCVJBJz2AmAhHrc3b9A7UtpCvjIUW6jgJYklQ3vw
ggEn4KEG99wEv4cv08B/lSCKfo6/qXUu+8gLyJrXSpTz6wmvXLzpJvbLM/eLWFld
ibQnhEPaKuA4epwj3U3uyx2a+YeUjoHxWWXwOTz3YmkuetyRzk5HkVA/ZwDeErut
zNdzDpJs11ZHZbT0gublGiqdQjNZ3rSEu7yTPtqmVIHemfMan4nxH+EJIFImXOVt
kdKygIeKMuXQwX07QCtO4zX7VC6nnlQf3I93KgU7eIL7lnkcdzBcDg/x/0pcxNY8
wE6mnKXkUCZGqg4CGvpcMtCpThwkeV1I/Jj7ZBP2PMkWtXjbV/fbIXaDfhh9HIMB
K+RV7g1JKiSd8crezel6s9KVhcEwZSTQz1ZlwVbzJ2GKECc+B9HzRPfJMaWG/6cd
gQ3ixUX/vOcKz3gSwpONgUGJxqXXGUxN6oqCOF3THPG+gl98/s/CUxdr+kqqPIS0
vyr033B+EDp3QfJ0X5OEtKSMU4/rWhA2NZjDYjRrdUQoYSnz+7knbdDzEpPXhx7P
NOpfp+NTMhOX8ADQt2aUf8UuelvHQxXmqVoHbagkuJrlSFmRZBXgHscQ6u25UmYO
JkC2HhAQhtleeWROqTaoFef0hbebOvmaBUuUdpPyoEzMeWAwk8rd+vWjEubUqS0Z
/skbimwOp4gwXt9QoMm2FyzRVP40jhk7/ZuS1cqx0FQKtSsZiBt3p12KjW4oi6BE
17/vBZG3FmICRhOYfJukJ/sR1hjlMM1oHrF6/Hebn2IHR2pmuSw9Rgvqxngliolk
pnhOeSDDtgmdSlphNZbit7MzY84teoaLo07SeyddsjxPhATAHXuFpZZ5WpIXJNiL
dr6RnR8QKUMoio6p5awUHVH9BwJhrV/0TocRsSF4rmOcdHzxxke7KoMV+DKnVSyX
x9yYcp8Hsry2lNM/OldQ2GNqEKTL4Uq12pkF6tpz+M2N4cHAN9aIcRRJTPcZLPFL
rWf7MV+f/GL5yNeELH7bJvc2GElyMTzYpL2cMLVahjvKC7/LB5sNUV4jt6VMZMnb
GJG7y9XRxiYvP9yXAtvS+Fyuwb15kDCPPZuLEwGRur2MLGzbilAHPpVFT4x36h+c
4fcMPMwb/2EobJ4ueJbFXSYIauND+sKpHP89KKZFLs0EtzzkykKYfQ+ZVAzX7Ara
Xcfd8G8AuNJh2NbQrZBxpnXn4qwVsNc9tt++ZSp3TRQpkruH5EG9D+Sr4FCh/DgZ
vFxv2uTSnheRpGBBks3C+a69Gv+cwlJ6J4GuVpJmfValJnpgo/zcs8G2s6pHfOOC
ngiOmXhOEjdEdYsdcoUXSha+KEfjHqFCrikH2uYj1xuaBgh0q57W0rokrvqel4p/
PheAocYFGaPL4F9UmEUCnhFkJAeQjfrhKpVHyqZ2t1qfy4wCtlpCGSi62RmWxNAP
tPXLQVUm4EVvagwz69fV0QdLPTLu6vHa+uGz05KmuMOOEJurI4DamjqveRr2Yxaw
l2qSCWtfJwX635TGDEKsT4XjYliUe6su3aLQ9uDu5SnnxJeyTFvSxa5M1CDnOK1Y
gZayCe7/G1UCnGAtxncd/xmX8fkxoVeEsrgotkFgANI42VWvphSY2Pjx/JxYCxXz
egX6M8YiuPrijgveu04OTw==
`protect END_PROTECTED
