`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O9o0O1ZuFm03eVr4YgcvrDExj7znP1XXLSDYHH1/vY0KBGmbsBc4Pj4cEix5yV/R
SM/81qLul6MBHnJ8kIT9Gs0qMry7fO/xk0ZzDu0T7W/oV6b0wNDeB8eBK9Utlrwp
f1Htrh+1knkP8alB9VBAZBfR6kqEMSvumQrO1FlUxF6h4B1jfLnHDkH26bT9zpyk
+nLKz23zRg0TNmvRI9W+zFy211RdTzINYW93SArAkNV9zmkwz/5hG94zOpAdaW9N
oEkPA+EMgJlNFGfCEkV4sw==
`protect END_PROTECTED
