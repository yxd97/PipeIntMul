`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFCGnQbjSkP3KiG3DM4lAmkbtyMCrrzC51DVotW2rzX3fME+DpjoI5wGlHSagBp6
RVjSp2LVy83chdkjJ8LGnRfBLa+t1if5yMdTxBuMdy04DWHfYIAkqrxOfnMHwc4c
i5/pfAIuNQnFaZQDbWbslsUzl4pm3L49IDSDGaYGP16sU5vBh8aMCWLhU4M/Zy8f
AtxlueP+g4NIlkrlJ2VFKBZFRwSsjOPHtiTqOy6gHox5KP65YmdDYpoKqCg1ua0H
riTvUwTRvWsnv8110VcFmQ==
`protect END_PROTECTED
