`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rh5y5niZIV7rX25zjwnme+nkMpf+gRyUz7bbaw+IBlFZFJPLltiQzjaaQUo/0RPU
d1t+Ka57APjioIWSu0FVJ//c7IxhWnIkHXjp0w5AzbStn7XlmFiN1evPKoKCJSoT
cJ01AOW5jQ+b2Rk/lAmtfFqfBtM7VTtGm5XuYXwOzvmhiN8U9ZxEQPq1bin9p5/n
5usmhpdHgv6ZmHrF+ut+jV/UZ6OMz5fnsHrqewWHW4d4oYjAahtHCrD9xhOcVkLt
swN/GwllrFtLotd2ksew90LHIuBVsI38RUf9kIraoeAzflg7iHsR4ZPNkGgqw4nr
3McRT5yj4sTt+kHG2TA7UzKZF4E6nX3sifKFQGKnqIoMr2qxoWZN1EanWXVOVRFP
C7H8+0xM0aZAeyY4pHodYXj98xBeRSg1IntP76thyOekwdsReHN0TjFc77qBXuyd
dF7xWSf8WW+3zRCcCP5Fqg1p/7LpQnoE+dIfc9UcyT0bHgTZs964SpDTRGZd4M1n
15KPWZ3MICPy6U5D7QxtKDsno55wQA5bgUlSlEpfjzI=
`protect END_PROTECTED
