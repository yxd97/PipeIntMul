`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1z1koRSeSkJAtwR0l+GM+vy1xVKPVVUthQ2Yqjp0Ns5ixt8Z+qoW1350topyp3YE
58/4r6KGgMsQc/mhnrWdwsMsRIV1uzEaPlOZ5QSaYpcBCf911ifzCUVEEXIBgyBT
E+bKIkZbFWG4NFldr26ome6FB1FdoiizYJBdrwrT1dVGruAQwXp9cuKngm9CxGwH
doq0d9nVncDAyRDXQv2q/fnT6GwVW0iLCyAPoF3FMnDbMqHTPtOmbSIrXzEjxc/i
Ppf7JyjvQYvDGd5f06BcfitDmsi7fu22/1VDiChHYAMaLT2M7jrrJBfSpTR1qgp7
RdOr2QPYyFfFjwfehwZCQY7GP0yUMBh1VxyD4O5oRpLz0xjAyzI4lp2/sZxCIe77
7ogI3TN1r8gNjS1xnMSbA//5d2OyDniAkVe6cKwmFs0yJC2eMHju6TrbdKF6aJCO
KBv45xsVXxXbldToS8lIvBSSlzWTzHIT4KlTt5wxgY1tH0tmLYHx73+1evZUf43H
M//I8D6A0giFwOzFkDxDHCt9UdxxFIKq85Z/zLWRvQyyHk0bsjLRg4sAkQIfE4GN
vwViIN9XDh0wfByVB5lQ8O0jbP1p1PrTL2uJqVLzlmft73kKz5DpuUbk/x0jueCV
5xtJovLLMS6OxydjT8lAFi8dTgdWQDLja+OGvww0EDOOsmCli24dmRrycyfmOldp
NoX29vg6Ks8FcmqFVklGYoLtWpFKNjH94z4PH+Ux39OI/kKEFz0OrQuoCIRVx/AW
5tp3PSUW7QRAUqENaR49E5UbZ7JTgxX48Z1kM0jFLhZgcVOGi5FFhwxBUxVyY/sI
yfrWv2AY300/3XMIy5CIZOUZMaHAOJnhvoU8oYB8XFg=
`protect END_PROTECTED
