`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H8zESWAhAri+s/IIYNef5XiZrlf1pGxipgVjALO5w3MqSEsVlsQ/Gk6WuCNABm4E
G1MDsjlxwedZ0g5lgyd/y/+4SggSicK5L1yEGUX/nmoZ4usflkWKq9KxqaV5NWtH
2P33lAbDadAp8EEXskQqslPqPeQAOwZnzA737k+RPlvIoRHGXN6XMaizocFqDdVE
jB0pSe3WB4gVGpXv8kX70nsw+9RUqiqS5CDwHVsDiSWtmniJSusUdg9b1N2kxMhU
ecgL2YBDoXj5PLlnIArTjE8FGWP7slY2NXArbZRTj61E4cqS1Pd1ytTdVugwAiN3
F3R5xyMd5yyAke1bqKyrzXsGO+qUPHxQd0draMWBVAtdhnHOMEDWPGxaN/AGuXoy
uMlns+lF3E0jBgezQ3yk8xK0a1P5NW7u44gDWidhdjQSCC7IdLYdUtGgHwKlLbDU
Mjk3G50f9elqqdYec7lOqkUkr+4GvWYqIqYchyQgwvvt2M9OdYEvYeqJakQkGeFX
hkJmx1I2dCTxa1RixZvft8GSEibX8GuunKYBg9YHVwsY8WBrad1yI6cJuXmOm5oR
rBgIXT3dHq5LSUkNl7kWwxj7EVmybnR204mRmeW5zU0=
`protect END_PROTECTED
