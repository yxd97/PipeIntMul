`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggh3WIpdqj76/Vqg3PUSt6laDHBtmE9r5boHd6qYcUrMkVS0fM0DDa0u2hCNWBtg
XzBqZ92tiTNpGk2lsnVLVTs+DEAGcE3L4mMkDitTWuNJduJhWJkASj7tZBQmFLel
vd/oYDv/vSAnfyOKf/bhO3Q0YT6wEi62hI4jk5M/zyp2pYLKx1bXLsm0JEDJdJCo
Jg52bKgDc18icDRupmvr1dSnJ/5RfAJUtgSMPrno5QBI6tljHj7wvfvfZA/Ef2zK
02ngbCl4R7YvDk+SlkTpIKi8237knr/09frGPUoCqWKUJuGb3Gx9ceMVjcOleKVr
WrLx1AAojejB7ComF2qlj9BHVzGt6QvX7O+yUutzK+dc8ZWP5eiHUV09sFYLW29Z
I8ueE0aaRVdctFG59vOlKNB9fH6VtAJUK5FOT9wJdIPhHjhedubVg0DFd1JqHl+U
+88eDfVjrPPBj4BzyC6Y+heisc3ircoJQuryka6NOUs=
`protect END_PROTECTED
