`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJ01YEu4Dhzprk0ZTPI5kpa8VCwGaQbtgLRgEMRc6V/2v8hOvgBvNeImO0Ua0ZTH
jsQ4erVv9EVtjT/vZUoxBjIV3aQ138FFs5u9K7qOkLVMdpdo6E8GwKChLom85JGZ
AVlen6T6Mc5aReilzqRj77NQIOMSruG2U6ffQ+EMsBISUYAT1ddPlx9UZsNGXbgz
dGXSa8aIuslTRNlN4nw3g4zkstWop8rhCgterjKLuKlFswceLG5kV0oWxvARS7G8
pQR1wP4s4QIovpF1/k+tPPi/04vA9SsNIl3uQDefJLRT3lIYaL5QbdAv6ijJ7FVA
yVWou7XairhvpN8u/GbMTq4jH5IQ+l8/59nIvTuK6vRzfrjRl4z5CLteC4AetXCq
uS7pOgxDdiKfnuL3IhWM2w==
`protect END_PROTECTED
