`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bxS0CM85YX8Wz4V9VPfejA/JzNpfgn4EXkNhhsxFoxvHw7+fzLbzwjcDJEX534Qs
3vL0E7jxg0aO21fkzTY9G8JIF0cada7EWSlwNPW2K5dn+qGWcPM7lkQhlPabJY0D
rOXMLVE6Ycow4iu0rVL6PI7RkAO3W1RjbQpPaFEmCyp+I5lP+28ebK0YXS3hl05d
Lz3dlx5L2cTZd2IbbB1AIGeJVEZenpn6iWXmgtArlEk7VQfTdQkNVbGWn2KRYP4Q
CZOqpT5KUD2TVu7dobS/nyVpSJlfZLZ2B0keJtoIGwjPSh0R3GGPifiwddyqzdd5
SzBJ4OzFI0e5wkXm4pSYRw==
`protect END_PROTECTED
