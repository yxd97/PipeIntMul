`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJ8YyK1JMJVLMOMTanDu2IgEhEjlux5sG2WKZebUCitOMdYGHB1u2ILa3vFiU1P1
uYIF3SphsuynDZgiohw6f6slLvFaIFKE7YS8DDxOlbUPYh+p26p/o0DBGZuDHkYf
PtE3GerWWJX1HT4X3VE7ZYOpC7Lgh/afZ92A9zWrRTBUFsqel88w0yOLMhsTMr33
QTfAwdgIfvVHmTS+4ebkEyRTiXwzkWQnp/uQqUaPOf7iUdWo1rSICE7tl6xuPI+w
ZqqNv/W7/cd80RKsnnipKul5aN/6JefvTTmlzcXV3ZccUFr6KfEN8XnuueY3wkBz
cuU57+KWUA9DV25gyc3C9VgLyPjIix9sIbzGFwBPrxKObadBdf8lFBUEIQrjJjrF
l4FiL8CFxEUcHX+S4xMc9tLbyr5mVaptqQClJ6D2p+CTZhkDvSwTz1mOd4Bb6fqI
1P+kWVo+kpKL2by62SMoqQH6uLzlKsmnGomywbglc7AmIpgDp9ZNNdIbwrw3Bqeh
sIQJshS5EmghlbkR7GzK1ACXGFLknxpFrDnfz7Hn6LL43LAdLfHAABevwWLPblUr
`protect END_PROTECTED
