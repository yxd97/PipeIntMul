`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vs3JpJ/JYV6jojv+WITaudSrm4N6n83f7bvW+sw5ZQSrZ3zfNYkT5zIX3cw1VfVJ
MVfmEdzIFulpSnD7vCVKwdMcFJeLUXOjZ0pj0BsDQkR3vp0ttpNkSfMpdNKhc2Tf
TDQniePNvVXmSwl0hhfJSqjBrxYnGfBmsXFbukBxsQeb5C4P0YO2UB0VaA8KSSdU
s2ogLI2gaWDKi60ZeVUYieCqMMjqpq5kbJOy0Q2ubXaJ0pI2yHMstB5+SnVrrb6C
PFrOW2ZTBRVvnVKeUaLe9LoseyAjbLlXDI31oOnC4KmLBsAfc57zi3JRQLkLOwv0
surjneB2eE/23D4oQnMLeE4PRdA+9Tjw165RB2J1xgpLZOsKlQXLNrTMhAU45vDw
P2qYgPtfQOry6Uuj/mPlxcLDlSwgQx6L9BN3nZE5m23iZop5+WhfNlYTyQWP6ljb
m3TguaU5rLLVxeTFzukFHhR/ZoPRyMJziP7HD+s6NM4p4t67jae/w32QZO8s5wFx
3+SQ+Lgjc5stSm+kPOgZveUs0JoQ77UYK+ya4ddoaS3NHie7fGzP6ddRQkOHimZO
Ynj2DxKDmGBYaMbexWFifNvJcXC7CiBxohS0qnJS0GgT8AxX0cFUDiC3uRazxApa
pAqq3sqD59GJk/QtfXWwpWanpHI5QeJywL+eUbBGWGA8JbuH9UeBEPiTrwGQjpkW
rSKmmu6Rc8dig9xU3Zj1gPjPTnWrDtTtyVAt83silBDH8RTpEHohodYJmCuzQyUV
L9YH9gCeH3sc3DIJrhQAE13vl9NNUNOt1qs4FiUN8nq7d1aNh56Qg04LsQq3bUeW
4tcci6A36boIhLeOsp5zjtwiLStBX0xVfrWJuowegGRIwRzxg0Tm2fkiSz74MWTO
9kfICvnWvI5Z1dLNYZymTvGgJNspuXhQLruQaa9YMbcK+0CVllbEF8bBsWN37taL
z5R6n0OtR/kL4f0pTEQXJ8SIGdOGWJaLlB3nxqcX5H/3xBb15/At/U31o2vwIc3i
dJoRZA3GN2S0a1k/2mNiw5BGAfXfSDmt9q9GHohxxCo227oe6dgXg3KRL0tYp5tP
NRhI22Yu/MMaYDEyVFcUVrTgTMK+SD/artuTZFjoRovpK74qeqS+6+o9KEGgWTKD
PbtF9462JRrU3nu6OXo36WUKqoRZLgKLs/6VQZ/PWVzGyTVNNN7y1l4PsRV6/awa
0wE+xyRXTOV7N1tpiZP5/vmKEzyt1wJsvGZwdaryb2nhW16vLdGrdyrdhNUI+rC0
3ATIPChpqcPBLydR7OwQnDHdyIZ5bOxVVDnf/h9skKSTwrJw/GvK/KkIpKi1A9Jr
z+6WY2Fkb7sZztZHVaGEbOoe233VRJhT7bzYCAwohf7HGLBLcKurWN48AtppmpPi
DYbeb2zbsRovWuzcoxb5tJ3RX1MXEV37tqCQMINIup8t9ECbXGErao9NgcbOsbsg
LVRjTsgPTu4DvkRalHPzFUcAqpgg486MTBAqqEDkEKLv+1XQMKhnZTLw5gqEOQs6
DEQ4JqYX8UmrfZGBfsnqnZhUcYB6ZaqPR4uKz7T4yMTv3AEIBXxpgzETHnhGPckf
gpCCxY2p/RlyG9FuMWNlg/xCoZq8Bt8EpOm+TuLU3rZRQ03eEeCprQvtEMBqJgDr
T1M2WG9DnO93mduVHjrgRQy1XhwQ6eqb6ngT8PRxiFF4LhQ7ETw9PTwqTqWUAk+N
Qm1HabByY0Kq98M+uQWNxFF+ZqVLlxvXPvE7pUQKBhfSs3iSppK/epGWqUbEGSBa
HMddtBlX2A8xqpWeI7iB9ooEEioU8Vzh/Jxq7etqN1lKTvTeXeuOwJ68NmfqQ197
PYgCM2OrD5Lpz7KdVP9kVuVa9rcMksmMwuRWz7BGD9FAWEaAgBi7ZeaeQa4umoyP
mokYimJ5Nib7UjNH75cV7CmqlWHHpfULj93eu+hBVDPEQPyptlTS+t2Dkk+t0Vp/
`protect END_PROTECTED
