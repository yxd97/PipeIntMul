`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qj2zIKNcxKCsHRhebH/olZoDvAjuaGqqMMeaNMY03QoAGQgixrzhD78LULK5JYU3
kaejMzgbRfDSUGbVwZlNFJ2XyUMYiQipMa0+uE+O4uyU44yuLnaQhVFFXFeBd774
30lXRxm8OI8PwN+XCRbHbLFgaC8xpHe4DZLgCTpJa8xw5Jc28DLi1yGyPmNBT2k7
WuX0/hr4tMd8KxSAEhtVaSRJ5hUgFKWqIFOssECuJYIf8f6k7l3yVUPCUPYON5nr
vfqCQvHXwQ0glGNzWkOVrXguS8CcfSTinhppcOFA3jwwYSaphYitXBxzPaAKTCAA
wimWRNSLmgFSsqnya6WctklSTndrnyNUnO/u5vqN2Z3bx5mrnCqmYHiR7FRGcwPM
4pwS+qDHCxMunfZXXzIs4yAdnztugoI7R2pKdQZ+WqKL+MSarPkr/6HVN1nHKsKM
kukxaCpLgOkMVRElg7taxU42TR8A7hkAvPk+hThU2ufa3BErl7TPr8BX+sONc8XP
1H8mBNm1pH6rCCQzkwyQs4W5YWQLFUi1LnzbBWgXQuoMaruVcC1U4vyOdCnP/ta5
q8R/7M8Ppvo91cPkBjoCeqRBB11wjt559lZK+3ElHPRTiMJ5Y3Dnjmb6F1twSNR/
ITryKtVwFZhI0tfjT41xdFc27+2DZuLYV/jSvVUR01mkS48866tvIWDcutEx875C
gt+6dgWLk905MRwxCF/7IRKIvRtfKGLlhEYvpm4kyjtNMZdb7z+n5r02XT3UhY+b
r9ShJflWFvWGOH49I35LY0Yx4l91QU/euNRrz5jO0v8RtZB1C8a5YC60runhSJhS
`protect END_PROTECTED
