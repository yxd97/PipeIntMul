`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t5nxYUWiVEr8XnmFXFIQjItXWLDNQWZV1+jcPKuzdnzr0Fk8ejjVBWc2oSA0AgHZ
83dUuCcVh6RQeOUOQPR4LUJ4k981KoA5QMoT9r8yVxOMT6O9evQsxuK0A6e3zOC3
85U4o9QCHK3I0ir9KMUf9b2C2BGtCF3Ju/Hj2kCwUtrXs5Xs7eN4STNTdWDHo99G
9UVpvvoKlaku7jUcBza31RyQZdvSZsY5VIa/wub4mHfS+kslwxPWjYh90kPD1/aO
NJTRQusNABH9cxe4NConNJV/0BOBEZ373mBSJB+zc0n7I6jmqqt3tD+XrlvOuOAS
vGjlts4uhA0BRsb4sWLOue9L0muHAwlExPcUi0rD8t0j2krl6cV/TZNB9CQbtJBD
ouliRgT6uWSoiJZqY9vnOv5ynbrek6YjLaZEjunIzoe9ZcfhMJQGb2+RpIVCDoaZ
N2HuFkjqG7PIq+JmtOM3GvLe3ckP0k3zuksDi1clLxk=
`protect END_PROTECTED
