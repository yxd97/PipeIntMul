`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
amY+pJebfD2Q9lz5RBXI8C9St2C23f6UileI30+DlHpSc71pd5+MpOBb76jc5j9N
bHDx0L5J/T6OsbIuRd9shPPitRWQT6dKPPqAjaGERkxf2cfVrGWtoMtkTNYGWcyn
Ze26o86tEosy1xkDtqgtag/qyfcnQol1qqVz59SGf2PNDbK/br2vn9pXQsLfpGge
T2yXnk3X9W4CEntvjMGgNBeOt7sANYGZOqzfqFDFURZ1nEaFBJ37YiWBrEzsYJLO
BDo8BOzRQJDuDxAzNGjv7udCSeb76VZTaUXmsI3PS8JB4UR4/boxJyz794GsAGP+
Z12upyCqih6a5K44e2GXcGhsH2UBgEjwwtglUh5xn2euaO1wKaBypfNvtT53VByZ
Nksovysn8gDF0bphJw3FOEhA+F1trKqyN8y0Ow73wKDClbpdmJf5icos8KI+xQ9Y
UO/4261Hrs61oRzVCx7ugALyZ2iZm5aAOnHGQsJxBf0=
`protect END_PROTECTED
