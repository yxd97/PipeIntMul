`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwvlxPjIWPNNukCVtdqmPyycj0G1c+xQMMxhWcOuB2McConJiH1N1a3N6BbVblft
gQJfL0omYg+CHZV2hXYz2f5upbKLny7nmMPK7p62bNLtpSFlrsvrXX0E3SyfXkcu
PTNjjn6SUS+N0f7IKBKnOeUSc1qH6TG15dMLwm9PYDDVJ5VJiG8sOndGGP1EwmMR
xJWexeYxcMywWIBTgGTdiAElziD/Fad7o7b5DkYvvHdflsJhpAP9QPqWJq1P76p+
uiKNHLHdUvUEJAMefXJ7eKb+KJj2NZi7o002VcHK/akUYdj0mitw0HXOYWpYJ1lD
HW8p7X+A4gdaeFiXAJ9h/gr5UjLBakKhZFfY0hfLX5cZ8jn+sz0LytFW9b/GERcZ
LopDgUIFX4c40oWjdguSlk9tRr1LrQz0LT6YFbuZzHygOeWVN83snSBDJt+DNqk9
Q/i5HsmcagqMs19hk9FNG3bfPA3ugxoiAKyVYb87qxKoU6U5seEw8XuNWwXoj7zQ
H5r/SgtTdm81QjyXeLQKvliDa4AqEHAvdAPkUGj33kk9c18Isrbckp3EiqU4HbOx
`protect END_PROTECTED
