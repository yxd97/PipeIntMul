`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XZOChJiqRUpY8QUKB2lbdbHDfaYD7yE+QCGlwKQ6MHEpuVCT3WUeVjGXdILQ0dm
FxD+eOsxfVqr4c7g7POjuBwHhjS8Qu3hLkgU+lSzKPLkYut0ShFShK/laiF2rkRG
grNQPTgpMU4+QI4vka+Z0StlvMtxP/nEp9pAX5Mxjnqw8xSqD3RVrVLhOk6/Sy02
wZ4g0/Rs/19PjcGAEHTAyJdzWsWBAFonDQboNdCXzkvICdnzAyWxt8sbMp9DWYQr
P/lboBGZTEyiJJTAsyNccIisbJBrMI1eYDHChP11ysN5OaizB9DcLwtHVAAxoB5I
DiJcxB6zOlC6q374djVTausT2EvK6ZvnyVlHHwMe1U//T9PIOx5K9kCb3IUdcJBM
B8WhuLerh9Yjc3k0/TR5jlq2/5MsP3zm3dpQNDSJjxgvLFXqVyF+8Mx/7zd1NiWm
Xp10BZ/3y6lXgoqWbEpLJqx5WPWCFZxGoR14DutnDAHC0OkEyyZG9GBxPC1gatNA
yWAXOhDmEMnpL5LYKx6vyJcx8QrAHf2IcntnaYStTpPf4TKGwZxXFIPflTPRpOF+
M3HIifmsRcJFnJZ4txBG0xkA+UD96H6fQtFZ+Izk//OLBBfitVxbarLoPKpuUwJd
6CjrNp2i6/bXMNsOIgN0UeQBqNNnaNjSzdncFi6iZgvPz4BsjRzhbhLe8tnVA1Mo
YDpwCJJsvzpuF7fEHc2z+HL3D62l38RxM+XgGgU0cOOrH+hLR8iBui51iXfH6FVP
+oUJ9tLYOqbL3N4jesqQca2HEYh2gdaATZlrGpdu5YtdF96U+e1CBy6r15ydJmoD
EX9STXLd9qXatEyb087Dl7ssQifFiSm+Jby5evaRTzoZmm5Y2L7RgK5Poxvog//u
mtlqFFYPevDEmaM/HQRVUdHXGjUkaaGp671bibtbqIczuNoPHxei+ImjvjO2P/wn
g4TDaS1baoTLmSQ4IpxGq9YfH6vFggkna0s4ANOlqv34X/po+FVFOhWMuNqGAgGP
7at64Vle0qbKMVtULWjzij53Gi32xKaKGDrX79kcm+DAzgrXBroHXn+QB5J8dH8C
RQ5EQ0BwT61tTUxPCsyjSo3aylIUEv3gfJUtXLjogaQsF5MjkhMWJPltsjiDuiRA
Wg1w3jv5gB7M8IaPX/AuBLzf+emi33DrwTjh3kpB0C/hltQHPU0SLynygqvsVSDN
LVpQWNU5fTK4M0IktvYutFWZjWTvPfJTfafPOd3MWHakaJM9+gvE+nFrzEFtHWcp
F8XxBBgUKYsLED30QjgJZtNXQwdh+9Pz8qDeH/g2D/aigyrpTFYZAzS5xRAY/KpW
c60yVmxfcU3O4uKjo0a2pYKQzNB6x4O3B6il9EdTF+UawnY3CMwTaduYB7Z2VbK6
ed7YKsOqUzMxYBQPB2DnXXnse0y8dlxI/ihrSzHmI3e+dZvKIVraOlZpdusiZykv
BOD7/nLwipzDPQoVZ9+Foj/yTJuqL2ljzPNyHvHByA+MB4nm9yVsLr480LKxhqee
S2nye/EISsw3GlDEQqL2WDXwZLIERBbRIZ24Vc9TF8mu7t7/Bs89HFW+E54U+Oeu
KWXhADzvvrOKIBDEt3sGbshM3Bl5vqhd5+nNzjDFxiE0i5kRY4ctKkWmpQ1LAt6I
lk6+A21g3WVtbX0nBbo3cPg090hSY/B1qv6pv9unNM68QrjeaU0jINRVzFxfUU5r
ibLLj1T8YBCLTQrFdDUU+JzwKqrbmCyUBzVqPcnhpdYRyx5IwGNY+fG7XRZvaQkc
W+YGZ8lZ5qOP/2eahdjYX+BDTj4rzWvbP37V2UN6iqS0VhPZbe2LAS5LSFMvvzLR
AO1D7Ic08pJMSWGh84AvJBzSKoDkZfYbOBnlJEEaB7uS2QWoc7Gj+3/7C9IEQMwt
pNYNCJfuAybPQMjq4eJI62FZbeenJ6dJ6TovYQ8cpJB3/H+OJum0EBJ2CSec8dEX
SesGPEgjfsK1bPq11fsnFCDvVQuLKIpJHkaE4RsayhNTlhzHkhOrQmmECM47zZtL
qmonLGTb29RorDJJSpiys0EGh+EPcKdWIcnDWfmbxhXXI3fv9DPI7B9U3yx05dzM
mwc8AYRQP/I3sjZHgrFZrkbwfM5Eo58vdhVabqfdBXTWP8zg5YrKpai5MoKhrV1G
8Dpby9zIJVJFEB/8CkHi1sZlhEuISzl+/hsgV6PSrrMKrEDqtxpIRgxdC+Liv4fw
kyAx5uMJ2i1pygBFaflOqmz0LkYz4CY9ctBKaEbi98oLyVtHmwK8UCY58n2XWEPa
FT5bwGI+MicA+mS52kQYzggKVfPA3CviA4FhYnChjyadSN8rL0o3nComSA7chkYO
L/LR7zCgZ0TmGgxrc62NGdoYo6qv8qDSaSZSrE4ps4r3BUGAi0pxOQWn/C5XXfOk
bCKaX99G9UsfAHCFc+14MYxx4STaYF5U6bxsrIifjpyqCuaYGfBgX5/F/w8rojtF
j0NOpEou6p5nZHYX/0g1Nt7XP10k4bAfRCYFsT8lSZs6DRgHSsJnaS2l1a2brGL9
E47Bvtj1YiQr2YlXDdNnU1PwzfNEJ8YgrV3uugVZJcxnGpPgkPFT8lj5TMGbppUh
EPdfNGu7rpO6C0vBEZQDOP2WMIYQo9e8D49NH0hIfWl6MrVmdcFNqdc/pHw95jxX
jVUTUCGhhkCiv4MZMW/5jndWSV6MQ9AG/eFJ+vQy0DUOw4aD+iHMDbEh3D/D9YyR
KicfUO4PPqQiNHaSyiNJ3dhHBweWHrrRjR1vTSVnlWhghavpw9TnlQOWD9guXxBL
RY1xI79EuYe23ZATyMH5zTAJzBApL5QaENusDKS4Kei36vvVtxE0MfbtsHWxgZkI
nZ2wUKfZHO2mpALIoN0gITFZ0KgWlRCfVptHVGIdLRPMo3MTLi6iRd0yL6e9W+8r
ZAem0WgGMpU0jGazYT2+U1l0LGSNZiGaRxOPCtoqi9ZKvjqT7oFBdA3b03Wu7zkf
HK0QystV5/snnz/ygZnLpu6qrwjD66dWMgBsWdtJfufSCqi65n/1vuIn0Nj8rEEt
QIzxs9BCjMEzwqQLOqEb4uR6MRW90N6uB7i0SIxWLBRcxbrGJQDqbHc/p0I2iIns
tAiOhT23fnJ5VLDVNlFB5aX22a0R7le35yMOClfjXde0aOD1jbb60oCkoOpYWiM4
jVzUPJDlM3wPLom8yWIooogQSJ8cGPm/S854ZXOmy6+MGYQRvD14sgv1Z5WZ+SH1
zIBvy1p+KWXhYexXqUhqLyztnSYSwAnH1Tbayo7m886PZsKdhn/wb71mrWdFnEQ4
QlKcx42Aeq5MiqNx71kLODW5luuYUD3lZDQ+9oIMzAq557zROzxQJUmHeYF8bkNN
LJhi8oGbuwXcgYXbaL7PZfk1wHshEEUd1EUs0QDWEqxEhCkcx3xXfYvnKC39eEz1
Vsn5FVBd9Ks3dFjOxXLaDEEI9H+p97ayDOvH0QqoBFbyQo28woB+ZTe00EllXAE8
XCMLuJP18EH2WkGWGdGign/VPfp3pqCOwX2oa8F9i57hlggUtmE4p3xsv0xmCzyO
KDpnvQhPe/UJPbw+tL+urxcQ7jPV5pMUnsIjE+xIwjW6gwrnnGMPKdiItVG2DTNN
4uOn8l/tfDlh8TBFez0q8YL+NmCIH2Q7RMkc1Rjb4t6D85lfTMnskfyrlR3AcY5A
KGFFGrWnSlIlggDt5HZv74y0cXL69DpFhG7cGEfQcq+4ANDE+5eJVia0FC86nitn
tSuoxEMNfqinDNIj+n+Op/KEo2yl81nsnckl+ZrQY3LQsuaLj6D+YVh8NFGFg7F3
HVeKLlptXC+5IzE47yx/pxYemHt1XPPx+h7CTBmQluzj0R4nzIOdW9YrbyV63E1/
xxJ30pGgllb2eJiSLI7VvGSRdTzmlWv6ppmmR8F5X7/5o33g/f31Ua3v7xDq+37K
Wtnl5Ay+INMZOVs1Ry41LNYNlmHXS6Rep1RaCbCW5iZSGCPugoltMLsr4xYXmGPF
q+I+ZjNloin9H/JzpGp16YCHNmOxOlhf/SvczBiXRdjv/EDeHjcdjPGUpK0C3BuR
sIBxf6pki47PuCB6kzUXRU88I9Eeoov4RWISQlUmnXgSscudK+6Lm6OwSF1iYowF
qN/XK00AAIZfHQbSDWck4H51YE+Ui/VesNuk7FP3OmRa+aVLwJRdZ0c50zC01oCV
X+7vXYx7IyM3Ss3tiItO6FhsvIqC2Fo4bEAzLZjt4luFAAX6qwCQ1XxlQUvwuto8
R1YtqTXiDGv2QE5G6zw4rW+3AWuVo0RkK4/89NRBaiGDiIJ+7ClUKsPN82S1HCR3
NKABeqkDHwJiKCsFQ09gr/+QFcnjR9bZCZZRdIqSDn6Tobc4CGiye9BTMW9M1otu
LzQootwHPI5/q1nQuCK7R/UsniS02vOYlkvbsEaiv6mhQ5tfi3NchycIxhr5GYH8
fYAktuHXW4F9QHFAG1mZqzqqyyh96scQChdwoQci4YBT9KdVyqTHC9pyRGkQ3WVP
uKH7rGaw2Xg0kABvrE717dDe9JHVpkPpk+83VmyhKmNKl7gaBo2ccMsMdM07/w6s
rLS0r2Vnx0UtUCK4QmLJLoYboUyW+QqKrUE4nqFLlzgjlALaLHJKSNxeUC3W/5Cl
Cxg3dM7/4huxD1uHw2wbZKNvHcEWB8wt70N6agxc1NjyoweEtccol9Nz86neLMho
/VNNNN6xeuGAPeh1PclA+o0hihPwHGA1vxtg2TfWk+QOSCqazRfP5i+kBu7QC4LC
lTjFb7mirc4Qs8/N/BtXtQ1mxP5m6OgIdUg2qNvf2u/sOQM7HXImi470d+qGtsxA
F/F1Tow+JiUFaVJ9/ulVR+Ca1gSBjPoYYFucP0uCRcOnH07lQpa0bVIN12NP4sn6
MtLMmSWlZIcPumJ0OXE6GA9bs2VpPhJMFHT+L5JmJCCjesZgsZs1H8pAUhixjEbQ
uiaFYMmABFahHmZtD5bbPPNE7x6xzp85cWzbyGrix4e+YAtZBF+DF5R3Hcr2x0Ti
TYdOcmpG50yTdlQTgqAXL48y5DdSl6bwQIsgYnZhTHxFevvYPs2YBhkXKpCYLljf
CZprk864o5jX1eHjft4oY1hCydoiabnFgD7D7wr8UwzNmXn5+3qDVosHGvfvaTJu
z78Eb8KPEK4AfMnT5ECXRQt3q6dKVc9+SLq81HtEl0CHVxBDbFr4YAXSuoyyKQKX
ZpB1PwYVoJlE4uvmUobeG5vDTzoX4KEOr3Kvw9MXl0oKlCRU8th7LAgClTtQmd6u
Ck0rsxOMhaTZvqUnyVuEEFDXEVuOKWFoPfeZx9+Il8eHMYzJJyTcycG+4zhOI2rj
ijQQqfpvAKnDsy2p4bjHUWyDEiS/oRw8KOO/OdzMVzXqF37co9pSUKFUNwGDW29h
8/YE6Uy+SYYuL3m4Y4z4hVhhmoo9rZzi2s8YWbwOTQkteFSGW2zchJ2B288KlicE
6g7CbZlP1ayLZiVcWW0gGv0SRZLFw8jw84TFdAdkp5a6A3/PymP3Nfm/6gYI3AzW
aiwo+HlOu42OsDui2NRaDOB6T7XYMBXMPz3Q46gXuX2EKsKWXCx6xaMJS4OdfXQa
7KAOBzczTZGpMC5W03qKcjayGVWLAMoEKLuvdI0Eb+nvUdJZohDuRu2yqcftEk6W
QSyW1J9HFnDWkT/iNJnvQgYgx/elDCxleZqbQPQUrYskF5n+mVSlg8nvQGA3QYsg
UF/FmSvEi4smiyPiBtpVji3tkT/yZeXFW75r6EhftaeJpdv5VChkvl34ZyUTw0EW
qiEN9j77dIzmsjlSbWT5xccIHUOY3kEOPOykJgJBjKSMTE6kzOY91dsJqyTzKMc4
UD5ZGh30qgmaTlV8J6AV0pLM3YJUcRkE63hJRWzUsibpdx2NlUPh2h53ekPqLoK/
s/8UkC3mYto8icGkFaQP0rgzIiFobrgOO1VD5y0tdq6KSLqT7EbJIGpDvE94vCpa
Mcou3xRyb/YVK26SqcoinIsBQxUk4ShUhXX2U8IgRu2nk7n01qjvDmG6mN9fSnVT
ZfVrT3pn01wc/vGTkb3YaaRcskuXDvlnCsL+pHIRi6/NSb+L7Y3l0F+kQUNYIPbv
zN9Akuwrpt8yW6zdTXbRMtBmfyoziuVK+agMvPf7NRLgKWWbQo6BWa2jSRXyfKAg
dTraWi8QZ33gSZNNjDYcPLhzKhhH38Hl0SznPV3c/erj4TGK3oGe+/a+ixC2q9KW
c/hAH1NdbxP8hYXBU9xguUHs22ZABBpZ0luwYv7OCmN1gt25gT1HdyWFZGlfCgIU
I3Qgg70vRbYEMAmQUdB9nWKCwFqhEkQHyXfxaYksOyUtOKeDtC95sVYenoZ/6dG/
lwIzYOrkpFQ42B9h1jbTUDdB7eDo5689Q1bh4E+hGmhs+FllNqWg+LWo7os9AGeo
Oblyv/mU2pzofwEcEIz9enZaxoDaZAKoOR/kI8zJTqwGXECsvd/UXYGxfFVVEdfn
dfpNJs1dbcj4wxVNPATrBHEiBJJMkm5CBHnIanszt1zFD/5GZeO3Mm39sUxoib68
X7AYOoIljU633NxUbZdXmWHKiDXwcH4KMKI87IOYz7YzHp+KuPTfgkuxuikFQPd/
u2ThNlT55ZD7SM2M2VWRiLoyrx1/ifPly2qUnMGAtLi0u5h6nfTI4xt8N1DM4H/z
4NHvfvEXMSIz6B8tiNFZOg2557wVxwJA5CPkzmCvRtbyUHc9CsD1mfOF+/kk6Ur1
lll8vFsdexkZaX4oPGLk682bFJsEk5iRGVdMFmZdIjJj+kZOuRIfUTiykpOR/77i
qjJ/HYghheeNonAi+8BDsAFVedByIJBRqM+TNHKYlK7xZhlXNhjthoFQyIX6e9dA
fGuVqDT2jGm1/MsqYjFtKC6rnJBkUaHkbh/jj8piP7MMI7jMdzNvYoT7B/tmHPEs
qk2HBIfK4KwwY2RIVlVTes9+M1O0stwOjwE83KzIfC+natqN4q7weyYwYQLFdiqL
di2nTWyUkaeDM5Zx2jIE4QIew2z/bj8KmOlfb21g8leB+0HAaMkNy5R5sQVdCGd5
6w4A4X/C3LzwRbu7xkNXolktK3X+B5u1LfcD0V2VbrAujsNRCfYgka6xaSiWEMD3
r1Re7JAr4oduLz+ulMRkX6IoZscuugGahBSXv2LDbHK787Neal3lAK78DdiW8YMB
HHBe03xMTGElWlD+RfY5UZOCTtb3PUxgFaIePb9UWVN6kRTTEIQYvTtqK3qhv4wN
KSwqU/Nasm1bWNaALSvMW38yiWy1g/KHBkfrvg9ya1pnQ+CD+KZyU6/9QkWyLcpc
ecjk3x66ravfk/LJHz9VWQeamYQzQLdD/Vjwr6ux2B25wbV7BYiX9n2DR6e6nqNQ
nzHCzmmWX/TWasO5Y1q4kzhMVgkUbCZ8tUhK9As4pp1li39IZp8G59krwGCWjnX7
5yW47AnLwLyyp1BKE3ul9zgRww044OmG/SXTJnsBgHQpbmIUO549nxUMzTg3/45l
bMan00Ge1G43a1eJ7BbfmSkuxHoMd0Ybxbb7VWKs04yS6rv96LtSn7x5nmeWNkZk
hzsYJOzSBXrM0ec2NI/lS/E6PO8uA8kxSKr/96LLNrd1h2lyPud8ou2ircDnU3DE
5Ti6Iu3ANbhHF/T5dauoGkFyybXIx6o3/62PqSuIR3aQEjZ15qnBBcgEUOprRNzc
3m9xoKesx94e7/IACVaiBscQdHtgojDkfqQNaKyT5j4h/wsNmRMcvCTp+XaQLxEI
WFgAVIdjJbnzf3q6+I7nDHOyk3jQ8aMY0JWR6CN0EzCzCdqBtlkk+QJLxsXwgzre
7iX2lvq6lAxdkXMJgUjPF1WpFp6hIUUHxPnPjp4DiL9UvuM6/GxuiRHX4b+HZwPk
nmfxwov6PdErSANBxAy0kPxsizymdl5ws5EtjG0zg7aPIhSbj9sQWVwl35xVPRBN
lgJL4s7io/7MVunTiqApH2Rd7H8mQ+tELHg33tY96jaPELecOgt//3sew0pDET4b
QLt1VHPFZ+3eFRjqJOAwmJAfj82BMWE+E3+6W4h39dkmDfwO+g3KH2KqZFnLAFl/
ThkhlKjmsCZtWTOXV9Ap69QN5e37/S8Vm6eFM/DKUsSCNofDXPQm2oGFUcjdSh2A
FYvz9a3NktSmDVvtI1Tu91LKr5w0uK8J/F7nbJoda7Pe3SiahhDyrWNeJQIxjLHz
jiQ/912CcNEm1jUWuTqbk5vUmItakY2R6apk9YKM8DOKxYVHuaM0Dlpnk4JlknzF
z2Qx/nkQcbcH8lZKZ1gW6stCHFPGDUy5WtABQf/GaOy/RWBxgObf278DhUyseDju
Ow51vKh27qsz4Wm6K809mmj0T7wdQWUNDPx2PyHUlmZWk6yD8aA4tjFBoY20c600
tuIXcGwRxWLXq0ocwGHmesv33Z2vWA9WkTppDushB/R6ewEyquIJAYt6scp3SLky
/gUHYbqbBoUjjV2rOIno7Z12ivQO+Zzo2rHIbkrpnT7UwmxP5anVpwSAUqO9tq3b
ITqfSRmRz0LQhwZyGIPYp0srleCXRhVE8Mb42sqVsZGMBglMZQkr1fPmdhprpY0P
vGhQJC+//KwL0iOYpSDswrbnleunv//qv8ETwxf+0P7WVpNz2+OuBkKlPfBIlNNy
iN0MNVVLrJ1/Lk7mvl2N7wF/KtR0gqx4KhA+3ZqHdouGZpIaUhYgpiCkYUuIUeNb
GPUYXGJkgEOXmQlIjCKnboFiPmxoPavp0+AeEzhUkg4vJBZwi6AUD8t0Z4RstX8T
`protect END_PROTECTED
