`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YrEtDMN1JUTlPH4XgCBCXH967Xekdgux73cFYxehFYOT7l2lJpHEytJCui4jc+eO
0Av6Dx/UzfgFTyKJUXfnQixBF77NvdIZOGlwy7ZKRkyIepdsXXWntySqXXXxQs6r
BhdlDeA3UgbSFRbDlfyYI+M8MqlMRKCWSc+hiLDufSPtRXjRcKR8iDX9P9Arf2nX
tqvntENwjfd/CgBk/EN6dVh0+Ml0aCQRJhhB9TY4CdhjY9HUzpZN6tqxn+Kb5Krr
FhhhmcX8bUcdC9UEXm1icT+T3EipOx/hgT7nZr4V+CdDwbGgsslCzPtyhznYp/bl
ezJmvkMZdJqXCozTNmmhAAOB8dY25bI4NxPJn2uE9DYfuGCN8nOUNYl0mzYvQGM4
uMsd7qJdsqHlwCQmC4eQL/fJuFWZ7w+P5qqzdsgMFCF2M/sjcNJAradZXQdYc8t0
qHCFOTAlhMePiUIRbfqQ005jfrYYgvCsaQvejL2kfrB/crlMhHNNutSyYwYUtu9O
VlIjuF5RyBLcM9ukpI/MWG88izJECWXMHnrsdjK+/XMshr9qDZMLHuY4VQPUNNUP
BmY9dQwFkMgxlxKk2BmZ84p9THBvyjbxP4FGkGAG16WuvV6ITbMYiQBNQsIa7igJ
ANMrGEYB7hUFUnYSfF3lJaj3AKaHm9tbaFTCDzTbZEAe+KMhK15QETsB9CaivdWs
M9kNlWQKuxP9J3aPohh2rjEOg1XzOtdVJYtIKRaTLEwb6ukyR4VOIQRgUJO/1fXi
qwRp2nqucrtBAEsWFgBQDnWtDmg2tfqRaHtoTj/y5cv+GNVQQBqpDULQ3DM0udue
oOPCz7THNY3kyZ+UhrbJsm/oUIesQE2UfyoZmwG4RUOQ/zXlkHfMxQkGcWmWUVps
ECKNJJ8w9g/0h90JtWtj+QYhKpr+t0lWwfV4TyFuLjxwgQB4ii0iJBpeqJzDY5AD
z7LqGcDkJaujlxtI8an3Q5EmqdiVGI7j/zDE4UNWZ8vfY+QPhhFe1hKUu35+pJdC
+vb6USKC4OLub3DKKUbXUH21TEqEGATNtafYVmgqmORqecupqX1MhMimxD8tdxZO
MgoHO+zOWidERnIBIJBxfbs0kU5Mn5x1WnFJjlOBoPDAkJmlVrVdWcSUXsR0XRrw
BkLC/1EFIlIPiNo46zwbu5aqecX3EIs8O3goZTedOJFYwD7YdVzNvb74OKO7/2Ac
SzdrwlM5Y6itDhb3oSldSUSe+mTaNKki5SUoMSvk3mQ=
`protect END_PROTECTED
