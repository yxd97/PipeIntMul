`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0aCnbo8QzDgM8vSQUdxB9soHOr+1XzljTo4di4Ng/P89a65q4Hyf5GJ7+leN4njp
z5MofA1mlq7WO2uDDUuJjMZw2Da2O8hpRv38KUTFDzOUwQ9mlZsMGH5dPBGbw0q0
1NJb9JB2xy9Xq1Eq4yh0CDrJQWkYaTb72QI0TU1xHbhY9mI3ucGmOeDWppTNIY3s
4iJiJmYS6R7JVlaBtUjEU0WTeQXpC6U2r2nzAog2873bnDLdq2iDasStc8U17/tA
5cjkqqeiSkKNAuejiR4iEDw43cll4K3NH9bXDs6uY2curPokiKyK1MHuSpMDUbtZ
JkwcQC8avZCjuUPVbErIzUzWIncur7xfJ5GtC2pEBUKAQ0opLp9o546cKqz0olsa
eVHfOtc7qW4L8nj8/GtFPhaGe+5d799ZLclDkrqdJy43ZauiI2W2HlhhaV9lyFIq
hQbWXhH6vkSogrntmoj6i3fV+GdL6r/bVVNWMb4mkrqVsqDk6X3GUjFvW0ExBNSX
uAf+jJj5TXAk3fVyLfDp3hxKp9g3K9GxwvLsMiwCYpiZNM4O9gq68DZiQ10a8oAG
OHdpedf3NmO7cMC6QwsL8txak8VB7Eo1b5eb7/IPuD67MlYfajh438B0shSSgynp
BOJXLDAi9lItBjA7K50/tlVGmSUaYLMeXcZbxzy3RGahvg35LU/dgXmoAd+RohTD
2u0y2lE29hcRyP4d+0/SNn4xjVPgrU5w9BqlARFg3FqmASO80+ojttmdVoJCpcVx
SJZsGofGIMShqa0BLR1rJY6/PAunOafspfA+vedDFioC/qW2MQiurSA1vD3YTjWc
CvGQv1nGN2gHLqloVlFZGvQqSXtWinkKFZkx39TLWWtLm6hWct190LQd/34liJWW
vjjFN9NUpC6MvDc2He7vNm2EeQ5GNDV+jfq3K5wnkgwAt3V1EbR+3id7Kvk6zI/M
wtsxQyqAkCrM+kamrwDKahJJoy+vlUGZiBlFUMlxtZlAIUsim2qSw+N1EP/9OWXz
B5yorpVgq+ObFb1msC9Sc/37hI4C/XoTW2dmqil/h3zkcKkt3dqbKYYvRIIgAEgS
ZTAeOxJVKLjd/WJ33QOOA+JwD7KRpHJDrkgJ8oYinEIfxloFZOVdMLOseq1wCSii
6eNfORZPw/b0RYEoa1rgbUM2a6VQhhD/3IkBAb9C78uSJO8O9ct5iixtUqPYKuxY
tIIAXNgOYpjugQ7GhOwSRDQNsRRkZdjPhO6Ugd3+yK6CsXFL0I4PbuqlHBoxVj6D
eCx1SyhW+0EUznlamlNfsr5Um+2lrnMhVSVOj7LXDOc1yV/0I80+F2+ivoo/TfDr
a0fWCA2dv+QNBGIVhDydZ5m/wPRXpvAxQTX7dtaWotc+BjU8Gy5o1Sr+pqE6gV0W
H/zuz+PnM/uUY6urDzfDq18R29lZNgcA3iZrXkAPIOO5rTtIvRLcYcpA9pMWukbS
2n47l8FGhwMqlCcI+PNZ6B84hgdwk+U4tBrL/9iy3Q62RDNWllRbTN9FhsblV+Dr
`protect END_PROTECTED
