`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4xXEY2Tcl/hGcDRTJkZaWA2g8Gy9e85UlB17eCP6NnQqlldFrPN9Xtc0lfYscU8
1B6z3FRHiy80l7qqPalcVeFfK6QP/kGRNksUt9tuR4V2sboE14Lqmp/+OxrAxMtz
sf//VLGNJ3cyMKY7wJzvIFgIdd6mUIFNuQ3EgG/5TqhQO32T8y4lFunhtHNBaXdd
WeS0WCjNr5eeT2xj1wuH/PzwtNQXL8p345rElXQLCmHU+WMRzie9AS8L/XcAB/Iq
8/RQHn4E0FjVSIymJZ2rnz87CMGfiBVx57USq7a/1K+la4De6zJSTwFHozVo/ow8
TtuJK7688LXlxypbfcgu0Q==
`protect END_PROTECTED
