`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBQJNP2WalCF7bBdWDU3j9dBQ2HoKNkp0+ywlmPL4zffvXobsHccjXGOsrJ8q1yQ
Rropo/j8Rnx09RuOZDtqmLAaYa2fNpQHVb2K07fqBZnw6G2RC+psdO9M5H7bUFfi
4J8CMpsNir2RnIwm9RhfuUEDHVOxqoSfNaZEtz/9S1o8/I7MMk6/wgtnom38lBQI
rsWOKKCbTGJexSK8ZflRz0/7JMUO0O53QD+ijTZpSf98qTuU8Pwgpiw4W3CocsNE
nPAnib+dfuWKaRBzr7e25h8PMJqfJOHAEQyx8sLf9J3riWq6xz5JpRBX2M9Z6/Fi
S+Pbssi3quPXpm0xep9oZGdAfQ5Gf8P4G2XVPHdug2LBadWaaV8xZmgwJVML2MlV
ZmWZz3gzyyL6LwpPjSPsmghL92mNxNr4w4bYoHStnd8cDZPseSu6PThplkKVri1S
8V0dpJn3QHL17X2oYPhAp7s8aRd0OnsQi3rlKf2l3MyT7V+6Z/Pc6o9+05ho7e3f
RRfj9zSgKhRZPP/AzQA9dVtmdsVTObrvbiJXbaHDsKshOpl2zEC2Lx3vYlxiVuSd
pjt471HvFZqd7TmGbTOPtnPaUc4Ugec+jaQS6GM2dmshDDekvmo5JA7cjtwyNnkf
UVbjYujZMIEpARfkqnYB04U/KCKRt0bMVOS3v2rQj44N6lfT6MLW7CXwEqy4LH0c
B/+sXhv2VxvjBFtr26YK9Qe6QycQW1To6urfW28UEFo0EirfkiVDjYM97E6bWPr/
ue7bIpmscbk//RtMFjWF+jUwjcR+PzrrvbWZtG7tPu02CGQMijvSfQZKYViam72P
l+5BbYw0X7Hnos0yKKRHukE9miksfbYVaxWORmBrbrEwC513J5VtjUxuSmszUXmP
DiY6fAtiLrBq7FGhrJ7tmxhUhKwhxA6c6UlRUHZDS+FS7p90C8bXSsfo0noKdtEN
cMLcgKpYEZ+C8eFcYJJEc5YKjkTnInZr2/IMAbvPU3C4eMKL73ZdFfOLpN1HuHtA
4VVM9Buogyjp6gANUDTBCAZDjqXqcF/ZTTex6Cc8qLUF8iXn0JIQfZZTtzKkphU/
a3sikgmz0jdbkhEI1o8O9L8PlHuqwoEVKrjj8/utcB/sHSdAxdobxAxgVfzLBysg
wFYfMLJ9lOyUWa9dRYj86PgS53e/OzDmJQ6HKm4X9PeXe7yXoVLXeyu1YgeFijhW
vgIuNL4D93pBy7Ehmr6ImH6PDR8wrS77eSd+P7beee1wL22O5bOAgMK4pXtDDoeK
EkSDH4I6qTrxM/u/McGrUcJ1pjASNUd+8ovXAEVgACdBFKpS6YJdXogBdgjWdM+3
iul8ypmEjj/+N6Pg6+c8E6f5OCAn/mHnGQZ5/+RLmaH8Vw4jYqUVr0XMipCZ62bT
CJdZi1eeY1SBQ2Ux+p2zVkHvzEwGGw7q98tt7iLKEBKOxQ1ZTq76n4/1UYaH9CIm
TodeTZwc2rK28lWAXrQ080vPZh4dqUEXPXVwAPKsxCcArclbYW57QHsjRqzwqJCk
djRJvJIdKiZutMsTH8qgwBoci/b6FfgYWwU+w967qD/ChNW41HZkdl4py0xjIsfe
wtq88r2m8KtB1yhNysPNY27yq2vwuPEsiRif6HQeVsa3TkXqFtLWdUfVBQTBR+TC
y/t8bNR9KcLs5UO/Rz7CdcQ1tLH05+oitZhOpw2dRPU0LpCOVHpMXau9hqZtzNGY
yraN2jpxJF+6Hu4XtFIs+ZViG/XZ98QnCET/iabZ3KZljAbGPcMuNC/YDey7x34l
S1/vuVsvts9YYZ+nFPb6YEzo45an2/D31iVdwVdrLz53tcad67NaBOxISHxjPLs8
usIp1m3XtLCn/+T7X1mEamJ0KA6+DgaK0zMqvIWHEvXv3l4znwWrRbhztCuDuUta
cI3/E6dVXfx/GGttPNEmOxG6BYZyA+9UA9uVuuT6rMZ2z5+hBBzsBOEOuEkM5CKD
u866NLWlZiv8FXNpacrZUO0XExkZe745OJvTzhQ6FB9K/VdZ5dwhJ0zJrmtE2NzB
7iAkJ4VmNOW0w6w4HxEPkSuvLmH4TW7uEOyD6IFHFnUWw3xZAchxvbPu5AiAkCdO
Ee+t9gZSkP9i6xUR1qHDd75TaCuZ8odMfJwiiGFs9Ml56S+MRs1qeBObzgvPoRGA
aBi8WQ5YnQ8u9BBxq4gFSL0CLMzUoxbfD4UiPGeqD4Du21UIz8vlwi2o6opa0s+F
rlTJzFTh3jBkITj0HrVgrSRFEIKGJYYx5uCfeMgfrIzuVbeZCa8YksxBSTy1nc0C
Ig1e0UdBgFmTmrdJdT8vvd94LxpgtPuMl5K5FTtwiOih16sbS0UVupSrSJDZ2V4t
gJJrVPZvJ2FPwgDsGPeCpouQGhzylQHV+tZaEinOn5IKsioInO6M74YOIKjwqh7d
6MsbhH0Hg++M2/ZRGxJ/p8I1tW8fTOEhdNMzzs7AER65psawHWiQOYIBd6t22eWm
LarERLg7rjdnrKqJyDK5phpB8V111Afhs9D7SITDg3c2dnkzFCzZ2TJCTb9yxTo/
fkhxg3tnvkbBvhVppsUtVY2OodHjcZ37e3UFN51NnjQ3T8wNYQiQijpsRvpBaL2k
m9AK8H5l/JUuQuA9CzCrT+P1ue/dDivfY1tIa/jLWIY3pzJvzRRoi0fJPDnXcFbV
67PhWXW4AtNteLWrqyu3MukRzN8LSgDPGn7ZugCCPQcu1r6QxyFV7vECDZsh9hmn
XqVL5zrgPPsK8DYnYrI6ie7L6QoawbkRXCpwc8tS40DaNpAnn2IoaBFybxWOn6A5
D+lm6PmKGU4PlrMfKsCN4ZNPp9SQ+khhlgqETQkziEkCsynWT7ga7PpTohaNfsgG
lkG89zWu//zrJajuNniutlwKQw0q2oy6TWCkj7b9NWwq1iZNntmQZcKRr+B/V4il
8DbIjwtebR3nYh00E3DOWjKwvdVLGSHAjdZnMCH+gGgE+/8dD6vev/Jf0esuMWV8
dFbWf9ffrUsx/oP8Oi8qsgoITGShWR0vXxx+vHh+42u9MhLV3ApETw5MOjZ3nTJ3
uR09v+JYXXyBAABs4sjm20+MeBKj+9qodFoPyIxmv3xjFCRmx/PjTdlOfTQkBrSp
j4fRRCnD2ug1vDL1SyVJP58TJaH5yq1nR8HDQJMHtTiMFcn3fLkrJFXxxsTAaKvD
P/gDzg87OUDMJ49ZWve125o83i3bVKA3Z51xNooUeBOD3xbhLBq/ic5VgsMBRHEM
TEWh7RdXli7fJDOluAiDI0F+RoTpy7lqiVpPbrLESAATSsYiWuUPWzlQa4ibOTwX
JwUvk5G+KEYKnENzTFD5iLuxaE1NK7Ij8tRALntvbGpQuGmU9GuFnl1XMudKAahI
xeiv55RFpWljt6dWdNh5LWI0Y5ptB7TaZMSIFCHald1jdW2Mgf+xZhFJRzag2BSD
iOkEwD/1eFDiQvSffir5Qc/jYZPD0u6B3qkd+DL3l6jPy0P/DI33dznQXYz+jH+d
1ncYD2pjva/ZuMAU1+MB2M7w26R9ZOI9ZQ4p5ee+UF/D4PuzO4r1ML+KShawXECU
UHmG9QbMXFW6spGpzCmNGcxGk/770oxWqSGtZAK650K9hfc1xZfiqq26L4h35UgW
UHZfrgi251271xB19bi+yhP2Z4+ox7xL3EV6QbHoH4DyZv35Kxo8Q8nVZOizTODB
rtusUHRysEy6oLx1x6oBZB3skTP+DEOA3Q0ucoYbncU32O/oRpw4S/q4eflrriYz
fDE0PVtAeO8ncDWCcNWlbgnJzSZ5a+M9kvZcaD3Bil6e5SQkK7kvZbnE2PwzC0H1
6OsizcckLFVG0tra3UnWP5+nVYFWc7UzJ6wpQ8cnam99M4jG7lpA/gF4UQU1KRtu
+AMLZITHOgNv/rSgLQ04K6zP6HA70c/Ra/0Z5QdLICaWrz1/pigUmVNz2ctECCk0
Og5yi4BPbWvKLjjweEzVJ6cBOdbrDAGbXrUI7vACMUY3+4YdRhmP1tZ0OIkFFObR
8hhqsVztUotHzmKPf+qW9tvFN+xJNZb+6HEq9vD+vW0mFMFGVhpCr0oNUYCRkvaS
8y6fcw83PTw6xbpovOjLlS1I9qYlwXJ+hpDCsozJjY8P+LuKjaqYcp0z0IyuPvyg
lo6T+hgKZWSygGBuon26WuTyM5PvjQp0N0IpxRUN2ObdFhvnVYcPkC0gm1zeiMuS
mMQt2aCND95njTc3hy5MoL51MgJg8CFN7+utFW8eUCroixVJdizp21+EK3wLouwo
BBWnmIkEbarUv5xMEAOv73lJm/PMlk8EUsj0I5u2cPX/UHQh0kznpEejgn+CgT8Y
W4jt4t9TBHThfNgcPvkL4FFrDP38+/d9ZQivhRNurrc9Eakygm0bbHREm0xZETy9
OhympgNXJPUlMu6TNmgjDdY9SYPRffQCOkr5fWw3tT9QcDVbuNz1qLPhNy8DGJLy
UoPJcvR2pg3DzA9jXYe14mfdh60oCcnxRVtosy+PQEqD8hyxIqje/jdTY9JTYAo/
FOVemOxYl3B3Qza0KLn4JaTM7dzk7DiYuXHPGSmzucEm+1QHxCLkX17RlIAWfUiY
CkQKvlN0piujIYJwKoNbXJoVI/2s1F7uv1Cb5RnuYV0PoYd1mxvHVSvXh4pvEQwJ
lgiwEz/21v3B1LwWCSqeaOmJVr6bDVg8X85QaWK0L0DqQ83zoJSYbDIN/GyzujTn
Ff0d0g50lVa8i6VY0mvdcFkkoUOM+btTDsZaoziaVhjVj52SbI4ISb3WqVjgWe1D
ImyrXggWgGK+wqgtHmVRCgGLc0aGfxYHCPpMRgoVR/rbZMcQ5J1bnT/LB3wpxcc9
uwpWY1p0ly1+4Ll/2qT+kGLt6iEWXkn3DIewrfde+VDNzUj/S+fUmmG+T4v/G+ps
2InbK+qxB6i94yQskLihfySE6DbDYB+7c1Avu/p4oTq+qaH5CDduZOJgvTQp/ImA
XnND3ZkI6m0A8P6Z7sCMm72xbAFWy6KY5QWJk9wikAZsuQ5Cl+f2GYF6Gjd8thqM
1QZP9tJcp7UMfcSzl0HdwQ8SZQ1PXwUecbRKRjnayhipUIXhfdQw90ZkZ3Mb+mOa
YhWahf/2tjfzSrop3A+zVoIseRiz19zyFSLR3RmY2ekyNFG0ydb1h7ZXmF34NndL
TocD1m4ryISad5WaXHIqEWG3XFaVQwOfMiCZvDeZdjOwD8YCGfudolalweUCO3T0
HhFAVze8ofD3SxZEq/gJ+MtGXzCeM1Xsf8yIdthXghZb58pJx1Bg6jROqyxtEeZ3
qOq0h2CohNJxR4U54Z0GW/cY9dFf9mMvCfaG7HqmJWepHFq+Bif1BtldQnnbgA28
U3dappuGjZ7i+/Hu6BEXZfYvbeWVRFtZFDGW0JB1oompXF5RTWLq7uZVaKgwkedS
pi21iUYN33p+I6txj1X8I0TioOP82s4jNOYw5g6qUk5BqQDBHEV37459CV5AIdpM
sBbXve5bNEk5StS0q9wcmu6qaeAKS8/y5OoI9/3nA9Wcq+oWTokt/1+BOFR37J8D
UHVfbl6GtpP+0WDO7reYUKO76isV5PxMaJ5skRLKH918Nl/VrN0ncqcJu2k7P7V+
3layOeN9CGYTMK4CrDFSBRp+uF5DnplT3xGKHk2O8eXi+kcANOV3eBxvdv+oWyWF
ZIYW0yVGx/qAP5CNYgWmyNW6i8lBUvegbgd3HgwI87GGG3NRTAWtpcw6kpwHE5KD
/UfMjp7/yhk3iginnVQ7Ub3jJj606tpAztMyj6ZAS621pVxCKnyJbrCm1bJ4QGtp
A+H3XLe932s7vbgsIBibQis0hd9hCbBJ7wV2oDEPIi2LEK3oZVIt0ATZRUawISTI
xNkalzHkDYZlxCLWQtqrqTf2fGGrIMrpri60PheWGqXS3Seu8h0NtzyLZ1YzMYmC
1QQd/GyZniJTn4qq0/EBTbkdelVe+dYsoH/cCOKh2BfX60clNTLziIhX7g7vxG5s
+ZlkA6bvOzuAqB2WZfrHhFF9pBzB2Fk5YyCHrLtfXaMCvl2jnyWS8X1sH2VS2A1y
4D89xD8NwZ7u+bGd2ILdhKcepPzuvu1cC8CJTAN+5i46W7XbI8kTmSqU7gUxACqG
duJ3GmYgtsijoJLVudORDlrtsIbTPX0h91SLHVRjmb3M4J4ulN7vj3tKLJqu4Amd
7zcUn+R+ArfTwmMF9pdJybsHd52umDYDNix9s+WbxXQ6zduSUItg6x2LSRjHhgQD
ensQfkZZ4l3az2TmrWLlwrB2S51+EKc2mbWgrMq0Zrs+3Zq5CTvRwQBiL5b8sLIC
RF10Ul1rCX33xs5fMKV7P95g0SZrkj9YiV/EcxXPrkfONbiS4GqaGs3IluScZKXs
I8APcp6z15GEGf2oW5jXXWHz+xLYuIO0aql5/gDT+6FF6bVxCUYH6rbYj1YEwPRn
c/VyDhgiXB3VxObubC1vKLlxla6s3s+UN6peNFU+GFi0KihaltumZndZ5u+LSFZr
I8d4vUo7Mfni48Eljp1rIeVt8dkOQj9wpD17L1oFl1Rf/mBph5QLl80fnTu5bUrD
fIVhhaoGG1hFsoV0S+/Rv9drYxAmXpesD+WYu3Mzcj1kP4eVLsIcyElLU2GT1RCS
f4XwHechjY1hTQDb1BjBjJVfheQ+E1JLlidCelvrAhBBFxzD1896yvKUFCGT2FQd
DMHCvQnv4epuxVlG5AIjaC26vNpidfuQIveKlz3WDqi60wJW1CkEJhCvBCenZqOM
Tj8Rg92ALT1Awq+pPPhczr5nT+oUyt1esXel4xV6YCZeRYWaV/t+sMhjztvCXbgs
Bq0+GdwV+FTkSWyzfMfaJNp3GodFijVpMMAVXpxZ3pOOi9OdJ/QDwhuz1bB+Sh/I
Ovxu4Nwnymwqc3ZCa/5VHbQaL09LXLzCID64BQTjt1y1gQ/i8527jkoNRoYp/gpg
32ZpRgFYVZ4V263VizXwlBYLcVLF25Wxe9C/LkpD7wFWJ+F7mRraRiIDFcUmlCSO
FZ8/3KovYGtMH55RmhrkN46AJ9mNm6wshj/miuZkkJyS/Mbnr9/WTNYJl4nXvP+p
E8nQsKi6tRWmkvrnQoGCK8k/WkQMkTCjn6U9iW+iql3ne/hyjkQOSIP83uEvOiis
d+M0gparwY4uN3EGHRuEwGPphAAw2UKFX8xfjEB0Atyre5m1bcklQl2L9hBc4ryF
j+aLgPGh5MEHyoTE9SrsVrEjakvCYemmRFjgftlOVRqWaxU1ExkKjyc/xx4Z/jqS
TQKRohgxilOz93t8+rVwcuTnwSLNu1ZaDjwX5V+v710FE+9cZyMR/uRbu9XC4UWq
2rB78mLxG4natm/R6EDhRDGD1xlGjGkBFrlRcaPOAFOIvO+ffMkM5gApet8n3Ugj
qyEunL0uZp9aRpzuQP0kf+qLX1HWnKsSrUFqEpe0wkxGcn6ZsVkZkcJAUT/Fka7g
l60FxWTxKJn1Cj40hqs9sQgGa+53BQa9JwYurzxMi0CgvTek3dqbTfXIgB47ayUE
gTQa0sm0yIEsRiZh2yG7prxfxn+IM529RRWvXx8NID167bsyKAeWeobTvBYG8I6K
5o3GSSa7UiOijxSMpEITggJw6+GN72601mlX7rLJgGiHgWnLfwbk2tdUKU84zjOa
yIsINyxlwPhRwKXWOFbtZCV7X8uBS82IGynwi9SSN+UvEQZ8JKOTXL+dKPnQ+FUn
Gq/+VVL/OMkHLKRZRyRWlAzg08UFaVWvZp9OGZyXnjTpJM04ARdRE/AETmlhwQsm
ury055dsJuNWMdKV+ZgDompBrCMgRDhkbTOZnkemylhiEghAB1l00r5Wq0NN+GC7
ezFxes8hktgpjXoLR7kgmLujx8N2QI+hp94YiR9U+BTuNy8aO/C7ALfONmkSJWc7
GrJbPXHvArDgtUvKA+j8NlRBoU6oKoXibAEA5fL5qISxLqQfgzpjLse5XW15/8vi
KdMDm+AR26ua6zx/Gfbchwz8E1xUWVoYJYcyO+1ZRuvuTsYkDWKOqKdhPNg5a2v0
MQE8hFl9SY4jDJhJW353YG0txWw86z3NV7r9a+DE9vcouU3u/Ni6ZRACBil2i6W4
2FGxwTGipaPTlg2Fxmdz5aFrBT7W9WaSzPK4pQu0/UhjA6995GGA/hcLMDFiKtyR
Yp1iH0412Ueep/lfjC2aLnweZPeE2Db3qP3SwYKuaafGO/hdf3rcpf0PrR48mGcw
pzQMIvlk9hxAxFUfq0CuW8QcQZTe8tCpDfLKl+fyj1TnPeuwzB5+wQEbzH4+4bt9
B8v3nI2emegyqvo505ZTiXLbaO4qp4fBuOOJhUPIjQiQ6awhFqi7C4qA5N+S4hza
8Cksf3aYGmps1Riylz6Hx2jqH1QpN3ZdflAmyR6XsGZijYwxHHM5Em2+xRtCKQVz
iy/XfPdnnJ5Ym7yc1dsgcsbznzvM9mi+yPCIMS0cVuYuhduYE0bY6Z1V52pcFlMl
nP9VXFAJLk8dy8QQdVrwpRPHgcdZzi/Yf/gk19ohycQ4diFzVsT//WhTB1o+YCno
0y9M+eefRbKZvJ7Bu2eKzku+aYIhNxeefr94K0o2UJ0iAAQFdxwXDuyN0eqp8vkO
OqA9hTqMk2gju7YRVJSwSvtFFsjwclY9wo3td+UfTbkfB3QGF5fUr9XB6+GO7LZR
9CvLNDU7Sz1BevgrivqMHGV/LivpBMPrerXqSty+5frSutDz83nStzpOKwUrt9ct
ppGODoczbGYZh1PPwwOWq6KF8CQIaAcVP7MBUbXuZ3W8Utqv83/tYcqdcn6gqXTv
xJrfPCFGoHDH1fDKUmEWcvxUF+qYd9EZCjliGUgZsECFL2i5ICDvIVZV/goegFWG
GZgFGd7nF8qif9jr/WG07VM0Lb84GHHedqxGjph8Umdoso7Pm8c6C/YSOsidPSic
seNX32ceyfgwXayYy6Mb+mrqeC5zvlK3W/IGNnHvyIYGVTd3VeKPGn7+CoIq4p3o
K5zZHGaRt+UkLl6dycHD7uyhgeJcb8a5TgcIEYHcl5p56T2EYYuPALKFXmM0mQ0P
qtr4/8sdnQWZwdokzQo3qgPWkANup5ujxYnkkjAU0iCGLtafYIBNjhQvDoOw4T1T
VdOrhZ9qwE8lpe/ZFOwB/gzrP58rEsSkeNcKinkwCOwxbeuK+4d1k/NSCOdIdY0u
znYPfjNKoCQsQsS2W8CCiYfN7YkmdnNGoGVkQ/8EcrzFND4/x/StGNF347VZcwDR
R/yEZokn3oXuLWO4MUzn0CM98UiMXIW48Vs4n9Llw+oKHe/wLc3AgRgO3J2wRsvW
ol+PKwiQhCnGs12K1KhUh57hBXhSK2fc+DA2qqNdsA66a+VA3jF3uQv5FqQK2kac
kWWf8QhAQ6MrwfhBPca2wZXRkH7wDRX1/3nX0LpvFKqmUp2ZrHyND0uL3Mg6++6x
FFe68t5NWsXqtbnZtdew25VdYRhxXP9FEUivp9GcNrt5OZOrE4xMAyRg05TX3Dcu
QDXpPrGbeG69koPBU9oJcN5SN/DmV7rCHnandaL5S55375c28lfFUHDlZNMK57J0
GT2kphebkYbE74dizqbNEKpmUSF7JPGKBsaiO2DebRU0Vt0VQIwetpOiYhjHytTF
ektOGdmyp1pwj4RcQGFIJG+9HZilrbTLejpW0UY4AVGxyR9Vpxd585fFyRnYb7pV
SSZwLetG1RfxrmtEU3fTNF2ss4j0Wg1XTadViJKrNpCwgMMboDkPnKet/B8C7fEY
JLS4+NpUlX5HNv66Lukc+DxQ8EvFiVFYQ4A1ovLoPEA6DkFl47mbVICKFG6busk2
urftHELYs7KX40q7BVG6km/P8CJ+tTXHk+SvrnhT+CIacgDipU22lR1XdGmI1Io+
nPbhGidNkuxHW7H8EygSoTpKgchOUxsmb1BTFoqiwRaxGGStnAqjqRRxydAEtXJ3
ttt0NA9M4QEF0hKg8h/YNwuwjyN02GR7idD2hU3InylSRnffswSUHFyOJnrF0hNh
75d8Y/AUJWaW9GgmZJvEHTV/fRuwbg/sRYCwJQhirk9YFG487sSstomgrn5VtxaY
MIcifDgCn9GnfwSCtJKopNm3Pn+989nS9xzcJixR+fCYOfBYxcpT9Ek2dZnJYJIT
1GeMtyIxuPiTeVLrdiMcd8mZ5vugMZqspamRe5wONs//lqPFjXZ7Pzg6lpocRr0U
v1jB67O2iIBXyzSwTWQaCI9PMT1T+Pnau6KM1HC5rK0V2/pR5Bm6xRXSDztKZpx0
/FGGmTCMy9KG/ppKFzsniOEfLa+SezIHcWzfSCwWX8nFT0GegIMFh+beXhx5VeHz
weEb4GR6SoQ7nxKOLEgKyZ/gxbZmCQyZqPORkGaCab6pSpYQLQxc+GlO+HjZ/rku
wqytOg5a4s3nLxJgAL1nev8TFWtjcmPxaoGrt0WQv10GrPJsGfbZWaxoweoIPXi0
2gKIoKivv45sAxxVHcKIDeFMcRSWH222iHZhQvq1Pfvr7Gyd8xlyluLZUxNg3UCN
3JbIWDIFuKWwLx4uRN6b3i6aiAdynhG6F0XwwKKX0Eb6m9Dny9XjZ57RmWQdd319
RUnUMfFfEehUTcz3suVOLBYfX2HUC66jkG8MZ6mvqvVIAjoigA53MBtO4vXw4RFY
CnzsGvCPbSlQnWBtsux835CLHnLlOLwkCnPzFbnGOj00nVW1soZveQ/LsjH0VI8l
hpTYARcqpdfkW/QJio1qGGuCZJiiPOq1rVLkxwvlHVIXzM/zKGWX2JSN3QYS7JD0
iz+loDB2dD5LYmVaU9nR2qdQ0EXbRC35c4th8blqu/2Q+oIw4RHvIT155qR+Uezr
rA+viiedpjd4QvwaaQZPmYhItX6mMDkVrJvGDYQ2JLona0bqqcL+k4C/vJCJWfb5
JWWUifa0u7G/WUMnImmjVXcm7kJ6k8kUm2oFGWswTgLOUmu+7o/SsHdDHm/nGgL2
yNYOKVqHCjzJZQp/fTKhfz71IHBVfNeDVs8a5Vt+UryXvgy6lbJzACc93PotJLSs
fRWi+/P5zgiU1MzPVfmtmqwrkYgmjHMPV3CORJ/TDJ1GOQW6G9yitz0tGmISAOKI
QXKic/n2RnFeQlZ5txXqF4ZY+QFE5kaDQrkCy5rjxbzz5K+KKbeKNYcLpSuWnwG8
G+UmbM5Lzxk2cFIw59bknerLcVh4PxWvyv8XK2lagGXN5LZoi2m/+ivOqkEF9jnC
WfLwTTfwvlgLbs4mYhcP29jNy3Qskqv4tEm5KXf/eV98yHkMjQ2EzgQ5Ul3ASmfh
rixMzhoxrIEMOpy5YN/MTSuqcDw1y3ZWgMaw3v0TTJfS0r4qzl+JUetzkia9IfDO
18mX0gmIGJgCVKv9QGenWvdKP3R9WP8kEopmbq5GxhwCSdPLnsVbosb81i2kT2GJ
A2otCb+C3/evdTAnoyRj4iA6Lb1i4uD5wjdPnqANHQlNHNRPsR3FrEw1Nv/QAfXk
Y0Ev4B9xCfR8eKEAljUVX27wHlrYyKBk7nOZQ5y0q0WtUSk8WM7sEffDQlCF3eHI
8nCyzp9LSDu1bXRXnaJojPaqN6ZkzvH018gCQC22+NVXbEwUqs8Qw2fzw3Ppaj4a
kGflsykzLiX/ohqi/SBINm291xe8wif4hOqRna7uI3k=
`protect END_PROTECTED
