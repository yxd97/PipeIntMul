`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FSn822ehCInpFUadc04VfFmJDNYn07pyHe1tLoVilXAWJa99ldU2Fh7dBmW3d6aH
2QRitAuWfYjzh/f1Y3QCJKGn3WttneDRDiawd1E39CacP1gniGWd7EzlpDhnPFOV
IQ0rvYHkm3MkrGbt5qI3rjqXZt5RoDsnk/sbLm1YTe9TXC3WmdiG4cvjpDo2JiHQ
jha/rfe/Acl0T/aZnIGz7hr2QbHTPUO+ms+46fiC3NwUAUmStMAXkx3F+FCqdS7I
kit1YE2CNxqWTHDc5w7R/xpT+wEYazVZHp/zvRDX4s91hpeFC0bfG7boF1+xx8fp
5s+3eB964yHSNSQKxaSH/z0Q1UGpRf8mEGlNj17uDeOuXwwEz/xITI0NTGm7jZol
oSPy3sdw2QT65YCkFiD63a8mUUiOM2n8oRKLnsuswGUbC6DeKkzVhmzspkO/Jj8T
O+p9jf+j6ucHUZP5lWJx7mkopE+D/S28Yz9MvtPb1HilZnCK5vv/eDHLumjUx5RT
0h3+NfpA5ndnXQn78mg49lrKCIeqSS9ILA/j9aQpGhzW+lrALuVuOcYVCRH3vBjO
09CR9ntk+k79GRdm2Z+f7CLuwN0jUzegAKWuAm98Np90jOL2t/LA83gqeJNc79I8
Zme5F120xjQkTXUqCFVZXOuuKl0Zvxhn2w48DP0lOskM0Z9cOwtDI6yOaLTf42zO
RtoFNz03bVJMcqhuLSlHyP3EZFfxg6QukTy2zSTQLJ0MOJI0Xg+/A0RFBmkBlVLn
inJxW4RSqkhRyCj75Ra3Sj9zDAHu8vDtUuJIppTotdoGVr0IYzkxDevJmII8wDd4
ye4z0/VfMZ/5e3Rc0CR707zvATjXnw+wvf+ZxR2Pfq3ZIvUgAaF81BQyaG5nNKWj
kcsHlXwIq/wVDThyFYl31wD8WCB0qLcd1BNwu942G2nGn7gh+i6HWIGSk1HACvL2
AIg133qLLTzq09OIIdsk0s5m+eklVSUdBC27pTVFp/Di08PdU107TQUaHHD5LVtd
DV90IWFh5WGMrnWRlSSOy+FS/mTXP4iwqZC0MXTHTOR72UImji/w3Dx3g0MvJHR4
H77hzGwyjPOCbhZvgjql+XU1ON1Jq4XyxTE773JVjHByjhN9EGbC2j3pryWyRRP+
DK7hRLOA6928bS1ZJQX9X47JRBVJskukobZnR9v7Gn2pLHw0ChBpWkz+zA96+UC1
ES7z8PQbZum72UK3fiAViG/gIembJRyF9/fCiPaJ94MB+SmpWGV1C7buMEqM7icM
azeyvqUKSnDOjTbSaCIVN2Sk9TiqvYL6WhGXbq2sgPeJZbF1QpECRs5VLCLVJ+iy
uG+o3ENBxzuMQFBTiNerfQpMRAicv3EEbL1NAYU0bYHlp4h+a9154UtVy4pUSkMH
GAlHy7OmmdgKyGH2AIaEpkvQdkOIzwo+43l1B9Y2U2IP+I8zoiFExihzTu6JiMuQ
2jbcGSnOCLU4mREaoTlmKHn/NgZTbPk2aG5uhhJANp5S1tgkZcJP0TCwo4Aj0tKs
UhU/9T/iViHovS3SI01pF+jWaQ22zaPvc6HOs3jJROa9uO+Bsx0eRv45X3ECyXQp
E2pYOOW5khruEWIkk2IbLyHWkDc1mOxUD/Tg8ZekHqsw1yj5N4+5wrVMRbOBkHWF
Dlw0zpDi4GAIo2WjmWPhZS5wVGefTg33oZPVd6o8ton47eOGPcLnwR0xjO5gHFbt
IWysBBNE6w6rX0h7cgv4CR/hexwO8ZyH6K29LHi7v7GZAJCvaHmATZjq1JwnR2/t
GhM21KPASanhWuWZ5hxGW42ikS0FB9mfMxS0eVomCIoRPH+AQBt9//7HnxJMGK0k
ddJ/uwvyF+OiF4v2It3YkRVhg++aSyXbw5OmtIDgDG0jRbONs7nDR+3lp6CVo+SI
047W8JpKFxEerWXk5Fr1ttAeLa1ZOyD69jtrbHaxC3H2M02UAptf6eBTUxf6uPLi
Zjhs+4H3QQ3BvD7de9At0FEuUXPiEJRgIc7DcvQYfwQd9oLfIIfUozntpXyNjQom
DLtgJZ39QOwyuZegb703hQzu+3jrmBakt7Gqo5Z0XDNyKFkZTE9+oz4NkbtK0sCz
ZOZiiwl4FkldUjJR69jn9PJfEf4NPjQnCHYNfQ3NmTg05/Wa4mWAMEbaDc7/qVYx
dgdj8QmeiQ8cd1784JMunqP4wB31znxbwjzKS22TmpD6qfg33c6Aq4PtQHwWRnEc
ZojG0xf1pGxTT6uZYOqtz9iB5Eu3pC43S8TUc7vhZ0kf4K3jzBq0bCr5eYekqq7z
PPyo6s+ioaxRMbbcsLeeSyieMrYVhk097YotzDh69wRrpqvwAaz63ivAnI9J97Pu
3qJvBkLWORa87CpHy9CuVvBeYzbggqSVWY3OYUBt0xXbezDNMdhGC7HMVXLCY2mO
DWsFoIa8f2cslXcpR7thSSeyeNWnlYa30wKj0uZYlSZ/V4f3Yr+xeW3k6LGM6fsL
bxxhUZ8jrSyIsQCq0kGY3tVqbGhgQNS1nd77D0q1+eCZ9p3iGBPLgjeLxote254L
yJUD7OZTv2C7jSOFrQe7xNHc3FkfOaehol+P82FWaJIG6cj7ax1EpVb4jB8rYv/a
V3++34pDwUpN24fEy/MKo2jJ4eGtiFx0YVf4v2y1v1t7jmo8wCv3nEf9sdtO29la
y0f7mPYrPvRskaGPpXbhdxmRkM1nmqE8w6hlOHtjstTAhKXtYWh5hvUFUn2ZWwZj
VB/jOZG8TStICbWCS2FMfGn+gZakma3eHCu6Fed+B1RSY4pD7BWFw4wqMABfZDCI
6wvsvz6XoTbtxZosUJpTt0q1kWNSWPDirhF+yMpsq8bJ5vq7ZHo7Qf/slErYH1jZ
g3VPpy3e9boF7qa6kkaCaBBTKq3524pUFZSGm7SJOFYSYaufDm+Gl2jAah40ZydV
ndHG1D9WD7D4ij6Co1D07S3+1YuvJlw65v2m3t9m2Uf7X+5QkcNGqq2NL0H/hOiR
bnsj9wwiCFj6LQqc25n3gj8ezjqCCnm4UOCU52rn2LakeEAiICDs3G92XHq+/zk4
z4/nfr+PjhzUTC2Jrp4f1V5yvwMagHylqCM+7mR05ox5FPE4pZZzrO4846TD880c
hs4KZM+PdYpjCxEwBHjz6ukB2cegdNUrjCXJUKeBQxlwXj+SJxow1CvpdWZ86oXQ
+X98VcQsqdH/6YX/QywfozVKyK9d/zGegE6Ypz+0RTKtIjEaw6PoHDJFLual3mSJ
CYk4jWUxlfoq937Rvo56LWHiUiHkQahSzV/Mw9F9SQe/D0/pj9cnjL89+mCBKyF1
Rr0T6GWN8oXq2dn9uePRLNbc7mzaeJeJ0dPpkMajCI1D9I6so0qIrBYB/2EAlChM
WWreVd5lOQ82xC6wwoHLC/sggHdBouw1LyaOlqTrShMkO0dbajaBtOVlVP/lYtUn
42iHuU1dJ1ywMfuTqasikZM7e2nKpVrNE734JjQZbM9bPWxCaPwWPXyTh5JgxbNW
hCuBGm7uAzYrnhG/e49TC8YCAEXbcUZ0ShNfhqFPcsYh2YfZ+ZIVAKwLF/GvUcTn
2cAQmJryWugyqvfni1yYtVGJMfGau6/Icps7a/4d8eovYVpYhrRMNyBgTilzEPMF
EFXLF9EbbuR+n8/KfK6iKneBd1NHS/QJjefeexmUO7JwvU/7DSZ9wQhi0Abkwr/w
te/xb4p6x5RhzS7rdWrOGgXF2YJuT4vn45McXF7rkP+2fLe3LoLeokHZGZStnREd
teXgmFZ6bZS8Q4/cvjOunZBzvQqxfie0fBCr5hSp2mjirIYt41m5EG/qB8QI/XsY
8eubEGhSHyusaVn7PBchk3+OuAWLHx2Nj5dWKNv5GH7lK0VVRbn/KmSd8cbSBLQE
fTLpZ+pN/hV+4Y/TJ5mJTcE3WyI5x6ZkMjMvfzaXjuKikb29AH+ThRLoq9ypXFBR
OC4QU/nOU1Jn8EM3soHY1FpN25vVSYK13/NGi2Znh4NvOFPwvvCQeQ41WZ56PbDq
HINUJKRZG1wYj9aedz5CWl9Ra1+W+GjhYZ7OSehFMP6gNnUk/wwbaTGXURURUWxh
d616Ei3DpXjNB95CtgPmHO7zXa9/Ad7LLFd5CvoDHwOmBtguDz3TBeyFH3p80J8s
flmuAsjufhy/Wd9hfU6JR098My5qSTQ2f04S3UdNwssaf3bmIN4JTstnzXCU9qXx
D+pQgSvXjt24pCcp/bAY5jDzxL3++jhZGYc88dhqOsES75tA06a1QfyHidyU0Rka
9WWikHjMf0h9nWTi0E67MGfBR991K2pBQ5Ys4S7ymFZk4HIrno9J5ZvoCCVmxPPQ
ySktbBceJkxLD8zg6APVQ4uJ4YCWJtw3/BovzIF7/mAN1igMCc+uZ+JCHc/AEiOk
H1kI3SbQyFd0QQ57u+f1mWrgilpGAmsJY72aGs8NhPN+yfotIYrvh9JoG9VZM88w
oh7mdhMFEJRPr29Wuc3fDDY6UBORYRJ6qz2qnWf1dMy3aPmyumWO/L7vEhMJCPtX
QsHdBaG6A7cUD85LxOYpXCM4GiKqZTjmq6Iap1RXWd/xJ4ohPG8O3fGQvry6aQ8t
TPQ0sHgdkT7jxve06NmMDSXGohaa7Ax8MMcdadP9Iqm0vvXpZdChRYSyKK65isjc
AZM8pyle0ACTyYidSmTVEP4YA7OtoV2ClKo7+QbMnAHMbMFxhnHYm6zbFUXyMINV
7A6t0jnVy6fqcugxqtJl/voaaNHhghQWMzesONL9FXxZXhNj2p+/Rm0CvoRzO2Hc
y63jmSOzbt2luK2I1EWFQqi0HdYc6VWYr3vuwwQukOWSqIeRosNPGCER5V6xz3cw
SjWw0/mmHVzQN6PITbL4z8kOIOJNeRzdhzokf/DYfdy1J5HcNCHuc7njaJxwaAjp
A0nGxu/fPEmqmfhmh/LzWH/aqehoH1TWHLW51z8datb8s3PqHbrURF+96GzfKD7r
skGeUv/1Ftk7BR9eXqFCJk7u5wFX/+e0k4J3OaYnoztYWJT8yZwaTLtVBtugEeEZ
YrEtg2JCSE3vwUk24qh2/A==
`protect END_PROTECTED
