`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iXG8g9zRKuH71hQuxxwDyAUNnZt9AQNM7Q4+CMMFbtUVsVKTQtr75wr3h/J3TLBE
yZsbgFE+oykGorM86Dz8geAj1Bfx28QILVJUSh8P9DqDYi2Tuw5wprzRP+66gk9Q
UiTC/9JR/nWdP6BnHbU8JyO7ZkP4STVW0qtA6H0EUQpL4TsmEFsmBLuNjpDEt4V4
fSiUQuUgTcKFmuocUHCD/4x/xi0n0dvkI2wgW4431LUPxlHBJfQQQDDgAXkA+mQU
pooXCZWRXXbjPv/hoMVIxR1vWG12BtEiPnAsdBRanQjZWQ0NQGdMTNBYjXuIdZge
GJ1/T3iLERpoCPrypDAZbfDwkKvvT+04YLaT2GODvPUUIpLzi/6kqxGSShSfLre9
C5WubRvHHvdy5fecI34oGKy4s8A7nxBJ+przIe4tDbT1sC7OMWiIJ8JIUUGFMzKv
Y2mDChyN+/MUSOJ4F6Y8wFMK49h+BOOh2xI2pZ8Es6ByqFpImr9+usJBV6kLbWb5
eqCaZ2FK9ySP7n72F0vUk2Mvbm7Or1b9Z8QgMFjE8Ak/n6ERu4vLdoliTHz9dFDn
lMFftdDfzkkjrWakugA5nh9Xm47AnyuaIzkgrNcy+hb5sAWrOrHx/CO4LhoPtgYw
YFnlpJxnzNcvcvGgu48vHA==
`protect END_PROTECTED
