`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zVAHiWilxfQbmGyn1y5VdfUmrJaPPr3ncW+b6PtseBlafr6zcrQCnmG6wrbeOOG
t9jY6v+H9CGnXz9qZtEn83feao5KA9rwOPCv1M07uTNSAqcz8zJIzQxTm4gyV65E
tg2OhukFps+W1fDP2MBJ7YagpMAVSdJOXtv9QmMx4R8/+djI5pCbAuAyXnvl8Pgf
18gbWtKBxVutGgAewTlXn0YoMFXAB90P/fU9/E5b1lE=
`protect END_PROTECTED
