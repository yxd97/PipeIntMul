`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tOlXQ0XULlvncRK3EE3TaLBVEv7XIQO0DTcx3a2Vs8hgiqJZ/sup9vxHta3MpZf
IqP7c3hf1zaoc1zQtWGSAkOGd53J6fCKbZ7XHqne0Dvme1ZAdESTmH/TiGajrxnP
SnOtRgdLpMXW+GZy64Ry4dXdM1BYILFNr6wYzKTlJlWNoBLsXjnRo/jgu/2R5eDw
C5qHLJcuMxKOSGcf3YupVhj6AmSg0s5ro4rFSic3T/5I35nkCBSQ1JjQ7NLL7/99
v5GzaaRvx+c+sToWrZSriykxmZEUZ83UaTQ69QmFQF9lVav3bxEhvBeUW+aqB4zk
Lv8FpOci7Ust1vbBJaO6sjG1NAMskH59cXtQcoS4C8K+fVSm6Up0GK877SRTMNgd
sRAIf7GWBuUXrwptKklmOzmFRgH45xM0cthisnw2+8XQwDuYeKREdiZfo00mvCFW
9rx0Ou4BUzGHhX3giK8wS2neXlmaxCfNRURtm30fMkE=
`protect END_PROTECTED
