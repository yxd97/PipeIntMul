`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vxzzXF9tyfBqI061N4GmCUa1hsOriHkjLHxynm8XJ4lLKzeM7Qn9QvRsw7Ay7dRW
UMv+BhatPlHXBLoxhhKmNn6SCs5e9z5AwPAyZ0+3BSUxkM3bIWApkOw1PDbLyJiX
rd2lMiBzh6Af89cT/PqEH1tmXoQIwiQa+zbmn8ffdAPpo5cROzttNrPOnzasWKpv
OOYadDuyzYJ6Z5YFf2nZFY+InxLHGiNBHix9ecB4l6CYV9SxL2AMIzsLgS7byc/q
kgBngbq97IPcR76u/kwNyTjkwdJ2XUSy3d15IyLFyvwkmPVQW0z2uwSSUIvBiiNx
SElVLJTGv63/r+2XTzCylJRLIkuIlxIbLS3XMCf4JBFEZwGZJZeCFC4wn8K9437T
jgewh7xx2O8mZP+sEmkQtItx+oqD+OecowCxdc/cuprT7ZCtIvOjOkarZfxQk0Uw
grlOHkPQ0La++sJjqRxUFo+GXlHwwki6rKaRRWwkoedD1HEn6s6HIns86EsZ+Z9i
vXnzQLWEPb0UJlDTxlPcMZlbDtmUzaUGT/u6s/rYQZGvgjUYP0P29GuzuxY1w6CI
WX1jYopvW64tirklgKlW/w==
`protect END_PROTECTED
