`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F/yLUpilSm8DHhNNHQ0XjBafy2h1zN5X294v/+fNiKiAyG/pCtNdDKCdm+6HOEyH
hIQ2WMmzpoRHLShIXpZ90hLXywU3lG+sjXVcUMZbXaE6sTSNpcZkGSMwnU217ult
SgUn27Wod6J6c/cWdVyo9RpAdI8KT0Jz98ydF0U8EIW15/FHhdUyEjfamOtkRi1s
pCwK4Yv1/IcoiTstBiOVhdeZhGyXRR+5bKQdUsjs0xakXL2TX4rGmYWtGUUcMcTF
77lW65z11hfLzqGY/ja2U9+2DxN3L7amJOuR1dZXDuPB9wWtL6PlsmH/Bjt/PZbG
+og29E5xUV+d+4V5JdQi+UQjh3zMx4XPWg3TNeAY+64kipuER50SdYVv3AoBNhQZ
NYgswZpNGcfDLLbaegfqXKGQESy6ZiKjVx3Eb+pVn0c8gGOXpsI57IOe3dpPPUP7
V2Gb6vHppfwKQNubYzE6FSVcPb9zqNd+V1Mt0CLOOX/ZQ9WqQ3VUMMmdfVgca5Bu
YWdhlniIz7PHDAeNTtNVRr+EG0X34/ap0W0VSqIO3qhcuFiQWftvXHR5LmR3rrRG
/l/5VgtvYQWAVT4PXw4ITCyAAfFz+QtXTzXcH+BiP0M=
`protect END_PROTECTED
