`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
msB305rT2q65Hvs/X/ablP5NPop6pmZ8cpbeVvVmNthgsd0ydKZg9obgEJO/V2O1
mkHPCtdLE/jfNOSM0p/ynNoiNYwlwcbqCvEn358Qs7N3/wZywRKqwCBlpfYwp5Wa
25zhmUQhzt7WTO+Kt9CBpW1UytCZkuBHMOg5b2Enmgn4L0UD3SxP1ZgL5OPTnWeJ
HK0DHc5lFATM9fDnsmj7TVcHjYHZDUaMgMs9HrfufrubyktAhSd7G6eV/ZM1IR0X
V/pkXNteQNEE1ByAzBhnvqpD1oURT8C/F4qK1E6WJj1Z2rEbQM0CYRsNPkepCrua
wdvtWq5s2Rg6c90BB6OAtn/SIVoXhIQ0QWPlMZpy/auoPA+PxgnD+j3z/l1B7VHr
2lnJpOwQrfELGA6jsEhoVm4NTKyssdgaoZ58jrxk3Qfb/8IYigC6R3UoFXIgciZg
aHTMu4GTdeaeeVym2x1aSpZy7HLIkYcHkJcM5i1a7adjZ2I0jkMDDJSgEKO/Sean
DtRkePvHF5VAZUWvysKZihUwAcwLDTZo5v6EXe+Kw9+OJbo6UHoZite6mnYwCFzq
uXPFP6ecK0xd96gH/7qVI9GFbL4ETyqFEbgTE8OBMNF1Y+nNJK2DDAS/RwMKWh7x
DtYJ8GaRI6Jx+HjsveUhSdlhWm1nW+yMxAxxXlMtZgE=
`protect END_PROTECTED
