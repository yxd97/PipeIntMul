`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lyTXq0QVuLDkManTB0XFOUlxNdAiRsr5vD4Uv/87cjO6TEGmAf6vclG7QRVEXgmY
aKORk4zCZkihqM0evyc973/PhwOc62uDocOohHsrXE5PvJU4QswqmBaq2WpWoPW/
EkUaqxSP3rJ1uNNNgC4zyJqiLpZmV6WzuYoQSj7u6MBrbXbIOve5ZDjmIXq56PS8
LUMtKSmvJSyx9sRaeNE1dydsBxx21Dab18DGUhHKt8KPEEglMINtXSoCRwqxa/Qo
aGHfLm3R1K7OR1gxCbrv/ZFLqQfIyCBFCSFiT+/wKIDGiqokLS3m4KNu3UeX0jHt
xBk0J6B/gZwlFmNUiDclyg00CsUumQdtYuV9k6s3CvBIBoEjZnti7vOrA0EPfROc
YEsQ0pCISGxm/FWW/af+kZYBHS9nc14jdlJ7o7Whj3CcupgK7zR3Own6vs1g//mq
5OrTr36s1L9ojZb2dMgMIhjbnjzvg2eXCGHlomXmQr1QfrNo7Ck9mBu+YPPRdE7A
/Ywuc2g+YQjGfG773RpCu4LfdiRt3GBy2vNnR6V27HR70IwG7935IUHV62KdW3m5
y2vDXDQSVXEWZg+X7WM48vbxSPtE0XaPx5i6e/pQ/SJ/UUivwMvQuYLNmc7Trb5/
UfaQ2/eV51Cnz65et+MNuhNP2FpT038UVThO0fCdOQVnuLIBFReWC15SKqyDo1HY
KugvDIKjWnHb2U4qFN3x9YkfA02lGPy/yde5hro98zlXTreLM8kCjIASFNd39SFL
`protect END_PROTECTED
