`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEQ1iCJtqrGCTk44nDEy9tf+jxb8L/KS11q6tU0U1xFq19AZGOO+67KgISZpg5dh
XiHf6erhcpcEr3DRdbmIIbeZZcP8ccot4wZeYQ8l0rbjPx8GmdnnURgq9tIHrG3R
x8yNwxXe0UJRThkD5KRnpLZ0qIY349lxF9i7oq5StQtrL3oJK0ThxF10HVS2/p6p
ovXM8218A/XTR7o8nvU73oM9iQVcxnNA3oKvpNF2Dpre1K7XOUhW+Uftla+JhdhE
G5YGpyPOr+LqZeIDY6jKPgC540D6c05KJ5zucNdjZy5DFbexLuisDsKs9rLWDfWB
W5mJ189/39+3FkoHBcwvH5q7fYvuV/LCcE0zIrvF9rvM5xpJG3s5ZpMEvNx2PhIF
Bz/BBWETspJBxmeDzN63pjUCQVFkopvg10v9wTHfrxK55IYozZHvp7G6TO2hg4kD
aEJ30HhwuguLOjGhQvgW2yP0D4sMY/QtPoAMLDfn7HJZhvdC1Wqbt8/Os4yu8FKr
Js2xE+GWO+VTkHGYw84xdXPz1b7DB19AegCiZGfJ2BV9hDvftMTxSdBXnfR2EDr4
hPwmYZU0p+tQv5LxYalGL4G2FPzyWJvaQuNSvQZp5WPWvmy00pECEcJ6pRKSd7x5
jy7q8IK2dhsHXi42WL+nMg==
`protect END_PROTECTED
