`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aih6bVD1FPwz+HUrJiH9GHferNpqfGtR/yeVOn+QJYRgoaElj99mDkBllxjYYawr
AevdmpXGG7acTAAT5M5t7DDdO7/2hLz/2Eeq0JVsQG5PKO5TUH3+golPhdai8DGj
4GHr/ceW8/YsEVNBBuAotU2ZH8cq/YKTmw922tLFvG/mPnMrJvNaMzjvxraG66EE
agDcAfjYHOSq+CRaytFwhLwYtt84Q6gKIKopEfxkacvC3xVOu8kwHqQ/kOsGJ3su
IrYIuqiQHdD4YYj5LV5ffQHVZ4/FcTVq6T3mmh/6jWNm6ZZ/mrnOvs3gQbpwLTPr
/IMnC+miEUeyTcQfPQmpv4pz+Xd6IdVpibeaCyiPmArQlmsduCh2FJF230+5UNGB
b6hbbFVxZ54t0wezGVZCDxSvGPMxIL7l1kKln86k6ZmYBHlXe0deH8Vg2td93lfP
VdjuDObLnMbn8gyvszHmmOru9m6HZYujy9WVHNhCtAJqWPDL5ahXkq8E1Octs6Eo
DLXxcaGktoYwSWQfZaV6pgWTo3RXe7p8YU4By8tNLMjd3zbPAAYdmTG+4pz6jR8y
W19amMoBSjiD5GP0kY3QEydrsLv6KPRnPbd0HY6a3JEi1aBpplyp9GyXBFk9OmBM
65yMkN3menwjNNw/3QBbZP7Q01mngRUUB51+BGW2qeYkSfrYfEjER0nQ/canDYuc
zEFUDXflcNxEr5TxD5bOXitYUb46HxdglzCLncIaQu1cP7CFAWnwJzopXDyxQPat
5NtzrMbuPpRNmLrPXkjyy74aLBEUgVyg2YDQzoiP3Wzo1y0vrjltOTPqIiebcfR7
4qANj2Bn/yt/VJkuR42C+YAF397uR90zTRx/wlLj0wE799XnaOfZV9Yb362lgTTN
ZIqwPkCmTtpm6rh7x2G+Sw==
`protect END_PROTECTED
