`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9PebO58YNonTysqSPj23d0AeZrgXM5r1ZZfPwYgm91s30E8pZTVcZu+DQd4obxbU
+UlmjDRBVqecN4Wcgx8wjOugHdGHX6rxz7zcjfhZ3ZkHzaOBY4FrjKf6gEAxCxEc
edrsGQ/BcHddtPIGOHaWopsmPOTALvw1CSWBgucr0PMtqGaTNA6PU12r4TAIvpEf
IC17VIoQLO6TxNJaabxzDNYFJ5mrwl6OZDuOXem7rYCI9supx+y+kIrWo7Wxivb0
5PxRfaTuQt5p1SDAtyBE1Fby0fBn4yf4TWoTGTXEPPEVFKzNvdBlIN8BdnuRVoTe
`protect END_PROTECTED
