`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HAsI2zKpownmFncH+7VF6aUrWKPAU8m+hPaTwnyOB69jrZD9hqVd0/rbFyHepllL
XFyouO3fQnBe6evsD4k0gPn7AikNiuKllOu1Pov5yXtAV0Brlwcz8srfgKgpQGOf
i+yX4xjICwOsQWMYUcEbCqgZhdFfCIWL+BHmLwpVS/7hZLiLoXWheffsvIaQe0HI
fnXYuSCYnmxC/qRF5hlGDgPoY2ZNyzOb3O2lOtdTP9eczebQIoup/02XxbW6+vBn
cSXOxiIVVV11YKSmx7QpqPPyLpSSeQ3BdcnnTCpxmTjMJEliNORsUwlurBQt7a+N
ALbs5ILEY5MioE15DT7ol8Tskidw2WMImO/Qc5Q7LOh4hCLqIVuBm6x0J7Euw4qO
Va55Yv61/2YdpHSygA7yDhBfd+LV2fLzzfj8O9RGZAsGhkXoCEJ8Tngk1BoWWtaB
+3XAgogCZMv9V4f36wdAz3PZUa4An5bkR0Sz7CW2K7+YaOZlCNu/WPyf27WyiLaC
yLY7pbIQFpJybp5GaWzXfKy7a7Ecjm9p1Sjc/PTmFzd3CetMLDZ5s7kg8kV/+EUj
`protect END_PROTECTED
