`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GP7oeexoIAq5pgavrbOSwdITciihEdeyRpRjLTpSPiyqdLURe79H/0pZq9lyNkFd
Qr8EM2btMiiE047XuMH32VIRXqd0Td2AiSvJnxjWETyQ2yhOL6Q4WQnESc2ttC5+
jYEHp4XVpFTAG4Ww5n0ZfsjN50qo/b41EVGMPh7gP9DI0kuF0P6H6QpNZILSy8B5
b0ZWTGIM2tCIv3BM/RVpAm6PkmFS+RnBmhiBMPKwbY3uOJiBiRSuBtm91Nq8f1HC
nlx2MSALTj/OVYms0GcS9N6lrtn179ryjlVasdO7+V8XqRg8JFZQ8vPIE12qX68B
hPijRWyqoGTGAGGUsw2CLU/qBKIJ/UBBfTgiJP5p3p20E1jVzpwoBuUkSOdAjYJ1
`protect END_PROTECTED
