`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AnDOfYwzc47VFnI4Z5CO2hRMDB/hEUNRzspBEy8dnJojbf56U6lkbtX3UR7Dnoc5
O9bN+vMa+2N5liPB3BD5UfFeK5kuO6SMwlXc0wTFJVIBPZ8R+/m97/5zjVhrggBj
8VgM3Fa/Z7vI8895FuA8+MUfPAJrExvfTP6kjt0Pv5PPOJLteGeNq7l65gW24Jlt
QWyxxhLgIjzJcWAfFfo9V7ONBPBKYYetx/xEhLDjiA1DPSL1ZyzAnnt+x2Btsf+V
7NtUc6NDwwynU68jKKJthYakz2o3xEhv3/+VTmLiOszGjopy1XDyrh1m7d9yDmzP
9Ed57CMdneqKeQ9p2pULNhXz/dR4ZkRDRioDZ2zsXxg0odH1fmlYD2Z0dsAL4z4n
4M1V9GFcqK2AgVRXVSfm/cLLMCcOZSkgTX+dkHvtfn4SDq3vzW5biKcHXHTMggug
`protect END_PROTECTED
