`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yX+uahAJVrfu4IaJvsddWC4ZHJOQj/8MirSEdVDzflfRg0S4ViOtXpewNE7UDQur
163ZxN2Xj+bhgnClYLpMTbNM/vA/ZO6bkJa8Oh0gBSYW39dRCsb+YNSSBKpoCv3S
mR7TCW+LImv0t15dRd8hCbKTvL0rPVuXcosdHgq0Lw+bCjVvgiAWIoHkMyZHpZ+h
ZCyx4FY8Z+t9lPfxxyykynr4nBUKP4H9/PgMtMmYbptj/76iZklBdCRHkQImpi9v
XJx71gyB8TSLXGL5+Nv3185WLKV7puw1BGv7C/2HmY8=
`protect END_PROTECTED
