`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qj0TaeUyo1qlrIyJpncwAqbn2WSUyYtceyME9GhabSx7y1/MQ4tbmP7FGX46PmzR
URWS1OImVjKQkqjKwg7+8Px/Xe0YcVH7RIPsBR6oilmkzdlx/uIi6pdzHiCZBsxL
ztx+0GvLT7A48pyOeDwlZl54PUWKSAXb65NpjivhXPl1O1+10IVl8ZuG9zYsc1Je
atekWqEV3mk2q0Eplr9QTrAKZiYfs55asa5pWq6ylWi5/DGyXKt4kudgTV053wbT
3ZekmFoCMEc2j1AC3NM+2g2HPA7wH6xCWusYRGkLnbtkmzMXGgMwxArySbNpyHcC
0b7qPfUC9YuFVFOjgqkw20Pgebfyh4xTrT5zfKLhI+Eey0+oUt//1BoO0FBD2qSZ
vLJXPXWrnkEtNuc4dPC4DUDFcHVfpfxDBlPOjFAiv5Gn2DnLx1DusNccqlo2cWFc
ZmV9ET9fuObyEvEEGCGKXA==
`protect END_PROTECTED
