`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yC7BMucC0/KX334VPk4rZmeQpksD/kI9KNSXcXZE1QT1Bi7RS9H0yLstk+qpgP8
hS+IOOVl9NntkdmLT21MosD9u42hR5eygp0l3lCC0yq0fMlUOmROgPNYXEoN5XBt
6GxIxoIAHmpJBWUhy0vYd4AcvCl1mRCIcGVoDEngFr7lJ3vNr4FBN1ZEU1+5I2Cp
m3Xu1QjB+vatg43LdDhoDGKLmphc1eZzdA9KVh4gWtDuHv5iMbeUVjnNkEKC7xQm
l2QdMYzddhyn1vUrs4CQC+G8kltP+5Kh7eHlSZGb9NYz1S9cOdSf7JnO5sA23MTe
OUmzPLhUcEM5EFsLmuhdWcgTOvic8VPTEyIrKJ+eAQD9XajakJitH4donCmRns8w
IScTnatLeKBbrT1yWEVTRqb53rbqVUfFqSfMCGSlkOM3tXmOHjZ9IxwKp/oZvZ+w
A+zuA1WyDoeeWvRjSkBSTovFK1oJhdlkP/xBuKvI6iGOmAvQ8cwBqrq0LermG0QT
PdHLseaaFRrngYJzRBqSssUm7rKnyzBHfO+owfXnNU11idGs2YG8wFvH3bdcRt5C
Eu0wxET1bGyVi1BCYCXCsuBLNay+c5rKD0549n7KrL6p5Vn6v9tPAAjdWav3blhA
G5Cjlq8qUN4QQf4SFqyYy5QcsDCeKDw2oGOy143pI9AczH/b912MBLhF4Vr+9qNq
Md89ncpdDWfL4amEG2yOdCvWZlJPae+sDxI0yZl1q+M84junlUJZMVdRzZPjBL9z
uFdejHRZzvaFDcZmJpzGT/RybW3jO1SB/Fx2Mufang6uHwTuQIVWmG0nX60waGPo
ZLmkvSXoJ3fh144a1lfC+VAeoTqrTHVlEOXDxZAxsVzfPGYeK8fgrLcAaaBO4lO+
E46cl4Rq/i+Bl7gVIji7dehybwUK7P/KIZmQggD3CoSMrasrISz3FfTkDd/pJO79
0OOhX2AWPWbd0oV2rWD5k7iMrQFb95enMRrbNW/LPcFMbOlDMqgwvQwLoE9oyvjt
MWT1RApHSAadNk4G8wBDgask+KKjgjq62AkSp49cc5MoMh8V0nwjKSyoi6TucPLu
vXpT0kdtOOnYT17KyKvG9P8F1tT7wm3ssMt4scdyRpIjWfGR1mM27KXldkI8ExyQ
AijD/Bv5YE43zWea9qVrJTujOTnoEvp3ImQ0P8WaSTunX+C04qR+P2Pa3u1tTzo0
vxl4KK8UHVUfxAgWZ8QoHzH6rrGfDpGxq1iZp50392Mt76H2JhCJ9rozSyFu7ZrI
xxisZV178VBoUObEQze1odJsElliPAE79qnsuiZPgRmIiJFB3qZRx2pTk+PXvkX/
wRw57MhHhuqPtBUB5ljy13y0PbEnWXsdeJ3CxBn2Sz+MbEttfa6qiOSRef1VsJBC
liIliuiYr3J4hECratFfKenLDNpSrBLCv/pAWtJEBiflKoQjpuAsRxOA0hsqUP0F
jqrk1A/p3FfQ/lvoadvcrP0KFU8zVwceBvkZLSnHclMqU319ZExDc2FMERDknwrm
3Gk2Sgi74rQiSAxoa0moFXsIxXacxCnCSkSDrPJv+KcLJRR5yNZGcFypAyxvMv4H
h6mXj15QWMCx8fffJrMZXUuvDS5mnGOFhZx0ERckgK27Z0X+iDZLnmitBZk1GfU+
lktH+mZpTfxi2YwcHhfitxXVUAc+jIckSsM/Pmq4rXXVEXCZjT/myLniphvH6zSC
C+5M+asT92NRcbrrIRfi5WHk8rUJlnX+uJBSeBULVBd6W4UN8B6GEXbZB76Pu7HB
n7Cfxh9tqUaRyUmtrj2fpTbRFGp9Va1lxtTHCXgU7iBzzQqEqwCpOrIjFdP2hTSZ
xOV5tZ6ZFTYoucDTyeZ0ifG5Q6tCE3d3ZLvv2SQ4KKwoNH1aP0uIi7xaTSNF8EGJ
lddfGfkwXb+oJYNGkLPzGnW9SPd/gj/2ETtv+ywCXwmkSsk2alQvSpZ2ysBvKHWO
i2NQyvCqDjkCofFYY6n7xw==
`protect END_PROTECTED
