`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K14wO8URXMK9EYg8SOCtTKKf/cQRfSBYU3dioLfVPgCKQvYpPqzCNE8oenSX6V3u
/JzzSp7FVmuJz2xiAWt31BvAIThg3tFNDcNvkiqmxvEeFJPYeGkBmt6hZwTGFwPK
aIsgtEi9POob932afJ8Z0lTniT0W6rEoT6+bfQ6GrwegqXH3GKvYEOHbvoP8iGOO
rQVTJZw7fF6mj6RB+mg6Q8Z0lbmxU+Sn2jWwWCqFFnIRxC/n0RMsychsy/cRK0yA
eiO+w+DNUJW3U+Kk1Uw9+Fgs9l4qHNc1gneEoLZxCbxDQFCYdfisns3VCzQcBXSr
`protect END_PROTECTED
