`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zEG5Ja3XQwDNJTZCh+TmlLGi14RgQpmpgf69TdwYqs34fdViXE8g7C3tD3baYTvq
k9SgbdW/7V6h0J4VC1+por80x1qsu/AmdUVJFItC/2lBDUVv+llM2buZQhqH+vEX
NQCfs3fohxqGNNmzKXmpcaGd66+dJ5O0s3bqhJjaHuc4OyKijHbdwBzzcVU8KQTZ
JIZoA4ndXrIiUnnYVtsYHPwG6nHOrBBiHUjvKhwwwdjRMWf39p6ayiz9eBpcq5Yc
y3PX34X5FNQv9/Os0kWC0noBY5X7iAi6VBsB9oDz3wEHf8CWq6Qd02RmlCkx/dC5
`protect END_PROTECTED
