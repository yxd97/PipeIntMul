`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4NgoM3jZr2hzDzL4u7m+/xXhh3WeMn1OXeM3ZamJNNF9/OzYvfTtXvN00zcFl+3
nsvlN8oHsKalcCSK2HxXQ0i0hWRcwWfhNtO8EDtb8imy33sVCcJXUql80qunG75D
nOYVxtP+NY2Q2Zaw8LPy3QRJfw6Ob/x7mw9O/eLlJ3DVP/r05IaFNNWmsyTDoSLX
+uTRcUjPGrIe+/h/YFBbU2TfGnYI4Dj5jZ43mimPgi/IgVtteEKWk8eGMnSzpBJu
Hwja9fdoO3Xda4I2CglmqSlC4IySbZJYFohVuZ4guiWkNMp3HXTzrlU0RZOxnvQd
b4l92wEym0RwOTXpnMaSVM//B3uBRYV62H9h3v6/bSEtwlNw/7DehQkUrA7PmWV1
DSKzme8U3psUW/Vz8+b74IbnYELQiKQnW0nCJV09t/RBJC7F/cV5RCOCH/RcOgk2
`protect END_PROTECTED
