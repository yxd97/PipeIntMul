`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjxqEQudXUhAfH0aUidklASs1sQnSEQuUzCCLjjsy4aUIKjp7DztekXxWlZ4UQ+4
EDVTYPKLq5Jaj7V3gP9nwB5isbvLC8c2bhEr9iMiLXCB69Ur4Qva8hACPVcffdOx
4Ej3880u/13fjqd+0AJVREfexid7C+8WWcQ6X4Quy93sS0P63Hqs9gFKTVe/TXcR
pt6ttt9v9npLBEvBbwpRxJ8IAK9yVwBHEUhpOz/iE0jTBx7fzfG6gBJ7a/3AZLmd
VtLasj3SB4O5hcZZAMn3+wl5WFS+28CAlditle23A9K1fyT4PbfwKbA++QoRtOwf
Wk6JMyPWISyL5lvVuLswAA==
`protect END_PROTECTED
