`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zm8GT6K4gT0WrTVBZGi76zrSoJoB3mvAbpgqyskDrvchuE0jzZs9KtCZEF+bBaQu
Szdvn4uXKSsQVekznv+kxugwFfNqepfcvXSr14XN8SwMsE4HQBAR2JbtpRCwYbc9
ddSf3FeU8Wat8hY9zP9+OpBrJpMiBl1zzmDBLqyjl5aBHibNhoVBPp5ghSSbTOEU
5sGdSCx8f9scsYriiqFxwASpvfdQ29XBHfN880ndLK3W4Kc0PmnH0381kBYFSzeN
duP3daL2GkLseZ9xZ3ZC7A==
`protect END_PROTECTED
