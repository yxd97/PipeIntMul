`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Lbh+tn5CZpyI1GQBhN0jCpCwF1OWvVszGnC5m3Cw9Y8IFqvk0VOBCzpMJF9A8j1
kxSYOt+5yMAwRnbe7RAbGz2voSHS59RFLHvmOGrBLH1JuUsLWOoowx3NrzeycI36
7xUalADPYy5AIrj+Tewj+sESEDAOeQrf00maC+VVpnMuUoORoamdqvcJAH0l80eA
bPiOEiVIX0zAPkhXf+1SFOZmPaXvdx4JL8rJYnX8b+oclKNq9pp3ATH9u2P3WHu4
ygrg1iQ0lWZJ+8KgqNYGnWETTz4PaO4IWRblY+ssrMw=
`protect END_PROTECTED
