`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
whZu/pztEmY1imGVqWJanjzFq3ASkz45F0Qj6DiFbumUjpNIMlEPDhZVont5ODD+
G74N+j5i87mWvzysBDsI9NSo2aBFZ25PPkrf7n589Kafjzw1oHoWqVcyawcXDM1Y
GbWKL8SgTNkz6LquzLS+4mrrlo3ipa0W5GrSq/5BVIgZ3T++9TWGSfBhb78aRuKy
F34dv+tkVeVZ8V6Ki0XhFOoDrTAg6O3Oy9Cmb9/sPX5wkG/Pt9Of0bG21PM16SKa
uqNMOBAzgxZzzex8SoMpp+xe3/y8rFPdYEHAXOXCwhaGocQPzFlPuSRLWGk8HpBW
p+jGwPpXg7oNUWan/hoXufcZxBZ9EFCtPoRjUUT8ZVDMSlFCxr0LW9WyvlmdV27H
DwShzSBnFcVLKS4hzBwRN/Elf+0/XBTV/dhl08xxqCLR0BgaSOg2PNlyzDumLOw+
kEBYar/uhvNb/tAoigpROexdSZB8xayP3t/+IN6RtpQco6ZgG/i+dCM5a8gbfINf
A4NtAoAHrAo8FTgat4Ct47zrM1MQ2EpuC+nhlOH6artMqGB/fCJEieIWOweMetjv
Uwfr+Jq2NN2xijGgyIImugB4ngWduScurUo4vl7FSrJwp494axJQ5itNXyzkgFWo
27JDwSevdUTDma3eSQNo162kveTSc6kAYo+eqwhIhY5BYBa3d6F+cTSxEIepfQ4J
FIbv1Vyx/YoMffe5wTdML93NnOfUSuv9CPe4OPuWnKgijjW9m2dEAb/DnmED8yeT
VztQ+0/sT0h3D9NxOwJTG7KBWpRasifOe1Tt66xHI+5f/6rcYjt8oNM1eiSDCc1x
4n/dOukRIdRteY5ujsT9EMm81WvpUtLKE/ef+8MGmM6Cp0V7lqUv9vTXUXAJetOo
tn/JSK+3VJ5sBFflvviDAajwTZlbVUcznVWSVR6G1LtbEzcyYUHzA6OLDSmgSo4L
`protect END_PROTECTED
