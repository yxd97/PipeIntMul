`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rcnd4m87OcOHn7njjo9KpcpDc207n4AzrXNMG1xyNk+PUwqpBJne3RYqUwfG2hRh
Ftkjk7bMF4EVHflCCTIBds+t8klm1i9yBLMpNu7WgXIbmqXJSC6kNY2y3Ir3fV5w
uscIa4ss5DaQT1hY9JY+HAZi3iYT0uHp0747+IwiOk8Z4Q5o6LqbzrnkhfyhStD8
JQuSvdTxnHH5h5BpWvPu8xi5s88XJeFGuUoONFVKp/JwufSQtJ6YSh20lDwAlvrO
9828rcH6mOWsxdxeMCBsf33hTwNldin1oJgMruBzMG13Fqi94I0ZhngP8y8f07qD
kSHM2vSkiHoogZHTl90m9wPtoO5/a53j84Ippfatc5L3gQYXQAQ/5w9Hc8MrJdId
MXA/iQrEq7KIZKHK+KmdYwohSNrWbSZTtlAd4k6rDSQrreXs28QC3vE7oU7YbnBH
9DMzXVAA9kjYRQ9Wp/9skFsv6vTrEZIAvvTSJ2WnAWIjbr8631mfnUfFPkutRhm8
hTs7Yv5GphfueFcSOnbIqcyIYRu3z0qVj6Nn7Di4hVNXaBYAixeiiM1BCuldYmv5
3fd/D3vILc1kybEYD6hcbj7MAYmSUHDjJQP/eU1MzEE3O6Z3l86wLZgfyq7OL0PS
oyJrO+j0FetwJu9AKH06oXbaskOGTTuQeF67Saqos3Fsww+SqlS79aSBcHCMZeS4
rxLWFQrVmLU20oU5pZdArA==
`protect END_PROTECTED
