`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bUq2LcV3qnEI2XsFwE/r4IFgyYoXLeLF5CGsFi7hDHbvmL457Ms9oWys1fw+dNKN
vJuTLDrKB7hu4cDXjve741VXtNG2dOGxbVyr3iYqsM03DHrZy61nWS3WMK7xutKz
IQPROGPvBpcCEiX4TRiHYW8obwSIKSPVbzTyifpgxWiBoFmbCrS//aiiNOdWSamj
uUBFVTzwoIvrertUfrv7PstQezDA/rQMIvpVif9qk8DUmE02DagSOUKCgTmQPbft
+hJNZRIbgaRngt6KNspNC7lg+B5hE853Bp8tTjoRV6FfhwqeLNDXrmYYDIdYCreH
c+3mSoi/VJ8epnEpb2V2lEvBEY0nG4QITS127+QGA4SjnAbQK7nKDzwpiyeN8mbM
Q2YzMuDA9uiXl/d6Kii9xdEMMvLV+UOu6X5RmauQLpHrR7hWig/0TVNxeXzfq3/j
zqHJ+lxEq3c231XED9h/gNXc8KqXW0zfpfOYYaIeJQ2LPkRL6dcysgZO65/Jlkbk
ulQH8uCmwuxQHXpkBWcI1hzlYVYhVhpemYy+78ls45P0K/KTGWuLvNbEkL8xClza
uG0Nqn2nmc1eNqjINl/qCVW0oWhR50k94cZ5R8PsM+Wc2NL4tCV5aZQvA+gHHIPL
JxhOEeaJqQ8D4szqe+i/IQ==
`protect END_PROTECTED
