`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6EMe/WGEYC+p0PcO2oODo6yV0luifxQnJZl2/+9ohM9yvic3opugn9NPGmqNjMaq
B+ISXLKNUux9MM32vsY+Y1k9/BvCpeM8h0oUqJQ5nJ4T/SlvAj6unbVO9CIsuyOQ
YdkRjQWrKCqFz3dVlmKazefFW0lajJVPH0Npim3yZfBK3GtJm1S+qWERfTZAOxaE
JsiUQr+/JPL0H71ZSZEsgrqQRCYOaN29KCDPBo+mZvMJupcP83kczidu5XDMQRpr
r9Jt5g4IKFmoEJoN2G9mRGIVQdQRU8OI0LC9VQlTYRkjDN44Kq3NODNN7XcCD4iX
OBqmv0IQLnuxJWYHiWmr9UO2RrYEH7qOnZ0uEpMGKmWtfF18qb0xs00qLOop7fpB
n+sFQgAiZJphMk57kx1C+IkMX8UPTyVm2t0HrMNCd3VwoDhaHezJkPA7bOMCV+ZO
wZF5mYSfxVVJRxwqoyThpvrHAfKfgaEobemZBH2EilcF/AMlaOzWsIydeSG6SGMP
qXlGtHBlPdF9SmqWHLrvw2JD/wAy00oBqnTJyn/FOKRtiY2/ViHm11JCPrQ1od46
dDj200t/oRQ2LHpSIz3s83Leluv79uk4zzqGKhO8h2j92x2pHf9M1g8zb+fqmoBk
RK4BDa7OKtx4Wr1HAJ/i3AYYnF4kEazUETSC23u0TLCnT+iCtT7r5p7cpghlLW3q
6exTbL9Uyeoe0ao16rrr3JWhFY5VNKhG0m1JpcSvFKqQQW8x2mwZwuyLKoBDZSQO
R5Qiow8qRFq7dVWRtRdWwX7hwbYC2GOJ6XEA+QLXZA9u+itm7lXUF/ZtetdIb/a7
/X0xzFZGBW/SB8arzpDrw9hggLisq6t9TAxoGLPtLoiK11/O5H7z0xLybP9tnWov
SZvSWCnU5Q8KiD849YbpOLzHVI9H0vv0Wmr5Y/8Mf0hbe33IIjaO3dRiHbNyIVkf
Y7L65e54jWouZrWLUQP0Kyddvn2I1riR+4H/gsFkJUcrGI5cyZi+s//u5vXs3bKK
uAn4IVW+v4E2JTUjzKcp8FIzatFvAHfFESXcyyT3La88NRiRU1P6YY6UnCKSyjv/
a21i0lIaQYTsq3roCVwijR2N+1d1g/KK9VA8cJTfB829/FptkWx5wxeWkn9zeCWs
NjILH6XCDXoXKdihCTlsxP7ST3RjvtFB+8HanLIty8XlcEHqGPKeslKEHf81FJ8p
PNJDoecpiL/RgrZFSPCXrG4mtBkP8mPXJg1omTQGGgtzne1HdnhHsM86FAOQIx7K
v9qrto3VlbEksFJuhViLfKeKKoRM3HOvNBwXnzNGAampYZFac5y3jCfDY0NJ3fJl
llpuafgMami7dwvTFO80BFbLsHNstVttnB6on5big0GOa0u+3v/oNL2di1LOGc1H
5/HowZ/aJ8ijMm3blbMn6wdv8eshE2SoFFnLHA0RQRCfHna/3PjlxEgtsPniY4zP
8OPzjMI3SM0ON4xL+3HkG8B5CK7XZZQORH5LCCXxn2SD+44GaR1QjFUPfx9H4mev
xCKHZCLDRwckw2WvBxLXmGt235VXd6tFfBOw5vI5gkFxW/c9u2mDFXlpVMLrK+ID
t2WV2IndKtgUGj47Fpoq00JDXJWwiC2y8a7WKeWx9lZJAH/6nQmVSR9+lkBETfrx
ljxSHEyRHv06zUecq+sNXt8PSuQzY63R2GQn1xFXiSHshyzOtgrMeQ8ymuL/kmSj
hMreSxChsUB5kchcEbU2VW33AecdGY8kkJOhZw37tz3+UnKs+Bybg4aS3WU30Mbw
TAN/D44ZQjJoHCsX8+R++WkfaIOb+nlE6LhTenyW4OA8w8b4zFNYfDiOvoW+rwQH
LBmM+2rVCYjnooy4Rvn4YXSGfbhE/d2JnVQSuJNotfdnzJErjaHosWc7F29/X7He
rMsrBNliZRs9ZYCRYhqty3VXqJ4qBHP23tc8loM4XUM7IGz7N/RP9n8LGk+zpA+d
o5mUDhdO6R3QTzr3evsJ+XYCN0spOicdUsdPfURPvRiEcjxK4zkhFALslL2KQ62F
y7SyJYo/E+gwRZFOLgG01FMDhZk2ll/G9m3gBzmmFIw=
`protect END_PROTECTED
