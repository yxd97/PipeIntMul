`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQbLfeqU1j9ZakxZdxUTpACf9ypFQg5pl/80KfApp8vvnnxz4TBd/tzP9mzROR9e
0Gw+vL2dxP3CnJSYnqXu7pFywbIKe1xYgfyKKmktAZJBqmNPg0sOHSSgOAi7ZZbU
Df4ZarjfswXEYScGE7aT8gAo6YtTJsUyp4dZwSN5xIB6zJ/lMJbZXi9qwxAz496T
SfoHYh4jf9PFw+s9XTgzhXwXsq/1pPnmR/SP3gYu44cJkx4/Qm40eOMl24gV2dmL
rINm7HfKhrrvHU/z3cCTITKyct8mpGrDSCRGpjOUn9u0SBYeUcfdl3tJMP5XrHxV
08NPG9V9vG6H/mX3ixEoDoVnXn3k2SyynhjKKfqHh7NG1ydkoRrSLreOyUU/pyaR
ktKWjfrL57rwA/7hmMPzsRO7IufNhxRgHstt++390Sz48DgOAtPSmGP/qXak28rV
1gxJYTNAkLhcoaUu9KnA9kmrG+MtqrtajnSVoQH86WCaehjT2b53BrjpOFMFpbtZ
+6B77ZcjiYrtFOCE8+ZqN7eo/3hjOwhB8ZCg5eFgYptNdo3Q4fMZhnCkix9/jA99
7Nd7QwK/hYY6J0t/rRYQKs27Z0/Nhwe0vP/DSrO/AaM70itOJuYDBJn/gPNaHaZp
jAaJSwtxkf4fQJ1u/KNtqQ==
`protect END_PROTECTED
