`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DcxcaohBSc6XRH6a2ft0IOCirbBgKYBNSdISN8SGsQld6f+1UsPPOVqZkw9U3TDD
nKEO9mfPykwQM12CjcLRvnRFbViCU03xDOFpKuzpokbgW1otngceUUzxI/YpyV1a
IVuA2tdxFIbcZOnv7eozwfhU6LXHs1xtyqc+txzUONYQOzIRvEZvknEkpWOCywGY
1109W7iV12Gxnxu3BYWEb3Ej3hSrb7cN+/7/hgArTfTvQZPOLHJeL/1/MacHbHkP
Nx8a6ftAR5QI4oQxeidrMXOlXhVQ4K775FqksdOP1kExSiyUDppYNk/+QXi7cp1P
i9sgsIk4vSsliBSn6TX8VRfJ8ZtRWG/N95jGOgWQtMtQ05GkYcXlhNAxwRnIbH54
F2Brgklob9CI+ZWeW4EzVmjz8usw8dUMdYmeI9Iqvw6vSxjNug9uNiZSamLncrda
afFqne8LaWvk4K6W2mqvQbLb3+qb9p/OFE9riRSiI7eJimf/TF5kUcIY4dHBrJBn
PeZDyTbsbUyEpRXEisTPR1rNgMiL4rUQvqwmivNySKHDCxhBWEONBzHRcf9rV7Mm
CiyCHK0DNCB0e+xviCundUd/S4zuXNszAh2kmm+UcR0ZmVevmQgolRbAI9QPNRmE
LAIG/Nftg08NPwMIhpq//nyIWM6T2VIrSLFjleKPyGkB8c/X5TmG+R5IdG5y647k
pTIE+Ls6fsGQZnxzQ5qWtnkRxQFcWNeJob6nEkq2so3vevk2kFKRN8GcMw9pIiZS
asYwigOyhqGP2jSNQ6tG8j95IcnLN+r0f4fWTa6+b0Y72PFiRL69/wHiThvbT9u1
9Ya7fT1Bb7b+0L04GOlDlqNF9dl5VOWiUwIWnA5d68aYEZTjsP8x7zdQKsk5HFMW
n3nEX0Sqy0RYhtKmiT7F6YRWrX+uquI5P82mgOPpgEqEMIL0rN+ABEBBq7F1PJQ1
pJmIW683Z+sezerUF2OKWn+2YRUzn8Z8ClsHjUGbSFspOKqYk2yb+S0AnNp9RiHu
s7wWzKoFTDahp8Gz+77MBY1xDo7qddT1A5stB5tLgnvrodYpylAypfczKV1tD+lv
qH0U6qG1xGP5q35UkiRUPSQ8dF5kFLFTzAdHjqvGUgHZAp2eVxUSc53KQm2i9GF/
j3QivqO+zcDMDXMVkUqHJUy3cqHiO+GOtMC08vsMg+zPiUzr2Ms3sISgrerponvP
7AetnBpBNz0vlkA0ILgL2RuOmQZLpeAmTZDt59jbR2jLAMi1nHRT6EpzHkZYHcHu
mE1Ip+4G+HOqq8COtUjOZt9OVanfp2kE1C9ELDo02FwsMN2GznmwthNMCGqm9md0
zqru3m0RxKj+s4JO3pe0NT6+kLUHMX4IHQUwdd88Vsd5XFs72HA60F3cpvBswjdU
hyTSmsTnm3tlc6zAs4B+/NRz8dudKF44ghoY4cnVAOfNQK01HssJu+OaVVDJ1ILb
I1gPfEn3l0EGyFEIC+9xgz2tvBbLD4jo6u1mHajBbtjlr2bsa0QtdpCTfTG+iQ38
F+bv3USAMmTe4VmelLiYcrmmtuCceqFrsU3R56ihyfgxWJ89zFql0z8RhwuZ713h
QEvO8Umi0IvR1oW7HHFg4wGK5PJQt3ih1m2vV1/yeyk9KjsbF8PPpRMMZzJk5LGK
gEtZwEMzpIJPArZT1iOzS1Ghd3HpgJBUGDwO7jJ/tx+9xCvUnpP+T/x0yebve/vG
Wnj9iNw7iYvoXX/cY1PwoT7omnJ/0djLuQlGfFatkfkUBMln10tMuoqQekDxOmY6
EUZDktJdB74zGoDMPobJqA==
`protect END_PROTECTED
