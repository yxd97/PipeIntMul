`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqlQClb3xduHfvZQuLEAuUBqtP7/dwt4hWcCuJ7Fs/kur+TqwzudcWwyqGA62myW
XOGK3LzLzFO53mY8lzSEzftviK4cx9ITXhx0m4N94oyBTPBdkHfO7sDlbwLRGUcd
4tvK8BqrwJmdA0ktPVo7xZFpi50X2YJaXYeTXDm/HNI++tSXGtR+hylrlTEdTeWn
T1J/IwWAveLDtE+AsoRb/YzhgSDmfOrsJ8b0cZ9VVkzXpIllv4w4vtUuAt4puMql
Q1vYWMUP0MJU897Dxl2IU7i9/VusZljY4HPphFlCWzuiXjHzchK7wVHs27kZFiOd
9ejEYJwdCfWVOJv205+B367l0QJYFiwi+XJIx8hclkFOaYwa461CZHrEOLn2Lfjb
0r9jSfjTJTARjrj3kHYD4j3xB3mlc4hs9S6pMUyZH0GQFF3rWpF11gxyN58xJrCv
ji2h+mI1kIPB9dWy0IYYjZGjfBtgFpVrmAa2CxaP+Ck=
`protect END_PROTECTED
