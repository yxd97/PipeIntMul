`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMIBs4fvu8RRGb9MSrr/idUCc76mGC6maeZFRezqeHKE1iBFZyuSElbrZoVzbF+t
RiRiJVlqiHvC331W9esirHYf+CVnl6XYHudT2UvkkgqEbMd89LvweCSnfxpG1bzA
5k1gtmVffrefhT31+siYEseu+1TBrtQd0bH6p+lAzSkm04RQX5P+ssAL5FGsj5Tx
6eEpuCmZ4kZKVp1Ukn5MyhanOCbB56zsZT7nLFdblSOnyGI8TGSYIadZALW9KhWS
6lXESZLo12E/0rcc+iyDREwSXTX/T2pNiY7PF4amWSSmcOOHgVy7r8Kv+DnzFDfB
ycFsEBR0bpp4+M/LqaVEAK9J2lHeA4K2n+ifP5AVj/QJ9nHJehdH8sgnowG8cEZi
gTiV5tsFzKpIWMq0wmsU01Jr/4KZxre3VS2z8LKYDBg2XgcFPawFDGRFKbpyAUwX
`protect END_PROTECTED
