`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1h7xj6KgVmDu84qqavjwHmuDkdvABuv9lPtb9HlcdT4H/vkbMlgFqeHv0D12xU3Q
fWvTGzsJ8RVTqAsIcnrVmTCMBtqCNYgJAQQUjHjxnO/yd7o1Inei/TM9bfJZkNaN
pTM+gXzIH2xnk6kKh6L7mfIruk+Mr3iXOqzeMP9kyQbBJJcyV7CaHeCYbRleF9Oy
AsPUbTY6w7g2k5VneIEbro3UwrogE3+1BcE7yKMFCXp0rGXfuYRyvA4QbVzflcU2
/8/vA4ePy2hIj0ftySiPw5colZJr0i+vM0xV8xaHfFWwVd+A2rzmVaJZi+aYn06J
znJC6FVdayc3MZMQyzyF7uyeNGgpkxt6R1KFeYw77gMy5Ko9BfrMthjAZa834+dI
zIVXtZoXfnPsnF8o5MUql/ne+rTh27YwqNEvcDiL6iR7ynNIO1sUISubAbMdoLQM
`protect END_PROTECTED
