`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6fn1RLKfjlHQvWz3RCDO5CTZVGstlJsQUpkgUp3PAiM3fMWkYAyA2M2scwR9B6s
RNCYcEdV4fVjope07sY1Idca8P4j9TyClPUTtS7GKVhCH/7o0TLjg2NerQJnNr+9
6Ef4pgG+5fhbGPK8V28wDME5OmYezi+qHz6QE6zN85KyUZePKaP5/Tp53L2FRf0C
wDCRmDqj325BU0n8CBXgTL63Ymdo3IDY1pm3188g6V3Q4VOO6hazPcrTjx/6XHKH
jOfQIAjiTGDAXkzwsXGcY5FjDjICM0ClGDf/dRDaB8A2lMTyG+jCT0/pbkARqgLx
l/IcuKhfTLa+1WTYT3LOJp5HKpY7K5lBNT1hkH+J5Q7fRIT0mGliOfX2zy+HSCwW
vLM0F1TSjLORXjcmJ283YWiyHMmu5uqoqjLfWK2GTA6TRZRO6IzccQ+5XlkXPxtP
`protect END_PROTECTED
