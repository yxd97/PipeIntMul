`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bInmfCusLO0yXm6NbF3rwIIrldAzJc8tHO6tZVtkWP/c2PPcEb3CCS2G7NYD0C/g
n8yHHrajB7sK450NQvEBC5jxQy962aSOxivFuFZiKRlhXjLgfSfvy25cUPK0tKXs
P05UyRnyBuIwXvlwY5mmKaDG2Z2XHNyL+vSlRp3iyxV7LYAwFCzzAwzAQTHLk7k8
C5zl1KdURtxxXaAiID0o0bv1Fu2VErIz1sBASifLGPngr57CqZY0ySfB+mGayLrH
LIw0MRCXNHlBj7zruM2q5oHz9g9aXu1ofswbQ8+ukxBQTNehp3nYkvu1jLeNF9Pw
cQrCTqkeaZs+n3/nWOhqkw==
`protect END_PROTECTED
