`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSkaCBGNsjFmsSmiYPG0VSurPQ/XxJRUxI8/PLYJR7nvmh7GohOi/yL5nYmNvK1t
LQWS3S725D4NyZWMkBl2okUuwdpifiTgHsDXcf3VuHzshy13/gybpdfWDalR3GBg
NxsO+gFVep6wWbqHmgOsaATu+JrY9VArqGXTBJvTSxP0098jEGmuBDzC6u0aYls6
9oq1M9YySG22o0DcpeFlT+1l9VrTjCoyYWxfdOp0zqeTOzbWha4GkgmXX+zeqKWW
7zzr9wiRY/XL+w4hThA8DyLN3aY9jk3JhINp/3N9Zg3WOVh3G425d7/grLp81/Dt
4L/7jI6PYTQMU4KrCmETxClO7xCsFqaxlGwRWgAC7NbADwQd2MiT36cmu25UnmLh
lAEDuJL1o0ECFaD9SfXrZgvpCt2Y9GGcy2veDMf4wR/XKUm/hEiRCRVvPIXdMEMV
3XPsr8ajQETMeljR18Qd1VLrZbxz0HuPzfmF0scFgh+BKY4fMf0Bj6KYFd+YLuNB
zYPAUhDNgNAOiEtPu/pGfAR0r3KbsMIEn32AuE9OpswITaGTSuu5N/lXr+BUejqd
JhqaFTQ7vuj2IeRWdfhMclGt7rlhh2PMFwccFisnxmtuL/p0gScyxhSP+11QfcOJ
Njc6ztrPkE7aAlg4YiCG8FPnjIgXtZ/d+9V8LztEVF/1iwi2NT0Pb1CokyFcvpBN
prKI5zBU5sKFl5fETweQ23+OdKMH8OigB5Fcivxh39U=
`protect END_PROTECTED
