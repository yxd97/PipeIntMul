`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3omKcb0xkzSKUpxjVs4b0MzY+0c1Ly/rOlDfnl4PPHzMsHlPKYB34IUd4P2DTnb
mhxyac2T0xOoLgeupKb8VvblZCWvpE7T+pK50il0r4yJrpXDslFKaf3frgkeDxyt
uLL+LqfHhCeDK9MejGBX38k5VTtvpKdI0/qIp1LmCEM+UvIMay1w/z38QUpvMsGU
YBa+JPLYHbkdHS1JCkAVe2meYg5kQG3lky4X9OWaLUoyRQbeha9KxhkJihzGvlBP
skbYOOcjBR2oPiuYjXycq09fSqPJG0pyMv3/rrjazkUpicH560eleGcFlMvVm/m6
OFqfmsD7DpljziFQ+Fsi8q6p3RXJlmXe4CbG6S+o1GJ2PC6ZWWaudE1qD7BlSCg8
JFnN+N+ZqluRI8Djgjn8Xp68kPetICNhEocKKltdIvIye8hHRbSDBuQj1IahtBtB
`protect END_PROTECTED
