`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mQ/QFD0MBfSBePY/7FmKD+kdt82FfAkPONUUevW4E8DZkyCHQRGDl8V6uyzEJmd6
/jWFGFCig94lBs2fORFtgJ0EPrUSRuu3qKIp+hvqX2ZV0YbbKnaO5NBJLho9Q8y/
y/SfGPnpZ8w8vFloWBT69oiTnoNZ0Gw+WS8/KNI8TcuohaSNYLxt6nfKmePBsLEW
atEmmLERa/t2ZWFubgzOAZrxzI5ygTvc8aHDT/H+F5+wnyaUK4xSZ1mPz7c3UxAM
vcGYb5k2s/r+4sRbD5MbbtJT/JflZmpMU5HHf8h/YR1LUrnvYksRvyDe+5YkyIoS
1CXeUO93TznfyeshNMW4Et9G/QWQ4Lxgu0VTkGXfw7AVFIm6yh/Mb7naLZvfgGFn
32uqPEJbiboN2Gib6hPOSJSlAGfSwwkrV8Jd4QO7g4QL+5pJy8hgCX40+3QkuHwI
`protect END_PROTECTED
