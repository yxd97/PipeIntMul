`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFBocGsxeOPH/EHAZRFfElGl8opgZMGJTIRM3e32/24AJBztP1lf66sLj02rf5/W
zhZ/iIolGHjQxGtkhBNyig0cUcUArDW4/SQ5lHWZsVWceKvPhUfZ/qZmslfywSMG
+N+c3Smdz7NFxbJuX3cCx1os7FjgKlsAti1mMZA2xbUGNBBSnOpLtQyLZQG9hJqu
2ezOaY1L4NCoW9LNoHJ9wziRlHKkPMLZmd4rV/94y1aFFlp8Ls7Fff31oCLd8MEx
nwskHoDaRlmR+n1aO/hiWyofoDqbh7sTv8fcTIRDVsWTydNfolFtSjdQEQBG/XVS
fsVEuizlBGGMcpaod+6zwc0Se96zk524JMcxIKOznYzAtDrJyoT60vguVm7JOFmI
Wj7WO9AINHIy3YFaweLxbEn0iYhXdRAkelRK5j4wieFDuxU8fPKltpZM4zT/pSHN
pPyo0AblPrEHo8g4TOR5FqAGY68fUPkWU6liunmH7z2JjloeSQDcy0eyCPdpetDd
or8g/eLh7zaQDZqFSRYWcJw2c9LeRNs7DHYa7cMxDXqmwLnSw+bcbAX1c9M4YARH
z7uJbwXUwIrRAOMVaNhuhLf7qB0kj6UZaa4QdE3E9BPr39a4WA7Ss03rnHspE5rj
x1L4NEMLFwyCT1Oqiw/S52RTjhV5aZn6Z98D+LIRuTFMGyJPYZQYWOrGj5wpKDjS
0z251dt4XSiggRnEE4lKnONlsT7Sq/svRUdJmDUzDb5TCxj0Gy+w338qqQAjVbrS
vuapTNbR14gGiEByA8wsXlI1qsIx22vgZil/cFsdFlQ55ZM70v8o9s0JG0oIrJmW
IKQV6WxFH9/JH5loB6nlp6gBYMnllGTGzGh+5bLyU1P27AD9c5gngXDG4CFf4OsU
5QfdK5zkbiBG0EQv2cLq5yzQJpzQtneo7IGB7/pLQjRoOW7fPf5OesGSzvlAEqem
7Z97iRNFhJ91AywpwKo18tT/zQxj5/1YPTkr+gcB/5Z5uCuFhsLtT8uTFbYQJvxE
CYaPhV0bYcTqVGiWKlYhm9tfz3t0SfiTRAdTW8J0+dQwNSzunoWsvQGij8wokANI
GlSmt0JI6SEFn7n2Cbo6shtbiGoaaollTOP9Er2gT7nhDcRjGuksGsANmr+/A6El
cmn2F//WK+8zcjCZfiDHwVQiBhDriAc8CenvsBIpMe4iO9gKTUwmKzXz37mOz8bP
a4vMsslreK1aHQKc+0xdGEuBs5+efvkkqnGHCnBQuFnLrGpEvPQ8e1Jq2H7CVyAm
vTN2kIq70XsUU83tOXi4anTCxTj94B/mmY5ZKie0u1WD+/vldk9bSNc0u9/fMjbl
l0s1bd0Ea2ruoKWSF9OoMQMFsxoKSpdUNut767854RGSOU9OnJEBNmfZ0ierwhbX
s/8c4XsHbQZKj8xLxL5HXSXWnh5NCh5nHAUX9vDSrAxC8pK4JJhGQgh3457cBjgH
jx6Q+yQHuyF2DYFNIobbexcdNDzAj+dE9iofiMWYIv5peSbVty/6hDZ57jkzA5Ae
8fEl7CSwcPw1jW4EWyleN20/sIdCbAWlOO1FkKKq69yB/I2sJXsI+R9nH5rbJEPq
TpGgNTfIUeU+LlXrzHCRmTkCOkKxozYsCUXmbbOJevxF8dCyCChb40YqMH5NjHFZ
YMDPwPwGNqE6167gblY/ZQnl6PnVHPLDKFPsn8SSvYi3fTDvK1EvQmPrh7MiHYdi
U08AlJVBqX0F/EwWW17Pg6LgdX7eF0xPzREsrQ/RQEeAp/0nA+gyFhRY2VsSQq8H
bs9hWr1iNMIKsYeuABP5RzuzTmK3hJY+434BC14jt10fsA16vTxXS/tfjlE+uZ7W
eDnRK4ynaAxDzIsoCmnEr9TmvA2eT9pamswnVHKnNBVhcp1E0mKggIUsw60nUIon
bHq+IwI8WuyA63q8o4H9PfsJcBvqSZgdu7h+Wn4WBiK/h9i+RTB4kF9e3UUUSGH3
LRickzDVQBLszerxtPU0DCSsCQRouk5Q0lMR7DRWU8zUNIrQEhR/EwU1jb70N/Ly
Gkzu1cIrLVg0VC9uglLQuNUcph6sZhyHqalR0RfM4EJFbAKY9CcXZ6OETpb+XGj8
0kapupbOvIfj5gRt33QV4OvRaORBz+cH40aV1RUnOI3kEqpbzXX760L29+9VCt10
+zrY2AqRO2JbzIkrJpBBSCNj5n7wOAh4WfK1j9zxpjcy3dPoEgUcG35IQiFyyVti
INM9M13Oq7g8mSbr85VhJMG1ZiB3mXBGsRl5bYBu5Mqot+f/hC2X+cHWpmeZN2aA
IGf56b58Qx3DYcMJBEQQszjCEsgMAVxiMBrNEQU1GIicmV8vCpemYwHgqTz51uvW
WTmfdCSMLyTyMsAc5RR3clEzFClOBgynsUQY2/XMyo9R8s7YDVm7DfhJEOCE+Gri
9DIp5meGkiAnH6ggaSUzCE6vPxd/if4T3fDTFnTxv+8LLTFDubfwXxv3Dbs4olg1
qrgkLAUONNmqwiRdr5ED8SLjSoHFbqr88/NmY5emfzY=
`protect END_PROTECTED
