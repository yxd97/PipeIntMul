`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZReQrGn+srhOS7cPzqwlHlII84eagTuqxGHsMh/laG3hHTVVvuvVf3S/FzfQ1wb
lqVDRqH9ljAsKHualizRvp2s0yYNYaW4BhMMaR3JYbqWs1I8dYIrCwsutDp/saWE
wka1J4lhlTrn/e3K3yS4dtuyUgwILmXSLSVHjkio+74L7qIXcR32hpVkaAC4Mcom
it7k+sNCt3hWiJo3RRvJyEx9y9e5hFEdtVX+0+4q/Zd7zYZauUPGy63r3LGgq9ip
XjU7NVGwgPh6gu9d7r8lM+yvOEur9eK4xGMUBP5w1zjKQdhjQDL4ZP31iQbAdo11
QmbFBTvUJGq7I+LtFk2bvdDf5qoq3BAG5mNO54RDAn+FZq/atM6BOpdUdTwjKgCy
f47TH6siZiXkFn2T1eGlnrrZsPpTyFo8neAr1/aUXHFLwgTv3YOz1w8+KuzMqvWX
k5c+/OnIf5chlLrVFMSXizn5O+BHlx+K8AL4QdA+gdyDO9Mxyk+Mfg6wHO1FNf1P
o1jJMVVZwDBtwKNpd2vBYjAz0gpAEWguQkLln75Hq95bj8CY//HQBXycgRF3Dm7K
MtsiF4Ofxihu+eZnE57n7CuoV5bwuczOUHMsOMGrtNFhs0Q29foRj+WymCRmpZZT
pBtp/AdRhiuQ1YaOctlzaQxmQmCReoNhWfJniZV/zWw=
`protect END_PROTECTED
