`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQf2ECu5evnlBwfnwckvtN9JBvN0UdKejX+rjPLuZpFRWZUl25dzFye4eXdN1Z98
G44s1JFQlKqNKH0tPDTUdqmmUJ/SCPU09dpRzo8amev+Oj/LSAlvl4r5stg58sMM
yUfhJOeQxAtNJ4NAnn7/bTuWuS8FmeWy97/+SCEQWbA5eRkeJtJZ8FHc8J0T8df0
qy4KRqGnMlRD+70Psj/CuKLWMEedsENg1YA2QA3be+2JaURlvGj0XCw24Do0Ej2x
xbynpyePPBgnLBIDRWzWzaXTEN2VO4wQtkOSNws0ChUGuEx9IlbaXo8DwiA1CqMO
sIjTuHyTsLw8M/L86BAHncOBa+2Qzy4VMNiSxTYHYgPwUs0eMDDVUtq1VYzaHywk
hb/JtyqW1ippcZGsSsPBOoBaK+Ahxo+jPQbRM5n7GtBJ/M/jWhudLNTDQRfuDaGx
Nra63fXxVh1DidApHhjwhoasU1QQG3cdGFFKaQzLwZzZE2qY05iRYJwFUhDwy6+l
i9eBM4pFt0RPUCEexOA5o26YCvZ4sXblia3Od0i2J0arLsBsJhQblmnE0qDPC6Iq
/wgD3h6ZPApf2FvklVhKFMY6b8mJnL6zcrZg12ar+HA1xh/KoZFGTbW/kc4CZk80
wHfxWyMYHJWzjufMtKx7Rv4O63m0hivX/gFk9Uz/hWnqfVTOCjDF56qF8KUjF396
9vvTAjQ0tXqIW/1WC3LgvwfCqOVmQV+fmVwpKRe61TAuLxjLMW/qYqIhUS6SzMJV
U+eV/pt6SjhGsIC8syQxEEy1eC1rkeubBEr/Vbk/LvXJdmVLymy1xyRVXqL6PYsX
gz+bkooh2hy7qIOR/10h/fECnOHzlVVra8+7JQ+5//pjIySwiqDpBSupRElSjcLG
rtEnA67OyAZTd6Mdq7RPDEpVS9gQUvW3fhNS0xpRET15XkdhrskW0nnDjEqoQUMj
yP7H2+8iZExwJy+HC5CR5A4wMJCxYdinqBDxfElWUewiVdSxUgHunOQOjVU7v3kD
5E4QdL6nhlYwLZmQa0A3wA==
`protect END_PROTECTED
