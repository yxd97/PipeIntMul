`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JO9o22nupPwOPfAnwNO1Axh7ib7JbiIFVPc899Bllp8P/nnIm6zytZsUehExjlhQ
c3iiSoMaVPtpyfmUgCuS9EXSWTso4xib5TRYB15amYJj0kjC1hAL4gCD/5UrloOL
BoSL3+s1LaK8RQ4K0Zqic9qMO5OlxdAoHTIUClekLNh7933I+KLC/f0PlqRK58Dw
s2+RICuiqmzu/7/2xgLHj83HmiR+7esotQiMEruslNgxN/UiYYbns1/4JuEc/3bt
TxSDxiew0DD67VdihHNicxiMKy5TZsTfLrDJa/b5yzvVSvE/L3TFAn2yQ0y7f9QY
0lDjAfKWOONdYVns32TBbiPFPRMMwNhea8iguHDou3UAY5y0werpk88pmlmSvfuV
zy+yqBfvFMM4YohZ7JvJAQob3G3LuAJCHMjc6aybTAx5bPISlk34NYg9SKQIPYv2
ImeP+ybJmEoZYV6bj4852ZbrHMOtaXnr5sReUFNvQnrD6KUUG7g8JI3p6/lfdwOn
lm1TBJFBP1XH7fA0sIZgRF82HfE+Q11Nttp9SwAeOcjeHLmTxiFKxD0yQWRO9rHl
CvPxHvNctU2IxeTSrTv0tNkeu9fzLXfWpPX67crLDVt/8TTwnVQ31brZtnlxk5EK
7vLavZe/cLwWYj18Q3g8u/RlIYnvnJnObCDpWzCEXoo=
`protect END_PROTECTED
