`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RyNx0K4M8WOUYruDyqBcP7c4VOtaCMW1zgkMXo9tnXx+OaQ3oNOP58m0k8ZqQhu/
o4ydarNo6Cc6txDwUvvbUjshaD7OCPXsRZsuK5m4PeZBmEb3yg9vDyeq6dK2mGlL
+1pzkp6vcouhRDpaJDbYGu2rEj3q2GDfoQnSMMqXU/fbhCYHIZlGFoA6Z6G9nC67
kosWjh5udQOg2Rq17gY5QvBNpBT65Ru5r7tYM7oIfdYp30eE0IUTMBtr4EuILuOG
S81F31zXH6OxdOsxMQ0vmgHPwX3Ag/no+vEJ21tVHvUlsGR3IdaSW16rZ2qogWDq
bFzUshLVcwNZuPhDBbsByeSfs3ri31fw/t+eElvlPC1tLndbEpgKoZXRdpahvszw
VGbcBHMGzDDwbFN4UlNdcRUDbMGzmEKyDY0urY8a/PaPoen691WOM2uxBvydCa9P
Wjx+5M13iXIEiE19NRu0Rxw5KkBP8grarr8sUuoGUGK6iagFeygJayBzIsoU/q0t
EKSqXMTrX9bHH7ZO5+I0z/KF7/fZNdqDFXpSZiXU5Yb8u30wvBekUjcEWYmPFsrv
O8/SumRx5YaBtWUGLy67KF5grCv1SRrzkXe9H/BHlEdU11Q/Z5WGh7iWCKx12wQf
YjSurkHyv5KXziSGDELJbntYK7wf45X3X/4vOxzz4kUaX5ImpQm9GLGptjXpPtMW
aar+rbPwpNHqyMrJgkIayw==
`protect END_PROTECTED
