`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwTnDYxilcd2GDPHrdLG9PPlE+ih5cT2eWjjebSGptQQw7B2wa3cNaVSioI26drM
fh5cWwGmDU72QAsE69UY2tphzfsClkGqOoqCZaabCViwQ23BVvrLgKRvH3adE5zh
TNMfzqXX08S3Qed91KGpcgHisZPmd2ZC8jdvUq4/1siQfC6UHcbBtisF6ovCLKDH
Zue3avqRyJcEJR0GIVtM4nLBzKxu/9hOCT+U6KEwXrGmFzeLEahfM/DPhul6en2t
AsTZXY+kHcK6Hwc8divgWDzhm7Tp6zubSTj6xG/IZde0KtR30KGnZtCtcS4p+i8W
SsqEVzd1/+ShK4s0YfVf130/HY68ErxRxxo6PbPcaoF0w2wyNYEmWdVKx35YZb0o
tUeWSMACmiaHcLGxmuZv1x+BWc1dq9yyJw4H6Aon6XiMWLkMEg1QYhChNzBP31Zo
5locWbM1idQ6r4GUAUda9AfyPW0fVyhMckK0YmzwLyJ+B7BJrFnkQfVoc1p/Q1bB
HwIsVCPlWhPj0WARU8cirH9McHr+UYaWrhB/AbyJQXgcb+c3Yos5+b5sl/0rj+wI
MHLS9xshQgD62QdThMPU7G1rCTJdrogIG9OPEjj+poqQ66Rm9voFXQkZHbFyk1Fo
uL1UCIEU3tmLGvYElSiov/vYTYHv6C8NcNY5rPUD9WGONAlwiJmjYZ8dqcdQQPuU
`protect END_PROTECTED
