`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kOrePM4SUP6YGT5Njyx5xI+bO/cyBRxmHrawrQg4RDoED/H3IjY0YjsPh+IA98s5
tUjGmhGEvDCCM1X1QoP95mcuhRFlwxnxF/gRiZSFp2L8PbSwoDctm17PBpE+/1bL
P46sn+u92eUKACHnetvFI5N2qFDkpCHJBOFzOgsm8tqpMsuZYj1wQJbKlIXZVaid
uTQI6HuBwG5/pMYaitFJoDYaV6lDZ2itqBAfVuqk/sxbnHhibO4w0XPtiuDBVs2L
ueQmTbRXlbyeNVVwg8CJcQnxRxi+P2M4bTvaUwdJwOlEUEwtwv3q4kfPfstzSo+f
0UJT1Brw8QF1htnYIgkMl1G3N3D+mRT7tJpc1w4y/0CmobWDs/imAZyOhJR4qN4x
T0DjlTm1GylbrpoWvsfyMYTjeh8+FVBZANJvkbdfLh/nB6AeTkoS1rXTJ2dXaVc/
p8YzkPxclhnSpSBLVpfukwEzMY3wI+7bMSmDCE7lG8NEQDIDBXyVL1KyIREc5BLY
2sZaXrdDEkQxEP0o4ML/GkmraQd9TV5ucgCwJYTkZW4qHxrRoFcCgQ+vIn+nd84g
FXIkM5AnO4E69cMySccSxLmC6U16oYWH/ZL3krZqvuKJSsvdWNMlWJoy6jTbkACD
PBldHNFcibJRZfXIz4qlIKPZcMWQpIiqXjAT6Nzrn1PGf+5P7s/lrpJPp65DtoPo
jg1/ffc5ur+/yL0nAvWgGSCc67N/xsYI4GvD4Ujfa3jaTmu38twe+hs5gicZCF8c
wpHzE6mwMvhA+J/EYkU0ONUB8GVsr7WjOCyTnUl+5uZmQ1U9mACYc6vkC5R6bpLe
Ebyrb+C4ljmGwSRJcWAbW29T5Eg0taxQumQqQ54GQJtvfsCphaPZJ7vpGk8BDoYL
6siBYlw+gEopFO80fDITSKYXljRs5jyIxXKmQbl7K7dLLCHd1ae7nKS7Do6xLBAW
LwpYsbmeeFgCj0rorb/XI/ZpI+1ULOyEU5n67W9CIpsIcwg/hyRvzkUExNO/+aw8
PuwBWvWzRDxmg1CSTB3GcttLzIDBgaNiqfUCg309UwljERfEAGo33hgBYdbqPGfp
pyS2x0V9pmIJg/v8HYeH7VLknV74Up+kZX8nkwMvPN2q7qvZs3GpR8Fnj2Nev4vH
q7NucJs7peiydH8PdaWhfjXEP3fPv6vJbdmcUa79IQVVMYQOOhnyGhoFSok0qOvh
J74KuO9E76iKXMr/zqIYi6mEgNDh+oUxwAdR5/JsV4x8vEIyCmCKK9JR8kGWrHNy
xjbdnr3KIElqQYKfLw6yk510nuaE4jVKFoViqlkjgGPv1K/+OFQ38b6B3DlpS8ww
ZEBMFIckrrG0/LqVPLUayTRpkILLOeiVvlpTBWX3vEMei2dgwFxsQFChzUEojDM7
+7ZpC7GBaiHgu278ypazkP3w4wbyBpyNfGjHhSKY+bDPlx5n3YSEuSEMqt/dy5NP
q3IX+DL3mXOmTf5f5dap+5NwuRgl7aBge5YJVwOusfikjanKauG0fLT6dqy/5J2t
gUZvKnlaORknCyzX6GgJYa32qXncWD32fOxgHTTZn+LlfwLE9J5udk4GixFnGcHK
2lFQqQzIEC+/ZiNk7Who2w9q95xLeKukJGAeywfRtcE2/SoZQbNEI9R1/q7nycbS
iodlBxSDmsnoxAMxxjPamyMmf7F/uc4jekBnPlSp8fTMXHJC8Ly/uNKFgRwHtsBe
qTO0IxbJF4nfytsPkJcG3a5Vx8OHccGP4YJwGunYhh6OV1U151wJJovw303dmWjm
`protect END_PROTECTED
