`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zazc1TnrM7By7KYwnhMgwWtHlWdCREg5QIg4Y17ZRGJcf7LaNOMMLcHsDbW4/o9k
YQlzPoc/2H+WhcGEHxFImgooYISVxhpS+UbAihqiOwqt/b6fkcW8au403Cj5lrGp
KIU6BBo8NXYMrEvBVkr6sVUMv0reMVCCdo2NdOI1D3lkEX0VKAgOa7d8sjMnK3u4
oEHcIoki876TUJFGsfGfoV3sGN7PdRnFbScjCLxNoIqMKS93Exgkd85CbWEik5+J
1XFZc4zc0ZFT5aFdqCKzOJ8WOZ9lEwA8XkmsiZaiDFCJ4wyGwp5zmaPJVXP1uskG
/YJzzMLWa5sp4JZrdqtJMhbaOCg8Dn2Vq8+ag6uVOMxg2B3QLEYI8hgh3ygerADj
Zzo1Ndwf7a8B+t00yKdFkWodDp/VmKBlIXoS++PzDkskvJJ4wgyRd0pjsiG3qZrw
TSLbDsPEhSx6a20WcG4qDI7IX2aYzgmImIB6ZjMoJNSzbVTl6ZOzm4geQpLKs7/s
NYr39avaW/5AYyhTkobGAkkxbJv41YLEWSyNi1VQbGP3uJklbNBwlHiV7lCbBVfB
hWeAfQbZKnxN6aIW6Ah3ryhQjoVdYbBVcD+JvyOeBBnsqSNfXZSyJ9TuF3YDoTqH
iGtO+Q0cjgSxRIiFQzQcj77PG999e3NzC9a0zGWCRFPmZPS9hIMlI4GJVP4FqcfE
f2MH7ux/3+0OpNXUMtDa5Hh7itB7ffDSdloCSJCgoXveHVd1EXF46jCGJ2f66MQL
XzHNeqEHK/zdFN83bw2rZEjTdVc1cxNJF3QgpO927vRdghbtv8NesgS4CqmWsfB4
dVfycivbZNNc4pXBpSN+ljuRY/K9SJU6WiDG49VxJfgUBf2L+clIgyLfRCrlIUUl
QwMM5GfiY8ocvU9ezV6NPELmwFSzlXQAjN3RmLpO5mq/hIgBeMV3BVc8hW2OWZRH
wUgAS36loU7r7qyFm6e8W1v/oiCyUUr4133L0SgKWYubz1sulKBu33vE7C9GnQl6
QkPLU2oZpvPlRibhHj3pm9a3P3EUg89W6S0vQANhi+KCYThQcgvv4gIIbFPL2vFQ
TOxEpvjWRCeBds8BJDmAseK8jQCaFC4gKw05OhlBMuKNLntwpHU8ken+bSojnMgq
EfGy3Ef7rVs3QKkHeoFK2J0EadHTw0knmtVIt8vJd6xStUNij64//a4nkXY4fmWZ
71ltdy/y/7l2nsMPEnp+oPTPrXoCxBvRt7EnkQlOC0myOx4RQZuMf2HrBe04ceZq
QYQrq6hrosJakBdh9B3Dikukt+6b9B4uLzXgJ1XKpeHz6eB+PMaNjTJ9QpSau00B
FLclggSucXcVls54/3UWB+MLPCoY3VFnMpPHVDjIbKnQCysgpNS0WKMTu0GkzI7M
oBsHyN+uS5FaW4DxbhLB77MB0+Wj/i6IlQci1ysPislzpDnNFGypuOmnTB98rLPw
OMuAPz3g5sHd5Ugk6sKG+7zNNsVgnnwXtRHosbHC9ejbDANxkuz2X69ir2DqHvC8
UtnRzNlpqMicJyhd9Vhwj2mECQLi6ZQkxLQEe7LPK+Z0Lq/vNb7VHfo4xTIduKd9
DVL8J7lzkQ5ZXemzg0cPoZvo/vdRS15vcCyGp1ETSlRJBx4rwBeb8s1i9/gXmo4U
ct6QxlKQhFC7oUAwg8zwIrx12fo7oIqXuvTlEEKaPSIFjdsEYk1bE0PJckeQx5Z+
L7VByoM6V/QgnUVcpm+E0h/EU36r/P8A6j0qWRTScO/jQhynBEwjQ3gZJPDD8pQ6
+GnptX+iNMH6r80qpdsPi1oqrn8/4+cAirJCU7JWOXb6qvt6aM/cUxVhCbig52qd
i9fGN01AVoYPFK5+CJSE0z6V3T0aZ866YCG3YzXF6oxT3tO/5MMWXG61/JsfW3wL
8AaoPD4YxDHspuODk+Mzjn/j/x291xj69v9duQv8FCnATY/6oLu6dIUj12SwRVIO
C64U3p74d1A9PNFk8wj3mEpZeJmohViIO26n1JerEpp+dXG3ehaV4fY17qruQYDO
9iAqcac1mBLUtU10bH3HhOvgMDe0WNx9ecs+shmj5xZM0PMNT0mHG5KP+F5QqtmC
CIcKS/DotioJOu4JuL+ZB/VUE1S2ij7WsBwzvtaWXfJDxmJsdSwnANYERfmvyQFP
xeho+DJDeWBSyXl86VbSklF2nxY3GI9V7IYSKtpMp7VF77DIrBo09htjdf+3rhg4
fDTsdbejvJAzYrY03uGusuJ9wF+X0lV9LZORNhkaIrf7qIzofHJMr6K3VwAyIvnV
KqnFUC8sPxMpwiDRrqdOVSsa3jr0cIh7Zt6LqzZk5Atp8cg+19miLopbdssWMTC2
qcHB71PZ6yaV2aXlv07H7FmRAKX7r6Nb7mO4CKEUgwmiKqRtaBZo0T/vwZUSYKej
qrS+bN7hQ6GKWAK0uJpUNS3GLwEPT9u70XPUnmM7fNJg1ePN0LVZ2ZReRwdmQ8v8
YBdUn9MU0CdXoptfwlNFeIyuZXkZuTgzTCJeSC5FMjQ855/PU5YdKBr054X2slxA
qI4wYRDQ3Ep3kURG0wY0PdSl7MV6d0xkQNn21bRYTFsT5FvYG5elEifLTP1xHLiC
gPhCQG4lXz6feDTmTqLbL+v8XLWjYyeXgG+mylW9Wn06fOY27jxJ/okBrXlCrUHG
Sh1wiuxa5xvB73T4SRuEJvf+4RlRIAt4TlHwVbPZZLPRR/lfdG3V5b3LL6ZU47AQ
TgDcJ9TDBQsuUEvhlEfECxvLi/K5Gsq0RkPH4wT5/ZpUktWRl16g/IcVIULotRWf
6smnqFEeXZoiqwM8mseYrR3mIuEapucegywLhJsnJiDdPmAoW88GqVa3up/7BIrg
CLbSxKLNBDL9tlDoBYRizyAgpm+XXXsyjJnrp0CXjRgcxSZN5iJtLFobtMuhCatM
5/N3X7Ee/pQzEeoht9fScXqlC/Wj0qBvtRZ8dJzyT6NE7CUy8DeVkfIEx7VpmFdK
29uzyKO9vbu9J4huVfIv+18aschloVHkkgSZg/2XWTawKSrZ6CJOcE2eolakMK48
pY9xP3D+NoW/45Sv/m6sVaCTi4gXjkBI6WGUOuyzjjz0IPtpvyj/M9e3pmHQtyAK
ceG6KqD800Tiy3t8Ai2CBsFr/DoYDtAcCQhmELR/7FBsoDZqnrAKG0mPAzUXg2qu
7t3WbkjzKHe14gAz/CNvBT323stl/GlJOdEbYYNo3+D8+G2A5WNSnwd4qFzfVvnI
Gr7tyrNX2sUc7w6Z0YXEdc0CbdzGJwlQd1fCFCBOKvidntXBwmwyi1PhrqnAHQXA
FqXQlO4mP+tv4BVTrB4McIM0JAXcMMCLd40Gy/sEyziYpKFSpOLhw2g6epbKOvEp
2Zs2s9Tp1nY/GYdcZBCPsRi9T/vMM5LRNOVohCoq1rGifsxWQiVMH8jU/DM0lLeN
ZGJv8A9J1xROlg2zT8BpG+fdXN8J5huDACVHWfGc8atlkHf/Sp7inpt4Ir+5RGUS
/oPNLOoFApqwY/tgsWghwQItlPrRmUOm6dLGyerlRi+BAnv7QZLlUyxXKADqf49W
XvJiXdvZINRgab2WMX2ssrfwrV5QAmT8Lxs9FI6abgnA3t0rpYhsWGnFJuXoN/6T
uUvDf1QIJMpddjNd/plXBnbJaFqg8Xq2WeC0gP65SDR2KstWEeXIwvbmP32k/yYC
dig8GbwPBkPK8KkgvfPSTMFJR6aTsKOxvHvCQ+S+zY2EC04jLCVUgaY1ThZDuyH+
UXfiBvbmd3lOP3zqhgrcRQutueyLA4FEzQH41uZ9qhUXXQFF532oln+zaXdlwOJc
bRoMi/carcn8ut6tPklpySAt89nVN2BMOSmZCxIAuwE/hWrR7ZIjUCJite4gZ7wv
ACJ0Mlb2CgSjDdOVntdgTZOwzMLHNoNnDm6pD3aePDV46MBPtz0AUxYlvkoNqBgF
LOwjqsH5gIA81NRNbYSS+rxB/6YIEwQ2kAuxhbQEIZT3mv7lGY1q7ObjmwW16Sm6
WbJMBMRVvO05XQx+PcKwQY3/s0lDoY/ualaqsQX5v8GKuk8vNBJMatqDfZaSrWOX
kJXjypuQPPXKJZYJa1/ZhxPXdHgelQZhICBvuTILDfk8qaPTYwkDpbt3fQT2VdHY
DpLfsMmI6/xZiYA0BC3J9grCwU/tNfyt9aBhfEM19D7b+1J5sqQGf6d3Pjvsawl0
LwkmkN4stW+KFf+LFjDs1SYIyt6TP17pRNxi/GEnUih4tVQMWj7L0X59pdXQJVbi
sU3idVTNAAz5zMFqf6gfCYoXMkVo4w/N1qbc6zxrc5v+3+lJBVelFm/B913VW3aj
9Db4WGdfJWCLeBhpW1VdenNxboxW2lzFB000rNxEAfCCP2BAy470VoK7WOS9oHdz
jTBkOBKBfPdQwWe/YMrjMDOyG8K2wbH1VpQozkq9pS9AMZcF/YcwZBcV+6InUYcV
aFwwV6OkMM/e1MjWrc7ljKxM4jGdoHzSD0Ed7OQyGKlF7gb1GqhLxIYLVX660r0O
fSiPLy30V69nu7lqnFpxfMgzRxmpjerAnryBuK82Xmtxc9aSzVkiTbCYXb39GnTB
2D9WoKM+RjBD3OLHOq17K8+WiC9N4nxZbsSq4KQyVZ+7hiqOKrDrCaCwJ/2WXK2X
+/D1lYilWA/tk3Neen65KTDgwq7hSEmq+YQ7UHCwljiwwikuB2zVKdSvlOLxtE1b
Cnpyu10aQZnZdSzHckVINATQ6If/mOtSC8e0V2ZTqzwSMhbviohEu0aX3eo+S3lo
VbxhWCNw+okSRHKGEBv5p+63F4hzoxC/03Y1EY2kGLDiOOavaxbhExH2PmzQjQzn
DjAL8nW0AOsU0puH1290LArWbG9V1m1LBqDB0joxxP7/U/Kpm+LxhaafXnlW5H8T
axi5csYsKyr6YqSD1rK0YV9PMiGinVZp/gneYXggv5FEKBGTbAhfdq1y3mewHDaY
JskpqnTqK98yj4JPbZzKikUQ+wcx04L3+s12HnRaQvi8HzWGLgPdOjUW6lynoECh
KRAs+S1QAIY9grT62ezyhcT0W0kKrfwFOcSBBQBjPpM3fn++ACsYodApGllWFOqi
f071xXPi3nqDgs08j6p7LjmnPfc0hL8xxaWSs7KqLjEFnFhxaIQIKiokKeD0dWtL
2tqkx2oD2XXeN2BfrIcnLR/MfLfRfBDduD0ZfuhJR/VX9x1qByyvkz/9jlhIPJXS
kPrglBQbasf3LhEVEHP/UDqqMXbTgRvJvfrMMzLLmQB4d3Vi0eMeJFfdZgwZG2+0
qwZKD7Sf6TQjNFuVHaCFl4TrQ7hXb4wnDwpRHtkQ32j1SzR31p/Kf53dkeOGXhxD
TMzH92L94yVYbevwRDTuA5r8zzXPt+iDA8cfcWb5PRYDqQjgKF6/0eY49SkVvpha
p3I9ANM5VP9EG7V4X/fm2NJRibvh2D4xmsx7UXoTGpIVzUgprBgyC1u2MVeNOYIC
s11jU5RLWLYnvRT3gvLLVb71rzwOnDaNpEsUl78m/MNgpZ/flo8Jwvqekn8VFTJL
WMdql5GbyH7ILeOpSxMu/tP/nMdxiEpVwx9jxXnDQ34Jx83OUNc87C4wgICNpFdG
vI0ezViWbTnIWkQkak9Po5jOnIAQWyE83Pd/LrfCVc0xV8QKEqw2sK1GXisHWXPR
dvVLournfTDpJVHmEMAHh0HaDOemKVCC75q24zEHADG4MeXLkIMla6AdBVd08gzZ
JC4gUSUMTrdgSFPQABUMNOctd0Oot0Xty8T+ekFuBjzQX8nh4/l4npAI0GyJPeLD
57AmaqaLN3Wq6hN92mWxGWwsJ9+9TwcWHsT9WjaB9/o30V30OaXWlTEobwgNGzgm
t/znJyseRR3rieQl2SKjTqEahUD1Sf1vYtGx0d+Ovh0TMOKcyjy2odXdcRH/oDL9
n9J857CO02Ev/wLDAr9K+awqi+INOvLl/2vhiBWUS14TNWYG8LlqlSZVgYCN9YvA
ina1Q9iiIztjP/ezv39DS+VITT/8Z9nnqfJI7X0LYY88d/PZ2X3Ku25v9+9QEc+Q
fk/pMVOdDjihtub/fl+7ZppOq2B/D6W4Hj8ngAX6w8U+CCopg28VcL8z/NtCYu4w
yy9E3BGR0i+4YH02n5eFNZGjG+ByquLUsSWfvnu9S5CU5B1U7f71XBy9N2blwcn7
K+/X+hw+burn9dLk0hH2O4/ykBDg2brQivSMU+IfpQiP+5SY4ciElPy7JF/IdulO
umUgGgVcd5EVCAy6HMCLBTyrY+/+hCOjzRmdUE1i5tx0x4YmCWOdqs12cxZ5N1S+
vgHl9YHwFspeQhMPqE1NQZX4XILTEwhsoDzB6e9pTora6s0tSvtvCHpKNZ1HvFQj
sphSHdfh3kij1dwxCve4nS5JztsRN3GBVKAiMMAZz+ZCrCbkS/7B+cgcfhtC7gxu
gsz5oE8ISj42IHgh1jfI8IZ4bjzWU82BMNReKalKdGRc+yilXH7TD775MztzrkEE
ktrskRRtjJWPZdXf1syot7nFghJHKYW1mPZNk9HE8nBCAIpTFUmMK8t+cks37un6
+Qx4OgF3fwG3zk7eTku7jBwReIdrEvFxhAOeRGoktq3Eel0PpKTMkg6YjR4jeWP0
rSmorU75NlAxSa3oSHM0HUwE7NNBJT4eeSLOkG5M3CaTbP8j+n98yGhyGnDu9TTR
NpajiTmnSykaK7kCBCHHCV34zyqQVs32RoecQdiRJP62pdMPf/+YlWZNFM3PA/dO
VHdHHlFP9EPdDoHAXXv/2/rS2Xr7LQHGc8egjqxT1e50yXrcgTedHi5lDNYrT/m8
4hrg4hVfiKAP22jn4afElFkLnNCBFU6ZMD9z2OwX1tYjCY18Yg03xWa9TL00dvM3
BUSanQipbHIE+/tqj08Z4B6phVb7cs7tCtJeBQ+NOcAwIs2Rgq8DjIxnBGHqlzC0
W4TYKXwmp8EPVYPNgvu8hVnWD940l6nJ9+1eKjlxZWKQhRjFfPAfC4ERK3mtKono
f+KhluHXVDxdX1CIaI/qaeaBpxXwP2IJh41RgHWLkJzQoZVEakF0pL6XIzxa5im+
kzzD64gsEh+zxKl9JJt6WTwPpNsj022AhlpjdJNy+4Sjy06KbrNnYJBf5ftI0Vs6
RA5LugvC+E4rEt2azZVdrL2KBSpWpd70CMLfhbABVG7YGVWRESIbmHFVli3kVsPf
hDCrRs7Uig3IUQPVGq5JfZ3XYMpz1aJJ3ayLiLC994pmY+CUyMCL27uvJLYUOTo4
ogXh8D2ayZI/oKnU903rjss3g7GZ+QMWGnXICx4XOBpSb1rix+MiQ4ARQMlDsQmP
S78awp5AJSjkfE+8SU9PgpdRA1hE195JbfpMAW6p+NCaPi8UIjpLBPRXLz/+Xd60
5VmWW2oat2e49ExbAhxJbJy0Myu3gpKsQUCCTw5RUmhs5rPdsKY+MWH3yDbb+/J+
w5Dlk2XdLAtnPeL0XzzPLEm8OsRNQ/r5aXKFOEL/VNA1W6ZW0+SmeZCBn+DhpWvD
5l0aTQqcfs4fO7XIyZTaffX2ZBsC9ZEyEq4n5W6l3iApkiLTjM43iSOrNeZ32jv1
jl38olzl+dCt/2bWD9Y+SPpAE3s0xYnVQycuGp4EX863HbZd+uJgnG82t73Q7sYn
THGhauUAPnJC+q98YDG1vXubY9eMLM9RllEsIeindSqK2FWeo4QKnUfsCleFlmPd
ADzyuX6rhzWEuaBgsuLVFstYF+2pUWgKzeYgNYlzJl8cYnHvuxCLO6dCbvM3BUIm
McsCB4+savIlmtXsCqy18yvBILBHSW6Sec5iFakRE83MwczCU0CJ7JHFv79WrqL7
KTTdtN7eO+9bUzms7Mj2C5u/qvKED0hoJRTtLU1e+w5iJuIInrydpVjB/UI9tYVI
cSzjq+N7hqeWddi4H0ZzE8v5f+DB7816NwXE5VMtt+KQ/XnZVYiG6hW1nB1zGi8I
NF6dEkwmjGuosdrjURQQ7AU7a68hB6lUn7swTZ0xfLsnGI70jJni4K32Vl2PIeFT
z2bsw6hbiL887KUTTgwnbPpBIUz5XA4H3aVxbVaQu7RnXQRnZhbNcHrGxA1+iQBq
638ZkX7G2YPrgkOJHTrCN47lMRBP8eOKU2kkJ/nI6qhnzn/bvtGZGKAkXqXJdKj5
yMtCpUMCYGhMBKPpkHGjmYREIv4I5TrR+PhOztjKtQvJcVVVwUILFFFrmScgJmO4
mfi8LCx56XSBjV00iMBIJDkdHzcDc9ou6VTQ7Txl1ok6BnZwYD2GhMlKdho3Iqnk
4Cl52tW3WuqCxEmBQqEDIvJsuS5yR1YJ56loYijlL/SrgVA4Vvtq0eSluXPY3vRt
v69nyr6S5eose3QM+UZRfUIRSX0V5Ec4FmzmpbyouCMHXdqGX/3GNSNzf8Ydn4/3
DLW3cT9SylNnsTvNt+afL+YDyEcS5AsChUqisyUOdqhjj/ZtpnwPy4HEmZ8Q+yGK
Eb9558KzJW0MexNG1R8SYcV4wKoSA0eZPUz5D2m5JPdf3mbfmIPBKt2zDDs1yhHZ
ijq4+bptLDrEyt57giaQroKxBq6Q18afFKyZ/2McrYzFPC9wRlP23O4Ue9rI1drh
xs1hubGLq4AqYxR5OqYvJbXovgVyZ3Az2p1P1Xht63lmrdFGwKUvBT0qbqbkBOGm
UEJpHCVwmVtEvKqKOl42c+STFP2ygHtIY5CyA5Fi0PdtPgECwBzffTP1ieqX02R8
WjBVLZk8ccZ1yAe3B+UNKt4hO4gT68EeZstH58Iq/znhpKAp+ffyJiUUesQMe2Oy
NKCxH0fUsJT4SWoJRQZzJ3+dE94c8nlbcOtTq/lGPjvf+l/UHL9zHilypbw4vsGB
RBpKgKpo5/VCGHLL5ke5gzSA16EA2Oc3m3t/MaFrNmA28ARNqzSmBPFqz85qgtBt
RnjQ3dwrqovLHsCCEtg6l1vfb6bgwj9ag0ZBUnT17reAX5CBEi9XN5UkhpohnT3L
bMMDnlnEOiDrdiUI+pXjK6iV9oqkBpruewq3yevuDCM7HtYAIk/lk2HPtLdHnPbj
Jc1CyIC0EUBmLuE0gOXgBkm8828k7KhSBwfsB+ocTx9uK5YZiWhyiRyWh+3TMUKt
AyA7v3tPkKCkrpMKetInsXiUcibz8v9nNn8rwXI71kiNckF7WGorI9qvM7TudLl5
JQg/PasD3scOy2pKrjXt4EDARq7ydZBc2Rx99jcoRNRAizeq/RiO/c+7mPgVMWhO
JQWhPOjFKmsdShhr5KtOWjx2c17s5I5bqkFPVYuErEDrq7gkUtoDd8eFoRTntffj
H3yvIidGOqTAR4rltKvQ5aoRhK4T8sEbsXSsVrqXpfaa3ehvtCrGjj7qdgS0CbDZ
bFx+ZFNTP+5v9X+7L09eXofAEFrT1ANdeQ9EKgJLULbyulwNgxQMySrdYv0oQ1GG
omeWGHZU66AAEq+D0jbaUjBuCpnmP4yhY+kVaF7aT3MeFbTR/nS2EIRmN6qwJqUx
Rp8N2a78Yxi9PiET1QY2ylNjRPuVb7Ln6W+FJSRysjkytEkXsnlqTV1+3wpq7Jz0
4lNZJuCf4pshxnnHIlWa4NZLzagzCtaHIo4XquWzo1MGU/smJ383EtiAr+6Zd+bs
im3D4BHSYTvFrGvBstuvrnmeqDfCe6f9kgSlEcTsCtTzBo3zNVFEutRxj8sIfnh/
2OCSS5foVbwDhf/YAKUSMFi1ygcAlUbSRfoq/uNagmaZ3jW5LaEsDrVHHT0pmOjr
EUBqQv8NoKvsY/EPK4C+u13Mk9utTM89NYCNf2236ZdlI7J7ZyRkTm/oamVd8B3G
PkCQ9D/BpDxvarhhaSbKNU2usEKANBFq36gRwGEyTw+ET/2ABcfq47LCJhBr8taQ
fw70fdHoRMdfL7DcoPlL+dyVjOU+Yssc3eX9Bvmn/LlIbXDp1tt2LIanEIXvlQem
HUmzJTB5VWcia6uiq6n6yDNR2oaLYvQaDjThfua+wZmsoEpNotEkNMAMLhgM0Cat
VCs5PB0yGsxw8rIk0QUd5OAeGlxVYcW70npC/YubidmVgpNvYsi1dx+SqUYGHSUk
LPpGLjs4BupHgam0xuMWyZHWq26zafwePMvpIRh6dK6zGUpj0zG9AIGtK4eZJ8kw
VYWbRVcXPwKV+s4zC5PHa9Gi/FyRR/XQToBgaCJcskZ25AxzgsW9AelJXNjzBq6g
6a3Gel/G10idO/hsXc0d6pk0kIvvq6r1Z82/H75IpDm0iovzYD0ko9iVjI3a+CpU
In6OSgXW3s9OQcwZj0iuHAfR+czHroxJOGqvJ/GKc+1dZwRxlQcae//TWtn27/UT
wQ5/9fVAXVaySiKswNNPW0FYA3b3RplMqCBZS+5UkRlO07sEGMC/J/Nr4S80AKTL
MGAUcYIBwOyQ/LtL9GyMWbkhSMGl8iDj/N/PiQoPxyNkEU/bCOXTX1DoeW9IJmJB
QC9ps+X8zZmesFEktkyk+DTL0/auwAR50Hjs2n96SFK36QV3h5/xwueJB6IIKhWq
aMO07tv+XYJWk0LP+RLvWnpHIkEyzJ7lNEtV2TICI7wjGuWFo1x4m6Rntp3u6f0v
BLZoPw7vR4/zFVltgY0zW+sbskASDGyfDIEClvexIYUIkWVqtdL79O5O3eNYih7l
w8bjl9MyHmYE8j3blaDXxQ7KcOXvoeMVVb10UGczK2JjGylShYZTLc1g2RU8ihzE
0kPEbMoOveFKy5Ofv0S+/bLEtsXc7DfxksJ6TDeyPyLmfC9ZKPUeIis5kPCQx8lo
pDuXCwSyP2/6oe2khnT5ChwGCHcCMVunyY5Gq2zsjwgWg9L8JYA3HqdNNih7/GPT
kSRoN22tO73cRiIgGqMMp4SWMuOnVQEvOKp59VF5GqlSuOC/KOK79BkOk5T6NCEX
`protect END_PROTECTED
