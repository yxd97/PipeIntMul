`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1886CEeMTJua9+I7+4siZaI/slI8IBKyHYhgAnRQAZ/pfFAKDRXWxEpyiCghGbc+
smmpEv30gkPLBL3OD9RhYu5KBKdb68LNWW99C2afBYIYLhMO587hbEEtmaqvmeRl
y8M0T9uDgr694BlwE0ARCcnzo0g29b8YG2CRVNkjv+JGGifepgw0jHDO3kFF+UGO
pQd9iUNvTs8dDv1IwHM4543Q1o72QWbpOY6wOO9IqBXj/7LMvlX3JB+riAwJqpwL
Yu1OGRm4uF2SZ89Kj/ZnHpU0PUAlh0GRqNQHHWajLhF1/wdCThZ8ak7e2k5lwLwC
YB7yBx/Zv3vP6kC20q0SeopAPH6cNPLAfpwufP3VbWpLYJPuAyFQsqq3GzXunxuG
2rgYnbYL2bymm99Ov1g0hBxp3ttT/AV+1f8v/nKYCDO/XqsZ10BAt77X0LE/2bPc
h9SUHK/ckrlkwIrcp5z1XBD8NBqYg1yrdSzJk/Xr1Uw=
`protect END_PROTECTED
