`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCv2PzPqU/edt1gf7XA2K1z5MVAbg/a8utCUd8GbOtEPv16iULRPJONzSdqc65YS
zfEs0MlbSAzNtlbfK4SxF1coGdMyV0p0vf4Vl4VdQ0KObK9O8d+5Bd7NXQLK1QWa
fk16vMtX4ajMIuEfZXYuPnQTDap/B4uXNF5Ls7V39oQHupWpsehUuRXmbpjeMgnh
a4mA1H4JbFNvMqxJi6aD6FxKlfQeBPTB1Pp5DkwF+edzU00W80AFjExe7HMMCJ8x
JlPYdogmsilvl3NsinHilEoh+fXjUac2zsZwVLplb459abhH1yXY8ebyljMECCjy
J+POC/FaGP9V+XFI4X60x1u9LSQecGrcLgaMuodfJtDz9qjLt3V4yOE6px21oDTB
Nx7jGSVDMaHckC+0oroyL9uMQVmr7HFgo4USCt+UiQMh4ARb4Yl6emjW62FPkMrY
axYQCq7cO+8xKD1zecIp5v2LEf3yqw5/X2V+YOoeXZReLFXJt+adJR8DjCgXoW8e
rHdnaZ2SinyAv8qHY7Do6bDxzmyG1oFyy9Pnmy5R5b0=
`protect END_PROTECTED
