`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IXRwDnjSwLVD/dD6CaDuag8LuhTobXtCq5y3WTiZMQKf0rL6QoFodT+v9He9Dcva
Zt13F+KuVtfFGjhHr61BuU1nv9+B6xxHkoCaDazMKKZP2kN9ArRW+LEjGb4mexgV
DW2uhFFzZl+mlLkz0oMY6z7iSBviHGg9uzEs8vnBMZ/X3RqL3HObNetDWHr1jvsb
1SAhXPD6TyUmBYGfLhRbDSOd6oBNvscGmJksB5QWA1eTiuuJf9B/AdUeiRuBGJmr
nx7jmXLDQQQdR3BrbEoSTwpqhT0xmpg0mO/vUt6smyXXMQepr+CKu5KgppbQXSCT
CPdTOjTdYxrds0B6XNz/GQ==
`protect END_PROTECTED
