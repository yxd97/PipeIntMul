`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BV3sQ55gtqLLnzF2KOWq4ESzOnNLEcmYQW646JX/V8uA6hbGwL8qK2ascKaufhMN
/+3axQLMdAUIgQyXHvBxKg+LRHxHDF7XWhjccwciT/Ecxo/GHBxrWEPSv/QLqFVO
jbwL5auEa+tbyL3XiTpqEuOZbAMpQC1GbOkXZC+tAb9aTheX8P+nOWk7A2QigVnI
ii5CbbFKI/nLzVzeXQRwuKEQlrvw4tRW3JXjkzSGIMnLpaBX4eOD2PEjrqQD8mYD
olqYTOBE3Ve5FSP2sDtxeCaOpxsx5C/hwgYY7wDVvRg=
`protect END_PROTECTED
