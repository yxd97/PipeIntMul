`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJP15I0/g8CraGmCCrEYZ9fjxuPOWa1y9nJmiPjQbrB8lQaFeK7IANisrrU6ryVw
3cAzYUgGiKxRioXbbT312WytOyrrVgi3b+yPf4JXMratp8DspqEl4zQdmy+p1EiZ
Go41cBM0m5tI7/hhqJQ3ANtT+ARYWEwvuYOdNA34x8ydg8k1fxZp8dABx/KYrHyz
2vQhRgCYS+BkfR1Vx/WKUW8QIwcMrAROFHtL7kY645nvfBdqsh/CkWyAEGSLdt2G
RoLV13Bilp70O/lBFsnSjtae5zFHbk77SxeuSURd/CPQu6aIFV5HOAbxZAdj4D74
3taKVZgRZhd/goDDQHN2wv8jua2MNlt3ovTUCY8L25sRAIx/3vhMdne3b+jQRO06
5XL2JxUvIfthkya29txae4ipNmgYsdItPw7vp4OhbyCCyEMvRGtnhvMzyAr15zbk
`protect END_PROTECTED
