`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAJnE+yIFzQVUImtj8rZz5ehoU9uWRYzJnBJf7OxHt5L/c+FA3lca7I1dUDjrzuu
FknMumb2p0IAnwym4r7HdqGspGSbcPRkbbV79X2Lc8eiiaUviLtAEfEOrDjYVojD
wyCqG5rN2+/EFXvRMJhfLLKVyURuvT43PaVl2HQ0yeGyHdpR7VDvxFS8UOVdonD+
UsoW/3PwKlSepru9Yl2F1sjgIQEkkjeXNflA3RkMxq0kT66SIpQTWZfpdq2uqUJb
8q2hUZiVxe7/nqeVJNHFzOehUuK5CqlWRFYLw0hm+GdLKcaxDoYqr5klnMC6F4B/
hBJ7iqmTr/zHApyxalHYAEovnxXQjHEmMRhU80+lvT44PspDGOXcNhRSMQWPoHWR
i3ZOOwTgqR4w/kewgeaiODy+3uof9juS/CkXwPVX9qtNymn13vomNIhW/VdG8h2n
a4avBpgFfgavDqwcRtzOLmqhaxT0B95C7Rnkxcks7SM63UnHOEtA0ysRN5rWjzfM
DlabzYgKCT2Qy3Z2LLkcx5fudC5Cn7PiaBcC6sfzbOxRNNfmNkB05KTuvSG4pdYX
EOJy1YbGsKtyvyJQ5WL/CaIWYQQHap7blhzKBXXbtrAoCEopMMBHgt1TFkWctrxb
KWkFkXtSLtCicDpla7nbPbUJ2VRdWOs16lsj+dTihkCrbpn/Ck00V4MWAyvW6CGo
8xg2MZBriEUkwVaCr9uFG19VrZbrZPOME/r+vwayKA4=
`protect END_PROTECTED
