`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MtR5M7WM5CXPp1LnHNslRi/polbOX7tK7ODoyeAm72aauKf31K1MqB56T6T2ZRCC
Jla9+9yw6i+97GH6Fq6jvz40nd+FgzxjScDsatS1lrnpIlqwjg/ukbNVSo/SRpc9
khSMAxEP85RGHA06WL+zon9TSNv3VYr5EXU/WnO2HDuR27xzQIOHuR/Mlv9JXurV
EorxBGCqz9Hj9/7kKgAfCjt03QosG9CShsko/aPZtL0gUn0i2B2TXPsjHS/vAKz7
yBEFkfFplAiqtQqyIFsw6IwZWZrt5dHzmSepjnzj9dTIcXiwPBb3Wo7t3wSwrylz
v5C8m3zq+iaK42dTBnDwTMV0Q4Hi8llbbJOH1HSqnN7yM+uFBO0NgQVzsRSUPg2H
RR1h639LA98GTrt3ev9aTLO39pOCFXrhA1Ftb0PFGbkB2bVatYHOIZ5iHssWqfc8
0TSD3dqkTObUMi5++gsJ0FZ0ro0p52RWU/O8VX4eEzIM84O6DXb4sxupWClPCMP0
pjOf3IIOEUdvp5KjQiNrcj/xdShEYy0VgbqI7c0yh8PQR28kE3tYYKvZcA6HctIR
rW8/Vba9Jpt0dIjKz2esr4Ny+YwKrcGUED/pvf5tjX2ZKQI2wipevPmDFuucbJ51
RfFxv3G5xR5Cj8SZpGy4H4oC1BA0EV/sgMMLc49bVN8j8IocLaGMeGiFRSncG9l5
+xCvzKlRmxULeelsJL1dj5F82hnhWIa6Az4C7uq8E3VhWTN42CL1W2lO1uekDGTV
bAZW93oFWwCdwycoOOVmzbQ3w0O7d1jZKZBccNT9Z251Yr3OrK6s3/6kUmc37so2
qN9QPUaTS+G1j5SEy0LSisYoWcWdiRdmOgMnFyegwZ2M3UYD/N9qXCiJoD2bIrF4
D2VNYMlZ+U53qM719HxarrQqwr01LBMiSJ4jGmE0ZURrsacTtwRORmrW9TVZkzrB
Atn+HuFbb1pO+G7MxG0s7wLiqP8xokJb6wvEhUfdA9Yx28M/djb4qzj1lymgTunk
6zk0ukDInLRSOqLnoRb21kHgvwMnLxUUTlv79bSEAIoExCLcaqRsFLHn/rtHAYvt
dTbqMFdh5JIgIVDHpXUcUpmFmGSL2JRw+O8iSg3ylIAImZ+xTJF/A8m6QVKCC0Jx
1H2FKbhFYqfyEBJ3qIhJbHyhWrEdCfBrsr2NBStv8jUQ/2ZSatheqD+jX8wedlQ4
L18LtC+HaCYmSTL5UaBH6dejEB6Sdk8xqHFX78DeL1LlPqWG7QXQzdtxWGygaQVY
tYRggH5PRs2gq0vJ252Vxf16PIwusD2Y29fX+kjF51cRkutBVOoL/IyBlw3MU/NS
9y+3R6fYmR/4L9wmwhdV1IvtAZ7uCo5mB/nL27TRktUs0hM3x95qIgEtNbIZlxro
fIv/MvDvr2G181ddIJ0vioA5lcIQ1cy9B0sW+fqI2ZVtDRKPeC6aSLZcq3pUPiCZ
B/ON1t7IwakbvEL1kleKGlJF/2q7JId9re2TX0roukECDuvtVyO2V4xRaJwK7+0R
KhAjS5GWpOup4Khwxg3qzsk2o1asWvVgMlbV5pTpZsEbGuSW3F2L1rlz2Ak403p5
ucNKIwRLd5QTGFumZks/yY3kdzFhb3CgE1nB1cEHPFEJtoHxEJjgakN5pR41gxGK
iJQT9IKxHAdrZXk/lSA3h5s8qxg4oibuPHihGM3vhcUp2W9FUwyCSVE0oXS2oLXa
186tyHs0nU1sWyclHHYCjNhnedU4H5Vrig2ix7vIPzeNb/Nbf5bpykJoD7d+XzeP
tf1nREBoUeJXFEJCG8tbB3nwjcGJh4u1hVZVWoA2m+lnLSzrZMsI5IWfqQtePHg5
kd29vHgTwDTvTixIsFDWoU7dICV6PYRZIoWdjdFoIV8nOIVYqMpeWvmfa0RXqMW1
PqtBk3VqW7gNi5X2CDPlVM9707Ci/K9QPS5pGWYbyJU5JefkwWuckDYWjK0HPG20
ra+BsnkPJEqWk/RcdZhrNcI7GnfOFj0NSXSGupLkUIJ0wXvPMQz+u5YYgz3Bb4XM
xxG/ntU9AR+2w51PojUbEqA2ZXVWpCz4Sq3iKogzmD/M/dBFoWJXqNRzNjvpm8lM
MIc9uow5e7AX53LfQMxYRipIUfrAdB8WhI24PBJlgHxuXPBLQ25Vqphw44aeGolM
UOK8Pw+mOE1ollVROiFk+InOI/R3/M/kAqFthDmJriOQSze/ZHAumAXFTLIQHCdf
EVcnIdD75pq6DnbhPhg0hWYzWKOdINv82B6jZ4Pzz0XdgRdB5ZqL2zxvVw5wEI/+
nRr+FI3r935jcjF3j0qujzGOU5s5/gYNS2vlpAugkTGR+cAEbkcMqSpZIC7BIDsK
rkN6K+X41Ewt9xZoi93DxjSKzYC20zHksNaAirfqBuLkE5zWcd9whu25O/9AHo1V
V0H4m63dwPFnl3pF+TjkTb9DIftv0xP3QWfgRWSefuwXtwSEKSZutc0pMYHmvvQ5
caVgg70NAXad9PezLz6WMGOyGNo/ceV6ZNgZlO8G3GRKRzZU6LC26vWANfjrdaHK
sTiBON/E+y5GV3A69esngtpr99lG0DRT2ZScSDCwyZYkQLVoMesbmr63ZAMObWt0
99+CjxcsrXczujNHtkd2xnFzcn57iEGKEjLJJtpr2AeAdhcJ4n3seXlsL9UBhNIm
KFg+bnBrJBwZtK95veNhiMbm9KzNFJ9RZndNK8yQdoip4IkuWVZ5cTh0CSZ9g2ic
Si5O+zIk7iN/1UOoU2eW8gbMYs3lfNX/s1lM5hx5v4zCA3JY/ByJ9dkqp+bqjz6S
/xIpxOsMgGctKHD/y7/tXG8wNntgObvbtkt3tZKb3ckb92ed8hYd8jyzpJYKhm82
PlM+Od+X25S6KVPIkTt1nCrrjELLuWLSNbq87ACSzln/PSucuQauAL+qJDisMyzv
HG22F0ARMtM5LxDToTzHlniG+CE+zFm2gIzd61IGeWZExQoIwocqL2hTwF7izKr6
qvZriW82U1ZVMGiZiPQLiW9w7lEke0PKXDynYo3RD2Y9uJi2EGzseA2F+hO+xN54
ubeThrfctG0CoXiZPKsEguWQUy5SIV+8b9WarhGY0gEX8XBZQxPVAT9rNwGk7VwY
ONQ+zUOelVq7kOFEvRq5Upwgw56lp2cIVzJFQLnR2RX8CWJDnciOAOf0od+9kmWq
yYRmColInIBv4IN1DEcqpQctnFWxaq1lezlfT9tWocWP4AM/JHkSB7Zjxj2dVSb1
lbMrM+lru5hzq3NABVtkkAHL3D0iEZXvXCy0MN5vzSLmT8U8/x9gjU3vlmPnlwAu
In6BlOmk2kRJ1dLFklP+f2xAI+CZtE6qwWiYNQnrrmgbcwsVid8+P920gFk176Q9
50nrJAIXoT625dwcgqearcqDlreNAvgRnx83BNH7DO+AsoE+WrMK21Yv9KIWKcuS
lv7nieqtq2I4Q2KbbwSVzfASmg8Vq8iqY2YqFzfvhQoZ5gAGDp2Lo2hYcQW06odr
pXXKbdRZ0rlVm1pZbRewIRPwzHKjyVOnD8de2P1IKGPH4iIvQMl10DhftlLYQRHy
qFZl6GjFvMYornva++Z+iq7S+RHXhuggTO04gqQ9ofoAgEJd3WsWuILPL9FgKtXm
YR57qKjOOocDO2IquNBUDCKK0R2Jw0sjb1B0C/3Euc3/COStcHafuk30ovPRylgS
vG2K+YHYEZ/TrVeRZDgPb/qPluwlq1xcOFh89BdnONfWo8JSuDNzeVCa/QoispAP
ZJYDVyK+1294Jvg0+jWkE9AuR+P8lb5kMnJAbqBxS7Piys1pGUDuY216pksI+Pz6
N5V5Sp0febeiVAzJvJvZNt2E0M/krF49WFT1nw1fXWrjAwyugsmS2MjbNk0joCdi
Vno5Hyubrhluvqvo0ho0QUMMwGC/DQZjex3JxyxjRz/IsWsX6UhsbWR31P+LKBoY
DY+zu5RSdE7bAAaLlGeFrFiFp0USNGjjCZ4Y6fXiHpSrDUXl9Yirs8huysXJd3XR
pcoYYRavfHcNm8XzksSbG2KlJSEhoKsLjr5BvbOyrfHHCvdCrky6zqWf3MIkxhKR
ut2MRs09jveGk392JTq/RhpgGCVz/ZG+JIcBURjKggC3vYi94CrvqHd1DQAcyIic
pHpYdj1NQS4TORxcVJ3ayq3cLHF0IBSIY7FH+Cx/mh4Ob2kz4O7ZjmDRmp+2sM/l
INjpqocY1lA7OiwD/7ADyfzGqz3B34vIeV8W6+4OfjeBNAxzv/vtmXVlCFk8TUtZ
7onW2n/LhDIAnwjC9Of6WhJ/QoPTKNbEwhAEV/3u8aNboYEGm7oc8MUhPOczXXpp
31rrq3rRXRVvnBJ1ckDtuHyUS9WP7OmfVas0Zo10HKV4PkfQXzSaqsN8Yr0QLvYJ
4lCYqKF8uzyD/GeoitHGkndVKVNnsBbipv3hZHYKuhx47o1/IysdfiLWAZ+VhQ+v
7eBVUSjIRuL86zC+1i2jWGoehiAOo+grPfc1hryJpbhmqXFwtbbLsuYf8R6xnHSm
Fs6FKVRfJWEBJsPvLeKdenolYeluO2AzpwvbnH/1+t+DtsyrnFYE5KbdpHlzOC8z
yMOiJzOMM1Vgwh9k0gQiyEUceNDTN95qpS/d/5ctFCbRMzg8xrBsI4NqRqv2S+7Y
VXPx0watf+do70pEIT2IfQPJ9ylWrbGt6pswk5uA+dlI8ZsPC4GbShGPGL0zT2uQ
IppgKh630PXnC+W8NYe/NwIHZ+uXSF5AQw+b2loHPy4Z2Rm4zgjmQQjObSTFxtdu
PkO6JrvZXB9oXqB9TgHZG/09VMbIcsUbaWIzqCJ6LcgL8v/ZqLZWSJZ0piJx/ros
PGkVHrr3gUahWQoSC1zpWbR0h/KigVNGhd8/6JnV8SjAISv8nMOAJ0E/I/xMlLFQ
OrIauRe903C6M4NNkdmDcBT/4wtxPX66E3FlVq67xRMXMLSeSKqMng9a75w09aJq
JsiSgwIN+dy8NT11Z4oSqzvt63SrXOCYRa+r8S1t9VP8mAgays0FM4WZZ0NUtG8w
A6JeZ9Cizlu0m8led+6AsHTqF5kB9FjnRNXltiQGaoCR6uj39ffJJnOu36fYGXzY
h/dzeBIOXS4E+gdR9V7Qp8J8gCLEA3r6iE4kCY6tT2D85EmvGouAv9unmyCyUBn0
1InWLT9+NQH9A4g/ZIAOWtNJMD34sT+W7cG+RV3Y3ES9BytZ30Lgj5aG65UyRgOy
FXeDhssxzVi6zSaNcmq4rSfctK4DOgZgeBkRgPgL8gCiklOerdfej8KVI8LiLo40
SDsAZkAb6Wm9MVAoT/ihbn9E2trawNWgj1H2H0H+dnpgZ409qt7yIj3tzVf2kRcH
qdJxLvm+R2wZ0wT02sJpVinN3kCbeFTCSuIs5WFGnILvX3GGmNKGhUH+IK/zDG22
04L8kHgEPOPeffNT4zmdk4lKyoeUJHjYfCi89Y8B+YqGnupMNoaD+rtlGA5vzkEo
zdX9sy+ZYytlaDG9Ra7/HTjXtv2L1Na01j7hdb/cgmYwLOnzcq+P7VvqSS9IgS6P
jEgcLDAcbwdw+5WkeRfhhGxcZNjE6kWjiiXwAwQvWV3mCRY14yhbCIvpBc4AUc3X
IlG73g6oDZ/Ex9ur6Mal92Sp3+tkmr3lSCP7wVbcToTuNq9fsotx6myqBjcgx7yT
yXB3vq2+X/hue4Jzzo2QoGh6XTF3rpW3sSuisqal/5z9Q6y1B8C5FL/5gQWYpmrR
F/SEXMKMUldBOX6gTXV1z5SzqT3j9TDEPxuhKa/U40iapBiz543h+cTBX8Y5FP9n
so2b8DBM7FBBo06JDT/pbUZgDHAH62YmNuiKgxhk56+ddLyreQqSUmCnPlkQTJ94
+x3G/ga9Tlezr20REC1czBj72Hqk4jKx1AUaXS3R9kugAznlFP95ujiBl5Ai0vBI
39/WiVUOTFuuajy2rxg4X2+7+x744aFSxtdrf0KsXAhpKrnDFs9VC//KJ9Kv1iCk
aT4ikfleek2eoXaQs7ksf6J639ecCXygSxfqVROAxSGMtbX/jskeN+Bby463fF0H
bZUvRE/0AUjMw1EuN7sqFuhrEsx32zxocuowAy2tt1iNq3HULVhAdxqj6kthjTM5
OAIgB/7K0qrIw5xRfGDhzbVqiDu8RHReOiS8XRZqJobVjPLtfb4mwHmjO+MZoRyH
zJ0S+D180WRl6mpTb30mWn334M6bx42sgMURLZ5kXOhpBbYGiNyXU0ncFv/iyiWO
qanrdNgky6VRXphVNoEl6W5ReA407z9Ox+QjcIsD+phfdIyrVnU8VggejhnYTLQh
/aun3cWCTm1RFkTrDGNUTS68siY+6mAel7Hqg9kZ3CuA+Yivo0zXT1+gVJ36ChTW
0YctyJls7CtLwNwwCqwYJLAfbOtEN6T1riY4hE2y0l85FSuPvcunPlZ/HOkFRFh9
9c5NWclkINwTdlppCTaZq3b+ODvVHxB+g1uI2j5eupFX4AvNrhBFRNTw2PMKWRdO
XHaCH7hgch2SZiG8dm5Cq4BnJJL+Xqrcoaj+Na3/CKgP4k/q2VyzhKli5lmWegay
TdmawJDV9p0Un5RhLBCVbQp4awvT2uG8LkwvcHlUSUOmyDgyEvNKKSYwOii6wkn8
t5OGKKxM1dXReaTN7mebY2g5iwKpaWJ9izWMApgs7m26f5/XFNl0fPqbGgn5JHUz
MEV1axkCSy8oUA0dk5DJwAZ4plFNW3A0hcZrC7of/wF6vuDmshm+4NdYevCRc7Gv
Ldb1U/lDpKZKWSmQBn0lBKKmjVqnkYIQa7sawV+DC7S7pwoZeTYWkB5UDjSSCNLs
oja+T2Dklw78PxshYeuQFlowAJ/n1tHz5kgQ4LtfuS3G9yh0WGMHjMNxNtQhmD3q
UcjYfTHUaolmealaenZm/Sj6orqYJV2LUpt85T4x3B3eRP3ArQjxMrE/JsJcSCvo
j4zzVGbrwEney8I1FfKtv1tXrhxr3WxF1dTu8TpGawuHpKqbO/arCcDv+L3NsrqR
2qTqF7aFnHJx6Ult1GMHF6C/HmHDvkVY8hnHgasfhsRSMyjk+Q07ljN8CUf9nJu/
p6piw+Ezv1k8qm+Fr1N24QmGEcsjkljkw7+yxIRbItb+cHX5VUgf+DFZc9HBlg9Z
eOGmxSMm0F4XGbSCE5esUHKNIiGTiJseQU0ifpR5K+ko8h5yiB9jaL/QNEmFy9XO
MkcMYr1OP1yEeoKMKjkjYfgDQlDIpgnnd903lafkHVNP7MRu7BAOlup+N5MPGaXt
VuMf0pZ+AdpgMYpaDfHV7zdOQySk+LtyRco+9Q1tG6SOYxAwOTo16Rk8yDVAfcYo
Qu/IEcWzvw/JVhTeJG9MH+/W8VEQiIo2/ClXizomJXIBauK8VhL2CtAURwf+l1EK
EjD4kTMqH/IWe7TFVNYK528FqzIR2vBx5Px1LJ3Rbd+e8yzL1whTuihxx6rEIUna
HmVbYdrHhJdPlv5xDWpmGLpBnQm7HcyVu+hWzOKCcwHxW/bgJFkK9iNL5yvzHBrn
qFTuicm5wgdHHSIOHzytipWbmZ1e9pKFNU4gvEfzJvC7ApRpvptQXQ6Dr4xVyN4v
z9oLfL004K633sRz6wusyYG+MP2+F2q9+oLIPMAqbFh6daBvjihX6nPKXDpCTGio
x9fe2uYn8LF/kAJnWKTQCvAOsZkvtrjAz4xxGxXxmWMp4itnoOPu4sn4NalMt1nD
yHVtmgTvwUFOV+JuO+TJpqpS/dH2MjHH/d3TARNlGavLRmmlGBMbPU1PeuA0vFJ7
QOBrI11efufTmde5VbM6ehWyPo2/Hb5zl2t42qgtKTj+FoyuYAHKNtReyD6AVpfd
b6iZyuEdJfLEA5Qjblhh8/YYwgr4goUyCrJKte0SDFjh0SyQ2wgkL5YTXRezivS8
5DGg3QNlROlp20jJlKlXiu+YYfkY+9/8suHjxp1QK3ZSA3Bkm0vsAZeEFApaiz8l
i0CgDaqgrlEoTx9O6K2w+lRW30TU7Bfr/Xx7jF7LKD7Tswoq7UVMH6O0hk2KVrwV
1PJjVI6PMQ+q+a6HPBZJxG0esrtHRSmG5lK27q5DG/kz4xwSKBEEsIjOsnlBQucv
0mgSuCDELqM2R2yWW9cB/Fh/AeuZRRUIR5t/qFMkCZ9CW33RFAWF7H9Z32tMY4P8
L/Kbe/1zcA2Kxe/ds07Vag7S6I6hEsO8byldWDXouCn/jLhyWa1IJueYxlgwb7Jc
JoMUH3pKf+867tglhfClo4GtE7V8w3NnOnpBQABj7PRhY8WJ5AgY6X4jkkN49VTx
8NhUXGJ7ecJcBrfPrtvvnGmCTBqeUCBdv86HvPch+DdRSo/RUciBXXCbVBFrsyby
I3H6jq8g6Xh3o2oWp4XUDPQnIEgY8jkYJRC8j54KK29ZJAFUjkGc4GTQzk2hV3d4
wrIZM7dY4d0wXVfiKHNKuBd4dxe9cbQK7V690ZTL1ZF9vI+aX7VKCEAqFBV+rirR
6+/mVHKEAJ0tBkBDPGmz6IJHbBAlnFhJ76iuNwCq9+H+9s3imrgrXj2fypSCuqoG
4BVMeh49MUhodA5EDn4vTcqOsyzQX+We4yQoV2eXj/pXzvr9JqB3LTciS2ghrVcO
wk6gQJeDU4dXUgCoKK54TCMRVw2+rfkBw16tdtT4C1CcEvPQeZvSpXzpeWc26xSi
dA7hic5NiYD/TAIeyRgi9Z5VkTf1yCHIASlx3IsIpwB+pybQ83aTAEEkzdNIbcy9
uivUS+Vnsso5rUaChiGnDYoVyX669P4GRTtsewHMZt53ATX3Hi321h8YYKOS33/S
bUBruRaGD6Cq93klGA8Ci4kivr5yFGQ6cWFEJkCL4DZLmJQMX62t5++evCi5640v
jtPuJZD/JXKgiaXiQMgSdoanBjB6KpY9mRtL9Ah7LvvlHsHb0sp53/HAI029/utB
Ha0bLNzS7LXpx6wwq37GWB+m+XTTD9QpbMDESKKe/QK3uyfV710xI3egV06m3M6A
fnLpRVHMef98GWlAnIvQEEliSDgbiuclqjw5Lnaiekok/Ltgsr86NtUoRrd6AFAD
+KtVBGEjoUQuxxhFRiFFnkJMoe7WSe1r61i971MeheEZaROQC6AZWN/wRA6u5L5b
KHjmIVYrwLL7tlpQTuHALYqjeto340EIwC6N+rhQU3k+4DgEKhe8ziSbW/P8dyAo
4j1k6YOFXjCcbDYYjo+IWSVcFysiNUZizX7kF5snInp9CkGSXtFiM0UOVxY0g5PW
w2TkzOSmHIOO14s8ld3Npvly9sxFj9/sIQhDf4xpr60bbYolSuNDfbOvAu/EBloi
eXthaeg/P+dXoZHd24fBRH2SH8rdXFhsc+AXYxVjT1ZGkDNFxVh/pEDwsVJyrwGX
W362+OMAeI/+814UA1vUP/r1lO1ry/lVmq1dr19iFz1YIQqfOkI3NZbU0bZSH4V8
fjCIVbAbqb7NYbGL1wKLs2i9vGlHidcdvy+Cv5t6TwEzeklguV2b+Xnxo9YvYiC4
PXPMFvyTD7EnSItjQhDdWBRJNusOWnYKbpR0MnHhr6egJzIM5/K0Ppv9WFgjCM2L
NOnHyeq6YFHGvw/x8/pBCgBZ17k6Ycxl/CdJBACmBwYzRHstn9CMW3sswHo505JX
N1evfPA91hz7+CWi5KsMfRCrJNw1DA8lDAcap9i793XHhhhh4lUe7So5q7p7aIbo
ZgmDK62Nmmx0s7atKPoRazuecDXz6yGbdStMrpPTETHxQ3yE5Yxy3WHiynlcIJ+F
aG4od+ZuHKcB/Tu2wWJ19fjfxOIt9v5JfB1tYeAAuSf4H3tLqDnYNbV6YXJJGNik
BKqebNWR5jyuJ4tlCM+w6JsOmUAZoaU/qfi93VCgryYl33lLHCbSlD8a5HaSNDkk
g/jFizYVOw5dHfowooF1BAGIqsmWaXS1MDH2dGY7owptY8kDmosPwkKfYf5AvVJn
qTy4aS7qqScq2WNnukk6FU0cJ4zNaVKrbDDWiAO/xEbQvoSRW3IPQNwHz+Xfz0Vw
tjr1IBKTefCZvpcufefIxPd2H0zd17sYjLUMFVZ1I0hVwtpPLyZfIwpSTtYcMoNN
hRqfL584volNp5zScOVyrM6UJREDchjSX+QnrNJ6DYDgheujgTweDNPKwz0PeWkJ
TzmdOG/uFHxDy3AH50sFU3JEhfxXIzlXuj/sz4Y7yy4OdghbYvg0pah+imEoEePf
W7/Q8fKTzGae52o1rOzKh8cFoD0CRWiNvGpB8iKQ/NVWR/NIKB72vxSwdCLhS3/s
mTsQhQlvk+/CxexKMO2x/fjp6CBS58zjUtnmG2lWNliqYuFKmsQ3h0LkvoQq0A8U
dg9SBGpIL59ulnjSDT7zuMl4YcytuJTTPG4XQfU6wwlnz3ajXQX5A2VkCxOVpRIN
gkt3roqI+RIHS8JKzRVwCdUEP9QZiDr06G6B4i/uwTOXpN0NiuXupjOJCBfHzBMS
OzpvIOEMzUrG52jqJ/6cDhb6B4gpMtm9BZWSgmArc1Vx1mddaV+44HF3Bqc7zntM
qYEoLv096r2nU87grJrnMuVPJD6gIJdJ/U0A/3x/DykXHarzqh2k00gTS07d5hN+
bIWA3mz88bxd0Bmd3TtHKep1g15hGzUxnGs2nIGFtMwcRZVpjzUaUeKnDncNkKjr
rYp99Wp8YzI0yghKf2gZHCSjP7N3WB4KzbpbdU8V6MoMqKZIjCEXhRE2rwRF5Vwv
V3E9lVs89Y7pdcXHBykmCP8/jRdfJu7GQn05uYb/shGjQ+F40bsQds9Fy3IWIN50
xJmzqSy/mOraxGXp8Szq1CMhSJtmO5EwVo9di7WSnE5hSoLzrS1dsvGrvQ/wB4Uk
KneVZ31IFK/KvWykRC3SUcjy40bSZD12jHLzZootoGLaq/sYxlANaLT7hxKfQoRh
8+oRT3KcnNT1LRyfF5EiJPbRfxj+43OQvXUECCoqqocg5rEEezF/p7QTZ3XXpq04
cn4I5k+L+fJr1HNYMBDeSSZJduhBZdfiJJC4rKF3Uh91pRghx9sVEtE3phl3PIHS
cue2ivQB2z9NDFJVRi7YsF0CgZM/bQKgpz0Ttkyif4PV6LtHrBcgq17ZfwLl/Wgt
fI0XCO+sx8URwRzezKOGeMcyzz3kt7EaJQGPDw6/mHYorVVgg0JyEQgPZ0gsO60R
JNhF9kcMBKz8lz5+89cRaqDFg/Y0c8AdrGjnLs3IUgqsTS7F4JI9uPlx1jMHhEQM
uQbEkcUc50Tbuy/J3H9tPW7uogAkWmimlVZ3PLFtz9kpU35dcByAXdTMPP36O6l0
L/pwAZnACzZ0u/3lP2Qv2ANtZvZBI+jK0N71UpqPsy3ihp2g2ks8CqTQYYUxD+bh
7LU7fSOLqdgJqL0aDeBhRfJObOef0kTAYWvLtSIisGu1nbG0TxdJsk0w+2tT3j/q
jzI7XoHb7tiL6mLnC0lT3wBx2yjuZlvYq279oHdahccKoDFZd35Rn6UMuGXMbCG+
mpVll9qrJDnXgvahHyRkiHEJ46Da0K3TxGdyDWmFQjdkMMtbjuxfi8ao+Lzc/Mqs
WWg9y8Uu9GJk0aOW0JRMo/cV/SEZ9L4Q96HghrHoZ++3cVIITkRv5aqqCi1hpP0i
8+zy4ovJtU193HipfhIMHBwIH9hrXMc8JyVqaje40ZqY3mYPYq104caBR191Wglt
pDwZFK+iREOPGm0Bh24gCTqISAfdmbFbsFHrkcuGPWY1qorXMBgSe8VxliFesP1y
yDt6J1S2l1+lJ0Gfzc54nS8TZxssXkLqKwqwDP6k4lO0oZvlGvuSB3FJpIx3SSZs
WJzJ7E5ST8e1iN++KPRoLjzj932SaB02YspkRN+Kr809h8PLxEadFHowHMwff/Sb
nGteFj/fFNnXeRz+bqLiIbCVtjZo6HE1DbbMbdvU3vAEaSMq5fRe2w8QWGj5J/Yu
S1p52d9psxw1c5hmsUnSDX5yoO63aFL/SH8PBf2O0vTmvit1PZu05KBE5q+vpU3F
MHGmMQjunp874O0nWS2Z1iHJrHxMvaJHLdMGH5f9FphnJqbQNk31noEkNo4Huz29
YjXCRgT5RaCwJc0RFjVg4v5M7SyRBGjknVlJSGgkYPPPq3Qd06ubkdW7befHzPbr
z5GQfjKKVyYu+5iCw9grumNmMffyNbFMBvFAsjY+yYO+KT3JQGhtETydfb7u/FgV
l9rk+VkJ43r7s97EGm2yq3GxIfEH+DOoS1WiuZoVeBOhwosGKEtdxwx9ZLVOh8Nq
281aG+QlJEobQsAhlYxa0KOg4cbqT4iLcjDH97wOm3KXjigNZbh3ofW6QokRyaU6
sbvOM8Ltq+c/8zm+jweDAR92vxRIWpt2XyqdI+Twqv4A4y00TAsaRbWq86SDO9aQ
qSxzJYmO/WtZQ5DmrAZ1M9+O7aJyc1EQImrW8bMnBNhCLf8p2QKKnyfXNZ0ORvcM
tYyqhblnkpMBCunRGsfj5GMw4jc+IaAdmsv4rg1hUhZAEB2k07fh3c3KJ2mH3Be9
PhwsZsShXdwGecsnDtdeimO/UrasxNNoeCLqsCzZnMIJ9NeSkQq6abDuBhKiItEU
/nMpxSsbPH2wiiQsjdAgR2wpKPwANUaRJSN6ijqLGmxIEeArx8FlU93TJUEiUb48
GPc5OBtiiExFjtaLarJbP87mWuEVI8TjsAHuGfQQgytHbQTy2lQEUlWHWJ9AwFOU
G0UBRNMbKkDR8sV8q49DtrwtHu2FdwhS3svi62alIq0iglR3fj4kUvrQERzTv6iw
5fmwaWfQMSinKyZGt1nHbVCFiLkJGPNx05z+nshBZpJZ49mdLn4IeqZzuDTecGXI
Hfv5Cb/njMl8HKLW7wx5nPukeaCudi1kMrX9D50CudLUUoH+u6l4P3K/kYGuBma5
uPgG+5pttYvj7y1LEtdQmy6Bjaxi/IV+pudEMvz4C4Y5uw+/HstJZWh0eFmTKAKK
SDv/JvZO/4iwLwR8Gx48Qr7VvSDJxnZaZO9NJ927v4AaoF/lJq7jSobVpOUiMPpo
eKo/j6en2xBzECUNF5R7k7/nfCmHD6HIzadhxnKZwlPWnnMxF9bCImMOxTBE73dQ
puleDvMu3e0ttVitZt/zS2vG0Z2DNIUypjijFOLp5aVM5qsdhrx45q1Zi9UO8gPf
tqcEHifjJn5L5qohWJK0sxMSV9EayM7eeAo79Ujq8yuPCK9gznGUdrZ+or/hPIAl
4iso3tjiADqCACpeKt+eDZuTP3P51wvDLDqwFu0nCqwPplTHXqIqLkHfhEbK5Y/M
x/jWNH7Ro2v96lEehBZltlVSSkyL+A7KIgkxc9e0TYtORIxDEbFw93RBHO97DxJn
izRQ3s4oC9JjcH9HIJnn3QozRX6zXdVbuzoQZTR5Ac2ToKq0oHxhxb5c6T90K/Ty
mGF/gnbPLGPm4byVA+qh6O6TmDalFSUNBvuFXCygHr0iVDmDx6fxMjfCuMrMSKPg
opYhNkDSF98oPg7Bky9czJkM0TvIHErDnPyT0kympwzN8vUPijcfqsOzWTQRuHI7
DAP7JbHWU+qxXzzRdAZch0X0Aw1cjK/sysVIBay+kjkfgrXcLCGh2h487DfPvVbu
1JsLBR4xevDJx11ogL5zzTK9iMZ8DrKFf/QjIYVziZL7bakB3yEH1ZNledkGCllC
MKWmqUCfSVqV9iBZJgjUxqxa1nkrCqzqbVQ4XMDIhfeNHtkc9ra7Z0InlDlTVnux
BGSv84SmXGNHqw/kax6bIRBa8DPLtkUe0OtCBXVqTmUCOT33p5rLM1V4BS2/mwJU
lPaIGdYZz7vlXZ++e+c78mGhWcOb2WHxFnEiS0tFcAgFl8XyxB5Kw1WA1wtD59r6
/6BWmsKejvPTjp5zIIYzdEF/YE3lZk0rKpU5rh0oO8mt+SFfAuSZXcf3k0q6x58x
5aIN02+cZvZ5oTDi5FBwlcup46f9Zd5SnIGWIDxkhbh9kS+ZU6rEEgQiDRhx+EH4
K8rbNKOydm7irWxEXftQgNpNi6ALJpKJ0qAXl9WigFYx18lkTNe9qY+Z9ggoxtWM
Eh89sI8J6rViC+IuE80YTHAEUr4XSF3s3Rq4iGD1VxMvqqTJ+EcMUJbbrPiSgPkT
mr3xjA/FJ1cgojjr8kCaZB1Msv77Rq3V0w/A36F6cjmz3njH6+GmBmHvQkFBR8nK
iL8ZE3QF6DBRWX36L+YbdxeNTRBO5c9GDihpZvWP/XoBoF1nHpwplAeMrDeao+3p
fC8dNBdDAoH0x60XCJNy8KSdrfkYMU8i2GYwBBbHf5hZ7P3QNrCrpCcfdhVepPfE
hmMl+NVhtQCSka039a6hQEyrmniiKVKQ7qpDMAcRTVN5CFUYHewZ0HDiX2ml3T9h
zPViEkIcxvBxxgv14Dw2Fe9ao5pOWVQ1t+i0P9hHevBcKk0DA9tdaZuFnA/Qj1RW
YAcl4P6jb+t9lz+igLJeInkEbkS3hkD/I1tvd84E5K/BQr1kJANtDp4nL6EFFsfC
RkO5BEfasXfzyhGPTpApZV/R9KJeiRnaun/KvIy59hg3L539ijZ1qPJb/4YOoEIh
TmKWsloX1wwh2u9sXqnssnRORf2cGxhjzwboPfMkHHY2NRJs6pBewvpmy4rd2eUR
g3/RukSeJBMVrxj92ioKvkhMihOcR4L+OqIHvdbdkzz400O4WebMH48adyl6KsH7
x9/1EO789E6baKKnRNelk8OY29dtTSuNkGY9GOMbr/cqgT62l5ksL7UQHLwX9NRy
6Cn5D4yR4gLd/tihdrmoAzGSWHDHiZzaES0IjsYVoK2/0LfBRLQL6i7Y5eM/MwQe
HWA2UzIygtkz71GF/6Cor9DC2mWJBo4RafQyUpHmujClyDki/LaDDP6cz9oJGBZg
Xza+Ek+wUABkPS4PeTNcYudYI3btkp8SeylibNSpnNnEGTGn6LCjLiveYGlGvJSQ
jttO+IIU7GiPMClUT+zEUDmzagZxNBffpG0xCWHgbEq+BPevrlipESnC0v+5jGMh
H7FbxqU0jauSWBkMeHF2ZahhNTu1OPr3kI6D9vTaBRLb7zOox0m8armPCb1K7B9S
a8vEcHecX16uKa3uDCLGZThLzE2J/P8mSaY0alG/zdPZkkkL8X5k7ViakqgxQLIR
d9kEwaK7BuTrc2vy6EfsabY9GaDduHiubhyECq65rbGTA42X9ekqDdPgzSq+xL1K
AOyRdyVDxxsNOXqyH01CmnxV0e2E8ljnsBtyY2GSvuOiZKKMWvCb/gzxdbs5e7kX
m9fa78x8I2XhF5VMEVF/mMyElYZsZZyCXz4j6zjSDFVmtlnpcrgsMMB7BnA6nWfk
FBS8MB+sQonf5Pyr0kFpSozng0emr7vX+mJVzr1l10SQ1EpeqH2XP5nT1PfF8yRa
SFPTsiQ/DCeUtgLGM1EgQS68pR8IV2HRD/y2gBDgQFSahsFP6QskUmXFAg2enkI5
Kav7kPH+6qclz+BDr7/60BmVggFvbPD3vUnPDzvLMzkDf3dqxeOa/B80IxtZAju9
y8bhiIieM2uiDufDiEjg4B4Gst8TPG+8fDT4sx8U4uyyW/1e4legj9NONcPPJT9A
F4AF9FcjRSvejWXmjShDavcef3a3/pN0n2rd4HlvmapPAznKmsF7jQ336Jzo8CRS
kxnrdZPRw1eT5odSZHovI9LwDmqpdtoGCGchwlK5u8S0xhywmt48VwPG2TAhS9E4
4Rgke8IlRXnckn449vlCa+sz+9LWzcHRGtJxBBRMF1MXd3Kth1In48vyOFd99zy9
5ANhMc8Jm0Rp4eg27ktHxnskyX5ex4yzp6aZE4pGK7xYqYsPmPKL5JVVCoVeSvGl
52ywoRqiMBcell73kbP2lJL+rwoD6DocWM+CncaPUQdo/VkzvzSiHirjdbHKxtY5
0UQCQS05mobqebwzNk2Yp3HusHFXG+z+LDLq1vaQNQo5sSQP+dWmJI9+KnNXb8ME
uudrW7oTcy3bDGAyRodPbmykb+/AlA4y4xWbBO5E4Jr8lEzgqduempjMH9cDCBWf
3nnlw2ouboY6kCe90kCXiBMbMdVP1SLTXAOi0NOam/skQm7xm9bRCLrYO0YlH1AK
/OepzkT15RdCByEYgDtzjhiWKpWWax7/H7zj5SsguLDVp4TZ/YWcgxKSd7pvYEYu
oTPQKKGiSfhQeJoTJXCwhs77W2pxDdNQWp9vmAKwY62mdklHqPIDwmIvyGmYJ1Kr
gqVxQCplry6SGuFtlwPPaB7dqeIo83jiqZGRMaxS6pUishJmk8Dxjp6S7KTga9by
+GXtm2/7cdcLi11D9rOz6X6tPZbNqwwJFv20T/icCZWRUzUTKkb+lmg5TRG+z42U
6aaPIzQKow0HKLhISGqmfxDP7Y91HVVazmg1z+INQt8cZ/ksZ0hNdohSc2CB+P19
c3GxoLYZA0UlxCankQjxU/JDqnPAXtYvXtz3inwLPr0dhx53pdmqTj1vxo4fMmQD
BGBmwKJhub2SfaxdMAJsua81SjOqm7AgGcF07lVmiL+WAGknYuYtvyoBOIHMr127
savwXqJqEJtjvWo1egkiDwXR3nxucDFe+gfQIa+NWTY2gSigHU0ykAq2a+oAHnDZ
2DNQHlzCeBnbYby1X4ZHDy7fmaGwHG9SLNhSol7zGQM62fjdVdnOVJMys9GsIV1l
KbxsMM13mkh9rE2ecknF1055Z+IC8O6rUYqk89pb62/ChPEks+yOatFAmLgZjxM8
f9n4jN5YscP7z2p6Rh9uuuQfRfYfBCIvQZkFb/IJm22uw4iYLjsjpFOEPvUuOLZC
bjIcQ9JcvioLjS/gcmiHDuX2Tb7wdrQhzqdEpMZTtmapIilgsJ66ZahvhTjkr0uh
O3/sX6d9Jtdfl4YVR3Voy2bIxnZMfVlIjrd6dD0JQhjX1QCEEIL7BL6Kkz46pIRh
X72sekOwTan8U413O2PtWvrYjQyRrEPWJ9XprG5iX6wZ5TjUSHa3SPaL2d+nEOKU
NYFxAne2FdA16nFlplGXaUGdbTCPJ1S/7Rc2vvFkKP9VxKNtdrWLBHKsrDkuzpJ5
Rg550XpB6wtoXWR5+XjJ1lvmwj3nB4HQ8ieRE0+763ojp7w9Q7mP8gTdhyQyQ44l
7Ik1qnjEjW0cndIe6c2HhOecBSt23V7L5SD6MAow37vn4PwKN5F5VafJGtactEbp
qStJ819PGqwEHQPpB9LS3FGHztByTBg02+FHCAWIOP4KJ/dfk5+eJts9OxIKj25Q
uynpVyX6GjEnwxIYAXVljaruLdVHBd5EuvqMRdof+cFAiCWXPb/rOeqEz6kY7ylX
6HjMkV8iFUCZDH94iIFsgKhG5NBpKhGJ8APnubNFdr1CKfo7Xfk3taLmu0zTSjKU
e6t95TncrGT+8l3AEh4uAP8Mwep9c2uw9XFHC1VaSSwT/95Cig5YXOFOjGsCBfoB
q4E/Sy6HWEqnZIxhS8zxHJawa+s8BsS6skXASZkPplqh4jnSyDCGNyHlVGNq6nuQ
BHPZGDzliPIIhwNRunRquvuoMCwEnokdV2sg3IKow9Wk/RWEJFF2AX4PbH1oAmNT
+POqRKl569EEnkajyVYsRFWD9R/UTucAj56ONNtZ+Og2YkUmnz50Bx99DE30vaTO
nX6wgeqgH+J5pD2vnyZLXNAMytIrjg3mdWidCj6ch4aF/L8AYc8WA1BSB9O/5L+A
fBWmIR3SUa4yn4KXtWeGn6VgcOpGkSmht+LCbkh+6l4=
`protect END_PROTECTED
