`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XS5b5OTAaam/BVMfLDZMUj0vrxefXLj5PZIIiLi4tY76pcrIQePjeKUtZ1YjU/Me
FekfibHCPKLN0ZA5zzvSXTWzpdsCjdylZLv7D1rIpABwh9fQyraayGZKJYIZvKPd
vEIbVrYoZgmSQpZ+yVB2HTkvyA071tZS38oLfRwtLwGvQpejkDq8UiFjZthygyTG
t5zVqYSRZEHXtbnSWYbwzCkO+si8+I79xQ99F9PSSuN1YgGQujDy/ekkilLvIHKJ
5yzGw/Yr5sb+brl7aCLNY2U/KIs20MwBr9qVWsLSxqPVdqM4J144rfhkPvT4Ly4e
514BPStqR+Eyg3T9AVl1U6gUBZ2Ll46dCSRQGkx2sU7IkcdL8+qPHbnReb6RtH7+
TKOkL0bE3tOEXvi7vSgYpy0eMRRfcN7sWJeEksacWdHZcR8rz7Lv65iF2gmW8ucw
/w6+Ps1UdEEIVOtzPwNbJVFzIiR1+pBm32HIERK4XTxNHBoWahjd+tO8HWfzyi8F
4p9YuaA51B1Hb4Q6KtZG9sj0n3pHCxvcwWZAhqkic3gd2s4rO+a66dND/ChB1N8K
qmFVNcwUdNsI1crfvCbG5Xj+UwjQ9DmHw01m5Klt0RC93JrX9KHYBcH8PKms84yM
Ps5ErdDSgIkEXPRBIaXSvKR1kwuzJiVRi4CWMlQoGfGM4L0OtwcezLlj84+Hexh6
eCNjTBdztEcLOnaRBp/Y0tey2pB05eg2xV8mnXZDhO17LI8SoRj274eQmM9ien7P
p5WKGS3g5VNwIY8OAkQr7HBwqHybaKW1/Md97xrdqeOrPqJ/RYqp25yOYNS/c8Eg
gxWMns/tuvvNYGr6oqpFe/apoz8ZDGZVWBb4T3xYBKezFt9vUI57FvTLiaroqN6l
QzPiqY5mq0nm76rXB+vAfoAajfe+pnUR55HZqKiNDUzesjXgMxcNyLZLNRReWsmu
NGrGZUdHv6O5zgzsLfLdJ9KX2UFZwjlgaX65N4zWBOIum7LAGmoWNWmfy9d/WaJu
q3/W03LDLmA0qjqwd0WRRi0wDFH7m0C38EsfBI/HFF3yk111XcMkfO5L3kJEs8YK
CjXI1sYhDIBa4G2uGYwrm1Y6TScRsstHooNX/6D5b5/Dq6/ULTfs4hQMuP/qPT5a
kgL36euYpJLdkfyiI5Iq+6C5VCZoSpGOXjkol2lcy1f3n2/L9CuEokTJZTSX/hPJ
ZS0wrYislAhVIVT4a8+de7O6PMc8m/iyByahX/U+BTIbpdKj2yrRAFeNymshKQuj
tBOMlQ9MoljrkEQMn0wu9Gw1XAezY038oSOC4/m3x4cAtdj6CT/RPU23eO6KCeY4
27MsUMXwkZJGigYFYerSj87QRJBhTAX0GJyvGQ9WLFp01JE8zkWX/zL56JVpCGC0
fg9ZBtbrmc40y5+dwujvTUOimZMFBwuRzVvvDkWhHJPKWpbKWriCWxuTKI5kwN1+
u49HOlDi6EELzC7w2ChJ2skk/+7i9ThXi3Cz4l1xDEnI3ZneJvcj9va/rH9CMFgK
x2ACHeT7o82NmATHUyiKEqh8WCMKWXzjFij16UQ338s6v+XjyJjp5vBPqHU4jm2h
rUq6/iIckVa4FOnZGz89cL20Y28OMwLY9kW8/QjtdaWCusHjbapQp0Fy9PH0+D0K
34uKd1lYR28l87DWUkJVFQdOQw9jDvqqG1tfrcFlc1XJDrGVemPoXug8h8HoWL2x
a07HYIflIxPBJPgtlPLv8U61ehiRsM7totmd5lKJXxNtn4eJn21VjLVW6AF/ZGOQ
N/1PlBAmFzM29ejo8LWouExOAjr+dgRRm7gno9KMpyFrsNOR5F9I4n8P6Q1Gw7jU
kVKl24mkFAmywvyh1vsrvtUET9Ch7clTRTHEU8feBCDmRE9dOMe59RNdCZGnco90
0LrVjyWW4HhKSsTejQxA+ESVzzwyzpTd6obQA2YyfBeuSsfW1SfDrmFdw1wMOpHd
iDOm29nP5IWg+lIdIW/nrAgOHTbUgvCcU0W7KurmTmyIr6EaObg+zs5Uj7zjeYHB
PB7S1FH+KoAzXH0aFtlB3KSgx+qHtIIeRGlgRWM9JsyV32FoIDmgPhDPFSJ6Yozw
S72r0yRwqAEBngd1YDMFfb/8p6jYgLq/+FI/mh+e3EXUPOQdxC6vPiZo6ori8C4g
ENTJxV8rmp6VkC1R21jGjshgmUdE6RPef1a03AgLpFMB/7sTirqLFVjAMm4kEu/h
9TfA9FcVAwdrdlQ12XRyzKgho3VNrN8bUYV/Ig/0hyq7HElBakOnR4ByYOt+qLCQ
iRernvGfngyHtUjH95evzGR/Z/HKc5Ef83zw8fswMKx+MmXJoCN1+KqDRKs8b4pk
XV8mObvFohjUs7UcvCEvOEXZjBKeEJajhm6RhZMPOaVDx2XIKFIZsIgQU6wNWecU
u93rckJGLsaxk6NXlgk61F4dcj5yzdC97rA66/siKy5IAiUO5iuDqO6s23imLAxQ
T0zmgnJxr8luYcY+H748hME7UgVfLq9TPHMtEzRI4P+J8l9haaRapn5ZCGCqNT67
CqiuVP37c28g04mR/ohpzXp0XYJVO/BfA3l52IB7eSVMcw9c8z3/mkjwXvbtSKB2
zWIQLArWDV4PMbp8S0/AVdXZ+lCGZySnvX/a4oexyRaAD62Tv/US06WL0fD5uJ41
SyU9xJv2JDnmCjcUP/k7+mtvoxk2zoprAzmTPiG7Dzubor2yjvI3JA6qwaUf7rgA
ffqNpqjd9NFcIunCWRfnhnDsOoEFe2uZh4I4Twb0bu4tnNhIn6Mz1dFmM+ggrdZy
5s/iJcqnAWJz4owah8IJ0hDuov9v7t1puhyuaiPrMvBdkDufsJltgFmyMmBzBzwT
cZNA5r/EhZSMHjZXTgpmGdlGNUivMTH3zZYFfmgoR9nSPFvS0qTGXg0Igem8Y1nf
pcDIVxE6w9I5HYh2YdEtSp7hPlT0IKUpU2jBUpdptXO/FhA1ftrPaqhELyLpn30F
V2KKMK82GSFtz24s3sidyf3MzvQJcaPp8s69pTE8geDRR1dLOMnvYN+iyG+MZMWN
bK/r5n5cWRk5erBMBif16tPe+LfIYaeHLaK1w3+10IhOwNY7HXnBaTOgyjID//ay
ER9s3jDNtvjzbKAn4q/AmdOM/UQL3oD0LB9kAVqZ+fIOPwomYG/RhtpTIhYHe88l
qqq93oSLP6wR9i71KkNGndg+F/qA3GL9lPJBeSgRmZUXpeWupJEmitasipdjrKtm
iqmU/w0NNnFvT9/U4OlHoC0FnLXtmYmAWEsi0m/kkhHUUwpqDydQHLC4KYF3SX1q
8cz4Z4VHlHdKrLuWLVVcKU4h2HXxTln9zkbQBVnq5C1Cv5XhCsXDhvCfBCDPOa4O
r+Z7YywdN3Fn1YP93Jxjjj9JU7vJN+NMY679AfBdfgWEbdtzBjm6UFNBu71IBZMd
qdQCFy8o/cy5Cvw1uHJDtHAln3BeXxJIg+qECiThGuzHvg1DFj4ETm7CbN9OWR5V
fFnD3In8Ww6AyezMATDQVWNpSkHvKKu9DwL6an0KdPI1qK9b0q3K8Zepn6bgAB5z
M53M7zxfyZu2C0/aOuJ3N9vVACJpS35UdTgORx8zH5/pZn/V7Ri8OW7IIW/4zQ8A
l6WXoz6YTVBzlaWqb4A0V5PWX1qIIm6V/Z07c9DGKOTOFTutTcn9lfBokNIgj4Vl
c/008FinIUbRoVsUrBfC5Q0UVZcf7f38CVimz+c923xLkAor6/mh2+oOWCPf6D6W
vCK+S28U6tm3bpY3WpO3aXIWxxFABF2OVTpNqOfiR2PtjCOoYD5+k3vOsFfcr06P
ILY/Xjzr749ZO/ghPijM6UYMkxC74HRKAuF180vC72rBqcmrbQG7GRkr7+ouHofH
CSDsPmzdhChi2BTcIMo5dSmlrE4l0E7y7W+Wi25CbnK7JalFyoKjz5a4NV5EYI1R
aoDVciAdvE2SZrLTGUrDLuTqCB5/KiJy6mlDPRrcdhujWu9MVxL5ooHyF2RHp8uW
ppMjll9XwTjEDv4zg0zC9AwOmXcEbyspwNAOlgLk4frHvIe8uiuVpU5El57MfOsD
hul80nc2nVRtgdYbOngqVIayJ9wWQFqbx1R5jNIqaD2MAt/AfBJ10QuCLIqM2lzt
MKYM65TAkvDaXi4mPlH2tTMZB2DMmOY9lyi2secPc54tyf7ZzIb3MQVD0DRGCrf9
pu8/JeSqJTuajAO090qEh2qbWCo1tuxdZJirsFehhEDpnnXUbxbcfWNZlxQ1XfXS
tnN/k8LWQm7Xx5IV7qhmGRj98igYxIbT+uM72mzFupLUaD24FCyxgI5eJcHzRz7E
l18lJcEJh+ldDdHztmg5n6xVy/ypwsFOiLASWfmfeo8qBVAYkLVT5GVQmCAomSvj
VdyAZyS0sknvbjc8+J10V2aCRtB0jFZqEzepIPOkh570WKYTIHuaweJiYlUAdtra
cgx6OMuyLggoY5EL28bhE6m73IfSiRqBJWXyLNberYua3U93VeG6mibLXQ50vc6F
bg1tJhysGMko1angtM0Epel6DqWhMr6h/8iKoy2/L8dmi7JrhPeIDN25PbBDpPAs
5Ec7axb+oQ+W6mDHdQIIxwEV3ZNWjy/qA4dUaEk5/DPM1YlxsrjDdS63BUmaBN8L
78fEfBNmVzCUUi+69mU7CMLAOhPs49FVEpPvuDw6pc1EmM05DTc9Ggl8CLXji2w4
U/9Hgx0rZBQ7ST+YtTyNP8gz2qGqa7WAXsoCKp3rMq3cqaCFpR2K3ldZktsdT3eI
6xGC2toHWolh0mqrTW5Z2PPB/nrkzqGSTursSVio21rdhMuyyPlCIJS7H7eXnXSf
wYBUl/0WMXqRd0F9lhQ+FUoN+05oJCXCtdrqANUv83A6QWzq1iBjRcclAoziWlf5
8EQFzh/KA2iqGBgzfb6P8OlLpISnNqhRzpa4SqKjLq9JbYWwMiiMe7StM4IwK8jo
fYDtLDVpICqV+0/wToLCOnfA8JGITHUt1tzcXdfSyMdWdisbIISpQixC3nV7PHYM
Jc4YVoDPMS/oi8qav4dn1rmuKGfmP64FyG3lnDckL5q55BdCbd07U6cgXjBU+njE
iHqAxtrHcPpj69mUUMvNVwU8bKsRp4xEOryfLBdVhjkIViVQ6xB4QHX/NzBSTyio
K6mSltsO50KUNccSdh5bGNmqa04qTwkTq5aHCKrimPfeLy45pjyje6tKt2IJIrxP
UkIYirypWS8b2cdFLBzrHMH2hcuFdaDmGs812RLBNXlje09J/WTkIhjtCa/pvA81
3COtFUkvhl6aiSKkfygBSz67f1USTK+vnPMWyuYl5CzjPPPdF1kVwjQm3d/Bdvwk
OTpCw7XQnmL7l67JyBGPdqWv7W3vAX17Gs7H4FJs6fpzzCI9aNNwJ5FpMK10CMsP
rFWgkpuoo4NukyLstK4tY0UFKjSo0F9nxaI0OS7XpE77kN+K/WRU9rriMZpUvNw0
c6xYDe9JUduX35/5vZXqb5fm8/AsxK5x+qP8ADFwjOr1fh+yTOco5yIl/LBa/zWR
i/8L0ZXPi70eyZKzIE0yRkJNWwrdNdCDP7rTi6LrSRePsim3K7GFLS7qmrQM6iMt
l6W8xd7pJE+xp3ocwZ6eHW7EU7mb4aJSwOdeM/no/Zd8BWPOLxPLC5n5Xm3mOXSp
LIBJcl3Voyyg3FLH6l1nV840Ll519gxgSoom5JdBcxTRFRgCNRH6EeQTThev8k7J
DHy+Us2b44/0k+E7a2V+/kZWOL6Qc+wEHedqkz6DVjiyNms8z9Bfz7ElQgemy4rM
H/Kiy5CO8F+ggZYnq6V80sQL/xJd96PBf2tWkVmSN6vLl7lpm8AXb6t6NJEZNPsP
ehyhZmmMh+6/NajEvMJUxXxwQZcnFekSVEhsf/qN6+EUCR3XmoEuMhXg1B4b8aAX
VdVyDPQwe2NaerhGpXzPPgql/cfgYPr6UcoJy2SZpnKz0hPh1tf4pQx8qpjnfRpi
f7YbRKSnh4qpLramZZA2ZxlvWl7r6/jxqQ7SukhUtIK8u5pgohqvoyyXiR2VJL4w
v6AwbmsfjGzwakF3PR/PJ0SXHyRUHb/F6dRp5V+D4UR1zuxIkDKRGctbTsjZrwxn
YcpxBs8c1NFOx0WS0PVe88zlV7Atk4Uc7w3fzqDmMDPruEicrdtyhPnoj8/g9HYG
rdELML9pcz1TZ26A/QPdefXRJnuoAz91U/7qka5Vl3YhNNonV8kH0KECl/RNIh1c
jDwpJO/90Q3ilvZmonwT5Tm81h1eNVrkLSOIKhltfzGNRJTVXvmP18cvyIjHTeSM
MIJoZ4ljeG6W8LeFXa9m3kvj/NwetQQuP2rxtITPAZc72ZiwQTm7/eBKgo5e9fXw
5ZMzj+c03QBUDbPRVdSrEZwqiH1OxPG/pU/uEx+mXETI+6GYpIIvCUIut78PZkYK
ZMos4TE0Gs0wyusO7xI7Bu82L6I5ZgMums6DGZh4GCtYj/ksZY7u3M0lFfMUstWs
qzc5tsbhyGhUp2M5BIxJkw1+4cCLeX5INAVfG0HCDfY7RMGjyPDSzQeLovzgXmRg
d34jAbgPXH+IJVS6aJzmV8UKktP7+BmNl6X/Y98KWsI+1Wumr+cfYu5MT4q7I1Cc
gyr1PjYTzBqkSP4+XBNuh+mEIqR+C/BYjsN+hhydHVmRwlmvuVXskj78rYGFBA5s
PP+LQTd+8RqeqdkobpmFqEs/Ivc96Y9Shygnt+8/bSJs723KqS4jwztnXIPa3roi
H11m+GDd7Jr1+S9YBLrMXe1De+jCoA/smblaHKlocC6BSsndPGNbAEXtHrUW4/7h
fvynCph2ALPYS7I6gbwusUCLPCUDYKS8fqkqI1nccJUzMxm2Pb5ZprQKtW31Sk9R
`protect END_PROTECTED
