`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6E9MWc63RcpYq8W+un5aofvXDkSOrDixXKm/XYG+Rr/xQn1/4WKIt3gNM9IT1P4
n/ctrrlWWvK9a449EYKTLp7DqrNdtNwU0MKv+9VNU6asmUH24qNqA+0KpyO/kw3o
XWhXog3h9YiZOV81tQHWLYpg4ZveF5hr4zqQSVEvuuiMAVnD1A0xSLXJwx4r6pU9
0loBgNka7dmXba6lu9+qz1ScT4P6/fhdaNU50GGOyWqj5M7dKE+h5VUwbOsQFO+h
jtzsExI+C34jgPK7Lk10On7Lm4lFidfd0Beowhxtc6Il+Js+oirIeNBkijd+QTR8
02X593Q441EGfHmbvxvCaRho3Y9qEieBNDNkpCcyJ2XNhielhBENUPCuCxN9ptXn
MJQD2Agn7yK2c5TpLKcrhSVROBE/8LQK/ezrjJ3Rq7SU4JGOGOAy5y+UDjcShofi
KeIqcZ/drKwwSC959mBvCL+wa2j9nl8M5wcd7DtNVCmj4EqoGtw9FWZ77S87qnWb
SuwwQYp/xoId2lwOAX+KLy7dIGU6JoWtEwKSVprOiYpPSmCrOsWReqxAVeb47IsX
45CvUiWOSidv6lSqHYWe9ZwikSFdb75JVgRNpnDxPSTJcw+ZQO3/Ejde8yb5gTmf
6bDKZvuDE9vRY0CEwJd3cnQRizgSdXy/ZAc95LOd711INsmr7homuEm+UNvS7ppp
1BR3/6tU++0+fNfKyfCsepnEYHu/ifwAzv1C1GZaw+QwQcmY6JjQOlsbuZHj5Q3/
6MWBX5P0vzm6ZKqoXL2oI9xP/QdHy4jur9zVjZCjCe2SsVNJ627rlsCeeBqyRDgj
FP0vquTkyCclajsfAZMqN9X6zwEIaW43yz/j0La1MIQ=
`protect END_PROTECTED
