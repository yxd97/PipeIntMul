`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ANb+P8ogh7UywfcuHQrUJfgHN6Y9zsUgFXjUFjiYbSHNh/aU8kRvCdfwL/oQ0Uhl
p+qm1FWfyFTTS8cHq3o/stpmZuDxTqsJL4IjUWN8ppw73r28HUD6yHEGktKCryYV
YTXwX43pP254YftlH2f70qqhGczTVhfvrEB2euPmmaVUleNWucEqchiDlP9UB8a8
VZo0G/c2by3NzVpFNOe/0Em2aTxBDOD7XdMf6mIrND/3MyGXu3s7+7IV6m4Ct1Lz
u7dihblMjSiJmOlvesXInoEcljOrD8gSuES9h1zxDgMWciUYGX5gFXjrsvXlw8jC
WX5w6dG6juXGuJ/FowGmMhxTyelh4jM+spuGIx0PGqybv/kuJBFhldnvVwDkM+g/
D/Pdj3bIp+g81EvL15G5ew==
`protect END_PROTECTED
