`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eoqxYMEwimhRqT6Dq12GLhij2C0hiamffTDlPoKy8B8c+6XHLoF6DTtgKHWpiIKM
h1xdM6fJFbSXBDl/a4giF0oUjRvVXtjPB5xTpPhQ8X/CvbQcvhZ9Nt8jS0ah41F7
s2+11DX4PIBplhPndL67yQtS53q/EA+Sj7yp8dng9SnqU5kY8cKjBKaxWT5gc103
FukAralxFDizyFc/1hivFdHOvuHxR4LY2YemyVO1d0/ZoL4h/oZYWSFbjWrbpY0B
Sde242Aph55ZuIjB/RvyjyGX+Nl59VDYa0QJLR4HsLz2jDCzjvXQ9l3fwSOPLtIr
TETtXWwXBPRuOa49oQ1xQPljoBh+YpsmbMDIf9SL0CV/SOclXnoYbKL4/U+Dp70D
uv9X88AuZ/pfschm++w3wrf5r9DS6joXBh9XOgCqV3n9BBBZb74BxaYUHRI/Boz0
zNVVnewFQCILkZVFhUdmLlyP0qXZhntVLvkPnrA4HTJc46hbqfSPCqTqrAvXPiVk
3FQ1tGfI7CvD1CZfOTrKt3Qc9rEigDfRGDPYQTXsH1C/nMJGV72yClv/OYqSERlJ
ViuESpSr2B2nt92C+oAnQ2gztlFUKaOJfYaD7PE9+IOrmdjkDcFXQeXluRO9CdW9
FP9eZZqjtyDGejyB3G8sS+31ReQa7LlyiX8il7HyiF0jjj6KUpOHQZh92uzBxZB5
8Qk0CLJ4IV13s7QbVMDI8w==
`protect END_PROTECTED
