`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dvkDgw+Xo6h56NVx0PvbMilRHGlyoqXLSZJk9pRQFj0S1AVAtUNcpJ3hahFoVk1x
bKH6smbOSevfAKv7kNug5P9z9czGnayKl+46skkALtOG0JYOaycflTIed38lMmeF
g1GNZI6uGh6pyPcUpvMnYxSwpZZPdf0khLBlv0ARQBtwe0vTObMaZhtQCCOsxmcH
5j0RA3b4qxQpcPmWEJiGLHddJRdIkqhU0bbFzU35gP6bpP/aLGjpdiDm1H8oKeHB
BscoohOba00ig2wWEgQ5G/dO7qdBUIZZQdFWkf/W3bVmUX3vlGY8WFtuDNAjcoxH
1EykkaIWmrHgLrIGnimWX3BN4bmpu4YACIZttHUMOPKT0GlD9oISsbXcOq0VbBo0
pKQzfknuyQa0tpPr8LAx7MJnA6yGVZFwDPTgY22clkrQ8AHNK3jFN7nOWRb6EOs4
DVqAh9uv6Bbsq6L/9jr8SSkaqAAxtbUsmtU8FnH+oM8QjKw9T6rLvQkv7/sVib6j
SFM+D98Q1/YOwAb/6wcsrKl6f4vK/yqxQwa85JhUH8pIEFbwG5xEu3GrpQEHX+gb
JqMmzOBr4meeA2qUSMctBRoOq1V2P7vIi5esSjwJc1iuf+/gBDXMxV+9Vvgah045
iDGylhXUiXTsvxnuT1M/kw==
`protect END_PROTECTED
