`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wU2AjeVCFHC/dH6QTDwol152J+Kk8hONqBOwH7CWw5C6mEuCgYBh0tZkdZTdQQf6
yrBm9BHqSF/0kmIeXAnsB3dF0+pQJdZt1i3QJRjCmc4XDYOSk0bI1z9WnxxPQ21c
1gNze0waXAePm8QWdcU8yDYqPsZmsJ9ZKV9je4jD2rq2+9tuAkgv7I9ghVn93oJn
22wInMbVmA9sogREhD7ualhvm2ix3QjAw2xpl8fohqk155VqJcvlklwtvlg098+1
r7hYXnwgM7ZZNqPJGz2eeZuk9xzkbluU17jW4KAfVzVRx24hGVn/5vE/k0DvRTkP
SjeWlKk8o5XjShHyQgOZaxgEyD55ff7UxDMXjKA3557ZSo39bACGBK7qtgiKRqB+
+QcBfup8bEG+PXpW6DIl3tmhV/4PvXk3wb2WOLmRR9RPeyMHwhhP1o48In9cNpp3
vZZWbxckSnZRBF0z2c3IIwsBlwmzeXhX3wXdNseFGrQTsY8t8M9ukdNM4s2WcQRN
OXT5IjmPC4SdR0YcoMYe+BoUzxpjl4zW6YyHQ635UBhnODl6C1QDrZo4yAiOaWQe
Nwk7boKbjCQVHXgh+1lK+saxTs3/ph6234p0Y9SAfQDsAs+ZlsnlUU/Kmhm9pP1/
z/BQIV/Wu4xhMYotLazx3DyKnMZC7aDo4R5sJnSJZ0RPZU/6INmb3vKQHbuugw4x
Fo62Gj0WQYFqVI8e6DYIxN71KEj/TTQ8cpzeW0x10XEXZVmlOtDVCngIGnD3Mtw5
CF1y+S3P0evQrPSnzI1h9vLZ4SPdwJ7Od87liDqDKyLXsdsFD8Abs/nweUSnFTkk
wiK2N91ac5EHPidmspiqovk2Uy283wU1/+MEhSqFi4694K94/jFPB6VG4PDq6FNi
3mpCffdXW4ihjAEsZ1OjMa2p6MXEQjm9t9iFqYbtw3tsASLLTIGrFX3R8dRywHkx
oWwphLweJoeaALip3O/7Vt6FSuZJrvbdz0peo1T/Na8eA30yrQNky6CIGw8iMkQx
52aUU3r0ZiNAANhOxA+pS9KLllxQ0nuvyRMB/utBA/8opwlQkbKl6T9bXOJdNkYB
VGeQC3cGcUUHjnKmNmmwbYYIjni2x+jBDK9SycAoj2dxYRx2snF6DSxif1coOmSV
tafnmvLABRcY3UPe9/huSgA1qIdEv5tZ3h/mVuFa3KZWdKDbS3rU+16GAFIQuqxa
czIwRwRb91aYu8fWpXINGtUYKh+VdyaskZj+8C/swdvaVfdcOj/+T2vmAYlcy9zE
hsCgDRlAWg86kl3+EbIxK/JLuBkSby8kHfOII0SuH6IUbss+sMkIebTBgvn25rgJ
MduQ++J7V6CKtru1mPPeQUZxiq6yXzj1hOVmIlDYiyu5e3IrPdgOUKlDBADqZG9K
4zAC7Bu8swstRB/fEAT/Fy8lAr9M8ChNqgCvhDJ9PRDoY98C/yQNB5bUoCBCyo8z
tz7qr9+4z1OGzA3eZUzavdl1LTnNtgOdYbmfbOfcnVDkMV08pxAXUeOn1Cs2ZKc+
DAp0VV1MznUCc8Gzv7CNYY8O9fO3t/6MhBIAqwUKDrTMAkWSqZhUskGtDkn/L88q
DfGzv277G9OZvp+81EuNSD0tQsLiVMD4CUR2BWDQXkQm+Y6UaC6gqgkbup0/Rz/z
jd11lLq4N3ukiTSz+SLFelrAnTWjmv2aot3K4LyimS+sFNUvfXd8RwbVIJQkRnzQ
R8PBfv2WhqbZxgcBeCO53PSPvbNkPi7abo88DOvqv298+HHUgXlRPGTen9sRvhdd
aJ1gK0Cgb+0O3m7UXhTl6r33FNYT8CWCDCinI7qdLwrF5QV9DmN8kam69SCq0Tui
`protect END_PROTECTED
