`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GmkU7hbposEDQ3ZlJfHVnfZlOvJWInxCZkN2bjPpQsPe0dReSyV+VBFesuywrXiS
xPQzFddOH1OuZ5DzFl/GhhxRKYXyByvkd1X00ufmZQkFmG3sD/GPo8tpsNfp8tJV
KNEfX946uTUr9RLAfKU1M6cL3IAjtZtf+zaHIpRZcriTXJFjQ5qFZquVtl4LpVlX
wGkGiC8rzRbM3G5/CK/WhoWpXcrH1E+kL75P8uvG9Krzw73HwPB3po8WrsNUZfri
JLsbiUDv9/8GJUuFRIvdHuLyUP2e/X/jKpn897kt8TNvQ0WwVAzxJv6BAdke3BLH
nMuSFWx/7wrsdhFLG4/enoSJ7wGlOba7hzUFrCZ8oTVhTVZFb9oGNXHjc/r4B/h7
gkhWniZcu8BYFxV8H44LcHphvRPWqMo8rtzaTSVQf3KWi4ZCFC6SJ4VaP0uxoPFi
N0/JwgxyYT+fcxaECmhPVfhxHXRvsLajNT4oYYZxprqFdTciWgFAwIGw5f8dspjB
z0y3xc6bksNGB5Qa37IFJJlHXJPA8jeBGEAIdMolhS9KOS8TyOBiFlC3UFtNLL6/
n9U8fTs2unwyydoTFDXta8MqaVXdjxA3iFl8CmgO/gHhZYF8e5B3WObKhI1bBJnc
Ow7JqAGtkxizACzU3I3JWarBLSE0uVGsyqkLAFgASNXMjL1szk/ev6FmkRFJYVzC
/7/stXVKkeRF58gAGpGaZDb2WpiYEPbmklAP9Bduv8qeJi+TXJe+b3u2U2YEc42j
kFhNGvYHQUe1uqZOWWDf3dmlRt3+5EAhQhJvhsfGvan3il5u/Qup44rjwtmDeb+i
3EtZoomdyThJ3JWJRpjXFbOuMt8WvcixZqttlKDq2cOdcG02eOzoeCBaXR2sSdXH
WfkIB+6Yijapnp1o+B5L+MNXHd1+A45TWrmVX1P+iVaoFcHBwuTGhTA7GxuUyTlD
CVcMzkSeITCcf2mQUxMmvoCGQbieLSlmkNAZL9N0OQKqLU9Iku3NDPH8752mEM33
rPykzKB6BSi4qpilEnfaOFSrWZeb2kh1HiCCGiVg8HdITTorzTBzLTOxWhzs76Np
jDbjY/riPyulEmVVN92jfYX0yzHgjwdrrCo/jJ5zL8W7xQstNokl7oTNgq+UYS0y
no1uF737FIjXM255UgDvLNwYHh3Hb0w1NNM0qqUABDRCkmbqTbEkAEH90d3ovPrL
RuT63xYFbHFv71eH81/M0wzacx03LN9ydmZy+xUEqzw0/oRYUyGAok64uZl1PfEH
`protect END_PROTECTED
