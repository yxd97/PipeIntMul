`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3NM1rkGWTPuxn3r46rWFaKLLjqYMICwVH+Dk63FUBEHz0JvI8cJpIRtjANXOf5p
6D+a3ci79DIdfdQhCJCBkm5B9fsQ5rUHvGKYx/FDN5pAYt03EU4cgMZib9i+SOhi
2Hb0BUSO+YKl1KWdBlzfeVQOHky7ztyu54zK0C6QE45thWxxIhhcG1S69pI+x5Ut
EIxUJ29AJt1d/iArVefIFA9fiFZ+fWSD5ajjtwCdwXl3IAyctlXiBssHz0rDOTmn
XyPOGsaAkE259hSOP9ht26FXWAQOK/9mtlVpJ+XMMahUhGa0l/uNBC8KiF0al/tv
LEqhP1sTPfcbhrz2w69vd5rnEMNBlSmUOCI4VE34fF5uOxjWsxK0rwa+XravRFZT
2dLG/bsmlT/mQXRogrpqztlni3AenxsoE66frNWaygii0HGuHXBI8Sd/sOsuYN8i
4E85i9ks6WyJA8No/NBWXiiJCWSB9Dz5HYQT7HFHvwrB5Jb/6EDsS21PmyzFDdtR
u4Jn3xyE7D2LEqKAiRJSa0rJBYmSSa7kZCAV8H2SlD1wquIg1DpiiFXSgNnGCmk2
QPtAm+vob5/xJaECMEetstJMESi2k5NtP4WyMiZghbJBlRZk5xzjaxwov3JunmnJ
`protect END_PROTECTED
