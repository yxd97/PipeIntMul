`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KkakU2I6dUyYYZbkzXHGFp/MQ3FBZNjIjwtob4NBhnX78pzrAGQK19YBkLMSfxVN
ARkdHzZelJRZ+d18KDU/S6SnrICdp01AMlsFLnKMbkzG/5Wt9VZuovWhsIY/4j+s
St4mUTQjru2xzdzFy6jpUWoVFWhgFULo2pdaEydXlz+tRn0bBZz0AoBqSWzlqBgO
kGxdjaa8p/ClK9RXtyMMnF6wvNi+aWtTIPNMPRtvN0Tb/bhK5ZcEzgFhl3x3GCgH
mpGBBUC3kMqWXAVaoLno0WVrc09lYkHzR84VjqPRSTz9XaLtA3V6RSWEMth8RyO7
py1Lhvc9Se7XA4qFG0XxuKlRYHkjAJCURBQQ/0ayvWro82KypPv01MucOKpI0+3C
6j82f5wShn2x3H2ZzOgLtxdQm+KHcOlZmmKsADPxRuhXCD9fco3IGiYtwGTSmkYf
aWaTLxVbYr/kOoV1l7iNTrR5gO0rQgQ2wFffhE4A24n2xPQsC94bR3hb6kSp4Ypz
Q2I16QZAzD7TRywMIxhZRwuXVckQFZVuKZEDkYruZZhSVWCnHrpCHuxR+Lc1Hnd2
hE/pWcyCj+muAsxyMScnUxGm4TFkEbe3teQTzefSniHquv7XBv8ieqXQVu+DmwrM
ygBW7p24EAr37unQV8/nDHMtOW3qs2GNXsA2BprWQ39Pij00cJWw5yKuISnf67le
hD1URmcsKqe8BTwzwyrFj8al3EjaHUpBgQzu7943MD73kKqsHtAIC3T+weMaOfvr
LVJ9gS68mJO0PD43pRO+G1/1z/R2HX1uH5f+bCehkw5og93JATf19gOJGoqUUsBO
lj2cO7Re6U29aOJNOkff/A==
`protect END_PROTECTED
