`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmlmenE6OqQ1lZ1Aw7dZqXrH/reQ5sUPPNb+cgfGlOIQAjRg7KbT5R2+zjToqh6e
lmbl+DJGGjIbv50Z9HaW/V7c6kqZ62seimvEPu/mfL3jv0swUt3WbHbVY0cpzjWm
hN+WGv2tRmGf0CMGXVCvIc7esVA6W3oOSfn9sOlO2yB5iNzynJIRhOFHozRzD6np
zK2/++7imrozDmTv4toDjqOInnUoUwBm9DLPr8s7FlF7MUE25hNSK0nzQ1wPQsju
+xiDRC8QalQ2UNHpQaQQavTAv9vsBg+ourRpIb9osb/A5NVLxFT89KJdiyBgb96a
roVRkrrh95p0ciHazg45yvSKN4lOXcbkHnxN7/hfI7viVZylOFKrmwhTXR4MLeJg
Kf5gve4BzP/dtTeryzrINdWZvoU6iksnuESHtl+bbNxHUd8bPPhxxFIH1cQ3Sh7O
C8cbkwtRXgD5q48e4hxuBI7Hr71IbabBkAiM25nrQXZbEuj22WMXdsIpIrFiYGVr
ZI2ctcJsGlNNTpAO4XOKWgBtF5oeNp8G7WB2Cjdiub12xbV+//y5GHkmlk8ortHU
7uQYeovCn77PBTWqqWKmlUdaWl/6Uc+KGWYvNTlBFOw=
`protect END_PROTECTED
