`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mf1RALQuYu50j5v05htpTAkNFsQ2+Otuwi/B+xWn0V5wzvfL03Qd8LrMMbyqmyJG
HYhFcyC9Lfr2NR2gCSkwGG2rJt+uioFGVfyLNWqfWP+tUHxWEGXhn8jmjJ1hJgBb
Ddtr3qxJ4rbGWIwV5asySqGHfJFkyJiq9/by5V13pQVCtFY54MGg/saZVvoG4f9s
iW3FQx2MLPHlL13o3oniNWPaBzLer0NUE5+y62L2xGSqgfIWo94dOeGAjzQ/nXAC
OrQ4q3nJi+PWFZVsZ72cLhBGmxcO6bwlN7PdTnPWrTeaQtM5uCeAidmNQ2hWxCvp
BhBid+JYDHyVCJNLwd4JOgXRYYmFoxlLbi/iDi5NvbS43zbfeLjKqK9uyBwTyAHh
cjpv8kYljBPkEx4rLFWEAmnaaZMMNehc8QUL75mtiNZcHoLwoV2fbQMN1g49JX2M
`protect END_PROTECTED
