`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fz+w29dqvD4wEk0lN/XJBwSFJjgN4WiunlI74Oaoi/8PM8pCxqtZxAhnk/gLcScH
A+j/aRdQyEwbcA7V9YXCWfXMNr5f2kXRs5oxcmzr6IWJZo+qqsev4C91E6U2OnQN
wUXrEFxRhY/vPOJY2hWzLMZ2gOOjPHc39an4+9d/5gsqS4y7cteFQtnTS1zPklHy
bF3twb7WySFlo3N8eCD3s3YJSyLUoBvyWrDq+D63SnrgqZoLhoagUXN5sNEUo2rg
nh7Hrj/WjMCHkBXk7MOvjkc/QyarB29pau9h5YdkhMYMQIcuMnz5dBlB/pxA8n4A
n+uMkCSQl/UfXarZBja5Ml819v9zfPichVjoqk9zQ6FtjC+Y3/GOur7Ht2axoVPe
uyWL6Zv+z6bjv6hzxy+yTAI032emv/hV4Tm7Mmuit4V9Gwe3nbQu2WTQnMSBzLnX
mO6/YCIlV9q+cr5yf0Z1SD0zDXLUa6sxNvR+i3SYyn6TWsfcB+GWbZCdyM8xpCEY
wTGqJu7+yFbRGIWItQaSEAo+vn4+/7fbGWDbBTQ0pKA=
`protect END_PROTECTED
