`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iSZ2V5dxJbLkiDYiLc+eNpBld70B2SF2wHxcpYOf9MXupAuIMuDH1Hx3nrrke6ch
h4UMmbJ3W4/SJ01nDnvwhPh+grlX4PnJNDlRhKH411yUcgKJ+hdO8P4rre44Rgpj
6m7Ev2LiOaDm2np1KJFzdbh6gpAiFRV+ztzB1Ewof1vdqoNIlzvdcXqQNxMXFxIR
B94H0/BhAFDndgDCQNPpY9D3AZuqvmyqJC08Px9pOJWliYBKpyIAolV12oIkkjlU
R6CxkZJI1aHthdh8Vxrxtg+YXBYDkCPENHdd9F5FMf0Nd7sZAG5Ub+Zg1pn8oIKF
efvb2o7pj1TDUSjaZTeJ5TQUBAG2HOhU9RSuECnhpsKsQYD1JXhTVOahpiWhsmcH
oFOKpEiRI/F2HM3vGVUInwRg18+2ikfjK2KLmUUywTL7SZTBAvfxGRUj0HiXyWCU
605/kBd/H0ahbwFhnmSRTKMAqeFZFpXjonnroLPhj+/XcmSjL7G3Pbzpvg15XsuR
/8Wx6uL6FC4R2mzkKRgdtl/vAPrMJVk2hvozeAxX0Po=
`protect END_PROTECTED
