`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jXWF0zoQ2zg/2sNAUXIT2WpaU8NLoGVlwghFVz1ns71V/D8IKjSpAZmObE3/MGnQ
wKaC4gAgRiDkfwc4ofFTrlK2c+qNuYhD907SFq0Z3hGsOLSBC/GyNYZi1BEKEk6F
jLpoN7AOxrB8EbLnHwp/ZocY+D2rK7xhNTeg+nolyTvW1O4+OIICz8VdPO1xCoFQ
vLJ5Fs5gR7Rb6dzZKnFhxTPB6UIzu0vrihI0Q2yl2uOpASbNWazx7sLaJWbJtbLJ
dLPeS31hjME08/NJM+yBkKbb0b3JHnkhcyVpGhtkpIQpGeROeTNElXWZsHLI/vbV
W6Mx6enQsZ+cIlb9hLEqhfhTZdC+ixXfn4DgQzIms4kXf/JTnH63lDHBTvAXme6U
`protect END_PROTECTED
