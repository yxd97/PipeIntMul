`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4jnv2FqCTjt8MatGLvD7RXJgQkA1OYaTX1IgmgWlxw6fR8E6/yJZpzdqIT3/dx1e
SbX5a7k1UJvLwOTzfTW4X9w1/m7FAkuJREDri1EKd68ttGvFbpWQasoKOuJITFHY
g1bT1/NwUzFOowuRMDx3xuSrSig1PH1p+ztWRkVIDf/XvEfLhcwTIY5ETPlLVstN
qFKwxwEIMzNZvTq0S8CilUyAeFeg1KFKiT2BJPWyX9ceJW7yX4jQMMHrPrARyNUX
l+9DQiZZJ6/emEN1tq1PfeRlOhNMxbdrvRmArniWDYHICr5Xp2v/8lJAvhN0qAeW
rPkcUSleYL1Wy/h1tnWGM0iPERSNVxaU1IFDHIjTWbIzHb1vf+TGwEO/6NuAlSTW
iWsokcKBoKQzb5IFUzC08UFQOL9Q/9AIZ7np3jrYWLJfgJoGgXcmTFzLkaeEFqyu
qJU9yUgWaw6P+bfpazWqChNYquFKMvsgfFUhKM4IMapm3hXjqYB2bJVXNmwDd3HO
`protect END_PROTECTED
