`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjuW+DaT/9i5vUt5GKQDqq1Qnuhm5gVTBXjEN5Z894FNAQcGf7Mm5Oofu3+ILd6u
Bgc/uau4w97tn/xQfB6ty9+q55CQI9oOW8Z0ZN7KiCfYyx5d7Evt0yjMGEa7YSOM
1cnu6skE4yM2pEGAAsIcasNcL9Awx2MAGtKzPnoy8kOJfgkMymzFHWBj0HDeTd/M
i6wXmZz8iBHDGE29voXKFGBB3IKE1k191fnw2wNMn41LC484epbDItpIQc+9UmHF
TSYKdeXPhkf4mx0FVa3P8jns77elzJKGFUzkRUdbN3URxnVdTS8YABYWBjvWcuDa
jFwo5TfDycviO6nAmMid6C+AtSBTKY+9WMdq7dSM6NIvZUJiDV9MztrFCeAbkJ43
bTF1C2JKfIo5LcK1NZsL5A8FrBm1gKeIKILI97TI1ONnj/NOJrX5G6w0rzOvVvXK
UJ0pBuqWLgRKC+cWWy8Q5ZtIYQfAuGG2/ThQh+q5nG8Ku6fn77Z6FoSr8yGGyHoT
S4uuSuWNob8c6r6Op3fsAfjOdgB+sNZio5pnHNZI3XLpQmDp4AsSszaiC2dU7eOE
Yi3eNSfL4XH0qhBtsUpSHC4n9mD1DSdDEEszTbHtPmaTx4rvk7A/Qh9gBjbTUMRH
8JEoY6xEQx/XtNWm7AodLBhak+d2F+5huFimNjZyu/0PlUXRGcVr7zyoVU1VtKm5
shWs/p1/qseFUtj3SWM2wz9sKZAdgftr4/P6OPJKL7/h/MchaLxKBS+tUQCeiui9
sxFJ/UxAgCotOu8Mx/5rNsweLVy4lnGbfmHbOEk/jfkAr90mUsVn4zjUwUKk7Nv8
1Cs2Pwcw8Ej7MEpONZUuJ2MaaOgLeMN0hqvezrlovInk+IkmC41Sr+X/+UB61bIC
BiMK68XT/ISyFB2zJLEXmrZs4xwNZQX8D3k5EG5RDPq/CsbF5hCBi+6plUZF4ET+
bkAXx8blAvH3QJM6OvqZibwpnn92FDdqyrlcDRX5f93t7A/n5dz03XLs6lPlRvs3
a4vLdhI2Tw14Jwddzm1oTwmJTdY0KIw7j40cAbglhabUvj1iAW+YD/FcLzoHiYfb
YkN07Xk0/vMBzZWeO7S3tYODVK9F/kjdf4CPOPOSPApjAHTQmmZpOIt0uU+00vye
4Y1U+kf8VjQtFj2mwAWQRNsjIIunpWPzlHFtd872iTO6VTuspqMetyx9DbkC9R+H
r7yZ9+5H41HnLfDR2/l062MmV7qSwmplXUKNn17s/DT/oOr4ukG1gq/ANTb8eYHP
h4UxPTIuN6nIwU0L0KoJbGJdQLlBMnz7IwIwIi3G5EfvGiCYyGwaOyXDNLvywoyR
wHTy0D4aUexgFaqubveCyGrlrQcMxvFoXL0M+fbyVUG0Ni1e8KcW7vXAiRIu+TQb
MNWc0VNVYysVDH7GVchqSJJWFPoIl03fLQSs3PDSqXomdov4feTHcn2BF+IGyBhq
QTHVR0MyevWZgLAe8a9LJD8rUpS40pY3Ih8OGjvdST/23K5WTCmAAs1VqMY9h3ph
kvUK8HRXOb+9Cl80PXxdQhmjuR4yR07JlTD/ckB1klhQSg9362+CCuB5rd8m3qN3
TLJYJ3CArJ8vvz7JQn49TYT7LFyJlN68Pl270DKIWpVr2cxQv3bYYYIHwOrMHsNQ
hLrBY5lLjXL/rh0ncZ7odWheb4xPhBFB9OW6CHRxJmtW7YE16yVPgaevfP0hlSqc
rKwz0LPvZAGZ1eRj6OU104I7H8XGY3uyOcirlpSFexm/8ZnEJx4AuHK33/6tk2fH
2s2FBDqDPxcUMDVrIMoE4AXBnNP0kb8Zw6uzTJxTX14bCZ4Vf43i5bI3WYyD1QyY
DQfycwfmikXlzoi7dMZnUZAQS0CZnc9Id+viTxdFrZ3pPMcLCvDxtfCYqe4tCgj5
h2vOMHasUYUxbDhxa/X4nZOtVb06hMKmqVswdcqHBT63E2o9eAYsCfZP2zV2UdoZ
Wh2TT40MXHpX/eu+Svy8PBKq/hT7iziBbMSn3ECXuztgiZaPCwZNcdjZwnkJSHuN
gAJ62FehRc/JZyAhzdu91r0wURRwwQ3kGXtU5Ygoen6VRi4d619UuLE47UXshiYs
eojmsGplu5weOZ6Gq84aZDCSoL9WjDsPFGgrifMKDT047Dx/FhgpIW8Vd/M3rY1/
wT9RwuyLlnTr9Fex3Isx6Z1iPZHpVxXR9yvKkj+M/4tHAtBDEqoVURo64+hgVqF6
/ft0d/5wDJSJ+qxDlmSJzK+WRQbIRgCgKrSoZwvPuG9Vg82Phwy4hso6WWDDg87f
nEujo3BMvbiOmBKz1qGaIdAOAZQ9wTOUe7sdT0VCFLHmjUtFlATfzHFW8PzAkrfI
nj89ALcKP/jfipflTAcvV8An+UV5sEY3cB8zCr81Tpk4Ptg9n4HGud3lln8Pkxpw
aVD3sELlbkss/Xb5ki8Dd7awRM4ukIozA9vmqtcDN3BK6AC/9fFCwaTBtxp1oOtM
ZIlsHZ5Ad2FetMGM/p7aKqyYI2GnMdMh8BUmxmz7ThZh5AYmeo5UE/nolS/pC1Jt
vPdrOla4FtAckwzWrr9PMERYrmreDbXTqh9ssnitulQlqrFSnOnluqsFaBKYMnd9
WZz2sIIhVPdhIyWkAetjg+VGxEJaVKUoREspke6lldKZkec8WXT6KvT5ix6j9zMe
GOwIdYv1/OrlKPmf7sdqu8brvECSJ0IhYh3HUXujKY9F47awPALXlDNHDrfpnBDe
ym6z44AdgYLd00cObiF0oj0kL+a81RdBjqZqmdn/uLe0sACGh1oqVy/SwkF2Y4wE
3lXMZg1oX0iVKEIphKCTf5ceGwQC3X3iIMlmRAz/lJaoZOeQ/hvwhf93aTH466P4
6DngCLuddTNYLxuLT+4ThLyYbDFXXaPpGtelxqn/yaDo4t/Gb/DI3A2ZCdQWrqwS
aAnMtKqlljw39GnQDhTHyVRveTsckb61C130mB1f/5WU0O5yPac+kO/OA+sv40qs
VUU17S05KWMNbDbhl8H3hyc0+elz1ojZgRWuMOQpW1vD+Z5b0NyP68gD1XXE66Ks
PbrLXpIxGdrDSsjwWYI8JxmKS3CHVZP1qEjcnRd2VTs47EXmt5QF79TRHjU1qpXj
rRyo10NnJKqPA0Ntanv8iINUI6UAX7cHESQvf02Tt39+Fcza5w0kjSurILr8Kn6P
yJYR92d08o0rtnr13LLeF8/XDMlvcX70d77i3dYvtYFUQzKCrCvhZrU4pjFJ/Wj0
fMq70K9YRL2UKBhibS2VCKgTZjE45fjCVa7BsD6bM1cwSZaN8LteuovCuMaN0yLc
W5Nna3v8nrOf3wGf/JpF1O43LDzHBAENjaqD5Maa8yRe/wrzC7bC4y9wYXlTx2mO
tf8JPKKVtE0r8pKoQsO9KV10LdSBtSLO2oSXk2s2JExu1hLqJVa/pn9AFiPgcSu2
MfLbgokyo5P1I2EAKoDvHiTEm2Rllpt1FvlSJO3f9lFlnc0PGkIfzlbKKiN7BalT
IqalTY1ez4cRzye+ank3dqaPY5KXZyuQIB36PIrAIBOX53iFoa0fB+o6jF215Ojj
YmDolaTYK3vGj3wckHAp0/FeKw6oyn0gD7w2WngEUNui4J95FjkAs1rmR/GBZ4BH
JMWgIWt/rMUirlhlIaO/mFw8npXcd1YDyRLqC3j5wI+4/uSnXrlhfTjBkVuCmHUt
XdJVorG3rt1iYJtoT0R+XbuQgJ+tjacay5WW7V07z7py/6oQZ9/YDPr4irTaQp4e
i/NDzMP6lnzbSntIeSZZC1kNMDCaae+KnaLN3zfQSlu1MMXPY/9eNEvkOYZdY6CJ
g0k+d88BH3I4CdBDrW/K6rs6Ye21dj0b3r5qWDb6WR7PDoPO1vWPTl1Qb9kXJbFj
Crt8V18Z8Pnarifw7wCJEkeGinkBS3d7La5xRv9V3ao+oIDxAQOjT2e3LxU4Iabf
aP8IDopf1B8XPx3o/E2F9bvovr4AmrxloYqgzjNGOttfLab321IZdVjmnHVlemUX
PXXkz/FOayTu5wYn1lWLCCP7CpnvMGq8dKyK3ikYZzllIRzTz5W7J9Ayn0SLVLA/
4mTEpgPkyGygvMeqyCKyJieDTc9iSfNHwfDgkktUbD6FRk8euLkUGEkQ6eCb6FFa
KkC+KcU24CqcgabmC757A5Vm/lANdsQos9h8YIRVkqwx0I6DrHTFEf4PrrUkEw++
SC7ORWf7Rk4y5j+cqNNXtJiBS/Y3NCqzyFcBARq3AZ18Vs83dEf8GKc8M02edrDH
tjXMnJ7SDyrde0OXOp8OFv66TQy/9cuBv5mBfJwTduAfzo/of84tYfY8i70e2+ug
NtOz4E2t8DJnTLgj3nloQEtDltBHQjpI3sM74DbGHirlggZ7WVV0Ik2+1zQq3EjE
0pZZ2VcdncMifsIWzYTEL3cFpFxSVhKzw8/gxTMOagntKyHYDX8neVWd9Z5SlNwz
9c9tVwkKv1NvgAaG3kPp65X74XDQijUQZHjKuJZEB3gqp37S0w0I3KX878sMjI3m
rspl7kzGrOax7OcFgNHfFmVdpSLY/+WnzEaX/x9a42EQu0G49ZAsjB/qOjB5roor
UUJQKnVbhsCykdMfMxcRXNA/pWlyJJR3Vu+DBNSnGjGH50w+6MnWwY8a2r94tR15
/6hI/b8GcGZUTodMKDyKcvdVuspLE3bZH9mQpQYrI22Tz0Myby8+Yqxk46rVLIF2
7/XYqnbybsBtbB7S8lOolimNEaRLgKjVgKFZ30ilStsW2gkVHlsSn7dyS47FNUBW
Er758/OjPeecs8OYR1CcK5Rhsda1dXGNQ9fjGYr+s7e2vuceE0fF0ydOZbsyaK1n
9VgifcXrfaqXPcKvRWPNV7+5/FG/qeG9IqkIn0ZlPRCdBThVPRe7aByBsZMCNvwP
RAzJ6N/MJUVMkKg73eO4GbuHQ4WJcg01DtA81fDvFRprPhLo7bcm5LkdoPK+y2WQ
esaHrRE01MxNbDYtwK42GYf4K9qxvxQbfmMIpa/TC8yIKOS3m829gW5R5ezZpVvm
8BR9QYt6tEWmy58mpNhn+rccuTSIWD5b7z4UWwBnmxsvB8NnUntHi8UpGD/5AcSa
ABGgbgadxrlOh2d1gn4o43U/VSPf52EpaHRrDu04MYzla/BIm3qEaL0s2qKXUWFv
egQWkMTd7vKksO9jizYmMDFWQgZ+8lD/V77DOsF9uL6Bd2G7ZFRiZ9/GmsM3w8qI
/TRbNhnC1Gt0lpYXXNdYOQOWOEY/04DhSct7j/1juIq2jktOjjDyjEc2bpzw6V/F
xM6/0hb4/vKDFLW9P4S1y6+V1UAKxFj6gX7z9wVbjOFKe+0JehdyWtbeZ2johf1S
vC8/5ikqm3LTcXEdBnn0cehbMunql+oWIrJnxhFSNXFQYIcnuOyKmExaiQ7v0EIt
1xIWg730klMyFRbSoJ/VVc+IAdYJmbraU9PtOgVIzsu2LtHDjsGUI7N/afKYCrEH
ibijmDZevlskqCqPmgmTYLuqnQghQALAXcLtvq28Au2/ddqG4KdsMUmqz3WP69ce
mQIOcyyPAtJub3lX1Vqpg4N+QI1PdZE23Te13PBCe/+8fLY2vvT+PbmrxEbA0jnP
ahIEB3QwumDJ0fr6SVxfJoPEUP4u7o00uo9a+itI2UMBun0WOvA7hq2nIqZR+8BS
3znTlPf9bTQwbw+U/1fM7Q62lf7uM8N6UCRkrg02VU1QZCKbix0rTv6gx1wxQ3sD
V8WY0VEGuunfiXncMRESrvUYcc1cgiQXo/IDWiB++RT/qYD96KGixSlettOzYitY
3xgbop+rRufx+bdbmUhv9JP9IDQ+8/cVIUOrgGPtim5q3fyE2/TeExgljgOUaQjj
aG9pylNx2XPZsp+zK1FoLlw2J/rS4w1MpPUXPA0Ejc2Mo+1pkVVrjLKh1SzbsgaH
vSJrXnE535yk6HCYJdiAKsbhZQUdAxFH8VriKJbiZCq2catgjCCAcQjTjdojQPfT
70MbdrupbrhhDQsNyv9F+hc3BKLzvBSZ2Aop6NEiaRafr/uS1bubJqAB9dzBQAmI
DQZb9FbSWhvRG7Damve1zFEAv2ts3XDCqaHiXiSYWN9PUY/JLAUZAS/pwbj2sBXl
GZuVQq7eLVpdFF5WbekFFseirSETfkTF0O/vdBEJ6yLz+oEv0OijKtPGcsUOVFnF
9Ar7Dmyqmlr1PT0Hl6f19qlSkDjkjqNAcee59Rc0WqpSpSMhOl9NxmxXNracR+bQ
FKy1ca9DN06DAwY90sz80aL1MobiM246YPgM+Ez5z+deidMJx06mdwnl9wzkyAAK
xxBuaHPzvyR4ZFk4Illc5ka/cgPKfutCGzVcjMy7bL0UMr6fpMB60MeMRlB0JtjJ
oX/H1UfdlHQm3XAnGUyykF2PGqzSHYiU2HS+Zc8mV7fVLbsz5Li0Aw9HP9G326UH
wf/caeoi8V+vOWbIlZLiJi1wCWN0v/ffQIF79ItnbMt/XXIjlkjvQtaRG6bU6pup
77EsriBnpIoacLgUO4zjnaBRfjZApawY3P6hO84JO9mx/+sI4fU5GgyK1BU4mdnm
c0ec4GN+5iCWB2ExVXGi2n7XG74+QgWRIxUjhg2XkSy9FZYLkce9Z4czWXo42NDU
SrCZWnw7npJReGe2ysK9ZvVCU8hrAjRF1/q9khJjoUHPuOqjUSovAyYkH9GyQaKn
fnV0bEId/vQ0Lo2liDVIA3dC1/Kq426wZf9QsA21+1LWI3xfG04R+qOHO5GOXBrT
9O4GcmnzAVeORquf4F/mGH46utM3/zBQ2g9OTHe5TOR5CtBSNc56ueZr2d/QL2U0
MTyW/Z1VY6W8ZEAAcT3md/8lqcuw40croXye2dWvK/17jUeWnm12MezO6r3VR5Lg
X2eAFsamBuXUlR5xqAdY6yqHzENBLsFXkAnWSHVV7XC/1LhatCZpDn0ssG7Q1wht
rF7licRp6f/+HFngqdzTaEAevIvGx/Nk+JDXTpcwTOYdIKUUgnaG1ugRoKv9OPMq
eCXtM1rgLSQqDxcHTHSppm/0eWxl6ATLT2r9dfAUSqqzTSd6B035nZtr6QkSTR+p
5COjHVu8EcstRmgah3AAkV2Mmn19I+8PsP3oleSZ5axWtHrMVy1flek68apt3fzc
+yBEEBY7/z6iCnddOxupY9NG6GrDrVYL1BcBWfDsOd+pHWykxiIsPBeUmKdJQhMp
5Fv2/PLzDJI8lhXdKmDYQkk88+hcOs+d27Qe0sQlVEfMqJnmS7011dQJhxt9s24+
9FLmH3Ye/5jEp4Cp+FSJdNYWurnd2wSxMJRlEAMTZSzIAArlaq8K4vXGnXnDVny8
N5ao3GeRMKXB4db5utM0pIw0sH3U6VPFQEyiMF9xq69fDQCPFUcosvpClzpVNhFn
01j7k8HN0O0Bl+H3mqH6SuQqP52zULL1UhbeRP/zOkgjNPsKMBsOYIIwEUnQQxOo
IqVTlAqU5zHtI6ftLoENJ28eCajKP0nmOZsv4SDZH08YbI46Aqyk08SQZzMTwpYi
fMqUvNZz/1vedG9cTjRyc2tjHHcWH4kX7sHP5Qh0dXzd67WM2RzkDubpbemna1yg
tfksXkSuf3232npmBQJHDarLCgNwyPR6z5LN671OTrT7TXg2CaRFLjSrmyOOxwQZ
9rwSV6Gue2j+a6K1A/Mt2ft1JJdXNZlllfBM/hUDoj5uA7V718WAjiXzObQVj4JC
eVwutheo/MV/7o60QC2/vnApLz54xED3zoaIBBgt0Q01ZgcjS+yso0ZfBdO9PQx/
Vyk/6zzuHRPWrDo1A4QYdEWs1ggIBaMkHD2D1FmbIhDWISV57lL8gL7Cg1hxmflz
oKCWKo29OJlv/5WzSfHbuiPpiksNlBnOjgGUcKQUfBIRCXUFOtOwMRY6zFANuBDL
N5bbrtEPh15VNTx2kRoJm7nN9hxxrfrU8vZeuxIw2YlDb0DC0C7XMuLPVJ8Zhy5h
4izj7zTAZZ+YWxtkNf8Qr1yTDxH4jiBP2VZEMo/5ou9gHYahmpLqjS7sNIlexCa1
B+E+UOLM6yw+q2c8ZvhXI8SjHcQ+Oowb9ntAH7i2BzyRUKzslKcVaoZurF+wX0Ps
DH0YA6n8snjasbpJu5rEFpftdYuLMNjmkv/FpSo+qXOToRSfT5y8zIvOuxvQXX27
xOY0xyjGCeEtqiNRM+uh8b3RZs4Yj5NFIW33LE41pCeljbclX79O7L8cldgkOba7
fq+8mr5YhW/gbnQ53Tn1RrIOo6jTu3932FaY1xtF0Yy/HDk7RMsffwHWNhqmJxSD
dbo4uq83SER0Pb1DNRU1FtQ7KIzRtMbzHAuiq8g7+9n9dAyeU1ZUxZoYSHXGsIs5
i0BhH8cSma+Gq5VAH7i6rOgYahr3mIicVboDFhJ0T/hcqqYxoGHzBWnh0C3idMhT
YVyYrbdNKgkS3VesY2WJ0qpOeFz6czibjCY4QDmeLilfOytsYOyZutjvNzRzB+QM
wFaVWJiyv/y7B/akH6pwsKtp4a5ZKH833uRTbxsauSIpL82vC/nRlcoFtlrnFGFI
3So688IWxuX/BhVaSRv0F+yNuyheD5x2qr0kVWceN5Rb3CPWGDFRbdT1OTJ/7WeA
IoY+7nJeErTl6xEjDYpOG+bZTnA+sgk2Ts7LH70F94nSEBR2ZLEyEHv9gSMkvWs9
SlYgxqkkcChs+D7eO98cDj0c1hh7iHa7lguyPB+epjJAbilw+MmC1t/NnerBghOj
HtkJdt3bgCW1DfL4vNHqUqV9Ex/nbASY9RNSWdRVop1oOszytsmRq83vpiRiqEob
0vKlgTdDpVR0aA0o/x6uEwmJEcppAWK6eHaZgppUZft61JdnIdYOiblFrSI2OKK6
QZoAE8VziCejxYHKY7sgTjARSywdrY3pIEGKwjURjpePhoUsBZOr8s9m/1/YX4de
rh9dOmht+Fb+bt83LJ/J/oKqpFBweOiIUNXfDun7CPzKsJu/aTtWnC03am3lTxYQ
cT9akdzrXYH2wk4kcb2KkXRBL/UR8GGE32CHHbbjuz7Fspzs7QNt0irirYJy1Jl3
ntsnt+xXzP+eqAPjDTfNoc9a2IG6AJ3MOj/wwMnZyqw0/UZDh3YnUOVJDtYzH0yn
RbNJZ8E2KdXD4oybyjCmiySsao9bWorNi8VDI61npwwjOvWdGCk5C/ng9OIb/xTS
Fq62kAvIqqRiUhkaVopXgoAuw0CUmNklwPZaG/GLtlAji8PH0Aa185tL08Ymo0Kz
mce/b/jNZkU5pksdGeY5zHattP2P4ShS94HvMdaBNAtyYQVQ9esd38BHz4xwznH3
gBWlXyy6QU5tzhBkYdUmrO7wTOhQrpeok5AWtfvwUT5fMoQaHDUtIFot4B1rahV1
UexViFnS56rhCT4EzmNpIcP71gozqbDPhw0u2fKC7ettsDKWmjfQX2pXCA2Ney2w
emUsWqsqaOjmBAIHd6X80pVfn/cZNXG3dQ6uri3vew5YnZat07DmIjOdK2M2LlH/
g2Md8JjHt4ILFnMjNbUuvmRupke33k47XqhBo3ZwiPktBUcxoRaIYvlHmYFVnRU8
cxM6Pqg5/fL1iTMcvKIsioDjTwSPYHOhe8U1I7uo1W8L8s0cqnAGoW7MXzK33jJc
RUf2EXaIhN+7qD7wk1QO5BLFeYOSw+hIERw0yYu0Qg3cL5jbCBdB/3rqnfkHG7PL
j6MFnm7nWC67AbzHuzMGyplPszZBRhD8Wxvvj23F68jd442LcJ2Id6nPCUIRvLK9
4clLHXSM8CG2iI5H4q1YP2301qAQsW1eSbYNOs929vFhL16Kg2NLwkYoui8g2uFQ
aTiQ8v8NSkLnyTaJQQ32vJ3AktAF8SuCrk7wrm7fdQCBOdkJNMw+2APbPDd44Gr/
WZ/6Tk97yfIBJHp6kU+bLMEvittJeR+EVSlTVExSR5HO9t5MBHwbeui+bL4PRJEC
ZfUDeln2wUUBYRlmmUTqa76AnQ8imud7JOWuR+hE+YOJcMO4OF1beAwN/S2KWGV3
Y6GPbHhQESc/wA5EVRyv6jPZ0zzCm9FVSuk/mgInVtuZ0HISHLd+EhgZ3MYeF8fH
6mwzzVQ3SO9LVQUyJQ0f7KfVvp8CVfIsTkjb5z/1RPuYZC3QEwdhQYTE7WXTlaFX
KisOPqRrwTn+MVHDdiSX2bSWPUb+cwYwRXQtfjv9FPr8hqQKp39pfotwBJMbow5b
z0oauwtfTpR/qtMF1+4Ra16QdtFvVtbje2gBDlD4glnnYENnxDkCKn7Ys0g1+UKM
kKkdsWfI/T/OS/QqR14Un6ipIYqu/KulPala1GOYVzgDQ6L0SP9HCEIwFw7+gce8
aWcsDrOgRi8ZqfY2qvJXxnNQfbQtO4vhQEPyUkE5MbB/hWdsIu9qgxGAnrp2T10r
OHgsvb6s7uTaGXtWtX+4x9xJL4d5tSEqKWkMd/cYJikbgBWdcfC54hrGoJLLrGTd
Utj3EGMW8iZS/H4JHL1yAwyJ7yOI/7pgvhUFdNAVzvsqQ6yo6GQp2/pCYwE8OdOo
ojjo8UiUzeKDBqNU2fJAl3RQws8ABs9r3FiJNB67X3wk/DrR9+bXQ9H6n+kevyVn
RZOWnXWjesGE7J92JYwaVX9flde1bUlGMYjyLAKAAGfzA9fwu1rvxG1qKiHPcSXs
f8g7D4YCVwRdKpEeHVnL+4hOnHN6OjY+a19tH5Z6Dxcrx5kQ09cZsKIzG/GFbbBg
0a6spw8JYhmK6Whyx8plgvaPFSZafz5byGerMia8ffPsnA/CtJHEcwoOWVN5ZNWw
nF93p76zW1k7YhOuSXjyoKVWe8YnXd5jD045hFfveHOjOrYfz30VRdPvXk5a/70w
JKwBJZWhe7TEpi4vJ+fk+9m1b6h9SqnVC9vPtS53STma0P9cokp9KRuX0cv5qQ/B
57t4ABhx8a4EPWIuf1pqyFD3x5wBJaYroFVrDlP7ChXP/tnWlBpGv2PdHC+WVpOW
NtVvIqGUzN005fFqljUPqMqBsd8QqcLECw1LVQJaMerLwmictoq36Qh1ibbq31yT
H7zlcqKeDcs6QIuXBE/NXbkHQIMV2WKwZO45pwoUa9Hs+K/9j5tgggm/7NER5fcw
bPg5AEI0IhApIA7l2VnIMK+ng//zx5vTP0/BWttBu/8ZxhTu0w1yhsbJfSolphDY
EZMlahwQRlx5Ew7Quvx7nQaMu7mVJzVRdtZrasw4j4aY9lqztQWvJ2aEu86iCxOx
qH7QwxdMD2EGLDouNhI0Y/WwoNDHqqb5E+a9tEqdWs2mDKP95XaoQ3535Wpc7XfB
DkY/YATuI++xzZNUVOqJYP00RMtBqx/yv5dxKJ7PTrUzqd1EN07/2eDRJEpFIpbA
0D5PtO5vSXEIbahDKZNRNmDit4MOJlL/UmuRM27IT2Q1c0thzymME+12x2nM+0x5
KnH5QGooozwKiixLE0a5Exgc8SL2up4zNjy8Vqof7ZvBiRGZ3hPOcZqRZ60BQKt7
37urhmrpWv2b8ceWAQkjHu2T/TQIOETKm+KtnxdzWaC+7/+QjDuKiL/UaqGSfqvT
jUTO7w7JwfWwE70Ffp4z1Bsd06rQU1HrgCYi7aE7XtxXcl6YdSA+dlZKlmqAUX9I
wRtz43BBFIrHDgFfLTB4inKjqQ7nhkQnSRb1HQ1ItE2GdsQ9Ji0Rhax+9sk2VRZt
tPy3o1toN4HbVvtq88aGxzpIN1IKnfrwDNLtNJe/xdUCyp01nNOpb0Kj4+KieT0J
b6S3cIMh/XBf5FodAi2E7wxRucdUC0mHGvAjD5vR+++qFi8ruF2y90MUV1r6wtdR
6DdmWoviQQqiZacs2SHCck8bngWiaxSCRecs/g5d6l/p7xPAblc4vypWvU4ZFg8/
UDvfpY9J+Y7r/fNkdT5SIzLELNshaKrH4W9jOvc3nBPmnPcERR9qERR6HGyDYaNq
iSGTtWHAMSsRhjjs00/aqMf49p1hv5YekqJgVYN9AISlEeabucqe5cp0XafEGV6Y
QJhlMK8ZeyU4lc5cmQBCsO19lMhLYd9mwR7r6rGHsEAb4AXoKfZkzI35het1DrED
akDbaE42e0Zyj/BaW0GdXXAhz0ecxbXc4q2U1dsBOsO3n/8rGP0r8vy2W2/QjCyw
I3xUKBfKAEvGE+wEyRrT4zLhVxV03L/zmtY71kfVGvF9zezWpU1k/t7wi2dd9Yid
vOV6xt4Tl3BtB8m5UggJulIctZpNvM05+HD2RQUMSXp7XetHr265UyL07k+KbVGa
+xh5IoMOU3wOgxm4JFxd481T8wEYdknf8u9KhsuNpQmPBPEHzUGEae9eLQj0ej0n
Td4mPylGbj95Q7Thac3/VoKHkNpeT6MZSma640xdYK1US3xL4k2Gar1QMvNjIqzy
3qbNFvK3IykfrMehPvzwlncQnS5vgJFKajAe/BDnkCxuS05TycvDbNP6JS8zwXKy
h9/UDBIJOoh78HK0ZAwlvszkn7qxX8tLXHSUldjQbCZWJvtV72V8006c5+63fQlS
1StjFj3NrTmj+2+sdJEO+5tg+pglR314ZLVmLFyRzJjtCn7uRG46sJPodgKrs+lQ
aqeIynBuAJdi03p4yAxvrXdgygcRcxmpffqvby7NasHUAWtrQsf4DrQ/QJOPuMak
B8b20MXsrrAEEKC1vfgfqP6e8ZSn5oHkqhW9EeDG7fpc+N5+dp8Ocb8YSkqEudPJ
j95RU6Log5C2FBskK9erWAr2lXXMf7WT+VifVwhTBeeWDlF/5kYZqPRG7zUrFBrY
sojGD8f1IpvDMJQ69Rw48N7hU9ImaWnAPN6qYxR6L5fgzw3peNRiZgOsf1yNqPi6
ev3Pmee3kU2YDs2l1Yl+sAhXZN+T4wA+ahRSAGrQ1tInh1osZBgxDZpTN7fBDNH3
Pw/+5RK/dLsdccxXAvYNUa3l03Ap8GQz2Y1RSVuO3Rk6sjrtKjx51i1tvbZND26B
ZCi97+sJLMXXc7DTFd1GKPYkJShxaCV3/UiPpdD9Efm0ByYYdpr9+SEbPG4xyS0Y
T6wezoxnaQYzfPOUZDN122m03uJ0ltgQYjoOmz8XhUvBDed1hbHoDoxuJnBXjol2
4SC8OoaHBy4Kt2qnY5XWRkh3S9Gcum3CTpYNZY9WM12T6dfmqJAlLWxMnD+k5A7i
2kFrM7MOxXwiOVVUXRWh6qZ+msiglwTa00bhkKHWR8r0Gmo8SOh7J0+8LaRZ9UOC
CMAEDXSEmwL18j55Szzum73rRWP9J+Ce4zF0JseQ+RkrQadQb72xSWAzBB58c9R/
fS6DmHN/VNb2tEAL3+hrSTXcev4DxH3QkpwogP4FJAQEQgMeF5MnBx9UlqmvI48k
TDlhG95GlhM1VdepuAahHoSpLmotyaGKdp/FguXyrzcMboPVlcTyswqb3Kdk9qAD
NZNGqj0y+evZrrbNWEwI4W5wi9c3oqytvbZ1TtFV3IfMFjYBWNkcMOM3meq+QKJz
+pCFU8onPWXsqPtNkUfdQ845GJvT39ouzO8VL/E1m177AS4BgZoVHMFH/bNvhtW2
alWzrcLGP6kR/HZxobr8/pLccpzzr/PBg4MJU/qkZAqJlddNXQuzA9FzQoPJSQcZ
nTnFdhO5k01XGJJDFHM4CZP2B++CGYcADL3iAeMiP+hdV0ylXS9B9Yo+RM5LMflU
EZfmqpr+EOQ9/YGiXtq5BPfaW4U7QWdNAbGuYtu+w6pot0BjjLYI4Fp0LFZ2xP/L
iD4R6Z64fkrdrTSCYFdp5dBGazT8H3zMeqp37VuohIne4mBOs3g1Cu9gV5Sf4P4c
z8/KH1VtTgn2xAgRDImZsbjgvGbwH2csAIIcUZE891GFIDhX92iHStlkXHiHxflb
Z3WdGi0nGoai5f1aWiP1T5moKXWjvaXVmr0V9sa+CDObcjIfPBug8luKJ0/x3z03
6bNCJ3bU01xNu0471+aYqdSxwdOXex6lqqiz2l6g21Qy0SjGjQ4qsT3QQ/4JxQme
n3rJwxTz3bFH8Mc0ClxLZ3IGKGZxD/XI0kW2fYtNUpSXW9gMw7mf8bUTlXzp5Kxc
FIuj4zXyhXuuw2YW/G4zY5pLPJCVaQ7agAOdj3XF4w5+FZAp1VD9evAjKB2UEpA5
xWDUgQnNPUrP8kV335M7mlRUKd+wHoc1ltCCOQYj8lLjMiapYa+KefH4enMdUSLI
/mB22c61GSTxnsPEjLoXNU1uMlt2NBu08gH6QMHwa6kaoX5Y6Z4PtJ3ga7ti13Ni
rpx72XFI60xILHuB7jSoEaOauN2CYaaHBane64ltXIqyuYI6fRKT6cn57WMFXAG/
d0vavWhS9Zr9+Ft/AtXLQD7ApkiGeuMvxNW5/MOY+56kV72Bfqa9NnpooxYbKcCo
MkswM28jkysp5twhlCdsa3wuXcDdmK6DNFHhacChdUY+0OcgwpHiSky6hDRYTnmV
jYLQ52v5BlEmEUx4Uncddaq4W3JKB1zfbFzNAlL23IQ6PCFZZuYxhf2Tfun+EfPG
yTfAqnvPLOh6yULPt6koPAgdGSh8+Y79/2Qgqsa2FrwzO3DwZzIS+wzRLcP/6nn7
UWnreMxaZm9gIuKagKeTyCwh88qD15vwFnTqwbCkIDUpK/KWkeFxhUK478+B98Wy
BfKGhmgN26au7Reu4l6FwauoMpjIsH6/3DXmTTXTDobr+bSeb4/bBtH91GnS30Ry
2HZcfh+6ri7pzO8AL4ygHEJsqdCMJPGeiDzjZqSO8qxuDPSGLEe4ARzfxUwPJ7CE
1xtu0lkYVJrE1KLCWZt0aS9ToSUQJF5cN9jaBwZ2V7QPBdAEDh1nFATfDX/NP4PZ
xesd/1kYD3AT7XOwL8OJI8lkEcUuhHbgPbPReHOrAAPZpFQmjK8xjWPLcnwL5huI
KV+aKEVSicY5+bt2STQFL14mrNJDNu6snfGOF2xlfbSYx+yyr7NWgYiA83LOJxie
iSYhvMKCxWLLeHIhLxv/Cos0+6VJhOVYldSd03hn8TGfhh25dsFG6AQVE84Zow2R
MQNPReOQehJ56FQyb/SgvDFHmUN5+tjXVEyMtib5F4gMm2u9blHdAzjKdmjLkKWy
ypnR5TsawmJ864fnA2h4QZvOTIp6m98RrD32z74by9MygOmToJejQlDCJXHPp6NW
s1t0nf2VAlbMzkybmBshjL22m0EX/pfq+mmfrI+pHNcWCBrVlOlsOcI2kqeBnTU9
miR6o5wdCRmhPdVnwAqv9NzShNUpX5CwDUnIOSsN2W0LPpepB1dZPTaaAxw5I+/E
WcCwqQLJzOpkgCx5k9B6aBlYksAiRLkU14TJ1v9PohMN4DDCt/94oFJhC7ABXFDJ
dRB+27vs27FksRuOA3MbcsExgS53QPIM2cszEcGRnowCchsVGnvjPZB4bJcNyOQ3
EbTW27H/2gtA8vBMDENZM56SCR3dAJqxbufvPsrtFHxXwATt978b5L7Fi2+ZkZsS
c9FOdm8SlEWP24j5hjreNkMiOej6ER4XM3fEdqX3pczFGJXENi7aZcueXSrBRHk4
vicPGDumx4I3ZMmjorucN5ggVBZTqopKol77vI/RkC8SJbWOBmMGipYYEd8fxV4V
`protect END_PROTECTED
