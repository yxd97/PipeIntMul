`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFLz3lzW+2PbPca6bzP3OxgcZ9RcbsqImm55DwGcf7cCxy5gXZvnEKcvIpB5VG0P
dqWCNYHNKsIc85hAB4n5QhqjRV/QFh2pjQSS8MM24+S1SP2xxIR5Agr1bhGA63s/
9b9fOaBvRFBg5Gk6Eq2huInOPBL2BLOZtIz/VWzzHFEBDHrZmyoGCCYT0d7j0Z09
6LlkMKqwJI4EuA4kuugbtBuVMEurtRVpuG6ZIAuHkApITjVYGhfNZWdmPYLOU39O
7ec5QVlh4CsL78MbO5oHF+d9SukhvfoNxVDwseuChDW375f4HQRmmicE0TJHVeI9
dH9eZtHsgJiJkyHPoZ2HFwg/zXHjGXTENlzZswycEwXNWKwYoHg8oTGLaiGUDhID
4jzkPAlhqbNUp+lqthE2nD0OrUcBOXlEdCscF8b5tZEE43CPRxkPiwNtVlq9P0nL
l8stSVx0nsihIAYQcPSW3iULdYVrtlupM6Nds/+J1AaEH4NTWFe7doIPH3ejWnnz
x5Of9foZS6Tiur3Gzyw3vjrIUsUDD69/kYDNvkgqqSQVVgvOJ+LppB5ipURYEYZR
nU1ZC9cSrkjbi4xcUgtdQ2WOgC84052siM+qWBEFoNk9MTzmXoakkIIQHCH/aD+q
qbVN0dlhwrQoFdte5XwLYwe1NzA6xCFJcc0Liu3Py/zJfZQ5dCku612KmSXWA3UB
HtzetlhKTcbxxav7c8SPuLZ4L5VerQjYynBjewoeYrKlI2M2cmY+2LG6LdyswQ3j
FQhh6BLExq+WV1mTgccCcxeg0it9GQz2QrYyAsAt0CS26Aj6QUDUUtOyheG+G3R1
IjooK1w+UNjxweAHvEi50UEL7Gp1z86qGpV+EjEih42QnOG4npPNn6FQwmzP9yZK
Sn1CVlM9DyKZhBCu8oYzBdUm86Whu+lYcL3+b2UwKTq53WFBcxMDsZB6NsoHwE8w
ZTWNjHHHMYosSh/P5yCka1jbuaA6v3dXH83jvapgxw5+DejrtfHxacyVm77eLJTI
CweWfRrrIcZHNXUX/TypzP8FMWsNLA69dREDzuG1qSn3L6AC5T4xSv1qCp+HBikd
W4mV2s5eKAib81Aj4M4aAsu8qrw65/eFrg+Fo7fBwS8APikoTysu6bWCiyiFHwgH
EpEEunyxQFDb5bB4SQkw2C13Nr9PbEyxh+NA5J0//CWStJSx1+mM9BBlXxKpsUWy
JfEbneBHuhpBvED4B/kdDVxq15KZOZMHAF27nKlpzD3MNlndDOTyPZUqVfGIzpgK
xtQGKQLoN5yIzK7kHw/42RTJAVEADx1l2OMyTIBS1aL9P+MSvOo7gCGdpq7Kr4M2
vm3Ucm4CeCJNPi5utckbzPp3G63NYScmaa1jiGh8E51Dhk2P0Bf2Q2yZE+UBKig2
T4lP9M6e2oO7I0qHabedTD1DQtDMGBtdImIMBI1GKVzFfuj8Freu6+ralXAWyl2b
xdHgm7dFHngH8488Q0SGdu5Gh/IwNWV0ScFbWvKt9LAWM1CwHpin3Shk7a9Aq5ER
0ZfO2TeUgdU7IBn6XdJcUGleD2devfYgt3UEjvQCyuKP+RkDMWFjQD8B8Kf1Pmmo
ICEm9lns3jQm+rRQ+pvhQteqffPfEz7J7thDrccwMe13ao5mbiWs/49Qr5ZZ5nCD
Mbde9d/9x/pS31aCrUpv7EpdlsuiaXvT3wxT+YvBYnASxluVgblFmhINCzBuQcKT
LecgLK4fp4fvPvFmHu/wV6cgB5GQzJ1gy4j1QvyI4jOhdZYvDJhdf7EsZGNVop6/
CtoYBdUbKTKeUI2FqteHGWtuD/Xh2hHeRxG81QVg2bKsMc8lvDpgRUlTQBvUCry0
R+umvwfiIf6bmbx+fSFm5RBsjiGDEHpfpNFRTGYKEgHirO3lFLdbWzohqMlRqGB/
mUQZpBvBZ9SaQttzAbfAZPEvBhzvioKLo/zXoVI+q/kJbghEdn9rOh3otGIRhEJJ
m4Bn2kH2AYw/1Fp7v+ejvD8HyEZ5aluTvlHmhHyQ3wS5ZiSMpXhEvz702CKIqmgZ
n3PQGZkXifrvg2wM6W77sm3U2EGJe6hsOsQ3TQxBzGmdYAQsjWXtl+581YK7voAr
KqqVkLRUv1JOtXJ6QvM9xLNEJftC6d1ZHX/hKOTy6ozR/i81yQbESdl8Y7E396Wl
4+QxVpnXCa9ZxsVFdiOrSfalPpQQAi2fpMOPJ8GLsKCFmKqjfwzzU3r30uq0KWHF
JDn/OmtiTwmJ+maroXXP3DZ7qG0RHawqJ9lUHWCYgUd5RM9StT6rJPVV05ofChvB
nSp7Lh0ZWaVpeb3lxgMyM3HLkfN24LJkf+TZlvrkLGklKqE3V9iATzaDC7Pyfkpl
9pwRydhj5MsgRRW98D0Krz2iMBXxVTFhMZugQR8pJSJ+RNSSQK3udjO4Do5alHeg
fRES/gS8mWB58wyOPZr2XMO7GkMATOlL6AYbkRRqfv/0JL77eYKYM+/GJ68gOuxq
rF191N1JsTyOIgdakWpOO2i+GdNHEpYlybQZZdTTU6RO9BKzAOxkogvydOpGMFud
EGa+Jo21JbYJH/UY1qS+grsUd9IJe/pkL/cirVhhpq9AKZzC0Xiir0jYAHUmpj4i
OH40lbgLDWloefqNlvVSuFmoJS1mktUTsfFduwoum3zS48h+KbtIrZdN3EELywd+
m0hOzBzHMCu10AxsB2aoFsaPpw32Jk9j+APc0qBt6tEeRT59KkpOkhdLTsWxUXZk
klT87PEq8M5KpjpezVvpuxUXCQBz+Sn8Kv4aAa/N9syu8lESSL7Ad/ysH6j/A37L
IzXUEuk5uko1yO0pgjTa6VUc2IhNel2vR1GNdNVsYt/2gdRGcGlV9zuvpbiUqvIC
tXnCYuaR7OXkw55dPFvWqOBwr53P469JuA+TL3K6TjNZtR7Ejhk9hZ+V4eAQEiSZ
uWmmsNcUGLzzOERBukR/uxJdz1/C/Zrc6zJIYWU/oO0=
`protect END_PROTECTED
