`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+uPppWVzEO21V8I3uNuOsbhCMvqRMVbBs1NLnYdeUzSSFMTUsry3mNG/qZstZE4
LIrM+mkiyhs3Ob2nrwGbhnlO7o2xvrXEXpvGHB+V6/m6xXjBb7uB9D8omRae0pxR
f1rXKhZqLdFl0CK+vcf1CYAQzXXGw+kqZyIhGv757RYYdOLqJoNBkt9l3lYLCkWC
wDRbieXCqDXfvnFsm6PnkDwIcJdwyXSlUrVUWUq+Yc1pmLszKiaatuRrA5KI5cB9
ZPOvkWxnVsoEXYYKADa5vMT7Gu0TdTK0yr1SwGf/GDVsmeZm7k/qZ2YHW4tDhGaf
vNapLdpPH+BTe/ApT/ZetyVCcZP8G8HiNn2M+rNQWTq5XovVbtQeKFnRqJQwGpeM
0d5jkZpGqUeAbOTDgKj0CRgOtLL5WN+gQ4D2XGHTLMOea8yXwRBfm+uDKFFABIJj
bUE9nLBW/clIaaSLWyoHpxmhqJC1rIgJTZFqd7NRe/l0u7P6vjsejKmCWvvFgo1a
ezUoK7CdTDXXhEmO/Mw+Y0hjwEAezsUPYE2sttABGUyhnUM9899VM9LIaV/GDfWv
tYXGQfF3ZY8XqeZXOi4RqVnYPOaDLBbBwm/BCBGm12J3WGKWZoh9hG/6BRWBn5bW
bY/Aqoe/BaWAmubgI09eTKLk5dyS4tjQaMfqZ1SILMulTl34pVmgNZDXwmleLkGQ
8lNcgjD4f/GHpkNHZa3w7fOKUQI0S1jvOAyHiX7JyrTDgpF3Mak36T16u79wNOqg
jcetix6rLo9jf2IMWRhavNJEtB8tuaZhXJpBfvd7gfc8mSjy3VjUTB6msrS3VR9f
e00k02iaSyjTzph4fDBKxUfGwI1mv7N4wmZVJ0QmNJX/ImXpl/5RpySH4JWju0kn
BBLdSb1twCUHqJvfnWjrTG4I502ujTOOw8fYLmMPm+yGAtm2n2FgcSzdFiUXevEe
ag9sR8NYjblClSnWf7lOdg1XLSwc3n55TjdKcSfUFye5CcrYvYdjl+iG/g865nbd
glOMShfoptklHN4kRoX6Z3Z6Wj0bYjCgqdcEW3fsysX1wfzk6Pi7jVCiA7SZ57A8
WmTL5Ypn0lYPnG0/Pxrf7TDnI22q/HKPHXOVRECRtYasxUV6UEld3rrAFAAYIXDN
YwGxj0f/jpheb5DNzsR9xErCYSDgGiyN2AscbkgnK6Qg+TNV5Xi2Rm5iYWa9GCyx
z7w6OuXGSbdX2bkV8ctFuscMZXtHVaF7NxB3hjJpJX20wxuOIrleJINWFI1rX9T5
5GmyLMFA91qYk7dEO7QYs7oaFpL1Mf8ym0n+zbab72cUEpmFWmJUZFNs+rjjJIOR
z8vy7/YEx+4xgte/OdZkHuuDlGMDXhTveuJaXGI6XdZQTxwSe9fHQHAWALfX14Mb
ObVfVwXRpBBx+p5V0pbvLHGNBl7r0+SShgGRdCIwXg8TQEiLH5NkQYCkBMM2K+Rl
lWumQvT4ovKN7OE85LiZJktnyVrFidXlhBdiA4GSzQeO2oUPavv2OKb4dJrdw30k
2KlHHemvtFwmI3Fm4viUWPy718jkYzZV9jaS9EDieT7u63w6Lr76KQTYt58mTpBQ
R04l+HY1736ueUFaZWNMV+kby9dckpEhPZHy6uDUkYseJNx+p3XGlp7HzNuHFbJ2
2C9ea0ai55WTswUwO9HVEKmMtmeC8TCGKw85voB4GV2VAzKMfLLDflS8lLME4Xso
riMSyGHu+Ws3yESngN1z8HV+vxA5VYMHICjWUvrjHhyVE4C7XeNYWWCwKbzDnvrE
LXYYnk0M8z8PW4tmvt2nHkdxHS3ELJYJd86G9rU56IaerZGF0rYE8xrjUtPpy5Rl
Ak0CR5apmzRuvU3N4E51pp+d28gq7rEWZAFGh1UG/ZHR4N86tisM7AS0RwEIBykJ
RVPW3P5Z/7No8ll+Ae3Eig==
`protect END_PROTECTED
