`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DURW7L93r7YT74BMS67lRB7Q+mYZ4s83x64Rq9xNdEeqiptjkxSNvbENCaXZvDW4
7nE6szIX/hFVtZklXzmb5ByutCvjbtrpuFcBN3rcBHpiE1MaGcxVMrHuCuySckeP
eLdOGYwC6XPKXtytiLoIZZhx+ycUQrSlu+wKi/vQN1APp097Djd94y90zpNCvX6V
F9ULEO8P6Qe/lKyL82XoTlUWEuGSQqL+0aQW8uMLyQNcQm6h8TfWHIhb5XbYhWGN
wYR4rkMcXXg2LlFXy1usyxfuUJdtosVdPM51/XroPGidinKeg2qLaWicrzn1A0mo
0YeMrKLh2nu7ksMawM+LzCRkrnxsCglYzyzxu5dtrQ951Xvv67h5ZIj4L2XjRBez
`protect END_PROTECTED
