`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fzhz9D/rO40LRsKu07Wdv+Xd5X4Dgr1SoIPnmMpaqTgasCVUes5H//n3BxpZe47R
jFohpm8XOSo0bbUJ9QGSpYYhDDbbRI5rnmab+RYNvcxsp2+eErOK1OAyVmBQ1P0A
B+IzCJdA0qmtdG4mKloFEAJagV/E60puTpKlcBDK1kx3S+mXOrZ5aQGhcFRXeO3I
hzyEyOMTtQ24SOKm1erlKg7/8tGauz4SgnARd0PXQK0GT1L43YlcVK86wJ656yhb
V51FzLnA37DCviP646pt1pg3o2viUdhhmnGmxJrGQEtOkw47HiKqu9NdH3U+MEW0
OMYXwSrB0qYWkXX+j16L7The9z0SdIaJEFi2z9Zu6lyD7l2uB8KSJIqpiywPChPX
ssytxKEzifeTsh+L1rj2JfxWbZzIUsFBrryITNAMMo7v4TjFF4SqtM9rU6fyCaMe
IorCTbqKeRm2PknWJOzGn6db/HP8PzrkyjOktPQaC5KocA3wi8dSnA8/2ClHbBFv
kGifmuKQHO6WLOzoXSWxlbV6bBerQWvAtROvV6XP5SzhQKkhg0Y4rEJWrIdIx13p
tE0/bht5q1y21yfLR/paLdtxKvs5IC9e0HBb2UikdEAvNHiDgjZe3kQY/33GkNuv
cuQfUX+E2/VK725RrrYiQzz/6JXF9RwJ2A/BdMDFFqOPncl9R3bO27xnryaUjyio
F1TSWgnbD6dJGwc83ZxkA9DjDvRnqEqf2Qdpv4tyVzE=
`protect END_PROTECTED
