`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WPY5eGQs8ZckL6g8vQSng3PHp+o2ZxMlPxQW8hwHSfUQdO2VTBvBajOzXw6gsB5g
hOf+L9xOvWdIkeN6EyVll5yYoJtcCTlIzKR+C1pHg2da3c8cWSlEg09Uo76cUst7
hdnSz7fNOFu2Ru6oXpIm2sEoAQOiL/N2r3HE49vdCTKwtvIZjvDwzAlWZ00oz2dg
tyoGpKa4DA6Wgb/qQQ07VrYpaFtJ49+VDHRANbNx8v0pnNLmoz3q/cOOKpcEcgDp
jF/XcsQXMQFGhXmEf7NuZ6uSj94pYoUJWsnEd1FmPy6lJrroza/DBkegyZvJDXHd
UTHlAeT7sBWpnF0p2oDIlpK/Vhb5AHTPR2zBWoLrA+0hBy/L0AV7hNz3KeClxc9P
jTviUUwhdcSxNOsMWQ7hND4i2uubsAsazuQ6hCBis08oErcQQm/p4THFCEmO4RNw
ODbGL0VY4/skg3HpGCl2UTPcak9V5/un0IUUG17R3CUzS9K3KG8g2HogDtSP84Pr
n7W8Y1Q6eZtASi18M9SBsT6VqOAF42s+7sW5yQ8DZHByFZYIx+c91wbUoZiwfYEY
HL9sW0C9+1eoQuvDwKmp47GzR04zpZzJeEL6Ww0y0uNrxCPUcm309Zrfu04DRZTu
BL3WbwQWjrGCSgZdJCi8514oIy7q03uIZ4I0Tw2lZZDDHuxFGKa5jbmoBeQfdx4h
jLlvp1C44r2JVfS17pcE7S4Z8LCXyLZjHURJoc9FzJnD5yz6qcoLd1OyK36b11+v
QodsmuWrTM+PGShGC+PU35UWhhfhUFyHwo66SoONNjxI8ZVcGw5prxwBl0CY635i
nyad67JcSOF2ZcoOcw4W+8Dw3eTecn5J6LzTB5KkhqAA3WvHqBhVbBXQHbZZubcs
Lntn1GUf3o0iQP9Nv4H+cUZJBFFOoPSOO2rAIuUpHEqEIKaHb34Ib/KiJAXHi8CJ
yoBKn0nr+y5VCc5eox8fdhvUDvGvU51lnt2x2zy2FYs/hT6YV1XK7/WbxhQTteyo
9JvWt6jNC9gt1bD0KBlih/BqIv1c9pVaerl8RaJ9H8PiCXmq+rYUkgSyc5GPMxoB
CJnbViupoCsgoyUVOWucVLHWAppMxyxH8hAdONZ5mLJ/kZ34igD3zbtNlqRK0G2/
1rBH3d2lbmSbret30XZL4O0R95vDFP9/4rNDVrvt+HiczeWYQTfHLwMqgWhetn4N
/EyBO8n0VL+KXVAVnQzcQXIdQ7p6nl3CNmpgfxBBIvUFPnENWhgMApIT/zyaylnL
RbSiOCcoxzVPKR8mcvCmS148tDUiESMeUvui8GvEvTzgccmL3EPv+DGWCr/QApXd
vS5Yp3Xn51Ro7yFE3mo1Vg/8+e1b3GPd7fNT7/MgNg0FZVL1kfpuIeX479+llJWJ
+01IDGqWIzKIB9E8lBvldpA5FvaKMVOPXij1sRaSyVy/teFsdG8bMk4hXJCINs+A
qNkdOFz8TbZmrzAkaSEz7RLUtAMdF/LINfLlivAf3p7mXYdXxMFymj0NP1SupFxm
CE626z7xeYDLjTv7lKkeA8znSfAUHNo700P+3QX4vIFp6KyhZUuvMomDyko8q9Od
mFfnhXkBQJNZGRMn5PyhRxB6tRm7Q85W06GvE0wj/zZoHPs5KLRYsLlcUv9jXw6e
9P2CPJFYQCGRkqWciAJ+iXdG/1VW9BeJ36iSxFeIfnEaHCit/+Si8BGTQLxGDYN7
/jXFvK4Pa1KOMb0WtSr/Vqx0vzODcdSWsxSVXXuFu7Kt8rVLm4QoAIV/G9v+lFWx
giGdaXJxjvxIx0wPnyXYa0z8SS3Zv/Kc+zdXAFMIaZLZIYYGULNniuZegbarUhI2
xAT5YgFochlZE4mIMBAHFy6pMVrDcEWzzik/byUn+w0X9+fIA3dNzoQK6UQ6kwms
VkT2QBCNu/v2X3vhCqseuvQwZlO77A/xXhHiPQ+wMxmm9wENiSQXaZjr7ll0rdoV
oyvrT4HD3tfc+dipOZ9qq4HvNEwNWJSqY6x/0jn8El5wPYiJZTfsnGiKtBitHrtg
Xjh/1qsLzRDsKBjj43PHs6qen+KPShC0I6CeHWGHbrCA1JkfwYY9Eh4d7SLbMV7n
fsf1UDjn0u0o6fmVDUvj5sO0D8f4JtksnztV0xN59/K09B2LZ2eBVGw//0ppZvRJ
PdHbEWPmewjPrXh2f8p9iLInS2pQogQksp7h7f1n52AXkO4T/KqOD22VoHdlmO4l
cMl2sEjTRvjIPhPnMdfXbt06AP95BEM8dRsTkxNSSLYDnNjKR0KlsZXEWsg1tUsn
wPaUqVrI/3qaHPzqnOJSw/CqfWNVTKVmrOt+e1USKtGZHsj5Sr+U8D4MBfmz0+T2
IAyunqxK1xbaMgX2TcnlbrOVaiH7gc6y4lzkCWdYRiubuxq68x2vMw6sCAiQXvnO
9aM56gftHVZjMApQmHsvzcgJbazVa9Wq0Q07kGGMno78TZHc1abHPFhfzTEQxYdL
xKZcGIRBAkscBtva4xskvSKnAuzN0xJXUH3nYG7Fq+TNY+hMZkVXT5y5smekSne+
zIsyDM3f808IShhCyj+23LEq4G7apmOPcDGGljabC0FBchAUUJtOphW2it9yIvLJ
M6i0GBl8ej3HlaX5Kz1GRhWbidfRQf/8pF1BDN+OTXSNLqXWxf/xAD4bKU9AIEtb
ysQCvvsyHB4rCiNWl+W/PnVJzGLq7nvVrZQgT7LhkiAmDdMDwg7UpBktHNhnrWBU
si5EEI5O2taj8INdS+VOSlThI45bEBZiOUDz8IFwus4VNzh+MOrhCr+DpRrNeGeC
KX1GTB/R2GtLUwLgB49dNIo7FUnkSlXOahuxfKItdaE9iBuUorrcxEJvsSTR8VvI
JGKlb6+puQA3PZlEeOhM6OBIsJXZnZ6ETyVhVLahf3eydqCvJxQiknXgAkk422J1
vC+gPDzIsdiStcpx0hPw1sEleTphl6XdJ8aHifwdkpWVN90Z0w4BPu7nCsV7HiXe
gc3rkgErHt2XKVYAwi4vYUvykomNgXtINNwjm+HZlJUzxGk9Yh74GM8huZsLR4jR
A+VDbWG+bFRGSmWcGrm/2TFDL4ZAvJO2zfoMqEcdgEzuwAYLghwF7wFY5QPsYLRt
Cy96yIypGnJHGXduJ2tKT/o7wITtcTSFagG6S6n/iWf3VBEj08GEP6+2hOVtOr+n
9Qlasy8F5fxtfxC3tQZYXTm/3DLiOExAlvwhtosXkTyPvvFMyWZFVtlwCrRsszJ5
BntU7d3TN73+X9bUInYDvj9188qqN4lNARVmMCAwCJ5xItYNlfy3zaAWsT3ZzOn6
X5Br3QZx/C8npzROqAvMNr8tBTMnfrGYPr6L7RPXBt/sckV+LJFHl/naw99n/SuX
Pfd1AIQDcUJIKJBAWRHJZEWspCAfNty/FESSmTBYKB/Dl+xSOhSt1AqkGD1orz6m
RmaiYIjLT/uIw+/k+M1cPLkB8nDDMbx3kr46+wfDZLV8ky7qw29EPK0Ex+WvSChH
jHS0qiCF2d0nSJABDJjlY67ecu8Hg29z4Xf7sGEvt8zW+7pfkCqbgdJx1u82lN5E
RRMVe1SQ7yLsYdJc1dRys7DA+DNm8LxBcp/Bz0GQNNj+8zaESvbKC3s4KsQGt2jo
gAEw4yg3LBqpPmRZCYEmjU2GbpHQr4rY/XF0HWX1V2e3Yt839AJgGV9TaAH9HiCb
yBFxuknQPv0vi2znVuCjBlRdKJiSvpnOx+4lxuljszUyJQMZbltivcmTJ6utjQ/O
Z4ZIXV2vL19kfUe47Tzv9AIkxq+obQYy4/PBJfJ8hIIJxgYkGKxjuaVKClg+Gawt
Bed+XQWGJUNBcH+RiawwL+HsEP+a8pP5PHZAfA/mzfAj8G0QpcVjbOyqoFstKJd5
v56HwAxsLrTLyn5np13tsEdbCBSs721nHXOiwJAvpXZfapd+WVp5jX2S8J9Lyhp8
ktF99aaSc+hd6yFiwRFk1AC207TiWiGcavqGelP4AHOAlIA6UjrL4cLuCleHk2nm
r1TGaWXgT3AWcLVtJxGCMIFUDODMm+zXUpStwT13D6h1v5b2AYv+Y79/RQaIBAT3
0l2a6RvGsxOARuFcmaotKepQLm3VvzoJoX3Cl7jAVqmRdo3cR0lSYtHylFgAu8a2
/Zupgv6TpKrIsjr4bb94G9C1jLmaEK8w1vBDDGBRxjN7D8Zucjh6VmVzPAF5j4vB
dLQ0Hl2F0YEZmX2e7U1bDsJuHm2c905PSgnegriiNIrOIuSMhm00i9/bgd+16KgE
7lYD4zi7Q0rc9szpBWK20KCu7U1kB9dDGlQ97bEZ2icJvizB7GffKu1lSqS0ytPp
6VhzeE4eHHz4P2VQ/murji846IH1Y4X1W+46dEijPsJmNlLTaSRI55X4AT1q26bD
uHg3NZCekHXfjy9XbixTzsPN3/NowdFUFDMPJbIIrPu+M0ii6zoDbbT7fHsIVXct
9c7Rz9lY6PaRg0Soe9mQeZqynNvqeFIVdj5jbk4T8CW0fTKJKyjM3/33zQnMH0HL
19AuZNer1FHhf+lGHP79hhaQleQiYH9xMHIRRqeuUt8vDEZMoR9ZP54I1pX7ROpj
tS8nUReBz4Kzd0SelTXEJTygC4cSRWCzKtlUxhQAPDqtjos3jbgGG3E0eytYU/3A
vXC3PDejVRLTFwNslmye3icepMI5D9/0QjlYOnrZ4ugcatO5ICExoYW8OxekONRZ
/5bOi2Xr0UFtlY6EyI9rsUkDEJgq32U4YwnvStI+ilLqSzl+fo2Nl4Kn//PFuH2K
lS/MPL4/+mcT3AktDP+EbxEfxkQVNHxBqOIMTTmR7Q6E9GK5hnKYdhmGBQ71cRc+
XAHacvVktvwKCcFz9a/t/1TbrC6PSe+QkwydhVFy61b9MPO8nHP6pEazF0UYvfXC
hNf7CxLMH2ynBmxzHowh5qx+ez6g02D4thBHZtwGw/435Qw59PrGMdrvuw4w6G0y
g1Wc3jW+ON0WOXQ1qDOzdqijpROJE9hMiHWly8QSygbcj5jwm/UkfhlnJCi4ZuOY
xUvEE/Y5irWw8gGXPkQcwMdjQjeihST4Y0B0RW+NQn3CovQM5FL/DCGkixF0vsHf
U/Mi4Z98Y+SIvuyFA3LVUYq7XquG7pJOu9CuEM0wpEKzKcj4vmKPms6jwczYiIpn
mUu3bagOtPSdV4jb+7dGXJsMDGWPjj2b8+k75UqPp57K5gOVXGmUMk0C5dqDy4jE
JDcKQpQWF0P/DxlN6NhD/KaXQNKM7ShNVbisFZZaVsLke0qdH4tfRCU0B2R/PY2l
HcFBUWRj0Gg0mZGoUNytMe3zbFDWovhdDI78gcRIbjoimR9fS4/wZB5WQShzi3O9
k6aJarwcDXdZII474YWzsiY4KkPhGhWV2tWZ/xK0xiW8HcMTG8qZb/KKUMU27Ne2
O0XwxKeHCJ+bJsKy2M15qGAKRN+0gd/fJ4PvT9VgXj/Trh0ypv5XenU3+82QKHos
D9NOgwyZEuSUT9a5apsF/06jWAdkdzqQQToaMaH8nu43cNbx33M22IK4RTxEl23O
k2yArzbQyoVxv9rxx7KSP69R2lnh4Sq9edFxSd+gp6g9I9QK8CdLncTYakaGhgrN
JJFi8H44en60DfMBHuzNddfpMnGCiSm5R+QbXqPcOu24fabyv1FJJi2I4Liw7Q+X
hrUQp44b5xFPlt4U0y+q5DhraXWq+I0qkiKUHZK8zYOYSQk02xM2Wo+2VPplaN4P
miFYdN9jxQuYooNbpuaOTzhcODotX9fYdlmYgFC5vAhhMv2Is3pLZtPoAB/Bp3pe
g/GoMiCvx93fCZlvSfx0Hm1rKXpcIOAeBucNdBljjRaP3NJEsjcgdrL5v15GChXs
H846Vs1L/fp/VaoJhU6xqDSXMnm4vGNeMqRSs0sZRF+GGUyRYFXqMo9uFqKmW4mq
DG479TbP4mxE0FMX8iAWfjy2Z4khQGXx9IrQLLiehuKMhTIDrXnvIg/INEvfgIff
mYoawWW9mxTx860QHPram0B1ByFidbzeNKXZ6lJLDT9kldpf+PJBiXuT6z1DzxIA
XlS41P8MODJwv/vkWOznErmDyabFgiw5u3GCsOc36DDrEtby/59GMpqzvAx3OouE
WNRiBydeIy/2hG+ed3YXMFLiucvzEqNkwd/RU6UHaLWwkAOKIsyHqlzpsYnCPuUp
zymvVSeVrzWp8/zF7jHdFwdOgbwhwTwfePjZ8mmn3+ArBFPLBauLTsp7hCGtlKIL
CDxOG2QnU1ou3DhYNvhf61ghOuj7/LPNQmjsoF/j2eqFtN58eemtqq94DwU8GUFZ
avE4nWIajqlEjhiIGnRW38o+RGybs5DSjGxotlxUYBmh84odt+WTPqZE6hJtuCJn
tZ0YPVgLKzuzn4xVZ7sU6ICfkymnFDD54KAMYkZzvtUnAWp2GbJnI34jp+Pnf+ab
EaCc2efyAtdn23ZVslwgZyKQ3GgdFt/b7FMadbGkAVO6uVlZrLfy7BK+lLx4o8N5
ikVrLB+jUbddMUIGwpNo9GNBLVDJFqxv+hGH/YkwNqbKuFg2RbztpoaWEJKwl248
WnaQa9l4tLMqomPlcU39RHdzlLaZ2A+zAvKDs79JCTTMEsCPeHHT3xbkMVo6EjFv
fY66dC9EmG2Znps9ABiQzUxltITYy2PbDzuhpOQ/Y/QOqyfXV4eT9l1ROpH6Dp6q
KWCKJ1D/0uaXH8clzZNzdEkfHl0QGBGcVKxklnCKVtVqAQGzCpBVMFlx7Xtsl2qf
E8uc6zuUN4jk9SxCcB4fTYESQsItOwotkqjggG4SsxZqaRbQuMMlOIzu2oWnSRXw
bZn8xbR06dH076XPRE37wv/BR/ol01WKqZrhhBiSX0fC2n3HS905YKgZMXcQktBe
dP+UywU3bQGWxGa+T7Q5C1Rove/oB6G5sUluDKA7g6WuzLXJpGUs/y3r2pNtHc18
yIH4me6ICQlI11XVTtI8yyUJvgoy2rMXnBPB4fPs/7U+yEe7SJDOif1y0lBGm7n5
YW2dZ9Q8hqKjpG0RATaG5uZxFMtmcMxT43Kn7ejrx9NTzyha+dudQ5blWjuiNKT7
Z5WOy7cpFH9cynhkC26hIZcic+shB9IZS87zocIqxpN+bgPj3duUffUbK6sPmPeo
gd9KSaeGSyeklk94wFgbySzbo+NojJtul9pOAUA5KXnAzsAS7tIBt4nY6B2aJp1/
d4RBk93OLrayEiJKPRLNvEB4lN7GfyOyhl11rumn6LxX/ChhgDJQ+UMFaUkuZ5B4
Qhrfh3nKGJaviHmlKJihT4yi/75pUovGWLdubpo9V3elZB+WC/NbMpoPg0Kv2nHb
wkVXk/AIM2vBSEJaG7Z47sOnZhsaaxk4N2g2Kh8IJGmjUkRhUcHDhBmCcdlQQDTB
/eIbj9wINoLldYq89ermg1eGsK/xB+qdYnNK9wBgCnVeZl+p1L9aCHgxoW3ioqk1
n37CrPPl2UsYCPQ0+iJZ0n2/ayUEQqho15BX7qzmE3OWlh73s/d9N1F/Ct2Dqzdt
sQ7LlSWGQk4FJUtbX4qhmgzMR7GSJqVrOjoqTChwFeM+EdoZNf2hUUp7z+EbdZsh
fEFLIg0J42fi8oPLyFTUIOXBRuBtGmO/XbLF9rfHihYU8p+uIpHlgEfO84aBV0mA
w5Fu54OGXJ4vgFJv8FjJnoFbcM7B07Qt2HIOko5MoFksKGI2Y0b6QAzc5oddnh5M
Jh/oYHULnEYU+Wm/3MeV+/9WcO/8E+7wTt1HRUHtHNe7BfaG+Un4XpSKrl7ztoFP
N0NmWxqbA21S/9W1+aEV+68vsQ9eKYqSPLVJZOXYg2N2DwdSmywgjTOHRKfEhIdU
bj1SffxUx/j2iNW5KN1C09plyBzz13kwaltd7UuMLjkefw4AiteNaHANfPLNbOCB
vA3Y9bWDxxgJ5HVrravQ0ayMGGQ9UF6ikqpQdwHjo8ZmsC3aKeM/Fs6JuVdA1E1m
PA03ZRm6CYPNER0nI9hcBk7v+GO2eJf+LEwshFj1XaoMm5j/l0h/8YpdNg3ImQFg
qL7OhBknL/YaBkbnTGrMhh7WRz+D0KCNUyDjVEFARvbiq36zCONnwqlamTkDZmJC
Teu6gXnIsUgSvHnFiOvTKHtFsnGIgYxCz6CPu4PjwF/IODHvnAEb3VyBlab/yriK
IOWG5JBsImSDlkC5Iy3tBd9efTATzXeCEM6EdW/45dNCOoKRD6UCsg9wGdn8ROWJ
EelxTbUpp5bIpcW8buLtkjzZqna6oUaC3Hj5V1VYyXMdJ9Xemd/VrdJHs8lMk6S0
8FkE9wP1n5FMhXp76DZ3ESSyfbA422V3kg9v29bi/nULusXOCK5ertraAJJLvO8f
MGb8NiccBPAMZqxOxYLFfws/YM4iyXpJf9pk5VZ1Cqxba2dbgXmBMw+/kVExdJ2X
MzyfsUkTVRPR6gFoGZqRH9R+Y7sU0w0FoYobTl7GHvSPtOL8s+xFlbX64a1TDPcJ
PexDqmRsadQ3Vx5yR0zRMZLsYz+Ux+HhPLgJQ4qcIxT90Uvb4jjietlsrdX5bWU8
4Z2qNGzAnAAKL6gY+zmbvCIEdsGIFJVPHk0HEmopNmVL8ZvYCgwY7IjbQRFUNGwq
Xr49CWsD5+s90+uWNFTTWtTfZK8gIAdBBo64zi8vd6SslLGCVPheXAXWGxYLZiH7
FlcVfmVpaOrYePV4ujxKc1Laeqcd4BeCbMpH/Cl+xFrZDzxGgFcKtvSXvIHsvDpe
OeLGJ0cs/fisdxpLpO4AJEyKi9s+v1cUv4K+oi3Xa/pLzWFUZO7kPP8emSVAKRwi
/+lh4/OYGIwp3DQVeqSTmbG6wqopmkALri3ojCwMKmjr9TCeNRzzPKSSmSuPapYy
qDL1fgLejiIZoERnB7djggbfSVRp4wFPciCj9JgxSuXLql70tbzWR4a4OiXqgQzJ
spqh+Q1hDsbGZ3iNXqhl3z6UnpgS+Fs79mCQxkOQySMuT144GOUl4TNm6RRAvJL6
lE3fR2MdQHkWcXOTmD6cxKiexj7eZl2ai4IbCLnptHK0Q2F+VUfTNQHFX2mbVUqS
oHIXwM82c/7hWgjHpmu23JJ5BL6dbAOzpCz2lF3xW5JFrUDvxERWXj9OOUxR6jYj
60P0hkdfPh1wfnpBfqVPS1ySaj4Ftjf7J3FDGmxVOesUYV09cSXDf0mLnN7t0Jai
OSmBsKJCV4dCVxvbbJXFV2m4AxX+imfzAiYAuyEyFSCuyut7x64FoBJXxCiGQTYr
9wiNzI9iLbB7xS5HYJlzAi2fppKCc1NNYghf0NT449DB0ryyRYOcvKEzsjH85fB7
AaAMvgBl1hvFj87FUsfQLLB439A27BvriUphWvFlzREJQevss92DFlZTBQ0jzRjk
MbvhhlM6nboE3fV05lO89LwIkv5zCAExzXXyZvK9f4O2w5Zu0apPMfGxqHukHkJn
jJz8fEel1ivq1VLtfi2vwCaPYPTpf9gIt2/dSC4bQNCsLQpQmZwG2WiZTt+vaWYY
bbCLZN63fgOlzk/t0wuNfT+s5gO3D5q1NxO1/EQ+UWdJuwJiokgTn6d9gx7DvyrR
t5BeELIOpk69J7WGPU0jf6bfVHFVfJyd1yDjag2dpk8WfCzeEUd7kNsfgHVXb5Zh
hRsHPuqMTJPpBeaH5gYx6g+d90BlILUODo6LeooBIWW65o2aUtnxQDvvapbEByB2
U63AEU55aTjoCpLO3uEj2cv1p0AMeg7g3anwnL0b9nmJtMrdeDCitWFvv/9ZixfL
kcVwG7HPFy2Xg1OuIYGfaPOGfGusaFJY5IgrMzGGlW63mqi1rs96gUWTKwMbdR1+
d2oIdk1ouB09CfnFwJIzcs+slA+zBPHvsWriAwcj6IEVyMZl74dQN3BswHBH3h63
lS/vjSXVv70rTEpJeSns0AAxweyXhrdjHjxEXBB/TetzyXI7b4AG5TN6p2Qw5K7R
mUSkDBdFIqtqFHEIBMzz9w/pDtuWs+1YH+KIYrHQUj6uR8otjzlRUujYHPb0Vrfp
o7MpVL6OWjCKumq5HnbT7GMMozGmL5Ael5BNb8cDyt0XTfM0WQ/DwXF0bpnf6Rta
4Onk5cK9spZrmvgBu3T/o6Acdj8Cp4vNdBlXayxP9Es4m602+QHLORtCJ8B0nGP2
TI64E4PxLNAHwoZyGshBAvaz92iiTGJV/DkEvmOBPgZU6q6dWKJg9AAJpxMPfL1Z
H78XAgEUD01WyWznoe2bZmOI4jmoWYqkKnQZIqziZ1N6H9P7zSvq7Q+NqVa/86iP
qwpE49b0x/nSzC+qLyWN9qFYD3S/2oAKMFC4Gj3GpdKlIIyFC5/+NeKE4wMKA/Bl
RyVuSXxtDi9HhIfhhp5RCuZpokn93drnWezS2JPSZC5KTh68zQxZ+xwbidpgQ+Ne
6G3uI0MKLrMhas/hOD30rwMU2FLWeZohBsoJVDB6kBpjpuXsGF6+ylxMJ1ePCwmI
8jh3eULH8qsBwvdiniwIyau9dhlUcfg1h6bD1aGnAt1CJDFx7/KV9n0WE7oVocZ6
RkXbCxY6FMRePvCCtHZZdrUme9OW9rEp6f3odlF83lzCxul1ptpv7wC/RPj8dQGJ
Ry0y56mU6D+odHGWR3XuuEUwl5y2tR1xeIoKcoj7qSJP5/4dbU68X+pJx/RcEC3N
/mh2klQenbNo17UXJPZNUl8gq2gu1BV6zHWEwoH0+eGy9gtSxCBtCdAKiQo6ehca
WP/acgXo/UcPc02Vbs6Cl2achHoaZiJu5n0AiROBgq8ZLYPI27qTVbMqif+NLL2k
qQFnREfBFAVAYHvOWv0NMevtNMHPxSdeL72edEwHmIr7uJ7uCDY0iB0E8MyFOFrp
k++D01xFd5wpphkrqkHwm6lywXBEft5L2BeFQN1S/BerKAONIpVdlcC95a9sCPkC
DL0ubMgXg2hz9SdIAZTtaz1MXSaGsI4H7wNPuKEF94y9p6uRj2pLFueH/MlDqGWx
v8w12Ah5uARksofpRsb3qdL25/sbTqYJSdqJnbzEkdHw3X4ti5EGqJIqC80N7n6l
Dd9hcQg2KFDgkK/3rm57UDGtksLOYSWIIZyDTHJRIQAYibtWGTVscw5q2R3u5w1h
GgwAxx67nvU8qoYATT+yNJpT+ZyFAY0D12X+mWY26hTAZnGgzDJMFDler/4po/d1
BCh23G5QBaAHT2Tn9FjQyaGNRINuzzI2NZ245vOMSPUXxou8nE2PS1l5jBh+Y7U+
87sX6gSB8Gu8r8JfNSwhSK70txCIUhA7JCC09YD8GxQaKKoeVbG/qY7fKJVZeOCs
PMEGD63BzV8J/Df3ta07xympXHghdpgxBap65fEEqa06ZeqmndDDG6yjmclXm8rO
5PX0DlNb6fYYrwI7oQGIV/AMAMkOBY0ssCAKH8P9IMDjDUqQsyd+TO+2T+m76M90
6Egs7QOZZMWp1xbTlmsOrM3chAqe2bc0nR5UwHtVchapEcu+4ZPGYIIgJrpHogPh
j5br6oSnq/c9I8PwPHyIK5EkFkna8/qy8hE0Sl0qgvHpuQBElklNDAjaMXTuMfb4
o/RMOtIbE6JzKSz7KXOBvHo5RjC6j0JK0vvRye+zNNhBHJsQKJPuatV4ACVKhyXO
Ef21mDE1NWBoa9SiZjVGcBmWLwdjVS8+Lxs6ogHslZH6CZWW8gbnYfXGlDfUzCxm
XAlDuelDNWtXySG2PTi8aLqoVf8eKnDPqxFT5dwlOsU5mXNZGM5shr5UY0Vh9mME
Xm/aRoe3vxu9cYZqqEbGbiCxVVc/mscniPncOVySV0wk8X0yImL0WIT1xogo+y9l
yopv8uoZRGhW73pf/TXb4qBkyBhLCPtBTOooOge/2kzb3dHT1A4Qs+OtxxATwDhp
mFMFPAvZI9Pj+/P3tzz6nMBiHhI5vAKKeCh6+BshSb4u+iOFdmYIb0HSwzAWoGIH
n0CTZkQPjUPyb0TAwAxBfXfdUqWRGQ7zl2ak7MJ25/YK4au3xpCKN0nlFwWCeOs/
aMmmxCiwirn4WIOdn/IrrVjaL6J7HfcjayqnqTsNY5tdsXQU/StazmEeQ2F4fzIV
WhwxEusvzQsfV0oBsXC/N7qwDt3SfmMvtBNmo8vfBFiJ8qMR4jX06I+TJh3JwtNZ
ciWyhJYV5Wtm+eizQEQi0VoBJ6FsB1ObtysbG10YFEi7vdE9eWcxckOlPbETau24
m0MlKbPyEHya50REpUJnh4MnvBUwCFUraZxwm4wvVfi5sQFlVXSiT+DAeXfecChm
bWExOEcKDmRHihc6sFW96kEJVHdrNKCr5J1JEP7SX2K1pAnsI8RuaJbn2ebdODP5
JB9D2uq8450GHrfvPi9d75Iflq1PIddsowVizuq/s5rDk2mXL4CJfKadsxkhZBFY
xW4etMBbMhEEDI3llK/uX8XUo3RWuxvVaJd3y3lzI/Rw1mOS6z9D5PrxITUn/iaw
1xjqaMQRl4mwa8eiasqe+cJRdD+5HRu1Gh+djODn3tY0Sxo/N79IBaUBEgK+yT4d
LYzFFaY8EJE8Z0Qb3BGo6c62QAnEer+NxH/zFukGUGsYB96TJN2NlRIOvfpsOw79
uzAoFeTb4lpCp7dLIIY8bNcPYT6QXOdY8bna4pA2ZM7W3rPZKqM6ojyFQsfdNr24
CFNLMMGBzjSc7vhB5DtQlf7yaJLVOmM3JbEl7K8svD2NRIJPcxWbHXcLaVSBMQn0
QPppVRiVAaWi0SrWyiu+d8mqt/ID4eutN/sQVaaRP1XBn4Abxp5UcIX2VXItJEpM
XmCcUpcD8bqGQDYzWRkMJvIUK1zNvmy65F+y8aoFvdeYt+iW5KDd6zMEQbylWNma
pG6x7NDcM34qxk5wJxMikzOewFoVgMne/XaKO6uc2cOhPKRu+0srFKvqQK5QAGWm
`protect END_PROTECTED
