`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
loKUt1uVZh5SIUyS0VgDoND1AdBEcvfMRsqJGIkpqTuhJu90fgHsdALx2tUtSPeY
KyrlHIJG9StAs2bE527A/3lUR2Jy1mj26WvTwhrMO7SSOynz8easZQoAztS+ip2S
gpcGpb17VmW91DGeUj4lAgSHg9hbVqktUSu4tFccH69H6+8WAip+xO7xvtwwqIzg
lTME5LrB1jEemLK/SdYA3BEiRu+qVkyHunOHcnYg0PeA5WTEFf5Jb30z8jqchurv
L4NVBBS5Hj9h5F8tbJrsT7Id77WkqmVoj8S86w43GS9mlINFEHAD+Xo2toCZxvFj
scvbqC8I5/D0LmEU6aCtCvGmR3sNXY29EBhkIkvGMVdV1+aYTifOrPUIPTNQjEuf
jsuuYDDAXBqc/2zlzpjvWqgL42BSszIchHy7B0gN7jtjfJoGqq+kHIfULEqVOsKa
QRwZ1E9Zff5LiL/2RFgGW2m3un/Cmd8l8ZSgm/TOsfYsNQmqQbmAtjA8dSMVvTPc
U+pCMIKhL++HcsPf22vVbMsBxbJklY19/cIzOzsVy0m5dNr5UM5C0HMCJcIkE4DM
+qEj1WtN07Q/G1e4rzS7x2kWvAz2Rwri09tSzh3LjXspH7zYV3Vre/b/wk7mC12S
PGRFDs+d62TpruftvVc+OLo1/6eJzwZQm+5bk1qKVPZLNWyNwAH5O1B0vAgGFPQS
NAdoRDVxfQXGYqgltn69AX13uOKry68l6s55b1+CALpGTsy6cz5jswjnqHiVbB05
fK5ygSlgWh/pXs3A08igpfGTlX38f5NgZsWSM8oBQtXfsTQW7+y1dU3H8kTUZIJp
tZXp5X4Z5XeWoNZCadfBKITFXOwV3W5SDeH4Q5/vj+7GVlzqcc57J+ChfUtylqmk
1cAqNlt19JDhKUbO/nrP/13Q/GYMHN1aTpXH5yZ/MsvdhVRpm+5pxE8r4gpP5d0S
xlaGFF1hLRVjjqwAUKFQj0jcMf6OPEmM0gTuIwgRSpLfNtldUFkOYAlnXNN/S0F/
G1o9iKjufl5skfQH9jklgzmT5K2uU62gH1JUf8EbmeHki9gi1CrBUfhjSHe2xd4d
pyffGBXgy6+nehrqaCNicrndtx612eYzc+HIrAaA/kXzOkt7L3YkmlREe8yLzZHy
26rHycQgX0tSiW4BrR7LMyRXldFymDtqAtWvF6Tv8IAw/uxJ/31ZnuY6Ltcs6fC7
2OUFWeKa/27+oYbjFeK9HEEQuQMS6VPRM1hyqzoIf9ct6qESzpjd/nX7mmS2u9RW
m+GHeK7Em5+Esrtty72v3E4BLih/Hdq5koi8HxFApbpdNqhkPvF/uQcZzmd5pL7D
zW/aIoTRoHEfPJCOq3b7L4OhIfAQbhA+KF/+lBKuhd3R0xKsxyYPFeFSGcGWZQDt
JIa+84XQrkqQs51dZjnJ+7K9QOvcH5ULDwJ8BfBfqfvqQZwcHXx8QgWH/ltaKzKl
+VLOLIq0WsphM++5dB1U6c5zixB6IdxJKavKT3URtQ6IdJMb8tInVpOyenO+pTQ3
frOqQIC3tWOMX22EOXUyyEUg3m14trySc7p/8/Ksq3WXFYsBbrepzM/LofQFwALu
7uo/q4V/mtENoYs+5kxiaAoX4IccAI/yTm5GfTIuWyCTGiLWBItKD0YnxKWwQstI
DRu0847S9Txu/j2wrrJ/a9QWPP4vfo1ptD7bEyb7oac57Cqyczc8s6TrulL3CMWZ
w9V8uFe4aVcZVHjz+VX3spGN7biPdHKzuuvKL3bRIv/Mk9bMmCfkLnf0sxjA60sT
A/o4pGxP23A6nxrhl5u5IQiyFlcoGbwKY4uErlMG+y+nkDMUL9V8qXA+axu/qTZH
T/OPV2r5pWgF9Fui1McPGC5qx37ftUwOyhR8RbXtdX6jyqveEWC/23R4LpkTa5eX
1aLoYc2neOpMgUYQW05/JtK03tO/B19N07nhLw2Cf/cWDIc7RhD57QFiaqJre5/4
8+m5QWn/yFh3AIDH8wbd2T24VtPbuf39Hbsd+PjlmS+nz1b53Jy45EF8XQx7aKT5
hQ15Vv97CSNQ5Il0Gwqtq/VzKAsffIOBLB352CABoMihm10gtpAAUPfN80n4S/BJ
9IfXFQS+455olRPGuyZXT8PsDdSr+UOCoMz2sp2LngN3ApJlGfvEM89AM+ZblqZL
ackbG9wVP+3R0iBw6vEEQvH9mBkwUioTvYZLV85ZlJXjxmqVz9su0oLidK2L73tm
7DPi8fjNBSXo8DZ7aOZmAN/x4e9N9NoRkLcN8YeIcVAF8ylxSuPKJJsoukClaWR8
WJevt31QHlcUFlOwSwQnCloluA/ZxxHOyrwvq2lJGglkdC4OnvxWPP40Clk8fWwy
KncmTIFMMrbEc3+tZrdqxgeZXc6B1L30a6YItS1/6WQOWlFEl8OamHcwyYQco7Jd
A0hpRF7LpZ8WX6lwLUWQsUAUFwAB9qcPPT1xtEcW6ZBNMYhFurgHzQLgjyAoK4dP
gFnH2Gk8z85JQuuaOPckeV56oEpOc+JJ5hprgQeWwVowHrfRl2gj0hv4HKCwNe/o
cpIrhcZB/PzRZQ3svRmn4/atlGsrHOPUY5oK8MFqMoCuWwAirnk5q7E6/ZnD5ZQ0
oYdM0bUe5kIEaIg4NUr6DkUFkxZEtO76soUpVe0A+8spQve1T7QgMSq0Z7K8Nhq8
1EQ5qt/jLvpCtgLLIkOIqGvyGFtInHufudwUNQp2DMcdqp73xPgYc1sjijda+Mx0
8yR3aWYbJKbLQmlBzGqU00C6cgXa64NtoAFlbInvUd16oDgIAuUPRjVvJlO0Lp5Z
uIttNO6+OMoulluHqf2JqX1sILkwSIuRzindVduqZzHm7SEZgA1yW579Hen5/UEV
5x8lXhUYnzKcyZWIMgfhGmWZ4aidJNEFMp+35AnVa07LMSmxkimTWy4PZN+7udHA
fY4RZDHsHJ+ilrZjdAMbcj+oVNe4HViNAagGtEnQx+pzx1AmnXE/ffFZDx+PoxxT
7FBsl7OS6UOyF+wq2MsvIG4dCTVL4I+BL7SLMEDG/ELmIOc/KdpsKlkT2c6XcBu2
jQ0J9AgAeaE7264ESlvY3DfC2SK260ZPs+4t7nWzfC8lumKEA90k1LyNW+k81NEE
n3w/3VnIe/aPsh1FWi8n1WO5WsNwNG1UBdG/6bJIvaaQ9Nr6AZnKPkFzOBV9+KYm
s0KcsUlGkZYjqz+PAW4lN6ovXAGScZX2CgzlzGW3CMN2c/rkJ8kx9XOItJ9dNhyb
d6humd0gWqpNYsUDpjJZtjcnCEN+ui2NeiXlm6HmfS0FvHdv69OB9GofVJUUxVa2
4r5XBTwgezjjBldqq8ny5TZzczBG2gRb8YsbnxYJ87ijle7JG9Jb84FjZFn46Wkl
9kPnXJUKGNW18hv/RLou+1pItpl4PGNrWjAzdnldu7VQTpmujaCxlG3CxumMFtOG
NqW1uXOdIb7LjLHk4hHZu03ZXUNd5Wnr6dGPSNE0yQ8/oGDG4bVPvORqshzFwUgp
G8zJVaQPKcNpBrQNcnW531BkkCdWZY5fRjEZqiv/7Y5TzAhLV6XlFE429wm2OJ0C
Br3WnhHXoa2TftS0CjmARu+B5rumOEcY0AuXjlkMUbHauLgzf1O6V4IFOfk3hByU
OfuP/sibzP3J7cIbfkHPfR8c8Pa7/sxXZuhEMiHw9wRI2e2Rz79D671bPNBj44or
qd/Y6pg5UGbscDtQorrD+oLK4IPcEDTrZRu8mwTYTYRw+C7b7wM2sXjb5cP1WQXz
VwKRqC/Y8/XDsBSU0PWb0A7n99bF1I7ZYOB0tWp8LQgIobPQXVUR0rnVQYmrfNFO
/wwknoFTRNTZkxE5NGMcxo0oO6r5TPj9dhQh18fIJNb0AR33CivTIfxAqUIc5ZqA
EmRVMBFUl1bZ0QRJv/+EiXHtuuxhlv35NKgsEeEavtRvHmzX1X9gio93bdAWhr+8
vhRKCMFbB6wgJuzknasaPJtsxa3925XDOJOwJ0VA0alPf/85Z6MjApQet+sZUjIA
/ot7iux4QZqsxno5AsbxiqLkJL5wPuNXhe2cCWBdQDTGMZgCyeInhtdIB1PoP6p3
qvTvCb4YFOJ9bvLyCwzhRGTCiNqQpZ2KN435IjWZJ50XSW/kLyJIwg6ZN0b48z4E
YF019Gyp5FVTLUBZiOJf0iEvj4s0EBcUmJau6AIRE+8uHZQ13yo2JeFEh95fZEvT
19ptF1Gj998hNXg9BSthfbxMO5KfZCOtMVp//ogoZQfh1tMzrfc94xM0r0pR2Qbg
oainYUkpqvjwPng648YwIegvWeATVtXASylDnLHosArQ/aIBMM5pmwBIlzWgoGca
qtUwuAyRAB6te5sKZ+pECtB1BzEFL1xN4R0YgozRJwLktCX5PC59WweoRAVERDPt
6kl5FwDhOLG2TCixnhb18XlLjuGrT2JqOq/pOoa6L97W2jO54xefOUxOo6knecT7
iCQCntU2f6M0rReArEyQe6HnAFH7OXJx0xKxr83TKlWdmyl+k9XMAMn5mhUyUuuE
WKPzPoLMyQmcU3+QTsnbMqjYYZKJthBX51XHxVW2MTQNVvS3yB+IuPMfu7FpA4fV
EjbxhdR5iouofy7WkDq50rtpeIbE7d9Y7Mliz6I9BvbRkGMQ0HwCDRctBog4kzQ8
QBD1pHyCUEe0KfpLcUs3QxjZ+avNGQj/JiVd8Tztnepm04OfOWHQnV/pIHEMZF0N
AvhJ9w2Yc+UtjoCOFpbs/AoYKq/61O56G/a3/T9oG1PcUreGvkgUDBj/Kb1orNo4
lVI2SKvPkg8PIcS6GyWQ4XM2Vr4D48t9oqoz37I0gyvQnpYyxmN+ncIY9u+V5bVB
hamE1Nmk/WbBtNmjFkhLwQZ7Fa1f9+CsALa+ipvmKyukMcT9yO/UYbnVEYmVJL4H
F9CEWhhUQ9GGpH+AUOL6qaaP2uQjUTGb2GTbWhTvFTsgUGIzrBLDtXgSDheYB85L
K+OzuK4uu+64xE2UlH42inV9CZAep+gmSRPUsmvTW3iRvu4TNaDyOznoX+H1Wkxe
gRFD99M1gA29tjFUcUAiP9R2ysLhA+qdWaL5vw92sMn7dmGtZJluIv+vE5VWKTWq
RITJ2FRRH2rejj7P81FjrBxvsYjDVltVYUyyTiiXgFJKq7F/igiCLFcr/nDK0tut
6vA9SM86vzkJ8KdZ25FWhPUVNrDoG5wVIPqLTKDzRHLV4Ob3t7UpNg/7ArlC9Vb/
b8YmGyO0o/qvZeXTJFX0C7gkG0RIKHSp7xv/OFaG6yScsLrG1i55K6e8luzlG89t
z3eB4qwVeNEoritUbAg2tiRgdogVOCy8UE7DxQXI8TaRNBXsC2Py/yGs5RcFYqWS
baAj4pYywFwTokNpOJyuOLlku+NzcS0ARyuHXqa2nM1Re2f8SsQBYQvtH3d1Yhdb
4sTjH6EXsoBvvGEHuIVchBin2lpOWEZS4uLENTzCs1tW9l2rOxUaK4KqeM7SNgIK
ZjHslmMrWQgZj3/p4loM8b1g5g3K+MAsC6WPPZ4wVtqgJ+z51X1+BZkFJfjEr6yK
UlXVjOkgEMFTX7EqL4NhzYQ+QUoVVfhCHZL/SqKygMcV/kQJgXIjIzXwSJ9VnR0X
bSnnpgrP86NLAS8XwXK8F55wIy9ZJqFwRZH8ItDy0nowGXdQJPI8r7IAJwg8ZxAi
4zojjV8BFMN0R8zO8c6kkj+7aHQyv0/oV2nH+6xU1u8+pmD/Ck5WH0IDj6ub6urX
+BoT+LhEMGv54OCNleFB5hzTDZVyFMf3UB+mh3eppaLUs0fNbUyBZ4EXSKExeqUE
eCKeoqf/wE9AkSfGQSdzIRv4gsM6Nx4hJ/qO9vPIfzm/sj3H/gSkq+eaKgnvb8lt
2LGH0XdYLWmSgL55VzO2DpAXcRA/EenRqVnfqyGRrKsvf7XU11PW7HdFyQkqNKno
WsvI7HjokhRdYTiEg4vccMY5khL4iubtliIwn2bcbhypsqvC2JVZeaa8Bzw9gpHU
Sb018lSuwKIY2zi1Br26Rfi/XnwIadJY/zJXySzgfg7wZ7r+5sRTwg8MNmNhBTVJ
Gw2kfmkXlN840Omgki4h/3dd14pnkx+KjdiRFl8r48JFpHDaFVB7w4eF+eZ20uD5
TJ1ztDYGbmY+yR0G7b+URpqnKFpV5oBXASFsnsAWSuJDIvZo3zDPXMbdPCuuMnqa
NsvXZvLpg6iOKA/gBG+J08A5+LmQl6HjWF4pFdZXCFX2fwu4D9l9DWLPvQYnxVzl
PAA1+VaCKf7MSLQ+nzeQDSIMIoTvqNqs+UEm7rUHLB2f4JMkwwchMK1ctYNrTIq1
PcDPYJPUoemZcwjdzjYtteckAVAcZu74GjOpiLhO+SRDfmgJscJfahSItO7UDW6K
9Gn1bFQT5jgYyESdr0YlJLtjfFqmJpwNV8Mv52yCXTRpTrYDOmVbpucBW1XnWtcp
Gc9JWTNeJjYyD3rLuxXZzqEPlcTLTflubJAsAc1uHOqLT83lZ8C8SdvVSCCnjJh8
YQjyCePOo1yFo6jS1j3J0BXSuFuCiRgm5YaDeurTZQ5FIDR56+u4wd2GSvfxwq/8
m1E6Pvmj8DXFVt64KLeuz/t0hAOBagUknWP/oJ30llY3QIaTQ+DPMOJdAkUJtxsT
/ptPia7u1tTOLlpsfxoT8mC0QX+DCidiV3BaO9Kw2uaMKVmh/W7p8A0gvlTm+O13
Z/Ex4sUJCWqKDF61zFPHUIg8fwg3gFizmDshmHu68bryAEIRVXokrPW00KKztvmm
HfD4NxEe9eICBqjWcaW4gTl+cv/mCvyEBWfq5yeVH5DJz83WewJfDLsSJ/ZbQzDt
3Q57HwIw7H6Nhy7rWRyB0PoyFUCToekL4euKjZRYLc0K2gBBwt7+yMOg5xriml8q
xLa+MVH4JFoosFOgCtMKlaKZS4aVTIFHP2v8fZlLyHCpcbYwBPHMqgIf2ZsITwxr
a909YVTzHpACy5fXBHhmnrg7nUzwp+o6lb+jMIvbjHlmV7ij/RKoChL9tC9AQlbb
NvtncTckMa5sh5+Nyeo87Yx412gnf13afEkPRUfaw/tjy+jRu1X9nJqF3b4inWaj
fpIQbKUTcT/cUJXrB/O5KP1o9qVmT3PrjXMxwo2dX1Qghos36xlPizKuKlHo2B0e
1clW6ZNViORvQTjmMTP5USL1mwu7KWNBk7K7aUNnOFTVc0av6QunW8dyKvqN/b+s
H53VxZLi+PxEOV3OnNVPbNCMHoUksM/r7Mkm3MP8xvnTtCzzhZeZ7dbMzMDYtXzl
u2M6eSbb5MvNsM7L/0s8sZpGOKoSVvf3Pe0lJpDioJ4TGcgh3yAIr5IiPzElBep8
UiBomaYYp+voRmmNR/8/gFQWa3QNwTzhw/lJpk3BSJQ7FUjlRUSiNPzs77SfFD28
HSMT5IGqPm3K14Hiqh4oxZRYJnXuLgokQUNEMpy4rlWCALFXUQcMKkKC4oc02R3g
ip32U795Hy0KcQKftT+/2KDqSRu+ZgQ6xFxcw1z4sS2e+0LNo+TLYwhvXoAj51mL
8LnYOEFEz4ap3JFwK2IDkodCZwxf+fEpPfLqyuiZBOm+qJyNnPnrhDRxTLZHg0XQ
et8x2wzjBXoihmI/LbTcUEGcKKk9Y1cAXzsbnhVxa74ok7MawAZizJv/LpZiFUpR
M/OrufbdHvqfwYse235QGUPaTsMUZi7EnAU2UuYYJv1XkA+f5opOTn+yfBmnkPdg
XkbgK7HcLWVK2JVaUdMmqlK6zbkNfUzGhYiM2Fl0yBqbDnxIYB+PworMaETpcX/8
rQ+l2Y26umHYOQaxM4QEXb+Wx4as4j0BAAH71VQZK5OgW8eBmF1E/zS8UUsZJim3
MdVJlKuIeHNQXec1oNtLcvImnO973rxcEWBeSdrnaqHmuzYWinoQvh/0afYKXxfK
ez4pxir4PAiPPFYJZhhor+YzGDvG1Xh9j4HGBoSLB1Yg5uj3sTQ26rOsW7vbveSL
mlKDBcFRXGcjUD4j4fLpNekdogUL/7t2VKtfgCzLnTaWAq9gDOES2yELzCayXt1T
ZL3zEVKBlo84AGTbrSRnjLiMfjutQWj/T9MIyxdRRAxG1wTOZewCuimzBZeumQ/O
I1qT0RRxC5xAVoqiQ0C3ej21dYj6BYo9juHaWIOzdesp8lFMnGdCf2apOdYQZ22h
xXx27ThgJIHcPvxOGv+eyuboNidimCqoCjoS8At/OELhwf7p3j9zIA/i3pzkuqDh
3RV4hJhwpsrojKhN2Sbh006pRFddmwbubQQaC2l/fyS24QjjSypOZ78wAOTV9RWD
4vhR+pqTdSmC7d2N2wz6PWdJZOyEV5D52IlWUZGRjVa/imRLhbhQLGgG72MC5XZ5
ypwOb722ZPu8ky9+Kf1wrz4qgC/J3iiSJ3KqTgHC1O0yKkfD9aqy/05jvUKAz3eT
vkzTIaJWk5NLXAt7e9u70RzRV+HrLYDRudvdbV4wxWeRnRnk5+26of4tHp9gj0fa
7CcBBlCV9P2c4OBV386EVVPUOBaZX5AyFvG2bSR7lnn0F5lZTSxG9JGXvCFc0xNd
ulq1EoSPDgp3j6+oLgrdp8Ch6Blq+gOzD4MbfE9qmauAqYoBy+BgnLcINJxCmU7i
7fYisn9lchBvamadFgOSCWP7RjrZygqTSboDSL+T9CbqepVQtHidSAcWijDh9kKj
mYFWj6P18OAf6njPWxaIIufe21WOXINTd3X8jBYy0cYA91y/7fMLvl/8zGi3YEKl
b41MIl6g2KZ6u6RmcpLeUgc8wZWSJpcmBT9YiFBr28FeiYd/m1DYnOO0328mlX10
84pp8Ldnx7c/mICAEZqipOxnPqW3KIZxng/LQLPFKrVF7HZThlLXeASBo/jvQnQi
KUk8ahBzp1lm9z0d4d4jV26b7VNZaDSBrcbsDCPLJexzNalrIMi+rhVATHvb3OmS
vR3RC+FSPcxEcK08gYSVXo8bLXYDzFkIlaTNIL+QVRvjU0pNClHIBAFT1uXPXYSj
qSvDXSXZns/cYAdnC4usxSjWyNiDdxTYtBp/33+7/V7q28Kc1a7m0ahaXDKLrac6
h8QBE/B08a7DtT7OafCUO/ywVxiVvsNT956Ycmy0RE+l9dFzmyQ2MRV0eRJkxIWo
Y5oAtwisLcpVksSbghggvaaf2eDwmzbPOyTkRmj7nFJ4/Lo3exBP2jrIluHcKghZ
0YE50rGWQ8udgbDqWcwAuLJjI34Dup6c4IleiweIq21KuBgOeQbkM+VtbW34YgZY
WxVUr7df/SZxg9W0mTYeY0+eW8h2TLaOLbSXOtvP3ZH7RCJx+6+GyIoHmDxLfiun
j1SHr9EtBmSMS6zmdYcPF77bqM5+qahFfEKbDygvfU0TV3HhOm8R/q4R3iiXCrt9
oh6G8XLHcsaq7+MVYWQHRR159+yPiM+RECR6I/2mbOZIbfWXdGfYstnyDP+izr+5
dl2yJT4WgEUHTQn4vR1lvYsiK0cA+xKCbo4aRp/vUh9//aeCOwvdl+BMjlDRST6Q
2bXT4HDUhQ/BmQQEoQPFczh4eXUEKZTmNANNQtMO/vX7KrhdWvT/cMM9hCc0ZtYS
iA1JYIql7KzLUYeCKSvinSnlkDOWbmMdujQ5hkACsLUlMBXe97lw1pgWaRVC7ss6
HyuEUAObpk1APxCP0uJ21whdtKevtA+rF50jO0Swx8/w0T9ppfMXtSvJ2FnuG8+N
yoFkr0OLMvwIh95/dDlXv2AR7abyD9XMOecJQZK0zo0yStNnWV8K0eLr8Lc7idwP
2vhfGpCK5ufnnL9KJWBMg7kzaEK3PkIQFfjwSgy7ATZ2JdTCgC3QxQKykVY9hGnO
cdk8exdhd1TuXdKoD7JhdTEtT5PrH0kWxqVeY/HhDTOcUUenjzx8pUYyMepsFGBv
O7m1tbjuxV93xee6b85pXz2hOPVg+mI+iQpyOVD09bKe1ryN5CQdZB6bHCth/FBi
//Odi83ccrOzjKgIi3N5AG1ZFrFZtro471Mrdl3dUZ6ncUmoNFOKS0pDllF+wBt2
4tBzdgYl2hP/NdMQ+iHsmPc3hImCzGFYrZ5VEU5sSyCuDwsVLbw+jmw9EbaTwbeE
9NRUprc2Tw8dneIXaTssvJhv4U81Cbhy38EC2K0a0XishPqXPrwFIpfi/LlkrNfp
2Hb/LkIH8v7fv/QaD9wcnHyPS+Cewae8VdN1/3itgTtFqb6QWP4W1gxyjHx6q9a6
T84xqqlnrgg89sgKCeACGjtupM3YDRr2R1OFAe802cI0iWHUMXdxDl7LVKRn04NF
sHQwy4K2mcEHvRBqQTLjmcXv6RGqyFKJn3pQqoS6I3LqL7pkzNUAv4i59YQ0lNfa
dPK9Hyq/Rl1rd3Gdj7fu44kQ20LLgWVHsBKMqAHWONs6/AUyawrJaFNAGUfHUpB/
66HiQBFN7voPPQ4hlOH9NrvGVNhMEuPW6l2zi1A31rywa9tEmUKiI5BpzdfiqpE8
hfUVW9NAT7sos1uwVOBdjVugzMJ0BqBjlkPJv2QNB1I5RR8luU2Os5yocaOQN6g/
plqEq890l/h3cY4Nm/GSNg==
`protect END_PROTECTED
