`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4K+l0GyogAUZ2M4UhlM97KIsorri51257DYtwb4MTgyLz4MppzUB9gqLKjWEldG/
xPpsIE9ZLa2e/cUhAIzCFoDZoHvneN3j+k/OPNINjO1ystsnk/FoUKGMfNDu7RdK
HOoruCwSeYicwHM6DmwxZTsyYwR2xge3se6PriuzBrahrrYrn9kpsfXXIgH2E/Af
BNbsXVplD/1nqqXraAse/U1Q5mo0lLNMVXq/nJu0zxbPqLl/E3vGN7xf2F7iLGbT
`protect END_PROTECTED
