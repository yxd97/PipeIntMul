`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/i30Hlp+Qqqkm1JmVVYRFLN3wydBmQ6wsCuDFhrQO51MKUMhH/FHcM2j5SZesjn
yGE7rq75QXRuJB1e0458+G1anGS9oQJ9Lh/WqTqPWXj4i5cIAWxzu04nAAF1oWsV
3tklgYgY87o71KA7loaVNQbUV/SkByHg961PZtVoqKXwjGffQ5rUJCHs63b2lm24
0yyjz25vhCPHuQnqoNuFnPvJ8NkkhBkHavuK3dO0PFm7z48p6k/b3VVVUWzOS7vR
l8J2oYh7nTH49I4PBwlkzS5BbLl0zS58zMK6iFFHqvGodT79Fe8Y0PnxaaawV3Ch
3bfY+YmSzpo85wyFSXNVtA==
`protect END_PROTECTED
