`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cIHsqtSgD9zvaQxu4JzrFE5gzmuZJtMj2N7EPwPRHs5sTGEsQShuwMefvzVJSbiQ
solbTe2AABfHtqrN7OXuHJZ3Gozvbv+hL2a/t3Rxs/XkgZFD2weJSNiBuAZ85d5M
mLYIarTB1YLeAzoUGbvUilGKcc3pxEb1b3o8Zqk/P9Y2wAhgo8zWEL9RXebplw+/
c11XyV4bhQ/WuEXoJdf8rlybyAeWURhWncDkKRVtNeNBSkW/7bDv4bhyShUpoKIS
p/ZHQ19v251NGyjC6WJ+K5okiKiEIDNQ9zzwkapXskt04GNXDf8f+3t/XSrZEDUl
J7rJ44bpJWucbujFhYLXpg==
`protect END_PROTECTED
