`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjWKVTl7BpoUyqfE4OSp7UzaJyPibzHrwXweVSx99XGZo73uT4fV8gf7n4S9p2G9
tu/3lGHzpi/g05YYwscoZqiIF0lXHwISOglnx1AXydj4jfD/la4CANICqTy4wwsm
D5ySmdjS/uIjnJcrTubkAfcZebcBZB/jk4GpIqGByQIyIWAjndi63sedIhJ1h453
58C06zt7LvK+FuLzX0WcLeJ9mw+dSLSe7c1gwAvAmN2bcrYOTyDEegSgvm1+SFNv
myN5tjYwDx/p/FKXWPk+dctoGSoPtCupCf3WNXRPJneXuKTAHzMVzjR+ZLKKt4iS
423r6e0fgAIo3YTQBCMYEkKAxbspjCQiFkZo6j9Cs5wIaA2WtT1sF77kBj4SKQy0
LKZegwA8yW9EmU5494oxxKc/VneikaVrDQ/X7q+FIYqqvvehDgUpMIxXSLJ5hrq7
Dw72EfXSIJ3A82WAjttE0T0SJ8yF2/Eeqp4WhRbogo/xWkOhLLfz118/1HDvuK1V
2kIOfZW0N3aJaIfOCUX5K20MrxS7tDvmoncLCvSmEFAHGKvtjg/pc33Ni0IQhB2Z
987izV+tWXQdi8exPRZXtp+9L0U5P9x/4/hg8eMN+WtI74tQhhzHIRYHltEgQbNB
NsJp6SSb/jLYxsiHa8LUUmbqoRrYHHRfBiLL83ZC9T/4lrTSojskpJ7DLDlnsnP7
phYoKq6B8bwso1YmZ6If8vn9WnGN3yWTqPXgs6Q1pgR3ktqA/G81TR9Quqkdla+i
SJJ5T2cyWyUh1QtoR2UEKLaTnzDptbEXfG3TvTm8S4Ek/uEZay8VVvCYwVBB//tu
TP1uHevF6606XgUCGdjFT62Mtn9Uebm+ZVo2pZeQKjM2H8xtLn+EC5hiGu9sM8jO
eu2cX5QjFJ5aXp/wdq5/x4f0IeIJnKSWCKw8I2N/TRq7M0CQlgeMRinjzkPCde3J
BpeKF+qr6c0BQW5EDckD7alduQugg7ARzJ4YNf8JUlMGKayZ9u2mY/n/TRmAa2me
tNy1JvMKEqtdn/T0khMrPSnDpFIJ7yBVU8fyMP7t1t/fOQURAyTict8wKUeZLrMN
IGqgfpH7mQNlFGwN8VDZ/xiD31WC5hNlOGbbg2lkQzJdyPmMwpJePAhe+84xa9kR
PMpIjqOV9tc5nEzMHnIj64FbqdLefdtaor2CHEiCLVGezbVCST8XrdC+fdZNH5AW
ebQdmbLr/ALz7SuYUMWiQPelsbwPTYbdcOsV0mRL+yTus6O7YGi3iYlniygHccae
jCGPbcgPUmFCYNuq28juR/XtwRYXQo2kCFbAoA7Xu4HTlMZg21SlcipaeQb1nmqD
w7J9sY0/fheN0yK7h5Qb0WzIEb6RpfAbv+AfdHxjjlk3zRimDAU3EBDsmhyWAtWV
BvlL466FePXBoUzuaqaDnJANrpfofiUsrTIzi4fJg4O28lvA9A/zYWRERegWu5fV
w5sLr+2PDE2V1oyyoLSDONHsZyXs0BUPoA07GRrGcEhqJcAPsTVhI6MKofQ44FTQ
JQ2ei7WZapfuc4M2ENPl+NJC5tZbQpdis6dHhk9lrtxTIpeUXt/X+AtGqS81ZhR1
nHA8Lta42RMS4szCiAgh2CMQ/FSE1NLwD1HD9FHIdVqnPwO3Uwflzv4xphEmj0hw
LMQrcgaaSgecesk//jK4gKcQfCRjcsE8ZENQLzfmcn7YRm7l9ZJ1muWOYJAujNe1
`protect END_PROTECTED
