`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9DJo5LDDfkVk3hOioXfuDgDsFFMbFMxZiXqDS792m3EFJxsdX72hLGMMMp4iYSWj
mbhEAEqKy91A0HeJY52yrj2eT2aPdIdUB6t8k/gB6QX9DO6F+AOyLKWkrRUmaM1W
d9mbdbA03o097FPMSt/SpJFS8tkijuW/OmomgJlSrqy9m2Bfm7E3FYxweOcU3TMl
6z1X7dtNLXSNwUOl0pPbtYKobReazGXXQyH1pMnikSGnF3G3kTDBFUI32MeimEzS
m3UXBDgIY74T2zulFwZ/0pe7agHWwob3XdoMOw9+eYifNXwNGYSyivpXa72sZzmv
`protect END_PROTECTED
