`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kBrZLh8udNcLAkRnXkHPYe8WwPEKGjUwr+gUXPsVJTbQ7KKd8JfVTzE5fdDa0leI
6EvE207iTlZ2SwlDiCfyMaMywGp0UhA6SJoJGfJN125CMOr0Ah5VgeM26rnL1Ctc
z9tmGVaBC+gaIN7TzrwTGs8MWm566JLasBUtzwOXj0CmOaVxGgbT7suk+flZUjua
Uj0I3KteBg8r0nDttJoXmF61qYcizWvtTKJZxRmy9h43dw2o0y/UUG3wYHKy1a0v
dOnpkgfLf70kqDxe/XZ1+DJ+Q2A1dbsSQjQkZd/Zw29kULkMAu3jiDhni+VM7MmY
qe/I6qW8e2YnjjHydIEmkWkbtQKDJ6qJa3OKFBirHXXWt4wwomeGWlofYa+hK7/l
6YaBgdn6mnfNmA6cnFrNIdndttuCwG4RTjaxssxlGxnlC3spCMmBfA5A0KUl5DyA
boaSASIzTgxcwDULx4HGo9k64vqR877eRYe0SYPgFGNWJ9PX3H0Dyqkv2ExFpI2M
JXiHscyPuPBR2mXqho5f5s1C8sh6VHkd1oh9VQIAfk7wE4LRwIfBlC5wB7iE9+mQ
Jbm5WNwqfCPoAG9Ngt/ZuGe3oxN6OGwBRXGLo2KNNgVlQIzHGgioXtjEUZdNXGIJ
odKwZXCPNTbmhfXIjAGYfuEaKlR/DEeqnbIdXGcvhqs=
`protect END_PROTECTED
