`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fpPY8AkpkCMKMDBfXRnxev2A8pNDu+v9C6ul1D9i3S+pwwDbI045XtcX6SJUYm3y
68hDEB614c5ZDyv3gjoYJkYSdPXCIvdZgggbSGI5HAmeW7RGnA8VJbcLvT6w22Iz
MnHEd+gHxOY/IlZgaTHlX3mx9cZrNqXWMfZ/RSBB0jSM3qNeYxjpyIVlU6c5jP8p
BMFvh/eq551ZsOxxXquJ5mwhpKmIEvjgs7KkfNDsFPGZcldohrGgCRI9Z/qw7yul
fWryiO34w+6Jt0cSb2pSfw==
`protect END_PROTECTED
