`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyHAx8oEae759TlWhEcVPjZDvWKggihPkTTz7l/dLHHQ8cLyhZxNi5rcSUeX7I/t
FzIT4/GoKV5i5WgadcIdhQJ/LbO66YPXSubbI9d2tE4rq/CJ5S3qUqHGixEvN1aX
xhNmehEoJE92NtZN3IJFaWSZ7U/gEltwtKCpzdRWJ32pYZakRqtzoVOkev6ftnxU
OYC5C1SCKuRw9KDzacpy56lMGDHwqLlbK2eF3AtHePG13GuLeAzhQRCgXnd3KWb0
yjyXhuE7cJjKgXHQ1ijjczhsZHkyT8ydJXZLPrjuJpCA1EDXgB0OKGnoNl1IEymm
OweXy+ZmMf0q2KRA8pI7nLGMltoE3LELeKHaL9xwmPcrMF1jJ+pdS9/xMa+EQEze
FcDE1pcVx40m8J40P0LmAQ8+i/e2Q71zQpofhG0Qq33+c4p/LXO+IT8KIlOaVtj2
z/wDUskpghxnI6aQHiE5I75BdU4yGCecD/OBHYPEbg8=
`protect END_PROTECTED
