`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PW2gIUNOLMU2tEB2KPP9jChJt+WtixMm956sNWZiSU9MzngpYEhE1UrYHUgAI+X2
z6Yys5pTr7Ex4LqEmCSlaJ3wQI/xq/R5XfrE5u5Kf9GJh3JqAV1Qibh9WoEsZV5F
XQRlBpNVxkNl0CtqQW21w4iRjS4M3TthVe8+GxXF8S7Xt7GLZhxFAikFW0o8cdba
Q/KciWAbWlXCmZLqg9tRjR+/pE1ch8uwZC/08pAFUdTnIPSUgH8Phjh0OrNWmIXf
e7n/Kgeyun7UqxxopkbvOfjub+ceT/OuG+0Cq1uJJ4O+6vKUSJt4pMIMvQ2lFlnj
VzaFQI9rB86hl8FshSC4W3bXTi0SauTKNtDjZZorCSqaslRP1BGiYBK8TjjYy3IS
3XxPZfDsmbCwRCH/cD/cTzrgxJIyS+w+SLfB2a8QQGH16Rs9k4MIwf6CYc15O7CQ
EhlFnh6gPr75XDhG30EwQKGZeW1DpHUlXdvzAy/YPQA=
`protect END_PROTECTED
