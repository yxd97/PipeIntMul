`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axDgZtXBnmiPKDK9fhgj2jJEmoqcnMYeUBFG1BnRcYSlWClwZBwNbwb0wMxqr6Hw
6ZONzhgLuEPeVNV03ju4gVUOCgcm7NIATQD++jIH3Y6jVnE2DvnnyUeZfkKfir80
2YQwLgIDsJ7lXjyhYlBMOHWcVVfNHaahZkRtj2yaO4tzXZ/s7AIEtRyGvf6CveZo
qfMpQuonUPfPpcVdh9B6Js4uWVDcHmTrWzdv8g/4Qf5E4aXR5NGXJxd2c1JlRFO5
WMyzscyJh0lrdvk5Mgwspj4LKqE4i4v82gWf6+5rfrMRME6VNnoywvHFC1jHv+OE
TkoDeF6NW5NydXnGtA0KkpwB07j4lY7ovLSZg2YZ1zBgvg0O4fpY3UbfFkjrZBPN
vg05HEhI8VYJzFAE2jo1v8dtGcsVVVCTkurTYeyy6O6aL/Ob0xIBp3iUdzjDxUO6
jorBIxCQ2lnSWz9pvZ17k91a+MeF0nFntzhU3OvJPKUF+uaQOLCTagq0+TVFM+07
pgp1ZShX0vZhwihBm8B8P0hLV+pttKUZan+rg7ZLY0fPc4eF25xqaLBy5v4l/IH7
Zc7HvlulsYBpaR2yfDABZhIPalFxkERmGw6f/BSI5zMikrTSrB4s2DBTX1ClBFaV
DIAzF4uzQoRPDCPd/ZfyNZ3GhWRDIz0gSXJ41OzlLGNcS6+05Uqd5URmLc1CUqCf
OplfgmmyVvir4MrdSl7iD5vUkzvM6fTJTvGpEpcX8ADg/ZRGw6hJe/19ON2A25Pt
yMH/43zExdvit+NqT90zzb5Zz0UkBqqpYivUyNIPCfRhr0usQirw3VW1Qqmu09y6
W+oroqLsvd2FPZe14oZ0Xpi7ajRv1Y8aNZHbJ6zxxDOx1I0MiZvDWs+cYoF6d3fk
nRfkbPdSBiwZHZayjqkZeilRDwR6JZkMswmqEC9OaCJESbV7XJLIjxVj2fqf+tJr
fYYw9CSXX7lw4ZET3UedH084CTGzV2Wf4LPqcHHFZedWR9pr2qH5pxevac9oEf7e
ngq/tUz10APkgyIwzvunPRvXa77c4IFcPY5f0+kM39GRryPST7mmhX4IwQgjDkIe
cuusmXwcJ4v+rUIJ7P9ilnKotkZ1qdAl6sJ401bWLL+rdbTvG4PhuBvqxsLUle2A
VSgQZrcxdYfV0hTHOYrmxp7LtUcsct2IiNN33hFiuXFsRPz/mV4Hsoj1vGjy/lLY
hQZ6Xu7RRYTj1P6MtF6VxSfrXtV6gbjRXwpuyBSQAhrbwttpX3mQqjvk7o4WOdlS
tZhynq2H/xH7VnwtmcfPzV83U7ziRP+VqoJYKW/vWCDXu8b7TQqu1CMy1IEF/t9p
tgjnGH4wQEHWLaIECpiZstTdcM1m/m4q6DgYQC4Hb+GSDjs1jHUaWGfzZNW68sOV
q0R5EX/h0C0sU0DXZz/8ihvtODS8D8nxEndwEP/3WkznRdPAm2oUID3vVEwBpBuJ
Ii/7s/QzGYSEAZoPmRTLnrIcvdcLjqFtfZ2nLbx3kBgMkVkv4snaCCLG82t7Apwi
AlJHTSK2wrxF9575BtBBuz/HBn1BulCULBNaim7DN6qyG46KqarBKcHoCQi81mmZ
eVJG5tE2p/5L/sLzsZaj4E0TtJyU3eeKshywTQA/cROcnsolhxzVolPJ5spPfvLH
ItcszjBQxeBvIuN7fggM8owlBLeqaWEHfpd7MYBXd1C/rPILzL2KRxdwuNYQwsnm
1KOyrB2wrtbtaMK9lj4gcxwYm+qJePzChGcYJctTPqktEfbOtUrUl7hrj5NB+4Kl
u3vi8PU4KR7xRq3wM6/75kZrb/hgS7f8/0MqQp6PZebsJHMeJ30lKA+CW7Bm0KiE
L0My5f49y6U6l5DRDZ1VuHoYXs3o4upG6m6L4W3kMDumuyaWnODMMRzGUQnbD7nt
3rzIU7H2KterRxuBsYFKXdco8idF9HcRKUy0H5j8iRY31Kyq4rGdxYp8NSTqlEIb
5ChRrg0Bl+kE782iGegbz/dEBPgSxYFkhMZ4deQdNt+pyVuI6fgnwyoxIWBx/vFL
SslTNSClAHz0CG1q7qT/lt6yrpPm/vC/dquUYWBjcAe83d7bhsuAS6BAio0fw7zj
Bn3oVjM4gmRJ1r61ENMDTD8ar1HbqGyu+PuVRYXZHY2R46TzeoQyrO1gRpiHFp9b
sv3DoM9JAJHXYEls/iSsWOk8KhiHGeQnzdXU4RUQnWiEgLNi8q5MkgPQCJxiIK3W
MUOsGzpzArsAPwLkgRkdKlUbtpTuRbq2FwzMHwznfknt2De9jJk5cDxXzofkYOMS
5VikjZEPaB0YTXYsNgejrR9f9V75RrL9na5CWvmKEsBjgQ09TBV1dLqRHYSoAVgh
XeVLuHiD1YJ9B0HtrWqaHWacgTqz0OqpgbWqSL4+N6a3j5XZLF6tNCrjcnP6faep
VF9Og+lIE6Boc8ATGIz7ofitkRxAa7A3YDTbPPZJ6e63RAZgLM+Zd1pXa/ZSnSGn
ujSFP7OtwDCZm9fs/iJf5sK1XM1TCojJwK68THw8n0qvyLZzW+7m73C1iGtpepNB
dt0neU3KGVMFsgc8NVjqJEkDwvXZBmO3ppEHAMRg3aWo3zWvrhDVeaHv2D44I1Jx
xknypYfCuyKF58nGwo1X0u2qeLTCA8iWFVso/+jSpQD+/KeBlV9z3ZbTSasDJtZB
BAuwvOuhxOMKoclZcsgIqhaRLdJrnwzKG4z0bK08tsmRkwQTIbESA7aN8cbh/dWs
AKHt6bGVZQFWOxCYgfjhZobLD9guuZy3iOt6AEK96xbtfjXNacr1KrxYX5DFEBIC
tQzLpmhtqiCK2YSycoV8pQH8jsY6WPq9JGZtAdEHaZIknyufqtyQVGKw9n7kAtlw
Ok3LvEpWQlQkx/HQ5NHXLEnvM7HdyUAzAfnr9Gai2yNPfRjfNJmU5WqgXh5gcRiD
rlG25xqNa/QlTDXHNyjHhQ18BBrX9S1L4mA31PH2RCBOm73M2xmjmjpuNvxqM9y0
+uEANe74336N+0XyhDPaMQj8dZYIXza09aUEjf2yE6MDr7v5LZnJU0MPtazJiRIQ
rID23GXr3Ni5MnC7B4sFXWGzq29rDoKuR9RigYw2uBZz1BsJhLkXC2UHOAUYP/Dn
4ZK2iuq8DE2mlMTDBOCeGHqMZGhEzYLoQSRqqotyk3ie2NoMrOGioT/WAPoxJi7u
QEh0IeH4pFtb+k43gF9ALDwvhXNQabtrAOS/iNvI/rpz4/EEECnky3y7WKQAkoSS
6kj2GJXp2gVbEQE5YJ+Z3n0bV7XMmDIv0ByC8eAbrQJoMAqwbvjB5plYFanCRiG2
E2e3/HpnPgk2O8OTyXbpAQ5STQaVWXuoakb6NywJD9N6I+C5KDH/cSSThEHyvJ2D
tddrehBNtyi9QS5V3KJ1ENyH0ru7RkRtbys+UoF9/fAsPAUqVmj8YhRXyuFrHj10
sHg/GYr97yzxsZEQgiQAKWsbroDu0op9RiMJeU4XdPfyrtEtdmhUMwGvZhTb5uaN
05UjnHxN3x8/sEO1q1YuGn8R4FrSBzYeuzIugAb3Ky1w1fsIzUBpheYfZg3OjZ3W
XoiwpQk2HMO7haK6LKBSEfUohSdOZ71x/Wuqw4YA6c5PWnUlnZ3fuL6yEX9PEigJ
FV66ZngemPC+vpmgH2XsSCCOhBEbTY+LvIL1L9Dhpfaox7gdJ/Iyp3P0XsIFuNXW
qczEgmR0cBHsp1ShRlrUcP1uE/lbNlRqWTUidbNa/dPX/gRoR+MkEdR/fnV4KW8O
t0X542mq5jhiI6pdaOqvH73CUKp/RtsLBNN3FBDgUqkQozuSZ9JSI/5Qi7JFH8KZ
JSr2znzSBd5NLN0oif63U6TeoBeeaQS8n42O0Ybtje1Q5HbWcAPBjy3k2ZFmcHbc
ghhkKCaf2NuL6yu3bQJBm1ILNcC8YykC+j7VxNDbdYX7BHuZJWi/G+nEEt/8QhD4
yCONsQ56ypq0omWgzcgrwq0vx7XADsWnJzfXAwtb2t9zpzP/DccJhC74AS2+NH8j
iP4eCmteEh2RZhyEn7jHSKfldyqyqOzbuT5eRs2+3xvjlW4m06Xo5+NAGDbiZUIU
TPjJJ2BvXdg1fhhaa/labHueWnxHxXDF9y62B9K2GMKOHtXcKFeR6HLnpf03Lh7J
Jptb7E13VuA3FTeKneM51B0Oo7mvougpfKzFJBallVenS4UWh9/OMMNUXDGkbGIV
2rttnBxOFBCWLtnvRoVwAkRTAJI821ytY5KUjU+s118UvBQ8qC79NfT7La+SO3iX
dHYcC5K1uoyiRoZgaugMVsblqFfY4rgotzXvxKK+wp2h7zDqEbxqMIYW3MLCFsT9
f0hHm8t+wHDul9wtjNxTgLJ3a9hJ01BNj+zeuKvz/H3TwVo+s7L/JEv1uYrIWUR7
nU42V0wNtw9L2S8ldHU9x3wAHkCtcA4cwm/BlfoW3yBxGekwGBl/K9S9yFgujfI8
y/gcVgFR8EerLzfNQYH0cZ7KIkSOihkFSTN6/IZXGAfnTzNC0Kg/VezJ4radqOM5
YCLTpxdhfxwKTC9KosLjEsqyBR6h/NH0+u478O8OPFEtuzDw4JJkuNn2/HdZduBD
CZWWu6crgWjYMaqQTAHqrJVkdcPMMnZVxEVn9br5ahoSHCWFh6/kYxzehfuTSbtr
A7kIkMHsBUJq0t+rLDJkzdAx35qGFU16w7RVjASXR5lFMqfO3rijn7UTRmnPvUwR
lKZX98J2IRQdc9QX4e/h9XnpswcH9hUNZf1uCs5PuHyZAtUHCWajWVTunH42bJ0i
Akufh+1O6brSoOpcM5aLDyMu0NiN2g/8W1c4JkyVDrGP3iHz8r2sPXOTemu6AbkU
gQEZpiW5PJFj6dpQUv6FV3ZVfzyxbTDCKhQiHCCAJtY+LCaci0vtUGikp6gkTMss
spMGi7x9FosladuniA7lIlbeNXCJxvTVG8xix7djsP2ClzDO4L7CC5QXMo8j7jlP
DenHpVMb+oc/VWlBssbPMaQnJqWOidTox/CgQLKCGAtOZwbleGyxMG6R5LUfqwML
e3lGQf5JZ/LKt8bMSVw11GEU2Nq9unRtjQvOOoFIoN+X5tdi5hWHZhqsB5HGkdv2
gIpurCBEGp07csqvn53EUJamTyhx+chjFvM7XnryS+FEp13e1A0qwOxJUg0ud4O0
XDwtuIPWpxZ6JVbrtWqPZNyL06xThgmX8oCjXolK1lR7UNMbjqRyLGeFywDjIaZk
fkl40Z3RouJpm24b7P0G54fYBkjKNm/tgo7JpVZP5QoBqBJnNTlU4Zw4XHnBE0Ke
cD0WCqHUSaFyGNJoUuqfkeAqLSQgkxBSHhdoQV2aHHM1B4CulDA04qCRz6gkpmnG
eLjaNaUU5U+61DgY+eEpg33xmFlBbeLAJRu5v34WIxo=
`protect END_PROTECTED
