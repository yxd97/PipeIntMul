`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meEMTO4m1dTt+aEj9iK/y5RcE1yG3Bdr8db+wYNycN6/Im2pBwfWrftnxIbbS156
83P4rzBjrIY45pitWSWvFZjJ82Dly5KnkrPJM54KbCf54KUkY4q5DGaRrEtPcWho
RCICOm1P6rj2ALqhWrfHm1NqCeW/xG2BEY8j3WU4TGAxL0nTiaMThZm4mVaSUhv6
toakb2oAMRqhf7Mx/mimsVTrxG4ZbnJvfIRotxZR7fybcYwPtuWZx337tsMKnvtH
/AD3gm6s/GKUiP31MA59iuiQx0mJ47HIIg3+KWA+40P2tJ8a+gdfJg9+4IcFJrgF
1JRS3Aa8PVV6ODTC35SlomZZ1LRV/N/PphFLFYBL9nGcb0+uf0sKajDXmFqSrxlH
hpsmEfNjJcePH3ZOXmaXm4NscDGUVDnhI78MosPEMLPoOfkjspMtno51w14QMaNo
mG+QUvfMThq+/UOwhrS+V5JA0dRBY7x8O180HUoEXacvON66T+JnuKHKOrPZlh+O
v6VNvBZD1NWq7yK0BQt52oPZHyTOm+UqHz+IS0G3+YNfL4dYtx6FIeeX9nMIXFQG
JPN2hrI7QX88rSV6Vwf/MPEaJom/Jl0C18DIhAC50SQRBvykwCbXS6ABP171wXFI
jFIb3GNuGCK9saxl5mMs+bES9swUC7w5MMc4NvIlMcHpuqoVvp4Pl7OMyY7ZRNKI
fGGzzSQP+cWhzYufLdKdRQWVPN9vJ5ddbqf3IXZN98kaaxHfyxBUjZYKlOgi/xym
AoKF/yCWAcCD9VivKxzQnXq6BcRIfdOpaE0V5mUcML6ocSmO0fppZLo3PNH8gO+5
PXyY4g5x56akzwH6MwzzwA==
`protect END_PROTECTED
