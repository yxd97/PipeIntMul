`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZzZCH6o2Jkq/7Es5tnKFRFX0YW4z5WqOjyDbtWIEezgW+Xs+E9lTKAt/pbnhAZUZ
C3hqeBfM28CVQdukVIAxYiIfNsEuVP05pusYwAW5q7r9O9pMBPILf+33ETndQru9
gDE2lDT4xVnUUyGKdEbPRLuKU8qCzsP2SqmhatgeqybF3qufWJpnXTSptEuQDz2F
WL6+4MRa+o0lpV7+049ztcE4ZDduzCnHnkT4T3ko3u7EGSFfsHMSiATi+dFI8rYm
WyqCjh8vYvF420uomnevMSdHI+PfFtb1RQwQKQdFjAL6/KGvVNiGw6/RFFFN0HY5
`protect END_PROTECTED
