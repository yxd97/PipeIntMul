`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J02GnOtu/vBw9Ls8MdvJU0Jh7prG2+roWs7cm6B+T70HnL/TDKaC6o1VOX9UeNJe
hp2sOxWcfvRP7dPpLzpWOtdWjOBg34rXS9Sz47x1XidQFb231cCoY+xiVkjDW8b1
UaNDsYS1fpT6hLJ31Beu+pEjetGDda+gnPV2vBBzWtLeuzMtZN4l2kf3FaJnovzb
DSdHIqrVAUbJ9cgtzilUoDZ4sqPdjnfopR9N4lBb0u0vBCB0RSBr7bj4R/EoqglI
4hofCWubKuYIZOfo5IvjLw==
`protect END_PROTECTED
