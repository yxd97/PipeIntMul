`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WLA5aKBdoRU82tcMw1v86pxw1G1hsz5cApBfriqMHnk7imhr2YnsPrRIoACw/rWV
v2mtVFLzmtrTjlwIyVIj0FiYtA8GGCJWyHBEC3g0XVZYS9wO91WpmNLJuX1I1D5b
2rAe1kjlrxQ/Pz+b2dHsiV51/yX99NpG/hIpMUMEOJRHwJSc3qwX1PsAC7xsoJpD
jjkJzE/0FNrUThqwZB2+HSdw4FZUoKJJFEg6PinfO1prYdbbB9RJAH1GCt6d2umc
wqsS5SjLEeq4bwdVJmplXoteG6O9SAak4BC+dlAj7R+1YicJFLsQVOFEd6EH9m1I
TOpDMQebQx4N7D55CC8duGGb9KvADN/peOu/CbjidkZejYYxu4V+oDjG9oU0Pv7q
OBGzXB73yLkEADh7RaHuYIxGuUUVhu5D+WlqlINiWDt53RfTD4S/dEbCaPH2QpyC
wmlPnNrC+FIFzmNLE/tuWP6plthj2J2KB1r1JmXgeUvqFPGWN/hAYehfSXiNrVkY
nov99nTJ2pFpg63gyVPiBg==
`protect END_PROTECTED
