`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5paiQWe6mN5GVNXMPTRSVkB5wDMR+YqoRuYSk++Ml4hVpJhc8sFgnPW+pCoWAG10
j1oxV6Vb7C6Ta1Fz8MlFwnlQ9D6P76DfvukhamRWRSUko8ZOwuA9pytAs8r28iX6
iN1mkLsXMdHkSjXfg3oDAdLd9X61GJp+t3IQWFXYMUPqX/AuAQerOQsV6Sfe6TRn
qv3GrQqKVaQlmzPeOf2lADz5lrfuCxHGUu9Mb0SmwTKKBNigHIQtHl6ufnuYw143
uUXJbvVI6LC3Tt6yhDOGTWl/dfrvfjMEms4/RqqOJg/slsAtOovW+eO6//gX4+m9
Vp1c18ID2FHrNxIhh1uiI0fDGZnYx0A4uhONcGj0bY33Sc8CkymGdnkyn+fI6oWj
PIRdQ8OdFiquwArEro9xDO+P7akjVPwvQw4V2+II8/+dErtjuz2AzKNX1nDE0er3
OGP1+DvJ/FwYeltTSv7y5aurQu0QkEtpQabbTuKN4cYJsWCujaXpm5KqiLz79RTS
ZPefDGYLLdFg0aYQVgLowbWeDyK1nHmxcSQgwRX1iaKIZrNx134UF7evL2piHDAU
T1lL+L0alHFC1USO18bl51O6RHW+ElstwTtpzxZ9fwInvCdWGlcxdQB4nPuZ/erz
tMqrdnzy339nSfwc/5v2L60vA9NXCUbokz+xgTMheW0StiEafqRjcD9QYE82Bs+1
bUMzy7aLrR0nlFODsHTFkQ==
`protect END_PROTECTED
