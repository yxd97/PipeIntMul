`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ndgoaw319u98UVPcbC7v66UeBRj5l/HiizeBCLN3SpWRbr4faEILlHkp/xGXXMn1
704vo+vAHrGWYizbPYkaR8zulFfrW5LWtCA+/da8Kwpz/YS9S7YxRWzVKeUZgAbJ
w7MEzSQBQHw7Z3TiyQVTZCMDOCE740FB0YywhNbN26HL8FBZnzxaH5L5U9RABqe8
iDJvjAJWYqAueo9vn5gYBJ823lWBBKVZBoPhKodYsrN0TTxABVGxp6+K7WLkRc/I
7ffquESecV1dOcQ4vVMyzXVMFa48jS/YbuPLWKNiw4IMI5rdlk7qZ/Dplya90fzK
l08Nlun+L+dOKve/3J7L2BhUSHRHRqSixEw/er8MFPhjWjIIFvLXr9mxluUGH26r
N5mcsi4aVDX4gfKCRgUM3OrLlI83kqKvJ/X5c/8bbPM+lISj3fuqNb3i9VqOpTz+
fcUBUUhAcu0EZYzGTdBEXXCaRG0itnikowQ7hePpLU1i+/cEG5AimPNBlHUaTtt9
4+YajzIaVhP+onX5NTVgB3wy9wsEir3U5W/WKFLel/IrMaqdcytsmXasxJnbPq+j
I3A1tp1ybpv4dEO/JEZbDv/zSByzsG1q11a4tRWpHKUB5IF5aO0QkxYvyGAdlmTs
/HyZWolRHmzqTup/t0AVrmtx9ZtHrU0E0C2WJBgMev7brb48PKdBq/WppySQSbxn
blG9+ueBOqEYqzHhYHzyJpjFBeZRX6jp7fEP7VBpoHyKHcTEfkKs5DZLIlMwLYHb
tXTYRThI8FpvBhEzfWKMJ0o1sUTrP7APWTk59NZSiaVT9F+H2Ez1yL6C4h59AQp1
T4uNTv3OSotfNOiqOKh3bpKMth/k325vixERVZMuNI7ZlColGtH8Gj0NJrUElAxM
JqbdSDSe8WGDQeTTtJmJi8bk+d6a0bUbZHUR1cIYHP4CWDEvs5BZn1VHjm9og6eE
MFL5/4U4rDdSepv8S2do7YSjMBOxdhLJylmYQG7ovM8pbv+hnJZ/hg2PfE/GzefA
Kk8/xf+IGlMAnpIHVUJHIXVXN3U18hmM5f08TJOZv1QL//TQatVBgR0tLhBdnJBd
MTzcpyy8JOJItM4e47A3Pi5V6GH3SXJtD33FpmOBBTSlwI0mCvkrPgPKhMuvXH0R
QLbAXDKQkGygj3fe7H+/Xez1vj27Iex5Szo/DmtG4Mpuq7r9mfwxxaSndBhZrI7D
LajDw6o/DqxTW661XJnMQziEnfBZ5H/dIHBLyNSj3lppK1Vo2wPHAT2lAciSivWO
QolEt60rnQSvHCBVeBsbMSe55QE+BkkNCAo3CGxcPr8Cpyz7xuBHmQX6iUFep8xF
iL5U+p6tYP/9Z4m6g/65qIDikT9/2KhtDDjqA7ONol8TbnYqmZtoaQVYGW7Z9yzK
udhx6/i0u+cqOzco/mmyQ0j5S2iSMbppqom/fIZGr1Be+YlkuaULQJ4Yoh2ErOpW
mwUdJ5u5ZcxKlXZSPLytjhdry1FKt0W4Qi2pizePq0yAhNu7Ma6peRZ1coeaGJgd
Ktw3YLpbuqQfXCha/cL2cSEdqnRSQV7bEiETUzZ8BLEr1APyB99Z8ylP6nO1mkfF
c55dGvLaE5dOIebCorjy5ttesSTgNYGxSyHTrzT+usGk0QDi1YeUig3kZsB33Chq
`protect END_PROTECTED
