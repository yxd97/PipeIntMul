`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PLbxThYKGvTG6sMMAPaNHEj8BLsruDmspL/fpbRlqqeGI17OTEe00gi/BfzEEMX8
EjrOjCSXF1bGtUpxWByCV/5qwgR4vRNuGjfkYk7DGuIvSBm7JObyyIBoTWyiMOAZ
nms5VafhaodRSJP/xiK0S29/D49ZVxoxQFkHoDkFkPHTALEr/W8nX2BO09L/7ZLK
YBssRFL4W2FBeJYCNCaG5F+J0W9rO4l+Rabru1kqhn1Q0edq7ww5gE/GLCwXchZb
h8eKltaKbWlG2LasZqiEsNUlAbdYGngHGIvaAQ3NM5o2hfgLXnO48K3YjagLTZCu
NcNtrszm42KiS2KaSlvhLbrB3CGQqslgKzybOckBBOlt+a7b/EKeXBNO7EDYFVbj
+D5xct2mgV6bgPD6DwNW4gBPVDYMchcjkS84yUZfz8fycS5YbpQzvg2oALFpIjTz
`protect END_PROTECTED
