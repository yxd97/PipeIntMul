`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKo9qOhM4iD0pw9ljFxWECy8Y5iXK4lZPj/NDmSs/7qgc5q8B7Pko//8IqJMOTAq
gYp6KdIlqUMZwf+JUQy0bGqRsGiXZhm8QZt5uGiDXZQ+icE25wgpiyMY40ctnLUu
MM1ZmPZh4ZGfeUcT6CDGmyO5EPK+2XtNULc0Tp8+8esZWNiaIJhPrxSmuVqkcH0d
EuXLZpt28o/D7P15Jah7nygbsI6JkpCTTZfiLaOiiy84S/37XBHdDlo0N7IwYDQu
gYSXnQ0HCjM5waw4tLbOBHGPVd3FotDLjtlrrprk3oQLMq+9mv5YdM1qXJSpmyyi
+u5LhUlF2d3YV5FhUcUV4ZBBIRO0oz37uFGgmO/Ewk3EuqkxmNzomofin0LHhSJs
OOTZQ93xbhp6Mgapa0L1Jkhl/jc9lnRTOta3dGyC+x1y7zHgGKaUGj1Cd2IcinPo
ciovFqFnzykHh/Urb00/8g==
`protect END_PROTECTED
