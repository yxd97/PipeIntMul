`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QkKnDD5/z2Qw5Xjtr1jdXS38IgDchFYTms2DcSvzE9cpkmOin1Qz4o9tBdMjxxj5
EG+RecFoWqQXAU4mav436rpuqLu+ITkvmHCvL8fpQkJcGNIDCflpjtbV2FUddoVd
FdjKhPSG04o4KenyOm3Yb0SZj9b9vE5pbafJai2KFwJVsEgOhVyVvakzsEgw0YpD
ec12OJkqNCf0hCXpFMsUYrggeSukiyHYWwib0QFsG/ghGYnsMkxNGHWMmTu5hE/T
/+c3Ao+iJyx+VXXmAvQvW7+xCSReemxyx0wgM+3nxlV8ovWEalV4UrdDoYBmpgq3
UjsWHtC+wtGVYpT7ssGOeBoPUDDlK9OrgZcLeMUZaEc5O3f5bgdbl7TSNWVLJKfi
pZH4gnF0Fun67TF4FRjRjJTztjx+doenhgv1tTGgf2MAT0AD9G4zU5ag/Lw7m4Y3
SeON3nDj3GeeOSWPJBZO7giVlp/jw8SXYQwdeg1vMxzXcPIA8+YrIOuHmEdn73eW
T94iVq1umy39Z8whBJ2K39Hn6sacaz8yZdTgMeFB2tn63pLDMrVoVlZmtFeRji9s
y5S5wXNMbx7UhN6ihNDILMOijaYRKRFXmtgZn710nik=
`protect END_PROTECTED
