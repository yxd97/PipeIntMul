`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gx6fxhcTDY2/JIKEG10/SMxnBNFEHg2cefQYyZKlcK9JWyzkOp7tP9Jwi2DpwEEe
ZULpTwSnY26lVdWuTP3PEOWEgjfDQNCVA2uwnFfGQstgmHzBBKNX3yvC/kvXS+Qm
xjBaasFHCEmcIncrGpsDAvMNXWO3qIDcmEM5B+YBxV3fgYqAv0wsC2gY8mzLEg7u
++HuVfKqnAQo0ZlIx8B2RFPyugkeFbSzS3FB+BVQguDh28c2jP+4OVi0Ivopgpgn
/Aej5iq24g1b8OpDn7lwdlKUIyhA6MntcJZq+kmzEzxAT3K+b+cZ4wqQE2iUhjO5
7U2kozMiGFV96l4TZ6KF5IewQ9e+WNpH34ZG2bqdWiEIehTXgP3CXY6lb8OG3vKE
wVV1LdGCZnp/Tx4bpWBtNYp0+2sFkvAWSacLCYEu1BxQ7vCwtIYqOV7olNe5fWyc
FaBuDIxyIUUJLvubmyhksqAMPHRLwEooElHAvkS+z0bAJ3iLzXtNFcoFAmk3n1X3
bz+WSpC86rfG7p3y5iq7UkD1HAEPR/yYD2qexk3JUWbX70mBH8gGxrYQVs6zyn1m
4BgdimwE2qvPpd0jZsKBhWWI0MsodtJuYITV2vYbFKV/tDHdO90ZoATixcYyOmul
0QePW5JDorlRN0tZsD7ihA==
`protect END_PROTECTED
