`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3UYSfKQjaaxTlF2XGsYtHIX5/dYASj5Y7GZ2kpM79eTzVBnN2mgsQOFIP+hycHvx
Ap8jITW9Sl+AHvfBVoHI1VfBeltRkD4mUcCk9J554q/2Lih5P09BfO52RrhHD1PL
pPWGUfai0eSnLiz6JAVOLOPrx0VLRRfAfEhGA6mbdSkHY1N7EMQEooBHFmQ936ve
Z7L9zRI7gBv1KqFNEQi12vaqyHys7TQYdEcSo9OEHjUWZ89DujWvrkiVza1NyGFw
29qdklfpLKqn6ft1FwA4yyzGFnIwQr+UFg9WOPlwwnwgEiTX+S8d2gnFqJRhX3uD
uKkA4iR+bepyryjlenKdv30qT9MnKnDFR7mlL0dz/mdtnwtKiqatkGSIkNf3mnCK
nPEm0dc1BHK7Oy5j0CiBYeQ3ZYK9h0VQBITxmtMRPEE5UzA/i4ah7/HsBu0TTTO5
Pq56Zfqh12rqUXElTp89ur8By++vXGMnJNF9WOnevGDdwr88BPJKcDBxAN0BDZp2
RLaHwRgB8AoOOdTj6yo1SrV6fdWzdOeUNeR4WOHWpTG1JgASe1aHUeKgIxv+RlAl
PfeZy1GBFyQQudveHSLRAq6KRm8QDVHgYdch2y95dv/GU3blyi8tFqqPKM828+RD
8AT1O6clYh01gEfjK4g5dm8WGR05ztQdNu0iKSgzHFKMoOxuHyKPg4PtYRbTiVHa
ZFAWqZN6iPCA8O+s9kU09gg7Mm1nAgDufQaboiV0f8bk+owuesTrwU/g7rLPejGE
XncejeCULJdZbqKynFZVYZupr7Q2/fLrVwPNJ6dL1vml4wNcuUpA5gxU2zQZNJpk
bPp7wPkEcAunSzb/Bd6gtobWNhy4DUKakRt9qmWbe/lEBnS7/pcdyhRRcGHSYG5I
y63ODHDuHAhZCS0lGt/Oxelx3rkPS37p0bWfRKRUsq2GGvBNx6a1NDS1TTKwupEw
6jajxwhyX0aKcb+Jezv/Ba0DBFUb1ZIBE2Ml/pqUZ8D+hhs1sJBl4Ni1BjW9rnr4
hmimpKz/oAhzvPgb1TuWIfJDwNLEU/sCF+P7gpulfnDzMN8mjUQJRLcZY7H0vmFY
Ij3Hcu1o1uxizmKfyWqVTs8QYrm2GQKCxWW3r6acXd7VV2+qzN8l0xDt3qedyeZI
n9QD9020zDeJh831hz4EG7Sr+OB/OcFyfdQ0fMdFDUAZEq0FhAeIrVblyas5MyXk
MNRQUtSsQXua7ZFBH2DTN/fGE0ye2VinUVCjF7LfO7F1aJ4A2Qp3MpF2B40cV/Rm
7VyvnuqSFX6iVlysUdClYJWXy1BzWLlON7WkKmhfluLdM6SQLrR6F4cP10o29CiZ
0GsE1Sc+jzkUa0VXYRNwlchTyTFxd1Z7DCWYVU3D1qQC+m6BbmCOc6bb+q034hAc
tj14ujeawE5QWG4IaTAL4aMLyI2Ekqiq3lQK5sUWop4Vt0dVqEgjU6puH9+1O+yA
z544CuNuGCA8mOTKP7ZWsTUVaBXT+xTKU1uYohvFaL3+ujbRBft4YGe/ue1FdxLW
LLl5apA9nSHmIcanb10m4AVPuv4Y480RVqG0cu/n47T31hGcX7Kz5Hy/GW7Qllwz
Td56sSOINQ9b7m+xbcpdaUozNbqyVyJlLtTvGcfxt0swK2UTxtMdf7ymfO7JL18d
VUnh0zk8f0cR3AfUqjSyKM3dRqLHDf/QqyFHgch04bISvmorPP6UdJiRTT7ej7s7
oIVUyV5O8rbSC2a+w/DRqVBft3cER7AjDBIVVUHIceQeT1gUOX4O+GnwtV3IiWoS
EFnlMoCcqJTu9sMg10Vru1ZKYNe9ZCsqL/wz+5lIVIw=
`protect END_PROTECTED
