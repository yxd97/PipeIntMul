`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QQx7ZNh4LIsApjUY2/ZUtSzQ21R2FtwzB/dUD8dWFAgpACohqVv2utaEtnl8zC1a
yOuMjk2ihkfuGbcJ/PJfv/YYNgMRvz0mWSRl9q6yTTd5sY0tY+11bWCa9lywxbnn
OU2z7GwyRjwERT+C1acc85EcHpR/jN50GF/HEJUWxnVsWY7uYo8Pgr5XF7yUYnId
At8OazysTWoL02uPK30/hqxJaqNTLWF++EyACuGM4XLcmwrh+MbVQvT8amOG76M7
z7c2z3u75//WyToHSwCDYxQy8HYXI0NVZ3koNAvTCrTNILUF1EXOT2dzfR9iwrbV
Orh6nR7rSnF5pa035pXIAkjKUGpP3XFZA0FsH7n06VDbgBbO145ZOTVkx/Q6Qd+b
Wd/9WCwWy6FbcSemQI+p25F8BJgS3RNOSh+eMpykhj7sfvC+MtH1nQbBH/V9jPAi
`protect END_PROTECTED
