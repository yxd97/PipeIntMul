`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRZjDC5BFD2J/JtibjqHaH9/+aJvP0PpCaifh/FMseaT7pDacOtK6dKkPWKq861z
Pk72+pRer8RNDu+lcTfeCZ/N+ADWji6ltsWcpZHgMbrvzOB6Vlp4vs+hljpygfZ6
Dj3rsxpkuVFgTYSOZOf2p5SgoA2QCvAZciX4hFl5lV+HbPvEH2AsznxPY71Ha/PM
wHoUlQ2hAMVEa7up46y/Ku8rrsSnbM8tyvo1sZ7pASawfY7IsAJWZGwV8zd9vF1i
hXIlOH9SrSI0wB8zt53A61vLPt/oWfkpGo1FGkA1MgE1GJ7p1AWS/4bH6gnq7qVr
FpzNJ4gp22KWSKdlvrwqS996XYE7f38X1nhIPOmHF8HoVNptmOwTAT5ZYmWYw7z7
V4AFg1+pa0+8hl7JoALuKdHiIxmNwAvd7+oEh/SQ2vFwr1UxgIgjeoEJD7LJlMlV
5cTj7NiDKkP93grM2mB5m/ph3K6YxEPclkn4TQ8ZolAw5prLjTyGf4Aj58rjYqv6
EVJ6EZP0Ok4GR0Ad3OaxlH5qy8dDSP5YEL+V41+Q6sa6yX+sbtgkypAhKWIoR72r
Ri9e42arlspWQruBgF6JdHNadv+bIHu+7IjvaWzj24EB3aGFfN4Ly3iq9tGdD3Qa
lZKJbt3OnMlUJQrcXVWsU/+aL4IiNJXQjgN/NfmyMOxD1NHJZFkTp1E0q3A12LEK
miKn/nxhXRIhukCb0te1HNcZ2/vEhIUdaQiIWz5oNTv1n9ZHJ0NbvxlG3j5y/YV7
IWOnE+35+CXuYdV/7H6U1jKlL7X3Z1cqbVPloF8UdJQQ2PLySu0euPxmw1ly6PCF
CATsKygb0i3cTIoWhHGgDaZRj4+MEDtHfCJWT0jpKWk=
`protect END_PROTECTED
