`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+bfB/WSEqiye/XXm8nGe4tJq8Rca/6AWSLHe1HSmpMnVx4RgcwOP23uBiqwN3l3
P8uf5tLysSj4a2GjxkCQI5uRlk0QOGAiij0Jk9OPAlwJitkUxQuTUUWbtIjOqidJ
+dR/dAk+hUShM+on2c1110G1bQNN8FrU0YC8dsjvncWhV2pJvTv8lY3RxLOsNykC
qhunY/h13/zU+8FAgY0P4sQixIVKcBvqnDmRkVNQ34G0HpqLh+X/QNyGesmJGrqA
hpUXQcdtaDsJ/wWofQbGUrMghes+x9eTKfFg2slSmBtFsD/A6vZWy3km4J5BAiB0
v0o4E9z0Hqy4+g5jHFC+1XuZLYmEtIupw9blN52NOKWpoz5x6Mh9Q1hnexwAxnkC
eIsKWiEMY2OT/BaLYoHYFIGPqvE+otNHg0uzUypAn3Ka4hTH06UKele6eIPhgd6L
6PoqmJSbI+vJVMuEGjTIC8lpz2axIzOCJacWws/La0pkoqU5cWOKjgOe+X/QDzf/
i3OXOO0Xaw8r3gDoyoBzxDsXZUQkCENLNtB2kUnFAMZr0UZii4XDUnCInaTmCVuV
sjlh8sRC8YJ+/gKkDE8NlArKht2na8bCPk4RcCVZ0xJ1A8gFQ1rgPSFx4QEjJ1Je
OwuSjGgYCFuS17tJ5TBpwovhkPikOCjZ25TLcqWpISn38TWD0i1dDM+AtJWOgbrm
w1jn+Vb9bGUk1Q9jq7R95ckm+nkBNroQqCHpq1r2XMUmQLwErruOPmAfFXwUs2P5
3J7/8srningSs+VZiQbH3g1ks19d36671Fbk1xhi33Er/ucWbtTFa9v5Xxcn3QMp
OwVQ6tnT4TD01qeplviSadHj/XxvdHKzGkYNoQTQNwNiJyZGYcmos6RB96oWrDit
DWSC4EucdvFUA98ChYQd/AOyf8r08RyFJrPJtkL98bkG5nBtNJ6SQ288mett+WEV
EyZBLUAZOS7tCk06NupQfH4jYBxfGl3eopiNHK5rm/BKBCeMJlFpw4Tc3V5zPQEF
AdUMzoqXh/cSLobi/UsLZSmT8McZtmU8V45TbLA3+9QeyLA2cdZ95oxFcYOsbCJp
S7sbHUkFHLAQZv/lMBevB2HscQRO+FCy5G76TNxfuGesGxhf5K5zmVdTgEkWYPG/
3mPWu1qgcx1Jn1UrOZT9ea2dKPjUnDu5D3ZiOgGLigH/+16/PQix30f931p0wvpO
nh9a2muvo260QK3acO6745N5NIe+O/fOr5gCTobj5/1gmIGr/IkjqWB+6DjsBppi
tLTXwmxzKlfXS0z7OzSJw470n4qbCjJ+CJ6f0tV2/Cjb1aRzm42HxP048NXrfVj+
H7rt8zkvMO09E1kob2QzC4o+/eiZJzNLpEu1ua+kKWbNSS8eSCik4luZ13N37fKA
il5FUtoVKShPq7sTSwshyzeXB1SA4tXQRDBtYnUPMT7cIROHqcNFhI5VabZR4QB1
WyBMxwQznItSP/LthWuGY8yq7zTq3eOPUobTa71E6z72fZupJ+WV8mvgluO1A+18
7txLGDSPAij2YkNhU/9M1LU6B2mbSlcVooo2rqYIrDGi8eCCyrQgUyUNrKmkehBD
8XdaVoe6uP7sKTZ5DUX2pDRmmvqbyc97CZ7FcT8cnXyRbr3jWcMEw6zEMFZ+/F51
AShCB2zdUAP+ix7i6UbSU+sfWnSMUMq6RNcVhh9cLo4jY4BaxN4/8GtVCCbvDDTl
No33dmxm3J6AO8Muhl3GxaEJxdaYMb6czB1dLX3twrXmflZur9xu11xRbM1gKQ9f
3DJ9Fdo1NNkWUZoiH0rIUNYFNtHK5E2jdxIgUizDDb5IUd2+G1UBEdIulKocCzHQ
rH+E94ctVYklWaNnSvks+56WoaoNCHFaLDe54M//8QWZaG4lyxc36pUP14BiZKtP
GOjHle0681MY5C8s1YivFZjwhjHOE9Xzj61ByYVSg6xki5fnhaEuDsl/PZSosNLp
0+lmhOC3KBSPFdhqk8dV+z4QysQ3kQPUIPVVhl0/seXcOWtdpHfVoFOVsqXYvsxo
K86+YKzVnYonRnxDt/veDSm4J/MgTjN8m7JaAZ8vRGGmpjMSjaBXOha57a+NitvC
UlqgvGiSdEi9gaN2EcZcCDIhn6ypMYB4XcIa6yjNMBzPnEWgBhk7YOcqEHBONjVk
7Yl6QOKQ5iXBztPufe5tl7XSM2ICSTkK6q7pooQfY1aSTOFuPRu34w9Xd8FgepAR
6GqksYxPZZonuItDnsAUYQChHjmbzTzfdvOOd9CSHs/IQTQ43DCmvX4pnA79Rprh
y18XCexikNKijepdY8YPz0JlkjTwmv1XHbZXVhaksDqT7idnv5DAHprtuNw4gE40
/WcEyG+2Wk8O9yfaQBjYjw2TL5o1GSCxuoYuUG2dlAXVgEW6ovSyvHN/K885BgiA
3lhWwSdItyNGVpk7z25zmt0NlMaV24WRGNzN+puEwDc5cpTrE6Vrov55/I6rSAkm
yZiqmOfCGjgFoHtMAs6OYbFJ8XqJ2IJzXdQepPED1GbW1xgXu8oNS/S2WOrsvCE/
f0IzFh+Q7TB5CwMthvHkZ1LzMrppNxyQDIj1BctNZz1hGZBsgEaUhEp8cdTh375D
aUKf7YgBrCfuKejJhBtfF9YTSFHoISYWFSuY9MtLd8cgprOol1MdUl8MjDOwdDT9
UIkkUopgRf/Sum/wkk7ieUgIfSJkM+YjxpHhDKkNOA9REJlf/dnWg/w/5virhuny
KCN6DdC9hE5sp9owCIA1IgHbosdxPNtZ7B+MrYd2qTgzpyMDtVBh3edr0mCpEYF8
5xy3ZzLCQEtQaA2R0dEzwfPeYduihPzP7tRCYg8ObPolfztZmpQuJg94zpkqh74c
xp/FzhRFwrOp+AAy5d23kMQe1UaJeNKXVNwv1UFVGMHCZJzrUVdYsM3RffHKs8Ol
i6PLO1uTWzDBdIjr/31uFmRHZ2EykNduOxBVNJnJ+go=
`protect END_PROTECTED
