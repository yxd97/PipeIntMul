`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MZPFWj7uVUgKIQuaNrU5Jaa72ET3/I5NBtuzTU1OrIULaWLoVDix0KYYL5gfjsQK
1ilYsJL3xrqwqC8Syze4h2k7fZXl0ejSlrfVwW512ThTpDsHnt9N0f8/0EtzpoqM
G9iofJocZggCd+Q1riXq6xvJQ5/yy2uOyl/iH4n3sJQPt/9sTyJe9+RtCmVXrXNW
wFat8D2POvTAlXSRNaz4VsJLXQvjiha59c4Oun1vF2KxzJEN79917EHSklEpaH8F
21HMxQzYHpN/eeMxl2ZM932dKg8IdOLzZuYihE2aC8B+9iuzKLcD3LLd12w6QYr2
mPIT0IrFWk7DdlDXndn52mJARauiAquWOIuOZAAQY5xcQm1GKeKmC54t2QW5RXUD
m3q5wmJWQdajgI5bYIljeKVSOyEZOsodV3tUDAjuK1pr5s3zBP1MYyftqJO5uEw+
InGJ3nlnrJkrYurHSbwF8wlSo4noVCwpFnhS0mTODYDijwEnaPlhF13wjw3SK68/
sIeO25FNPKk8dDJsFvpo/qRzbK1LQR1qp5HwFNBot4i5g8Bh2eWHzoVHzrCYAnp7
tcL2IO0KXD0Z+qEZPfH4e6QYhhd+aL+hvEWBBxE5xiiTLR9CPc8YmDvgpQf9hedz
b9g3pW2Lq39wWkyUYJDV1Hmqb+giRcHuOFtpa7/BiRApxA4Xaljyic8MHLfBUVrn
XuLKJzHpDOUiQrCmAnlIUrXCBG3B41Kv4X1ACqa4e8Ey4mOh8sSEV7Tbs9xwi1BA
79ufpGcuwwVEmuJQKB2VBrqEBGxDfCKNCbVG3Zn7+NoGhkpd/JZV+AnrTfQ1bWd6
uSsjfy4BZUdJALv0rNTg5tL7AL3k00f/3rctqOZR+49ZnzbK0hzriXYNFgKRY8rh
DVePu2uSieTso78mLkNW952ktwQ6Sxh7yqksNCqotnaDn7Kp4JfSMSd+B7kjbCQu
SRL/FmI74c5Ck9bIqAJoftVIbe1jva+enrWiJwRB0UpHmP7MadO271oZieWKzNLp
30zBhB9JITonqyTLMAUnC/PNHMWCeP2VBKzFao5rnI5Aquvix3lTZi1695OZQLFy
XcM2qjwpJSatuiT48Qh29MUH23O2qc6KJKVwr6SK3VrB/s6mrSLv7AjOqh+uOXDh
ETjfAbSlQU+7Y92+dhiUIlL84VgW2JbnuzogUW1bWl3a9l8Ve0fkZw14uLda6QhN
lYu6THtImu8sKiJnRmBe8dMLgXbaJBGSmIrdYu+C63l5mt4xjqDk71if6z2nbrmo
PQtRunfDIhUMtdUJFaiOEupKZBzHTH7JZJmioYc2msKMpwZbE1fUrb3FITtRNajx
YaDyFsjw90/fO72fdbCYsfAZ3xMdNdyxLfdmUL7u9sqh0v5I5DIxGDoe2t+j2jjm
3VM/hGS0P+rQ6FA4B+qnmoksdr/5emkqX33AZkV6TNoAwITDVxf86a/SwPKrY06c
iaTfCwQa4aeLp7A+kAO5uFxCpVcZuYqWFIXhQDOtSJlY7f/B34b+AC/y3mXRFvAq
FvxqreelfyaSYc46UyXqih2293VgIYfj2VPL+xgiApAeaUbneEjRSQs01Jx9zKO+
7LHByhgsAYBJSXJMQyb/nNUPyoSNpB5RlHpKwVXjSQ9yN5hb8mqkNh4u1fJZPRfy
WFkSuh5WPYY9jvil9odnH8RTNia2+yW9MPwGJCGUUw1hj7xK14GqfuOHs6/P5p2A
PZXUTSXUrEGjcaxJQdfvXsLrcb1OkI9MbwjYcn0wvX/0sXJlrokPLtKFp/QQIZay
DFv3vuE0jDE2JDVYpy3ZeQ2q5sC60XIqh8j8egroE700nR0hpSQmckGDW1+3QnZs
8v0kk6M4OOqBDq6kBvMOWIYE+qqb3ovDhNyf/rADmOECfjUegmo48ZTQSOdEGG8K
G0OmFzpvBt9QepuFV+ExgfOlGvhSE03W1CuAYIO6zc0Wo64o1ZKuvzny5d5WlIda
PGfqTezIBKyN61KQH0xCum/fdb1E1JZGn6c7AzPO+yNaPNVWq08bNPfaQofPy8BG
jaF0KnRevqBABO7xZ+rMHGzpA4D1TQ/6ePtTOBzacYu5F/Y/RcgUjgreH0tzh/yu
wDy0WXninnTgGkAx+w2zj4Yjoal8jaXanMBZ8EcmiPyuIzMnOgafWSR9z00fWQ/v
7i5l33Las1kcmAtDV08EhZwnUOaLMqjN3k3WufICcvKsLn9cI58vytvNpIB63ulM
jZhdzrXkINGGZbZQ4eLsnF3ncs+pnwH/+0GKLlFP26P8+Sd9nzdjPFGc9LA1s72G
j7xBXII3vcgQasFJmNZ4RLmn23Arx++Q5AHWy6YBMkornEDoD/CZbVl9EET3ozJQ
LPhWLUGJKKA7gU+aGssU/pw+R7LTDTHouME3GXot4Ztuvxm4jA6svR0qoUWOX+Jw
zCI9z8UtfjG2z2662xeb04w2eNZd7eVmGqRXihMV4i0V7NwMPkP9MPqTBkgYkvGe
gEIVujC+Tzwgsa+X5Z5sN7XQRNW5DD2zse35JCaJ0GKfoe/rFlIB3xazmt0eLTNx
BjIPcO+9Lq3he7JdacVVhcgCdQFfW0oeUK6MeLX9Qf79umxah/I5F4VaKw9aoOws
Sx/VE46UUDe7E7CEijhN7l0zzr5tVyTem7UycmBbdG/C7gnKV3JCpUBGMuHN7XgC
i7eoBli/K6D8yuGAfnNhzSMKKCaH5n9RD0mYNgiWR1EAgLDnPidc47aL1W245hr3
AkhWuuH6Wc/eQk77fufq8EFoSWFAEHddqQZROWHUwhWRxdYvuXEKKL6W7FNBjqSI
I6pLgJvRlmM4FMDZIYcSWsfY75WzkVoKJfFxso+rEPzcAMm2HIIxN630UR7iNVhj
UvCo0gGofnu2iGGKdiX6Ai3cHzx1JXwJRnzglOYbnV+IbXyCzVZwKM1SArA+LffN
UM5ev1bXwph0Vstumk1D6J905CR0ECnjZUOrktFMgHzi5fJdiS3yjP8Xd0DVwvAz
zmt1hYbbcT3HjNPy5f3n6XUk1lwWoDXHCmTVc89wFtTfOcjLfNA0KJO1fS9npBYD
Rb7NmFbOBvCvrlMe4FWkgKOWRubKT0DwxU3gIzfdhNBdNip13YtLUBVFArWu8iLb
Brvm6KWEFM+mbk3s6xQogMkiyTVQ2TxDw3gyFZJ95JfIYJi7WaHRfz3KLT+6rKgs
LkrHlGm5la3qE18O1HvoG/Eptr5NWRcjtECsxeeke8YoCuChVyxZhDEmo6nAoyNt
5tqrkkXe51DJBHfQWq3BOhcjxoPv6Ea9EHl2gIrc+XKqfwGe0Wa25ydkJ0JqdvXp
d8NyHYPuaRoJCPwkB1FROv65CJfpgcgFC7VZz77CrK4w9zgNR/aFWbK0QDpqMnQn
uNaBVkE0kGpf87LP7XBs4w4ZPVy0kkUo8CFAm/i5BZ/WbEmsjHNq9AI+nHn/ekbi
DmEhneZyth7Q5Sn34ygGYgiDHL/6ARSnB69kSzZ7D4BM/Z2EETtLAuzLpJhXiSRB
bzkX5Gv68pfdOx/HqdlXAc8p/Lnw9iiTO1FD3PDI3nmQQtyXFmGtL6yvxMlRVgOz
isXCQ+vYDkSWhjv5u342ICJbK/6lyKT+bGEOlCfTpIDCtLNct67bj1jORdzrXX8t
diiM9dYAhut/zxdcUGohraZfYjQfm5015A8HHdTzFwpgrVFkrU8K6Ly/0nyOFz3j
6IGhmOaRXZluJaHu7ip+7ictqWWcdKJutr2dM4qePtz2eshYPKJ73HzX4KHm4bnp
`protect END_PROTECTED
