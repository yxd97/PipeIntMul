`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tvpwrLWJk0F6OgPhGgfMw45NZace3eVkMo2xMDbkSjMgxzEkRk/zLZr3dTSNV66o
tTBSti+P7/e3+tNOZfYqrcS4NlrGfwsTKBHDlzw/18X4l82doYM8c0IcXxnNnbku
sV6X13YhsXBLyFl7RfDIAbiQ8FxkqAFuCo+4Bggx9mbhFOd0pWvYm9qV5bI6/dc4
muq9E2YI52Xckq2kI7KIhSLiwSdhEJELqcF/poZ29JE=
`protect END_PROTECTED
