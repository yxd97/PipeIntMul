`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z0YoNXuT88aUXSLLVGcJ5uqwV8c5v9vIJ6TnWLVGF26HgOt6U2tX+cFsnG8Lv4Bb
SCt59RgTTb6PwakVnRQkE18svo+en1Rtf/NlpJVgCysYP5bjITiWvre0YaSza3KH
GUEin3aWJs5l/Keey6b1Kdgu2E66oyuxkcRhWxt77NerRjZq11F6SkFwStQsWQx3
dQKET1QmOiu9S6Ae1SmbLYWNiOtckGv9Xvj16XglDCEUn05pgNUoA8Dnp6CWf1pX
fl/YtNxNsQWcEP3uW3mud3vjLYCncQN1U1GitHduPyE=
`protect END_PROTECTED
