`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/dKexT+GvpqMhvIE/ByGFtpIgJfm8lkkBPQdaQpkd2LRfA0DWda9mYGcp01Rgft
qDc+wcTemFpiBJh3ijIvOMvwoktjaB39PDrxJ+FWG2jAyVRLKMr6KbAsNYRyDYlx
CoJJJF/6CFaLod1QVVeXxzn0lHGhG0QqZjExcBVmW6fWmAUZ9SLT3YOY665L80bZ
PwNnv1JmhhJ21C8jXQBu88VTFs482u8VbZXmxbr/dsNlsZNU6UhmpNggYK4Z//p3
vAYwX8gSyfXVxIs3/nGxim1JUh7ePbVJhzc09pvFlEjepY8+p1ekA/bN+WsgFNUk
LibBPWDP+qHoT7NgCexteawEesr1AKpn3eUhW8sO4t5qbDqEiDluMQQ7RFC6GL3V
4+mggzJ2xKIGWn/c4NtoTcmbdmZXnsU70ZkCs37X+t1BYZGnCywBwRvPiiffDbBJ
sAlH8IRhagDaPLc1qUo/r6IdNjIvaNc5vAbKWrB06Me6ie8SKV42mZu2ZaYz9igF
InQ0SAVWrw0g9ZcT8oT/l/gG/FH7FsePhvw2IXbOSM1LM6+ofeKKSSzHmCgWFBsF
yUkSW36jSo5W8+YDTaFS2bj+RpuMpDvAanJz5kS8A0zs9kTuFx/Mk3F+srHShLJ9
+01z1Yonk6im3fEzUYUC9MEgwyrXQWg52RNFVfBKfgQXsqhClE8K4LgAipY+9qYT
k77K6K54Q9pmwdCYvptI3UOwYomfAD/pL+hmm/7dD1ikESAtDfUOigv2sztLYRd3
H4gEwzfJL6QkRYWKsYt5lxglPmqmZj9iIFNk4g2RZeJVncHxFuImbMTUJ9ea0Bty
TcQoLLxwDDGJF3tkJrRouV0dMOG0ZBNCZK5HBO0bCIWzmbFFesMETXi6fH5I9P5u
DzaU5JUVQLarkzgN7PfEBeAtndEXVyeQgh39HM9YaPYHQBGToif2fMr8MgKtHaDJ
l/EBXUJ4yMllYzSi7a7PMJbAj3cm7Ad5afpx5tKnpHDD3vx5iT816D6eMToV7Aee
24ZNjfTFZrwe7ui2rQAWphcDP/kNTFQv4XHzZCKWsJ6UR4Cd4z2LVUO9ewOYRJAY
271OCem15fUOEySR85G15V1p7J7rCWQ3eqPFHpmIm+N7oznvOfr9oUr/gsn62NIw
y+ARY8NguuIZjevkEfVAOh6oq93I/tJGqU7oFnHmxRwvNY/ROEtsWVX+T9+xUDj7
xb9budkmrn5H8G1wWzAklTPtktD93BZ1RaDBct9hNOk8m5jykUHCA54oDWif72zW
TT1ejhL1QROTQEahuG6TwCCLUkMAsrHt+cgdQJ38R2kXT09BqUMBsp4Q8/HBrPNm
Fw3EDaajXIUN1nMoHrXUUQzBD1FRpnqgy6tZCx7QMB7SwIBShN34EvAKtgDfy8VM
pUyfZpIfd22qUdo0AwTH2M2kreOEp5ggqzJ3t+WCkurlkFlFCNqjncxrhQ3Qq0jg
mtiZlOXHfJfjxCN9DNXNhGEIeJZOAOhIyaZ+ys3a4Q4zfoYj9XY3dZeXIsqSSRJQ
CMyWVJ3OM1YfAHPBp/Ydia9nBvdQl6lvQbCeojv8elD6ISpu37PJ4llyf103jGXe
QBeDi1hAK+xDPQonFanwfZP+RVUA72UaLvctzKWJZohEiS0q9D/fJtOfWmAAzKKX
W+mc+uj5Ce3jU7AoYwhVIsm8CnvGDWZD6Ut9I3jnQpBzrnu2I4rzPDwmAJ/wvFrW
ycc5lh/c9Cmc6Gz/YnihKJgipvPZSyFuBP8ozmo05aDpkqGyCZHGD7Y494vYHTR3
xkX3YhiZHiYBdj1XGNGYLvoCZFpfctWNedryGF/fCdDFg2U/1Wpitq5sogOfk36s
/fsPhUElHQSqoBQuxcnlNkz0xuAWIo8nIqKKnU8MoeKgllKGR/5dvh/w1nU1Gdha
xNUBc/UdtN5W0JBLoOPlmbO6BWCBEs6pkwwsqXQKpK3zJ38u7OH/VnHFkJh+yHqk
9nEVOGm2Rtwrr+5TcO5RDQ4WUjNtW9bxqoqXdm1YZYK90KysSbHjM/tSfWe8LMoB
bBJk9McQ86usySOsdkfGrCvrMQihJJcSciR5iECzkMxcBNrPO/iAmXp94e/cdX20
4LcWUQueTGxuthlhxEg72Dia68mGhnu8RUAJdemy/r0vR1R0Q3Bsloar1x5Htzzp
07q+LV8EubUPPYN41ExmPcJf+78p6TasY7fHFb7J0C3FYZXiqu3sSKbWGd0DghOf
xDrvOh9+dmI3p5X866zuE/qx2tiTEOWYui18AFKDbBwQDAuV6heoF16g5Ag/9Wtk
/BiPd0oY1TbfLMYaOBrGMIjCM+HFwpV9PvsnNy9iGgFMlzWlabh+pZy18m7kP0/b
RKzjYUfJFXOG4lBh5DQx4E/eeAi/agITRAPtgjNV64Nry5ZIl4VmbDB541jC1w9B
maHF6D70fs2XJY10Se78c4QwR1hcvaKoPtZGiLglyvBi/K298DvfdeT8TQDPNLIg
e1BMSI5BDQ4f98UNDRP46kq1r3O0qvxpotaPlGAqiwuT+Xfli+09fxVGThJcaFN2
17USJv+uG5CJ6iA+xRLqcnjZ0ww1f97kuoZYSOb83X+PMJhgfo6I8sgLVfI6YXKR
d/f8fknDACyKVajCSWUnxIAxhGPYYZBjkISG+7qaDseGToPjDWF06OxErxijSCvX
1xBhYj5xS1RBTvw73hUKHlBqsAEOMjFwkv/jWSev3XrKgDFo9WHoPQP331MVyhS+
rELKXuAX7at3YWCsXbSNx+OC9M5LgbdUeDwOgfZ2yzaYLNLljMAMeeDOytPp2wud
9S9rKVQVAtSB1S+4+KKfo8V78yEfqZZvMomuPiyQg5TsmeD0mXOimozuoXcGPQY4
x272Iu7Qr5dAo0Z6gXw3wBRWJ5sL1mXsBhD00U6QpbWbStFR1DWyOx6dbllIFPXG
9MzbQ1oOr1o78jeRFrb/o2nGYe1Cop/IR9riPoQfcTE8ryKNeq+Wn24AxhQpLLH2
XWmOpGpCUd4Fn0znYJNzj+ccydMoaftJNbNaEl+kqa00Cj/xr593JGVesUixom0t
13w7a1E/FO/BxPiM/nMBl/8Eqjk8i7GWbGqmN3b/quTtuYHkxB586mUxkUQPXGYf
kq2Fn4bwLmgVUkKodLPmgv/dxovY/KdoEROG+godb5w7Az+XTbYUfg9ZRx12kC4E
Dkyvbs6Ojzu7RbZj6qTlkYfH4g247kcHVBi+unNzLYmc5VsJpViXbHXNnipwujSo
12sH0XzAjA87xmqU3a2iJY4jna216Pj6Ll6M/1mPLJz9XJl1WXtNSCfwBQtuScHJ
+s1G/WdBiQwszh1I5yhvThY1dZ+4k08UAWKmJAD0cykVXPX2pvfvgBaoFrEar53d
J72m5tMeoisvB2K7H8aUZd7H0iOdsDiOLjZhOTk4S0anYRnK5qczHVQ1vH44q6Kr
tH2BzQ79mQNZipz4urDZYSHgEoXiMugFHC7p9xEO440EyfqfVJm+Ju3dh0E5KhUJ
zwlhg0zGkpaMjuVBmktO70y3+vPUyrtY4SoDRjYIRbp8Z3mJ/L8+/w8wgD+zjFrP
VZfsoFv35WEas7RVOElyFM8A2TvDle9LiJ/+vSbOeq5EIEP3LYeXHIIIF6T/Ghlj
wqC++QtPl1GVnrWnaYSNUP1pk2n16nGRGp62Bq6NR/KkNEe3rc2ISw6G2HWqH+wO
ZkCmqCtQ/oOAn5v0B2E1b15eYHjT+kKFucHodYsPCpJDFsondcEnDvKT9q2u6iJC
La5oV1+PedPLzlPZT7Knl7rXJeMP11uQC9HyjJ0qrrO+St/pSkEZoodzujCzvUMN
mo9JMlI0TBFbTWGdscmXf6kfYH/oAWi8427yKogySZFRmvjHZDHrKjtKS9CaEmRx
r64BLxNhjvaV+sHu9ZSzDi9ApdiHqtrDUqmfUbW/h07HH4bYx6vW0QsDbNuOvkyf
HOvFil//1vKvxLZEoHA+Wkt0IEeYRYcfcOq/jHFGwucNod9jXR2rm8ww3xX+HGES
cct9D8ZgtOXzGFcLcSlwL2gs8JysyRzO3mx1MaErGvvwexocccu1ce8DV+rFvaAN
DYg9SRmvl+Pj1t4r6w9LhGb0MJFRaX1vPkzMHwL2La9eaGRu4RN0Dz/SpZNKhoTf
S0eWdln3IHEMYlo3nnyJpumTNMBlbCKlKi/fkrIeACIJ6+bL4ZyTWfFShkgZPvp9
yp8uAuPI8r0wNYuxqXA04i3i0IVlhw1UMU4orYrJ71OL4bfvEVWy4yvUEaYzt0xF
VuWdfPpZX9zov0m0FphlQF5s7AEB9W11Wuz49bPvjtuRProslO15a7VNM3/6ZZDv
Baik1dPvvYh+ZDX1G+C1IaUBDMmkx9/i7dcFKBI9mloqUUOxLwU0bFBYHi1AiV6P
Lll3LkHl0oE0b2IggmGwe8YHE/jkYo0svD9cf1gLAB0iBqWeQQUCLNdeCR8EV9T+
0MI1gqVEp6y3XTww8sPPftLiIkgNNUD/lUTAW+/aGUGG4qqV/IGyQvGDAygppd4F
SbCQUBAtYP1diON7YWC5Lvq50ZZb8zm3lOyeUrk/BF4DLZoTeMoU/l28jvJJw5w2
rOix+j0HQG62jgRUzAgspV1mhokRE6d45T8cPkDxymf6sKp/d9BpGr1o4t3GWKoh
UK+dAY+MZPtNOuJ7/+esJRfMwoJarZstRidcZhHYvuM76g2UafHTdY09lJAWUswl
ZUVJV1KdYZoNYFXjzoZtRg==
`protect END_PROTECTED
