`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YbG4XHNbVtN/C5+WqJSqDxSywdvCfFT5qZMS8suNI6DKH8yATfXBo7yil9hzG0Gb
oRuYWvoU3BmmtUNKiWbHNATzk/0e/9nsZDHJ9SNK6T5qRQw04Y3+mlmQdLK+69qk
zgy07Y0MbYwcX2f2V4HG/o9jq3ATa3O53wKzCHWdLTfUnXG9pVHNPO4TEq34EpqL
Yxt2f/sMxjU88sg9RQOiIg+ARUNYuMFN43RXZYeiib9iB3pmE11x2yoHQ/t56yDg
38dxjv4iGcz2vEthEblGkIFEYnfm55nDAFy3T9/AKkbN/9Sl0s0P1eXwAJeOA+Lz
8UrGJBkIdOWnsiodD1+nHPrOi8AEXpbUJhJmj1kVn23JcgI+QYnwUFxMXrYohDWF
R8jAwJjzUOIJ5A6EvbP7s/MZHxMjlEbQPhhdQ0799nO3f12jhNkvmJuariImcWUI
Ngjo3ffyxbzJmk+0SZnHpueMfv/N0MAOr0I5wECgOCkmkKR16/rjRiBqedCENasz
cn7dgMAEmzY2te2TyCDKbFDVxtvAdNDq4dTT1r18dU5Aa/3MdB3koCfSrUqXF/62
EAAWSujgtX1py18yYquulWvWpJ2Sql2PWtqUb0Y40NIW2ZYl0/o1XAfhtOEG5wKA
3qSuDuSNAvsVYGaH96KXNMMDYrEdB0kcuL2sRbfLaDtEwBBvAjDCQrd+shgqLTkc
AmIwxcpSM+9udx3fUGxkcwoZt98JRIy/0flC0LbvyiEFLnsIoLZ3u+YkVv2Tcllx
xuss3CO7CklY9Zb6sbR1g8H27h3jdFnm03g6lKGA5kIVW/PvzOPnp59F+ulT6i2X
WUkkKHZGK2J49WsY4qBZFl7n64gf/TpatrCIG8xqTtxXXVsyVdGLUnIeFVUa1+iK
hB2Y6GAbRVbUtmwzESxl2TjMwQLeNoMzZhBGWpvs43U8DqOu6JHta5Q8yTRcnqxw
KkyVnJ26KplhxOsV9qVo7xuzwuExPJ7UCMcqnIeMiiIuWI4A6N5lvcWoJlkzvp19
QKxaISjUr8wpg4Mvoxiad5+541NEJCf62akE9I8LpSUW7skH45YswXo+ymgtAQXQ
mFtVwBG/aN67TG0LD/ZBhisT8HXf4YOYf0R1b1eJalL01fP0KkDnjfsIpSAyvER2
8ooHF5JtdOil3k2lQzdI45Tcll1w6CC9fY/fXTrrtLJsYdYRGcAFQ3iAxIrYSE8z
`protect END_PROTECTED
