`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QobS3A+4QW+sKVUUrvFES1nQHmxxA8Lhb+1XazMH4QwJOy2uxWvLeFwc/5k+khgY
xsNSYze/pcak7v4wlktwuhCSpbb2I6F8ZbTWQ6n44KnXMR5bANIdm1v+BP2zkxme
tpqc7Q8YsO5Pt+htI2EjAvkPzfEzRq4/ukcvnTj7yEYf6xqUTqmneqxB08Ul5nh5
tKUEpvSHvqTyvd8M6t44epkOTB5kBrqZDpLIshvSCs7VC7FYbqJY7Mt24YwomOGX
l73NnqKPaiMDamgmBT3U9bLDomRGDtRz0Xkle1mvCgZaw6zgVJ7nvNNmIa8MFozs
nfTBerbHyMeKaGcRjlCrUOq5gZN7elSI1avAGyAb0hhfORRLmgdF6fyNenXiFo9V
HmISYeuvBzQMnfnTI9QMZkijtKxSr5TRi1Pz3f3O7mM3qIcgZ7QFcvHMUKitWXaW
zpMHZG8Owm6Dkz+21ZVhocVXJCfSxj6KALeRX+lu7o3mlpswgg7TfiUTsVq/250x
moW5YNq3NyWEd3gr2WCDadX85RiCglQ4WunG4nCOTqaOTPFTXpW35vAnoT2QWH8v
ZXge1lCc2O9JkPf/akNOpA==
`protect END_PROTECTED
