`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0RDt95WVE4jtrLyPF/VXXArRQgt61Gohli4ox9I4NVC+fy/YeR81jh5vng80Ezy
TX1wjtOFrunfOyeXzYtWkMZNT1v10jWo7petchmuX4qaCerJJY2fAryB+mDxRZLn
KDDibaQeZmz87LTURn6YoydlEpR2T67Tk/LYOdp0IQZH+jXESoX0qbxmVCiZJ1Nu
8ANgq3IyKjiuc57jG9HvYQldA6Rmc0IfshG6fD3Dxw0Hx0TLEObwwtOQY52RCXFT
t96MlYPjPggr1eTK/qsOAvlyEWFhDdsimBHCrcBZ4zCuyf+B0kjpEpgIim4dm6SB
GLY7dHixk0aQlb44xq6qCyx3CSd/SKbe+epNihE0eryutst9vGJ+FK5FHkNMSLwY
VOFDdDkT6Iuv20k5jOqRa5Eql83H2H0fQPHeqbrTPFeOlU4AvFzrUrYwrMGNLmQr
NrYM9kyF/g/YY/AtqZsggGBF0BTnrJ+cJBD9wLUsOjOI0ERmwjCs/6y4RqbCnxDH
ZPEcxUcGi1ac6MMHosYzHnfqTx1b4LJ8G913Be6OALYgOvoEdmd7sgduXxVd4deb
T0la4He2sXySqwC4lGvvHb/ImXgbSp6sC3zgstOcMkGZM1e3hOAMlafszMEvHSFo
0R5jFy7L+TRKaJXrJ8rtVn+S89oWuzwslzPCPFM/0gulJJWO0hSWtrMYu8WuQGR0
NnkBRFcUiVm4KkMX8SRg3XnbC9Q7uuc+b620DxsQWVz70dCYxp1KRU+QXUEAxKwW
StRbz9oiEybrkAL9iaM14jihGN3QRr744zPdhE+0+nDEHhUGNPf7zqHmW56Y4dib
3dWVteAd4y4nAo3AH5d3qMkx4d01mJiiFuFid72iucScZyI7UAmlLO+I9Fn2VshX
3cgiLU6ZYBgOX+UkBD2G6vRU2VrXoKvpC2DTLeGM+lQMVtnWAI1OZQcWIylPNNMk
TSazIOCatAL5Ss0bib4zjg95OiENAIviZqO2IOKyke/hoZOAJo6YWZsHW28ijN6P
YHzQDgtP1SGetLTmbfMBbtrbIZB425xh5hhuHzhqEDjNP9n8Ho7ioHUMjtwp9986
QAO+H8Wm5eRXJDJl6itIXFB6RgePU3jatsZ2iEDOqwUNiMXEJpPNnJn6RJbvC2iA
PyO9kDsz5UGAjvUlTDdFyhzgkO374ucihsMlCkMmfSlb3j9bcX4Aqt3MtJI5XX5E
RAOJhBuz2hcFwMu9GlUO0NCN8SLhrTwVDFALEUwcGbPxaxxwAa4EAnAFJa1Qz8am
wYP+xvsWAfsfxHt01pS5qLgNZG/yOGL+zxvnZBMv2DXyqzDm51rEeFQ70mNXhGaz
P3nOCILaFrb+ag8kfgOS7HcQr/J1hdZ2NpJlqdCTyiiXpKeAbw4M+I8ndrk1O2kH
qL3hsz37Qhe5IoxZhPyIcAgGUxrRqxgX56MaB6G8C9e456kOuDHe2E9S41C85DeV
hWH2VmBhZ3HgPkEyau8xWLobajwrafiOKgmwG1vJ31oXYPyTbIBCaw7rbq0tzloW
NBgsDOAvd1C90XwIq7K83mJhLQegdKCQyhvlFzT99vy6JjtoZu85JKklYhM8ioZ0
XK5Ol8a+yzd12/QxipLC8qM7nPjPPsUaBDcoIlVJGzmg7tM2Mz+UdltKt7AlgujC
giw83EsLLaHR0dmQ9JG7mlMURn1mQVDGz8LXmDGo+38q3CFZmf8+dBCCvIktq3Q0
gKwl6c8mjcb2A+5eBpqZyTWrQ2F77p7uncmFMp8lzFr+08hs3yxK3VJg98oA6bYL
Ry4fBM9ozL6xkm36FWk+bMhpxon1jd+BelENwXQECZytsjQF0EWz2NtwyUTZoP0c
G1ihyk4P5BIWTFsA518TXzI2hXcMPRlbCnrrYKGjKUn61/kdXsTd7Gb6fqtKZekQ
VsPg4CugQBg4kJNUPi5rplrc6AFbjyRREf0tXFJbE2n7ZdRVnYFWwBaU/0zlbZJ1
CAHZciLS77j+lLWP/AAh/MP7Nk/sq3cej89rcIWdM0bGspnQZKEVNaKGNyeFwHkU
tTIusOPBqBvwHobLWvi6wA06JW9RS1MdRq3qW+HtrSI+u4ztsLiK8Do3gDz8Wcb0
UHpAXHoZTDcn+l0sIuafRW35JCtghsyTDmnBA8IyxxM/DunV+CCXPINAWOlc6Bk6
l6cgM6WBZOnBFGJY1Mqk7IRgz1fYpSSWQ0NHbyOJmfw78Gj0Yi10Z/dXw2wWQn8o
O3HDvC4/qBb9VcVjnCkJz200/aAYcyMaDzXDyuGh24M/IWprC8LAaekePM2dpR24
VNu3xOJi/TUwSMT9F3Uhm5Pve2lUhaQOzAyp34FCZHu7vloqHPbXx0NyIoSqk5KQ
zraIXsTI3nyVrv4Fa2Gd7tYVaKl//QOBj4pG2h8pghoJW+s49unygCBx+TD9CPlN
24gM95OLlPrXIjCKUUEArKapNHIzMG6iorlGT47N52Z/yTS6Jn7g6ZpfjnJ+m642
x3hZgK1cN/RrOvJaeUtEOQ==
`protect END_PROTECTED
