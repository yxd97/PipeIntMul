`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwTKZZEjRkphBI8tfgitYlcIoEFeZbjTP34HmokF5pcvf5+hlZirgbnQIEPzS2vM
vyaMWmEwX0nWyoWAPNbW+ywusMrj+9K4XOfvEIbcF/QgHKfn0qDQqT9BZ2Hqmcjh
3aUNEWT2jJh+HKTrSRtPkSTwlgW0ED1dvab64MbW3qtHj43wHSgg+C1pVFdnZiFJ
O31qyQUQ/68nC+Bv9H7Tg3G87H7Z68dwI40hCoXQ5P25VInRJ6k8b0giau1whAEJ
`protect END_PROTECTED
