`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1GUreBtcKSRr24qrJ+Qix8epqihL0s359L1kOEWL4IMkqnIhVqit65R4tKftCkJR
CXjPf+iPQ77LHzaPgRM4mt1l8aHGTtcnllbF0lZG8Oaf5PikDd2Kb1OroHeMyTa2
EeimrnBFKzv9peXvS4AdqWrGLEAwswUT3IUVRzytSYoxI3pgzlG3spqJMs3u5BDA
X9Lczh/5Xn4Oon4NJqksTZZ5QXwI6GJ0UDlP7mPEiX8XlbKC7Ty1TDgmz+l8mYj0
H4cKtn0Rpn2TE1+9eHMnN/TCA1AZED0dshs6SvqPd46zpTHxueUc3vpWAki6KNh3
iKjy2rTizjjmt9cEF1/UZpb20/+n1v/fi6BsvaCmwLg0heIN7n4Yn5iu3f5yc9zf
ZO/OJvKB9uKmvCi2DldMKfDpSmU81USuQ1wycP95F8umwt8bq8TZWhesGOln091k
iwgEWf7n8yNNTe88YVOdQ/mkEiUpm43wdzMxXcezRrYscOykoj0LIkPwAQO69pD5
IEJCwdTGlF0ysyVDMXk32D7IedEos3ktcfDb6N+5l+HjHeuYGKr+FNx3GrpGhxzX
k9z+NSumkpQ/D0lWnp+gR0fFxrhmkBx4m2n5AXjakPbDEhhgiQLJVr1O9IeW7SwS
8m/6h2/VDgQAaBdhQ8yHPkO+69f96xsr3aPS9E4sPF8GVyrQHO+4093l9VWmGDWD
PLmnSeyVo04FrSzPhwaxWXd8robxehtJw4YEPmSN7yP8611oW0wehlQvUy5x+7OB
FCXrM9aNimWVDAMzDayWjRwINf3YoHGQFiDtOUKYbx1uAi2wxqaKHtpO/3PXkAdH
AFTFwqszWmBc4ym3WWPdzYY/QGNfuEEaMtpX94/YrpugaW8w15xMJDqEv1MLSQOS
h4Mivs5OGIH8YksdRqJUr+L8sIqigpglt7jTn9oEYvlxoUEA/uQoR8GXfAxvgB9O
IUz4hjZjknfPo7HVN2WzFn9tq3s1oKT7YrHalyRJQP5LJksBrNS8EW6PjpDq5sMA
t+ba35vQYNKI8pvHERR/LrzZMgFmW/ZIjNybblrda2l9Wbc6D8GnXDAOlL4bSjWs
tzkZChNbKqjVYb8OMH3js2xLsWfd3LFjfP/JbVlIPOfOOfFe0PeeMa/4Xcw/crul
Uyi1I0+go0tVDzmPCyiUXgJcBbwX89JBvs1unsjQUDf4rhH2YAt7IvD2bAjydqcH
oBHObXZ236AGtgJezudXVaxewvReafM7J0NzP9YIQL0ULrvv7kGow6J9ZsT+g9su
l2BPuZ4lb3QJpYcuRWdVoTKa+/ez889PfOOKpg4S7TDjClrygn8poqq6AbpHp5D1
xunn2gVSqQ0K3xcHQYm95VcSn+UtnREdiXI6PSpBWbFQZQ5tYvVJHGKLiVc1NzY6
bqzSLzEqE4YgY61l0dzZiNWxNLWlKv0jcxw5Tx96UvpHR4RFDVtvL8MU9OGSziek
4iWtRReAx/sXzSnBOFEf3sZ984O4rPpUpjczFSOExmJ/6O2us+5STN4mwy9/yKl5
ca/zcdY8YjB+WPDL2s6Ps0lo1yeuidPVvd8DpvJtIzy6cS52b9zXVaexOts9cDOG
jb7pT5OhyQd+5ZbUgWPsVTX3hQh1I30evFLNwvZe+hLEvQk1jRq52Ow4PAja6KUs
yVYlYla91fMtdefrOC4Cz9yC+0SscHVV5U6GKIssezo2TNZzTcPebsXIXxgqL0P/
qRYY0GwoB/FegQD+uctxycG2gepiDVw7xuP4N8R3PXlHGvjDXHuAXpBpZbMSK+3f
nCH1VmxGWC4mkT7SBCt/Fp61BEqxycIwDM438A05W8XFgDMvEXmfXtaOymWp1lQS
ypiGRc+gSuXt4T0vbO64jk77JeYvhXsotOPKm502Qwt7ow7DT65jOCFumvUTYnLz
Oldi8UnK8oQwbzMABKW3NHXoRySyIBkgX+4GDGuS8Is0gMLdBHTHk+FWpglDeSZ2
hLNss3sFKoOIEZa+jl92YjVShz/XXVYUcEdPhk43fDcGSFm+oZUC+N1fimGlAtvG
43/uKlMhaUXCTIH9nlxv1ZDKnfhWI7KNUisT3OTIHBGLeO5BCuE04QOXK7S402qc
rNUiaoxGhsGNmeRu/Xeu7xnzkryY18AHfir0ZV7x1ZNM/FNWn2eelz++sXXlYGnW
KeQspAqtBhEF6OvxCJjUZMBCZPRJxakxvNxygWVHePdrVJfPGdDLgxNBicOpjwA5
2GjiepqHIQRib9rqYvYPq8+YfkwSMsazT+8RVupTkyV4gXbLMwVNRwp6vBkfl/W7
0WyS3FOqR82snp3wqBion5Om9Em+VxSaj3Co2kYFDsXOATRnOhaVnx14zOufZt4O
it7oL7CIteO9hXU6a2fRWTzoyp1A/P+wogVKFN+CxpoVEIqPpgxuY8IzRu3BS7sq
a1yk0L8NvTUWQ3y9pr8fnFGEXdgqKNDYxAirrBINQu3D5GF2FrLWdj1st2ar/Jpy
F3HjS2WC/QtsiCCNP55VLDhxhwpSnFsg/cF5m3kHBrAHZnYi3AbXTrYkYQNnVd84
TntcGle11vHnXNm7vI7JxU5WWTbHWzbBWXdIfjyA5yaZkejeVzOSirE//DcigOFG
1XPKuOtNp6NY4LcpwCfwLEdqwtlrOrTR/44kJi6HJ3txvnVRxYzI8JWDAEcOl5ld
6Lqqpil0exggGvNoBIZOaCWLSnHZ2tTDUvc2WlA0bvwhno4P3hmofcEJYyHyE9Iu
VwJ638XsPICQTKX9ejipPeTWBpwfhIosFAhoiPnKfkBlzI9WCtZA81+zhCFbj7by
RNgv9q36vBSpg+jsrEJ2thrvAxyb2A4Dvv3XZEhGXTJWcuRa97acE8Wdkg4Rd0ev
toeeJVkmlj9ZRloTLPPs83kXm3EDYTqSYdofW/b/osygg1UbozFFYjsS8nRs6+ft
SXbY/5MkFO1UaYbyxyKHTFvwKPfHJwZyguyrL17QMCUT5V2qzvP3foKEQEE5XDYp
5Q4gbbZ/ByNvOhONl8sK0oaded95IB0aHG1wJZfXklJW/n4yyA35QR/eARHOKzrk
6fezPhfOpHq2vsygL8vfA6ZYGe0tsB3EXvXF4UfwKYTtCxAaHncnqhpZ9HBHRsJZ
qm8PxeoU0aIiWkgW80ErklQY6Q07MLmaUa34JE/9AS2AZIlNcTFW99aRn4rTKP24
s8TX6YXse6QSAPxnCHFk9HFX1tfQcLuuiX8hjJuEzmMSGVQLsDA2ygZuXbtPRYj2
ROB0aflxBexzynGHWe87HSEBwKdhupRODC8ZFdNVjjQMFtxCp93EaIkhajeyGw+N
awa9qo7mq6PyWqjY4Ktntd9fALrGYz/nKG/uwTeBiu6OiFCmVH3YhWVcNQZYX4w9
SYdjJRTpX4qm1wWc1cxQbwQEkDbyfrsfpubt4wefMTUZQorgg9m8pYTUZt1/45pE
iJu/TUFFMQuZbg3xbfxBCv71vcjFp/naY+YMbv3KTmJSH8O423XvcfcQLA2mrP70
wPgeHtnZHCfdIGArhW+zWnthgvUcKHjieerfPGtWWlPXdKsZUr63x6IiNTAo6gGn
iMmaVv0cYaju6fcWyiK20/u0x7uGVZOJPAiJ/RlgsuKqSp25h3ogtKHWAYaw0Bli
lfdAkb/pq98JNPRB2jLEM9UMyMWYsCyP5V8NrD1i13/2wscetoFDcZBjBpZsVyFo
3S54eIVDYle4ZJWVRxJsOMitUfxKUT2EeBITkaygYrErxgpP/tkJd6U53XyavXNj
oQlGb3aTUP/EAUvAwAGr6wotTj0sX/9SyLlqPCXWDeAOdYRm7lqCpc4csQ4CUD85
KddL1t/h/IhzDYEmcWos/ceKpLtSfsdA8KPBrNKA6EmDGqySFQkFLWDg05fqzhgv
jPCqnvgjjjlimxW3ViATPLmoQeVDhcPxiaVwQterPN0V9OAe69NV1R34N0OKvkAY
6Nb0TdY04H2Jatxer7XUMmK5C6T0GkrgU0iIOUvDPYDpiy6QCXJzQofcqoV8Eiuz
r5xUynilVwK5tAp6mk1gsQCyPgoZaNGNHyjKR2m1FozlObxzFRGlo5fTZFufPieQ
G4tcXvWkWlzHsvETw2YAKv56uRZxJHQlqWjiIV0a7RAhzLo2QChJPoO4vtqIXppj
NUpfDfGWlukKBq/pwCnEUdZHWHRqGsu9vVwCvCY11THKTMGfQZQoWY16Nnwqq9I1
xNmK0rKz/rpcs3W/sUCWIBeVEnrjlbDNWnnzF+Cfegqudo1Ypn6gFThvINCYdr1o
5W2zZWUsI0rc6/BoiksNQDgeULoqReFiYNvWa5As2X6qNHPyLdvqJ29kvsSIiF/J
gy5dbSUuHGTN4zbGxDMFKJ0Q/vnLxtdZrnYw3r6MBtBFgRJ/bciz5tTx5dKqkTew
iZuVyEaWFiNjPR/028j/HtW8BGfOUgQ8I9mNWcfXcBKOmhjcOiLacFn+AbPR8cyO
xVr332gB+BD0eC/K/ZumS7D/cXQIul0Jkcbf0hgThtsjoiO1mxJ8S2ubg2Ex1rCN
bfNwjHiAfYgW7W+7r+ROXbRlyEjmEejWldB8fOZavqTzmMXkKmizINDgPrQAfzAE
BY8mJ93vPbO30wwFaSUBnG9bO/0Dd/ILD6D2tgUrazo5soGYRPKYpQdt5UB/2LAZ
6uG1B4mBwTITrhA0LBUrtc+UszW88NRJAXtx952acQ1RXsLb9pQiwPZdyw8s4YYK
dVwFu2RQM5WRzg8uPbOL2k5kzYUVB7hdIp3UiVRYJjhByW+Pnq9+8PlHoX/2MjM7
aBCDLHfXMNmh654C+or1GsHzvV91bze4QZDqKeNT2lbOQU+4FjwOf9vPMMBiy+kC
yMrGNq9BI97UCl/O2eTsE8oXtBvtMvHUZrUndThBt30XyD8KXVa2W+CUstvE3zNV
YAnyw+YaE3IfwdrTMF3fXcKNw0KHCnu48GJKaKRY1r1yNSQBoX8MhGFu76qQnEax
NbTU6+b47wuCguIfIoVjO17XvBEPiE6aGNdoZDM3QYqZcG1ps1z58NOSgwvSNP+j
c+zqzTDlRg8PyO0+USH8Mw/ByQQOMvPr9IhuyVg9GI/frJDLpR8oqOcTDrkTlKX9
XX4VSG6CV83GPBQ4ntUoN2d8cgeFbbE0Q1yv3eLgCSLR0JxJbXpsheOIQpXHUtma
HIHLEZSlNafq/nzWic6jq5hNEdtHVAyPSgKUqqt2VxeqOXqXLfSa7SUEs+bAuiHQ
N6uRjFVFt4F03mLLV9fZUhXqvSIPu4sih0KAArvOHCzC0YH86rzCQe2gDq6vBbGr
WkKEWs3VCGeb0hJZO3+4A2x+F/q3i2H9hVvChA4fQNyPXIdWshu/pBKXMamllMr3
ZiBAIQnk4vMHfgSiUUQZgfMt1vrOIsId1jt3IrqJ3vW/O6fWRvIqx6fQDspCuStd
CSSZwiylb8FI+gAwxlN/puP8iQHeuUUS4itMjHBTseZ0IHBwpw72qKqsmAPttnR4
Yn0zupgdFIu5dZbpJbJiINgc+OmXrlYbXxrwK6rdfTbEa4efbZdzLpkM1HLPUQdJ
D9QBW021Y+wUVsB8bw9olvMxUgU+oA245MDzfCiAkQ7gOo6Toqykxq1o9tnF9rhg
8AUBTa1a/ZfEKFbNwcbYjZXk7G2bTpD1D8V/DW4EJ6Kj/hj6vj8yKZQvx1GA8q7t
pfV5/+rp9A6uy9GT56BKz8Iv8m8TiRICGEEkP9tGgnWUXv3UEVJxVgnuLk2QBOiS
Mp6ixF9d86okSMqcCRSlASFIp2lSAeSH0XdA5uaIWkd2o0NTxLnsdXj6Y/ZAMqwP
AAQLtQ18NeSfYMkx07hmPdEs33y0Ut+3zGcKOg72Ksbd8aLh4orH24bU2UXMsngD
+ra7jzmBjri1tYqbP/3IdgXp3qy3DEm/Aw02xMnXggwa5nDH70uA5coKewyn/fWw
EMhJpxKabDE/iJgRygwHiCBhiX+lpi2r4OQ53VP5Zk7A7Zwv/rxosUv8YgrPQ8Sj
yGTHhjMRyO+vOc7H3JLMjVG0Cunj/Fo9yQ38XptozDx6qEmRyFBTzPVVnFJkH8JU
UFWBILz5/f9sLJbAgNW+5L6sbtoONmx6aGkgogvasuy8U1TEIKsLFe+ciLWLzE1n
ol7h5tahJ/bQxlcovLy7sE5WI0xY5wy+yDxNswT/t95W+cdiw1NJqWbXLtAwRWUi
LxqUDzsan1Z3PGZ6LmeIjHcu7Bcttt2fCmHoZYo56hUC6FIsLTJSiHkf6vC9uDzd
VrwH/fyd3zDMYuWxLShZviQgrOHMLsLPTKMQzMOozSj6RKY335/ETmdmMyTI1l+X
N5N45M0QifmJnnPKsi2dnMkAgCHsMHa5VZVKwXDGrJOO0EP5PO1bg7808utpr6QC
quWmFOJuO7SWgE5lJxO3zuMcxkFlCA8qi6Ux1U6A7QEoLwWurD6FuUgPEk44jKdn
5lt88K0dynN23NzTcjaY2uR81W/QSqawtT9JWePCBg2B6wKRpu5+jiFp//PeCRMZ
9TGqoXZG9ekbaaj7L4/LY6T4bFxqqYk36TsUj1mAa4T2+qRtckcpwkrjBbvB+f2u
ZTiBBBoTtGkvMxnUVrklHskLVhQ6rkxzn7Dwf1ygOCP7a+2JxXRSgyiRnkjNYyGD
BZ3VUS+FvbaNtgUnggeIkBbnNFngDOTWK4LT6pjA4MdNrsDpyIKecY19qRZWLM3k
cPLwIebPXv6MNfLT1LrBCMP+b9JnRdsuUmrh/EATB7XBCGhu2WyQ0xFD+liKi9mo
fDc2YIkvaEfjDwAEatVbP0u0oN4/TA7qJkYXVyE250nkF+1aHLqbpgNBrXQhr6Vt
hbGYSB5E6nCfDaZWEeAYNhWUI4FYxmTfiMBAv7O5H7ZFPg/65cQOYN7UcSwnilbO
wmIqH3l0AJeSgxn/yEu8UIW1ntBxCGDoLLBfMhYpzV7cVLlv9zKUvhxQ5tENHw1h
SXbl3g8oRFtuCTfBDeUN7DX9fanGfxScSxnWGZn3fEF84YQ1t4IAgIhDf/TVLnSF
8o9orP/YCzpzVCGpYN/Ha0tSXIyFq5vRW/WrEKPqvbcDy/+RetzIdocG5gOh68NT
wqlK+eXjgMsED7p7kWX6JYbTKBLmuWRbe0rhUvHB/hdvjhYvjAsLreNNbNbQjX56
Hsnl6iv/rUtKlWXkyQ0Uui7CTESOM72eG3IwbSNFpPgiweKcLx/iHOEnb71piHnI
8g+aGO/leQ4MyVSm3Rjusoc9LKAPB5xDH02dDjc5fpJ5Qodh5oWhutXy5luZ9uhf
AFDUNABYH6LE3PWC5lqev02jO6z4cKH5kL3JVR0usi/9P38qUhHIaY5saaz4OlAx
rgMnIqqJZYvMFNo3TqHfTpVcrfrjD4Xx72H31v6bYmnnAMP2+J0hRjNAxTEMQZkJ
MXKoJ6zPL5oY8TaUoVR8hKkNVnMgucAUtedn3DAS7TtZChZM5YilS+v1YB6vVaD4
+Xcj5Y+jSBbQfXVeQV1CFpIqP/HdRY07gYBQ+v/NDdPnPr4n/vQn9t66EocIgxgI
d4NRqYHsAM35qH9wbi+/s/q8n+gY5rwQUFWOVPYXX05WfDnGAUvXXZkPaFsDMFAk
98E9kP+toizDxExGF3ZzpB8wi3nbuVUzwr2lYX7UfuDDEsXqPTMwy9yHRtmRzMw4
TUdP0JOMG6b73YYhfm4HUiv1SDuZRCNjtddcnhBWLL7BET93VU7Mf4ilCl4tiXpE
SjktyxthkTH/3l2Yk6vNnMjhThzJz6/KxlDaFs3I08xIKnTGMsEa6aq/kya6b7A3
KEO33lpl6tJ/hOkvyOC/ulU+9bTn7qWNAWZWYfbZSlzRTfX/YtGayrwutN1sFLOH
p+wREuo9+1WW/WVxBo5Xq/sWUfj2NNYEqvrhIXDzdnMsZ5+RxAEDHGSyco1yKajL
9hcOBADsopU5odS/+kXigiRXk28QAUR0TedCa3uYrILgdgwEKYZ/+l/AcE2FjhkD
4qZvBfXdnbZPh4QhIMRNbPHKjl5kBxoAxUqf4OtVn0Ga6+VLgrHuBOtQBX68kRAx
HCuKrALRhTmKF/7BaODuBuJndSnYKc3IGdzJdg7LBrwuKbnxGzeRfCngIfHFTIHW
a3r4eCVMKXpA8qB6QOMnkE7CziZuMqakHQDTcxa4rGkf6EQ/q5ldmYWI1KR+qOka
HSvk69GGNH8Liw+tQyq/0L3FGP6PAOYMq/5XdDH9cKAX7qfZ1qrSTHDw80d+5TF/
UScjwtqGJHtVHg/wqXF9L6SPPevEIUoNDnJangkTdMmNdZ57eUh8r2nVBVjVCuS5
yD8+oeMMxkkO1UKTiayiuZdMCCfLjtvPqPRQrc+wR1R8Eg6y6/DDnPMx49FlYdQf
1w0VFtYvJ2WTlSqx0P62g4RU4mBLh8Yl5oxNtRig++guMI2zczLXKAEG0bOm95sa
RaVqXIVUKGAqFhU0xqxFnS4T2/PVg0HdVkQHg4i/+FI8gdfI7oXcjACt/xPkZoTJ
02Hmw+5qf9FrNcg+cpxJVEDQIGVlP3qwnAVgsmJgKcuZku/DD0KassAFmuDCkxyH
bMo/JwvZsp27Fol+5+D6C3cUwFYsiExyE+OdwZYUdEqr7ZjNda5pt9X0IdP6pvqq
5oUn34jb1Z3ePHO6gFuGjff2vkn1qClj0qlUKhLOfjEsQW26XZxds0RvI4sec1nf
7MYZ1xfsEkdpg8yk+Mr6AOgZamoDAxc4qwDLVfae1pdxMXTncwNEVblf2CGl6g63
SWe57Udkm5NvVATg8p42ZvGHFRy66MAFG/D2SyEDq+p+dsKkynZh0sRMbTNmUd7G
tq00PIxeBwajJ5/bU3OnUorxq8s7erixAhNMpBj8kSxPUGJ1L6I54xrb+aIMCoY4
haOq8tjBhWqwoizs/s7W0J0DWo4hN8gtxPNqEs1FwL0Mjwb02veKTSQtbvSLsWPp
t0hyWJIU5RaYRywh18Iu2agQBjJMTXb+Z0NVc0iWps64bFY69Dy9JocB29JmCTu5
A1sf+K/WH3Q0MZI1kHXEKptffYt02Ji6aCUsHylGXQPjW8wBvfD2a8F3Dc4bTsfL
tAOwuDE5+HcaXZhb1CrfWtfepr22i1s8MrsGTIDRTGeGl8mcyO76glvm8R42gdl6
ZTBfkZqPwKP5yWnVKnUOZ0bdXkpzkULCirEQB3P9s2e0VDkGqUWo1TKY3AZWpmLT
7dYx83KVgfUExL+XaQIptt4BWJjObut1CZCbuBzm+SJqnWcWtMIjGTzHbXFI6mqk
Et4AOuPvfYhUjUxa/o5ZvhuW7eumCAC2PmefrN8MOBTLWotUk6O0x8ZfPUqrqypS
kyzXjUurIxkpK1LNFHzOAaNOJxCEVt17sj36d3zvlz8mrN/J38aRVcOCGdB+sIEs
b5cd97OB7mIf/QtPW8UXxBgdFrIG/SclkkrNBoXbcFRpnc291jUsTFI0aFNG3rfU
VfLhmMNnFR8BjJuapfV2+mm17rdSIcHJu/u7zr6jUceF9w1xXswGu4Wjz6Z1k2E5
l3LGYLIzqHgF34w8AgHtMG/Kfuspc5q93xr0z+zFPxn8vWug472EImapvGkX/e2z
OTnXTLcQ4taoe/K5nmFNaDt2CCBKK/Cb6lzOFpTfEYz12ft7T3CIhwCmcJ3V+G2D
f/kMLie2b8El4yjOAMKgZ5UtExpLyl4UoJV5LQLtnAfFk7+65o1MAD6P5Zcxcvyn
PnTNR+sA0r4Ljp2gh0Mdx+/I3WyZyzULK/nneAxvw0/6l+F7O1Qs5A3NXbMq98r8
PZ+Oh8LOv+et8+Eg7xxNZVRAC0FOZ4353W1Jc250QoaYPzAfIB5iQwoYjNhEQx9a
rAlai2v8ry+V5FuPdP/v86WpCjez8o9z4XO5gW9oiEk+6jwAK4UTK+YODscnIVY5
u9egO6nLAT6VdM+0C14ds8D+SJ8lf6XoZSFvSMPm9x7WeAKm074YMUUVn7zD5YG9
VVXwrPGNZP7JkbtFIZojhUDVL59jNlz45y5y5Q17ZMrCaDMKMPPtt3d7CoX3V+4K
reSyjpjgN/IhBTAQ8JIdQcb++0dI+MdiA0YOso2Kie+6YnqpP6uzBv5+dVhUb1Os
Hkl23rqLMKYqR2+l4ZvuvXXgkxONELuiF5Kzi1zQxqhafOO7Wx57IZkt7XRoVxxS
JmfNVfd2Z1iJDkjlrMp5+bn9H7DpttRmPa53/R4ccq18Y6LdW5pzV94H1lc1U5TI
DfsfWspGEksyav6NiiVLUWT8uZCr0/kYE83px/nQhnVwDYEbXvLzOnRDGkOCElAz
P26pONkkplb5/mMlbmauZ23PnSdcfWDtXk9aG4wK/qi0tgblGml5r0szo11Ov0XN
77wQjcSWddiLYHvJb9xgqhxw57G43mJ0vWrgT6yOteR0lDy/ekfy96HSvUqk/dMt
1/2va5me0uLoskzCQ+cKvdt6MaHIoBOknQOz9Bq0UCCBw8FFK2mijwCgInnoOlom
q2dp9dKXG5wSN2bliDU/ds8J3OuXPaxToILej4LjH6RkN5c5WBbG9tOSWdbJwwTx
yTYA6KzkeMpwwaS9A6NipyDCILMsVb6Zs2yZ6HRCBQpUOTXsDjLTiN7XmJ/2tQFI
7S7XFU9zvtpnugr1sOFq+1757J/4Fnn6hGdRmSf4EHThJKYMTmbHE5X2AZ1wUWwt
/hghXFGTnx7wzKUo8GSdG7aLAmmHbvGg1QgSPXgRWsqo/E/b1tGtiawhGd4Dwpw0
hTrwg1kAFp95EsNsPS5gp6yYN/z2jZPzLh2CbI3KEQC509xT9pJzS7xirV5c+zwi
hgvg3a0hU1YYiVdwn5XTexQLzDLsNupMdfOA9ZCrVRhSxcHDZ7KMgWFfnrqLHH7Y
5B29yAinfmdk12ZH7nyntYuh1vvHFAIXNDVfKj9lMb2/tII/M1n9hpPw1C7zy+ZI
LTIUHNLVX8+UpUS322Igdo+mZcSshALDSM+pbv1rx0NntAluR9dnWb5nWwPoiDAw
t/DxawP33xwae51mhY5BM/Rm9GPkuLmrcsWYN9VtRDDkBQuiVcnD2Tqddj6m8efj
sD7ms3/VVTwc5UVXOCNBzvEM5t3xbQPhFqEQ8PvvNjiQjUVXfZlRf+lGOeUidKR/
UwAt7z+HqlKdtx8zCvUKqPbzWFG3HKtgH8PW/PpLU39vSfnwrP9gU6fFWjPJR01D
G13JDgTZEk2ZQeIBFmTGLrM3yGZoPkzV3UttalzFn9r0Djbig8phvuzu2yd9KDxR
CkDOwAOQrqI6GLgBd/2cjmovZiIryRhHYcxOcg4bPBXhMuNa6LIBhvynjTsQkals
Q8fK7cOoHnrrYh6fyXLTnnUAQSZODbK7EPcBD7eqB+tfcYn67O6UBlOQPOaU/tu1
S66SD1uMzGqK0n+RqzLdALjM7sUwiglCMuNnfZHhtGFKxWgvzblLspEg6N/9QtHw
TenW+lK85fIoUROL9nHoW49uUXcC6In/oU1KZ8FOLsVhkiUoTt6PllwXNQb9u2Q6
ObEpSi1rQ8PBpQPZRbmJwFAvcbpKrgMPVT6CiZND2jYBFUgEK/1MHUWorYgpmIx8
AGNlGntGaNWSgPnhR/E7+nwgkxGFxQfC0VnxvlrvJyxRE/JyxSoA5Bnds2u6RF08
+7eFCqyDvHdYWcqVIqvhtEMuBL+ce1NkGXGqKZxd9ZFC4M/dOGgTOuDkcM76W7tS
NwBrJULNfMXixRPriyrva2UYZJ2f0zoNoJYt0+qVVJetnFpM7QrtBQ6ckGcDeMUr
KqqbzTapySNQQiTC0Uei2MlY0GznCrSME9bZ9FxxOKXlbmjbf1vhdePpEvlaQpjC
/itYr2ARjrYKpz34BCjLkhWDOGmw/sRxk+T+iGvjAsf2kwIlyBeRJYZFDK8Kvm3P
SvXxwICg1QZHUQ2nhHJUOWEvqKy2PgcaafCJkCdjP63Y5KfXo1OwlRwPWUpIwi8r
W28NAxDVfQTCM+Xqo/UpvZMu5wePYNJVCYu36mIJHAIxDRrzJiZshimN5hqz7e3h
XAEUMYsW+DGxnUBrr2eY4P0BxfBWhxcX010FU+8RE16+WZORL8RqO0TrwLtA49hN
ZDBGczVJSG87nbkLQsaRMA+FkzXBeRfZmpmoieDlfaVMo5J83jBTtv8B5OXa5wFT
dyMgQBjmmePwsEg3vpRIKoKNjB0By+VtUuz51e13tTPB1ZW1IB7kS158NutTGpuT
et4moLV1RtW9LREXcaFV43nO9Fl67W3uSpljOZvRCR9b3/Kw9zUYXNBYHs5lb+gO
ODyk21vVjpJkqSYyIeyKrDotaPa5M+JHrZJU6x8wEaNJTXewwVYckARXybYuRhM9
ZlFk3JZTLeFg9/qWT9Yc/MK2dX9nO/qYCBmWkkLJYX0SXtdaWgP4cKynA+Z33haV
nPABGZZ2Cj5V78Sj8u4waXHujKnHDQkPsB2pqLd23WwDRffvNKjWfdnZiuPpFU0T
X0cH96XqtgKk2mHC+3VNS5t40vwxkVQ+EPMPV380+Xaddrwym/cREGgipgqpDkHS
vUebB9kZN3ZvfPEUmTUl3rvMGfzPHIi8OAcCb7ED0vaAPcihUdwVwE6nrWPaLSez
PtsjBYMNMOy23p6tZgSVtR2rO6G7WnKIWMwjWTKvekC0lNGtbfRF04+e+JHd4u/9
ZkxcSbILrOigdfx0LCGks0cBwvgWbiAGdnPN2tJSVsUon94rEqJ9h9KUKx4XXwzK
XoKSWxZR0AWGonAd8scSn8d9Hca2ZrEOPXjWkyBsUt+gY0NiJp5TAMuXtEdZKALs
fsfxTq+l0w+yLQZRjFVEQluuA7PVEl+mj2My3RBJ/ao07XdgdS0oVoqo4TKxidcu
TaN02C2ORooY9mJd3y2Xpn4RlskSrOwrxoDxBDBqlUVwwzyoymgsYyaP7xAzMP43
kYdb2/08PVlPTqr9aFn8ilU+L7qm3n3NqbuqQD4Gi183ZRvkffmuJej8Jrb1+YYg
bPtP8Mi875qFeVBP0Erzlrzj6+PbzOnyg5x+27iWB10zbV3/fGCakVec5UWZJacg
oOlisZaQq3jCYSXrHIwPDzb7ZwBQJo03dOStHOimkGg4fG/X3GQybh36T7ELciY1
PX/3l2uuSnUjRRIIv2d0K3quj23vfoyYQnfR6IIwJPHSYbTe0QUEVYhQp4K/W5F5
O0xqw14ton2ZsN0h3sz4NuDfoRM6ZiPWbwOU47rSEF3rzk9RcbndANFwKZnUroaY
2KoCpdCaTxJaIgv49jzrdFaZjqo1g1iIEdMCu/3/Laosn8crSkaPELaOmLCIOsuj
iCVlRPxxwtInS+wXJIeR2Rugb5xVgb6gA5CoRAax2KwFcF/BtnyHB+ZhKxIg622i
Ro2xmBtyNuclOp7fERWd54ZOOIj8QJijUjmWRS201GLjq2nBN1/gzIqn+aiQWRts
d7duzm4ODXguSyk2QkXFzmlifp4a6VHAKREZ2Rch2+mgrNHfVi7U84sGD+cz3KeU
CH302bNzoGPQ/dkmzTmC6vRbk7iIy6gA00sBWhKPFK4+cW8XuBf0IE3FdiQoT9co
6i2XOZp3oRe/ly2aPpZbl0IHyoF21I+/FoXt6EBaFrZZFPmkZhJHK7algRWN4FGn
NOOadKDtSy8FUU1O00HwDx2Q3X4dGDls+BlXKiEZV3UhTsTaH8c76lL1OCeI/yZO
2W3jw7KDlwuPuM6JflyZWpAkRxSyqJR1t4ZCVWf3CyfOM6PfFKj9hI3ZFGCy+ula
YyTpPGqdoF8dBjQu2nBebCWtbHoM0iJOyFt1Lv3yZVLEG9HSF+yyD2boEAZmje5L
VPNm+qBvs4t4vlyvOXedCZBdT/168+JWRniojNCbqvFgYogtCxkcr2wWH4+IegWd
rjL2xix9KxBe7htePIYiJs8guF92TxX5hG4mtF3zn98m2YpvgNdnJDMZh1hRmG0t
yG8YIrtR+s47oHyu6rYARupIhFJYyngXvfanvf+4GPmpZlNZVmY71XZ/gg1qP0lT
NT/5+DRtuv556apZUXBAiBoSHBJTLStOvOd4hlYhIXy56zM1lB4vDqw/4VRkOOwm
OzmY1/JSgor2upKAq96gT3wqCU3iTMW1g5y1GeTFGM2eK53BpIa/QpS6USZrafUS
koTSgwwXYmjo/r5rNZGBUPlOAyNPNcTrt1CKI1zTUPos7tdrzsnoU8lRnPVYBXCs
na6nTCsFPFY5Z2JUhglCWVDSjM0ToPTymeTgHAl4no6HJqTiWhSyF4X/bZAN+IHJ
0VSbTUukBpceYXHKIMWFbtXNjbNZEf9gVR39VdmSIetgSkwV1MBBicpEwy3dgAFH
cMWNpaOIaiHap2Tp7mjQjVUhyHjDxospnBU+2ttz9Jn6I1bMJw1Bx0ntmgLpapU9
EQOh/+dY2NDKJL2CeQ0ptHUFR9xJh6movLKzDzIpZ3gYnZq+HUbyUuAmQJ0AkO70
ZA+K8rRyZeHk0SttjEq8RP8KRzxUmFBS8sPuekymo4OudTp0wi7FLWNMiYQf8zhn
fNjJpKOWiPHv7wPP/nvnuwrOGlRR39MpbW6N16rATgjetXnkPfTyvo74gkD5u2iT
QqgMA4LRVJP53lZZblqfKmh+JnBLWDuxZ70UBUwHgV7zGjLS5I+/nVo5tXVBerMx
TBFF8Q4KJrOjJma0uEz8ebbC/GXSASohQbpDZX+bpfWd16JX6q/H5f/JbrJv9TmE
42rYChyn84xwptyxhExH1T3FOd4b/HFG/FCDRG4haEcJKSNbSml2BtSPwdzEMZJ8
D2/Wh3k28r+XjJNLRWZydJp9UQhmq2yWr5Y9s7Cl1t7i/qjlrOpqK6mSvLATBbjH
KsHz7Hm/hecSZjAfQGJPP09bIY8m4aA/DXqul8UEEC+raxku+NmrpQO+7ENuo0a/
k1nwg1lB59EGLAt4caTbh3BBO1zPk5euVdiHwQvEgb0k9UUemAhEyWLEBq3/VkMe
Dg3KjxLN3WQXMG0oxFtpqhnTXzbX/WS/BM/ix3FujjfFpDhCsNpl9UG+/gIwl72u
nbdUmmSt9MFUpF/dQghY5VKArHJ0gIaSq/jY5h98Z0g903EUmYNq8Tg5TUYLmX/U
XwbBIiULedcwx5Mk4o3J9WqpNE+McE1zcm6txgWUeRhpxfHDC1OBTng/c2SeMh1a
sElHzvPh+7fj9QIvKBoTyA6mfqGRD/Xpw+sq/c+30DHe/IDmkerfTpks6J4iPM3B
foLV7UkeFu9PA0aRiwJKjbomXvlHG/nNyQ9imbdGroJnx00LWIwJFbRDl4/Lpqm/
5Jjd7cG4V2URY9TEDXozHYkrRN8A7VQ/FAuPwcxUgur58SQ6X0rxnPQYg2YW6G4U
iV43iyXL7oPfjFGvOkkGikE5pCYYl23+lLSU3xzZy4GVXqc1qWOFNOesDrP778b8
SN2Dn3pc0Upx0sA7Xwk4ei/C55lopBmqswEuOwTO3OaYAhuJFag2OItMRuMn9NoN
ge4cyMIoNhkM/qZPP4dj0qtith4aHHgfoBqPpIkLfn79Js/luMjPu6S39+Mi2WuK
NXzg8z1RuLkFu+nFP8HgaJvG4iEXb/C9T+NR1/HjAQyb/ZLTe4s2jF2JWKL6djtN
Tkjs+FWaChq+nCyAObYy95K+Yco+y6HVzQICaYp2qZlDI1QbjNTHetGu+inBPeHz
zAbVKN2p2zcb/LGaLo4U3xSxniAFVdzT9nrxAUdcwZdnHgaGlttbFR/QSIoHTX37
mJxG0yCuxPtNWHRzR0JXjiPVlTH78uGTc/g3CEM9dcAL403ejTbdKocimELywQ2Y
b4cAlvpewT9q62hhxiavp099+s4BxC4/nZP9mWAC/31VbOCPIsfJdg+ukfQutBhx
yz623KOhOuuElhL3rAQdK+DIBm5uarBdUhOo4gwthqJ4SkFV9QIvqPmCA/z7gfbZ
no7mjZgL3O79NwJOxGwbfszhjxkYUiQBI9m6BT1D+zWkdtCxV9HnwoQXcU52HTog
cMi659iqo6BOPhdb0FGIeYK0LEA2e5CusmSHF/1+DJvs/DZNiH8BtyGmBFpJRiZ3
Y+8WeTVJKahSmkTnUnhRhsmLegYH294n6eqamLaW3ma4TMj9xOiHPSrV7K/4gOlx
sm6o6+6mFmgdkv1JajjJkgDHJpZWq0aYDbdHcawqSt3uxXGTzsa8RicTplq5FjCb
vL6S7LojnZWrAJPaOvU3T27h/ZBNvHm3tvjUHMzaKhlHLwtq6Kg7nIY0kpF2IlXG
WZVkdjmXUkSP0+vHQq7qIMyiLnz113EV0jehi1T+uu1IWipA+2x/Q3dTHPG4qeoL
Qe7dUxs5TiQCvbmh2BVkfBDQ7zfW31V6RIKDKaAmZVDdGChnmMtNAcudpcdaZENK
+kIup8XwY0074PwKiL7Z1Klbj0UFuXWtiNsyiSboZNhrPIs0tbSZfMTMsa6Vlema
5FuR20aT86YRaT6kbHbfch+ZwvmGuYnJU+D0Ik8QEl45SiO+iZSFvYASYR8QQnVy
wN1rmvirDKLaMx/Zj5ZCZldK0vBZAM3cddQMmlV9YJizIZZsWz44R5rpkSCbYFxC
eSCLVcT+fdciOVdb+04QDteARFWFmsyNFNzjSCGpdV4G7Jqo3sCYeQAMdfUeov59
1wADV0KTTPa12+HnyhO+Sn9iTy97We5sy0RT75KB5edBVD/EfKQfB7RocCoD27UM
VOZndPzwnQ8hhy1FOK5uW55Aw7Z1E5aB+kX0lNgfoFNOWRfBy1uRkVukERCfsJ/X
KwlZDNun7OHfPugDu40siwmKy5/bgOoVxFl4rc26ySvPZg7FOHekVQfVsz/mzwUP
vG2YeFEMCoJ7OpyWF+phq288cY7/fLKJhUYnGxVjZKbCXoNwRaENekd/Y5i7EuTG
UHYiE+vCXDu/DAYPgIFuRuL1zw+FA9S3pPKwHMAmXHj/lLknZVL96O6Ee2dVf3QO
uAIR4ms5BwJhsZnWm0q4MBvnRJUHVFhc6S5X4ghxLU0dA9V6wwzP0HofhJmAh0JT
zXRP1R30RfYSo9VVpH0bqaWURTznI3knA9ZRje0/HHFG8TjYuEB+XoZ4r89c/OmH
lHwEurARaTFCypTaEd4HKpO8z8Ffi/ST4YKRmjhMcbvlDVlJ7nqXQA07fp78e0zJ
kAjucBIT3pqTxeDCeLR+x4EMkpcJqWpn0lsq4hliloM37H6bQbUxWl8rdfjBFFUb
1O0Emg7vXXJBMi8VIL/b/0Rr4CkElmpbDCgH5hnlNdanJtGmCU6eAnRPT7xRW0Am
xjv9ld32pBy0pwC1g2XRRo3G5WDbhi44pWlGlC2qPa9h/b+KxJuQoXwaPZZ5vytH
UYxlaxjEyn4LLTiBYe+vVvWQ2gdfKAo3jMnBd7wnPJWl6ow3zKFY5bC50iYZ48kz
yw8a5sJlwJi2433b/dvJea5t6wmxPet5jDyow8fTiyUrPAHX0evQbDHTUESPvkoO
mcYzCpxSVJWyHz41fZPmdChOnHdd1YZTmUIHbAAglycMHqJuYDIt3L7riI2yTqHn
g2HTTHp7/mpXawgZ355HS22qCU5MF+qP4QviL5YMyfQ8eHlTTIrRip+9DTRYZzqx
jTnxxOK6TqBRQudvEad3djll6xkWtTVig66fdZdxLa3hsLy3zmHqwemsWnrl4gWc
GiJVrOJ3Sg+iV7oZg0KFP8uLJs6cjM8b8VsCdWwQxfZIiOn7CSQGxAkU7W9UG9+2
iy49pjpLcy1uvye3tQ7BOZhiu2vJMm9IUHPklDwNEIWSqToWPWnZDo0SWL+gWsWQ
Cix89VxnuQJcDRzhZOhuks7+Oje5RRudID21hzg7KFrUx/308PRZEqOvoar9vTYb
4nRqOthvASgIClVirtX1OnVAV5JoECMIK3dLd4kWT3PMBCX5yd8uua2v8/XbuW3G
xe2tY9bJvyFPbHpY8vQ5xqn6k4w7+xIa4rHCGuUaz9YImHhtFzeswhbInnl7WC/2
evQeWIkWe0vZIUUCWWB13DNB08kAXmO/NuNvkO43Y4ObtxH9LO6mwtReJTRslkX+
7BuLYxfuvoSzIehCOqhmWBMoHlEgN3ouqEwTNmFjAi9Y7SNmvU1RAutycW+coTlz
aZgJ0EYqQAiBFN9pRMGJxNFXJ2O6rLHKL0c/enc+26BLuqfSJ3oy7rijf6RmJxIV
QeQ9TLo3i84BGyIttb13kjvxzlfBlcnJpFHEg8mCdtH/eU/MkScwzPkGPX6JQ1c1
d/NJdWPUEKAp5XxesaqLrqAtVKt3uogufy9OqKuFmxUHJtkI+j8vea/pDnyxkPtH
oULGaGz4Bd5fnAvhScFdE6DzWKrNt+w3zLh2Ru4nFVs=
`protect END_PROTECTED
