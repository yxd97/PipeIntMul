`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6r7gFtceAIauXbuRZokUaPZwj8GefheEoj7RQDLQnpMFhghu8gTAOSSYSZDpXSs
0VIgd04XomE5NMUDZyDTd/ujNuuhwRMn+BxQf7uiUL9vzR6NV21RHbk2CYBqh/SY
yF4WmuOGN3dNXqM3JRdvHc0oSPSsnPdsJZJuIhgcA/k7flqMBto5A0L0LoMF8+Js
3znZVT0OOZsT0xgDdeBkna2V3QbKSPjr7+9OiR3NXj/wtgQQKvRKx4svqn++AGaD
o9IsoKkHvwiFCO9b5ujFfaOHSfGjZRav7vcadfrtT0A0pNK3clCiOMTWGSB26ANa
z3/veA8UgUK4y5mHvtjaybJlVpZ3NwPqbsYJNuKHHal7H+CjwqTxK3SyimVoQII2
imk6sZzQGFnqw6hCdd+9zpxQPgIk8DYSY8Jq7SUx5JveCb869Zq7QRRIpKG1T/Ki
HZxto6lnLnD19iR91iEyZivssSgv2qG+231P6p5Dzzi2SS5X5YP3oDOWmnPGjpVx
m3MvtaxFFngAvxCI9ywCRysJ6Zi+ypOiekH6HLo0mfM=
`protect END_PROTECTED
