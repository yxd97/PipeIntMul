`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBKgOOfa7o+0+lin7ME+uyeCRz4ygUcz2RVze9aVjZp73XRpU0URfwk3a3nDV+uI
mX/iuTcykDcDm8HWIjOiB423C2twvSzBreiWRRP2KPbYLGUt28/dLw1siqU4EJDt
88FdcHSAs8OoYqXpMv7LHBB3Y9nSMyMmt4AXSTuF8hyXY41zfJZO2hCF3i8uJ+rF
HuVuq97rsdMYCzFIECk/FrKSxgzb3mgzfVxBft5T8nzpXmk1YUvDwxwSZswaxIyp
EXOHnAgrVIl0XZ26U+91LHjqhbfAo8mHjhRb4iQ8OP/9MK4dfuAVFHgNcHdrcGSP
cFt1bX+RtP3DU++P9HICwzMuvdbZmTJQYH3ulweEeO1F5Xclb6jX+Ns2pkvq+6GE
/qUnWxptKHPmaTjLiRs7n8xHiY9gLiHKTIwwGQ08fXHPx8OxuqiqTi+fMXy5CaFB
xkBsQGriOMqHhmBwnlsca0ni5X3zjVYrFuFETEvX7sUSH9blIS66xa3lmfI41ZRK
+WzQu4hPVs1yXNVFaF5/lOSZ727IEyFR04nvqNjXaTFucuF/pJAY2NP3nHsg4FMD
35R8cotfzK5lO8I9vxj4ODHMMDbJsBFSTOeTCgKK1+mm1rhG1JToGn238ju1gbSJ
ftsGH5wB2JWHsCi9AOv3a/VqIwYC6090nh3dNQuQHBSbGCunm+/bB7tTCxiJ4FVj
hS1t7mbCgGgJsYIVJX25OwIk4flGcn4lvqVKo8Q5kYhLbkwO3FQwYB1tAVBDy7AM
VS6SH4Jc2E3ShNfw/sw9DulwTi06qQoz2iG4zPRBjs3bFk6ETIKtFdwNRLNzBj6I
DOTb76ypS+9oAXqzFtbtpJItdq5PwHbtebsCtJDCfaFjYrh4NkJ1rpTZaAY1DZq3
oCObl70sub+OOtPB2fZSntNlGtcgA2tbjL8tngOcOaz/o2xKetDHuURHFXGqmMIP
veiaQhqHMdl8LVk0zqnDsLyqu43Q6OjV2+4NfpTCzmPytCL4S8+wgQX6FolhHDLf
hrk9uYCBA2/2rFXOaKnxqyc2oBhlVoe1YO3Og71KRCPtD4CfPRj3htaNY5oDeQUO
QhjHql6eaCU/vVZAVcw6gP/qXnLzMrs8oE2dWt4yM8D9hpbOn92D6n/9iU4w9QBD
ZZ3MpxaE0UuvtYVB/wYXRH4uAWNQdN5SRTuPq2aZ7UbQgf1FBlf0TwgoQ9sN3FDM
Pnjc0NxsfhtCuZ21fHYTDAdvbQl5BBopaeizubgbKro=
`protect END_PROTECTED
