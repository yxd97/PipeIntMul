`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCtUD7jtA/kE9I5ZBuXy5aURd0YtW1U5Z4VZrl8B0HWMZo+nqfPpVFTSckmNci32
+UWZYV1XDdsoiNPCflmIIYKaEJyMSoHutS+/vV6bUJge0r4p3GSBamtX6gt6Mntb
oO/LE9vJl+UqaMUawUMMUWo02St7N+n+KlESgeSHyD6HRS31ljBTA4Owmf8S+vuD
gDCsaa0VjbmS+1ndUEg6Tb+JF98gJJURKQYKhwfWc+LvU3XjIKKqs7JErgfP04Y4
MEJMVbejRJbBpjKliUBkC3Dq/gWoexkHQuFmjJF6kzOP3dGcDUZkem2WhwlwIBMP
CZaPzNoZJKATQiuHeoXTX57X4rSuSH+FFWzO4f/EVvpSPQ2v0dw9B1C+ywA2CUoq
jZDNhJazvvXnahNrIQWB5CrPKLAkWb9UBmq600/JzUsBwGPPIkfgwqPB63pT9CpZ
ePvHD9SNDetYq5+1lfCISw==
`protect END_PROTECTED
