`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zze3XzOfHFuKOrpHXBhOoY1tUWIrbyLe/v+/Qrwr/eYhaLx1mi5nA9Nzf6nXJUGg
9v+B+T+q06Bh3Qjnn/ryeSi27RcqnSx8jMKlqv1F9vMuKHGhLoEl1YofU1j36uz3
MAKS4YUVgnIrbWw4tnx3/yhsqwCCVovIWKghau00zrNXJUwGvCcsNnDnVsOuna7b
/5A6g+HAXfLWi6tLkDLcYi2nm3pAxkfOFTsjUek+IgyfTRRL8JnCE60NkfIiKr+4
A6TkiCIUwXUZb869GqqQgHtvs3ZNl2JwaqgYJxqMN/2W01QH4E+59oF8VUNDT0o9
h58MOoioR8m3HcMae8fa8lFkaDzztBMQU8nqFJ5j4c8ylfDdYIJk6rkDkmynxFct
b5Os5uy+8zBl+KDVGxCRnA==
`protect END_PROTECTED
