`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6ynzYolBnjQXyMeOaU/dmkq9GMzrThHEscBtG8RA75smwzpq4JUA8MWL7/Ugxsb
IN90tS8eGm++bMO5LbtT2q7Bj+nBtVX6J7znzLEuFx6BabOXsSgl+1WtZt0qLhfx
H1F8VhaoNco/ShInW8EszH8daLqlnsZsVcOhSd36AJtOHg16z5sOmTm5z3acU8bq
/6nouy43OgGWSzHtSKqnGDwqazgmUKvw6NkzBbcGWRrQ9jirVzrESU4fNyibDldm
pX0iFMZ1Vnt2TQk0jST3GWJe0xFrEgpC/uAkURtWRZcqp4zZAjZ/ndc1Z5/Ho32U
2n9SPKV2vws3QRiABFBWeBZEpvVKZNOy/GN/IXVYEwc=
`protect END_PROTECTED
