`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umefRdGG9X++nto/fEwSOa0bXSILSwVzKxPOYYkS35kOcSXKg03D1jqGl4w+b46P
bEWVlF0semRfhrJvvZsXim9wSJ6Ss1BWEtMBIVsSLQ02mu3r1n4vUocttj5WphGk
mh6K5HVMmTag9aUFTp/8r0BYH7Zlw2VS+IweGHytJ0QSmrWDNE92ZOjoEbf/NCR0
OMDF5PKQPEhojm5NsPVBQQq0EuEz4vdvKr5xD/a4TyN8l8nXDT1pGKATWxEWR6dh
j87yqSLaksgpc5lgIqYgzDU/QxXgKohz4ZRsX68mQpDpIhqvPbSoHXPmAQNTewKe
O31EV1Iz17PelRRVLmerOqY+s44juQMciNDQuF+oquOsEHSasF08XxG4I/tcaBaI
ArsWjZYZsh6wC4TdEvN6SVwep+CtIgrlrB2UZOmnqnFpqU+FcNyb9Nn7b/J7wnep
BzLuViSTJwB//wJy8M7ePug6mLIG/13qXHQuA6b2jxuBpm9XlwbTym4E+GXn6L1l
R09eg2p7QisxvWwhle2oRK7d/UUgFpImreO2chd6dr14ykY5qdag/SAUkb+SSfe6
za1N1uEw9gtAT6Tb4nLH5udGSoglt5FMBO/CGXSUhM0peVP98fwfkMxxvbLWabQQ
XZhOlWrweBmsJQgIueqpbp06M4SAS666/GTr8iuW4Ns7paqaod+/9UTtfHZ88oVO
fQmWOlP6Vez9vxqUYYK9EjY3mx4oWJsvWJAYmtN+sHxFcJoweNIf/1APRrUgTDqV
dpMBWzbgamITXV3sY5JaZ2aQxzlsVJMgcJkDy3OAFoRPmeKyQmaRsBKWwh64hCxt
ULGwktb75UTyhSZCGrOs4BT2RKvg16+WonaMRZOEYyrGP2rxAqr+SooUJbLBgiJT
q0bMM8QSzP9flWtKT3SfqHyXbGMKMvk779JdpJP0zcI=
`protect END_PROTECTED
