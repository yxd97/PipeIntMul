library verilog;
use verilog.vl_types.all;
entity IBUF_HSTL_II_18 is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUF_HSTL_II_18;
