`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FJVFZ2qiuZf0iyEfWpj82qxg9V8lRBsyQ3buULJ0Y3+RqYvNizTp7bmgGuh3p9iU
ma3x2rpiTbNMKgaYAfNZQ8Y7BQrJbyIuqa/iaKajeFdEf75JNiIxHp0r20S1OXMJ
W/W+Wf3r2fJnCxfhIBTxxFLQMC5oKlHqOvgHmGkNX/N854d0VBpuPM2pe6FQp3LL
tJnablG7v9lAdcn3zrAYUSgDHtx1pze8XrUHQveB2KuqPjlRWiGxEL8oHZ0ZQBAb
LQNF9EXtGeveqXT4/7rHZJMkAx+p1Ml+yU2EbjCOKGu3HXw/AYQUbaPA82xEhn4T
e8bAexYslCt2aQTezUrsfM0iTem9obSRX+kX08KjZPc6NvXurbZh3IILHzgrrFxy
GR84MnFQeRgEtLMuk5MAcITsf20EhuuCK/rV9Nt2zL0flPymjHDsazAEFoZqzPRK
gahk10M/6zDoCyMWa9tuLj3ZlMLuHZpkbYKUNRiXhdJfiEr/1Rr2MU8YuGirGEPP
8veTzbCxb8W+x2sjr4AZLtXsRjC2zdyN3JxVM7Eqd6o=
`protect END_PROTECTED
