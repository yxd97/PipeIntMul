`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OsHayTO6KZSkWmia/hc4F7QHUqK9VqXWgz6z4sNJeqkO8mTWhIQpcGW2MOrlVtZe
gyjRtEF39zTWog6AqXWwjGddmIfU8naSuZAOnKN46S+xyowhUwa9WwH3NS88Zahu
E3YRPHnU4I5xLfveY/hoAgMXa0lbaKvG53FGHIm0Cw3sRBaWbbEj+Tkx/b2+QaeH
Q3Z2Ih4eNtCjxogfjv2agEU6EHv6V/5PNCKfbaNs2OOuPGXHNTwuSSxTwPYMi6Ez
qTvIN7GdtRJYLyvgL3s08anPoJBb5J/8BS1EqZe5QLf6HiBY2oQsCi3f/Q+JCDTl
htCDN3awzfZVh3MZF+quMZqMZBoRYVw9B9aTQGSe4QS9PJisLl76kG9fp332yibT
SOu2Xxa+0Qvm9Tnl5Q/CaG1EQvIXNrnD7envlRfk4TgYNaMzu1V/qhUncsVy8nXb
IY8/k5FLth91UNx5XvmkUpkjEMsY5/d3+L0OANylBhkDlhIQf2LknBLbtymY50Xz
il71knXXc0UIpigFdC3ViXEzrVF/Ewa3OVnA+DDCmMZ+zDjKJLSs7h5qZexEfMHM
yoFGpiUZuDHhFxFoGn0W8eAz+G5FJKasXGPyDsLs4PUiVZ5MrITJDEapi8z54hYY
ap2WbkN2C1druFgexzOHyWC8OlDvjR5r5S/Et2lNQ3txuIksBoNkXFN3Q3ixvLZr
4WQHt5vGkyjVGE4svA6zfo3GWi3Jg2hxv4GQuiaceQbxG8cuX1kansZ/k32amrKp
66c7LMm/cvLB8UqTPQTCQRDuM4qq6mt9jQgD6RBliYsO6PzzYfepoLOZS7Iw53mX
mn4evyub9yLYqPOaK1ClTm1UxM8CKoXn74YL6FvX5XgipUPJTRFnyX5Iw/vVXBqn
xoNrGzfjXqaPubtWP7fWndiwOyqnW1/w3mWkJQL7aQUvpXlKDsXFVfvD55yhAdD6
ZBJHuJtNhl5lIeAh7gDzG06nL7nqIyjv3VN0vlTOSR0S5m2JPzWUcgCsYjA1PAjO
Ev1a6RM8tQ7nMxBl34ytfNXpSI0vxSXCZWXzwXe6Tn/CDLqfpVLQuLoFQfK3CHF0
4aSmhN8ukg7SQFuJXnqtb/TIcnAwMLFHfwW0TIT8bI+HjlmHLs+l55+pNcMEMwQB
OKvS8Rn3qkBnL3kuH2/+sbqqnfNAt3BWSPxuBuVbo1sGy2mBk7kQUGttdceXRbjD
nGpQ6ITLq5sLjzqJovGIEOFDJEzT8t791ilslnZNrSYGkm2ZBMuNR6xU9tR4/lK/
NJVNvaYx9tZllzKrLnlY+CIqjniyAwCdaIl7VBF0BHl4lyzfp5LRN6GyXM+dTL5g
L9NiAKWeK7lzkQD9VqN0DUXVmot4ZT8xIwNi1v7XK9wbzkepaA1uXSgZVprLxkg3
LRKfrAvNeHzRaIveO5aog7YxslGyyNvvYugD3QFkfGFs/r1h5ljPQYC+erkCUrkB
l2a3bOQQDG6e8vf5NZmWyBuYnUnMtEI2OgEjlHS+d65qJ29NNIswFifi4AM4xohA
vmahIQRLsiaacJoQPbwwLDduqXgHtXHDensI/cJxLubwW/zSXLgyZXRfyT4xyRzX
y0vlGTsSniBLccr3AM/GBw==
`protect END_PROTECTED
