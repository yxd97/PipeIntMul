`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MzySreKoZXzOqxx7Lj5MtQTRJ5rhqy/PvQUPRH4ieJAsaUPn+X61Qpjc2mEWF+1Z
i0vA5VR43Ci3dV6w63FKpPvhOv3mowbzs5p8RHISttTi/ZDSE8OGEgFhi8HkrtNU
tgYV7+CM9BmIYicwX5LKI3iDJziXxFQnRd9f6BGFlsWOu/mgJHk68bn/t0II4knV
P1TaIf8iVUr8bVQtwUR6sHRAtwp17LbF0a7LdmZsiJfyplTADjrhNQgXvhehL26f
THKI9B6KLeAXNHV5LaCED5lkX+rDhR3/70wq6t09I1lixsLnZ2xXhRishsvovSvG
B8SWJZYyl26+vwqK9xLW09V9EphnmNodG6G0MeU8ymB6LB8sdNXd4tAeV/6kZm3j
nye++YEAruG3Fs2rDTp2b8MglKIWJrLrguWlRAxg8kbULwX5plCE28uCdP8eZRou
BNIXgy/0Bl6lUqLjtzvFfpS8fHajkbyVxBFYd1VFGtXjkylVPFoaZ5kqyWfRnFEF
eQ3MWnOnIB/MdX1INZEjO74NQMSSUAvwCUbRBvtp00KBZtKk1RuoWGASr7tyDMY9
x6t/E2TuqoDZkFMTL8QhUo53dbAp8tWPylLO4gUNIA3IUTrsj/CZedeTUwaoFXX2
Zlq2WWeGAn/aKYukjdQQthATvJKCLVYHpAE9H5uVxx4=
`protect END_PROTECTED
