`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YqGSa6yNLLAyEo1pn8lmwETfU7UMkBmP9+QOItxBhaTZgtd1LQOP/gMmT1yFWvj/
K9HoWo73J5K9MNoTsiyBu5t/3Y3cUz3SstIh6zNNTItqcZlka8up5LZh/vVQAA+l
HJpwhqwABJubsaxY+g0u7UGUwIk2C5Hh2v0tmaIM4Kjx0kiFX4MKk5TMLVfs1KNw
/NF3NseQ/8sU3J3MfwZA7CUXuKD8xuZPBIePILJrUrvbcDr5EGO+ECAS1PDX29mH
VP+GAHgszZIsZ0AYIKvRkq2yERwqD21yECDp2BHTfBhMOZ/7/kOocDOhCvT9k8TD
6CTwgPE/EPMCCYQ90GeSk4X3OiP/Kr97NZk0kGAbTqFFgjCtRpTlrYYgt/3/c6Av
OGUz4/PoeL6WmgJq3gV8vIJ5eDFZe/huBtnMhby490ijWa/jpj22fXLElSGABfui
rpLkzEoR1+zsdX/ABeUyWNshyZgK5Iw1BAmp0O9kQZwVKMwfMQEdKCQwBb8YSOYR
G93NU8NYEm4m0BrY/ogT70KjxE3Nc2ZoPYf+GgFpDTqWoenSLfbGXL5lvb9JD0gb
eZYI2n8ti7THwVYvy+qyuqXiXMRykWYzu06Atc/E1MBiVD0B+biGnZ7pm+0rBXbZ
pFpA29O4RKRDnLotRltQf6CeWCrKCRXXoyqqbOZ17wacgRpp5P9okLfmGxU2HqlQ
+R52RkqenUXnmM0zEibwZiaQ7dIdOkfC1sVUOvR+ZU6LZKNceObTdXef3air3Fq8
FcUrCeDnlO93tTJILoxZ9utt0RSLsMoCBcHQkmxm9FUBEk8eAqqki9cM/5f7lEFO
4Kp+4dH03zrpEMPGsNd4dekPIjQHg+7tySKRRa3Lbe+PV8XOgsguH/palNHQA1rw
lNneIgDt5SSoSBSCcPcAJ9iP/fzniJZLq1KAdGRkQm1kK4idO+LnMtTHOBbijDa8
`protect END_PROTECTED
