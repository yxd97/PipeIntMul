`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yytvsOaSi2h3HlUFyIIeW38c+cFGrNiZS08mcw+c8koGT5FWwRPxwWR755jDFn5O
xkzdBpJqf+8+UqegT24LbJknW9DNu8vlviJJwtjezr9q4sCr06uC9ROQI82I/i/+
JdlvcI7DCVCgQQxs9BE4ScHzV3RgU6cPlFi/vjA5ZahwEkAJpN10s6ZX/Ea/FzWn
3aao+a5vPIhDt/eSX/H2TS7vZTvAKFENWUhH7BRxKSxWgW2wWUWARCsWa9WvlMnV
HmCvAPRRRR3M2iLFL1r/1W9j32f8mFvQa7gxz4E9VMzvrd7E9LrFmoD3608tOrS2
lVKYy8d1jtehMJQrxPKW0hJo0NWgvHFRwFIJPBbxXwRMj7IKJsFR6EUCV+3tAsIh
xNZkGgjjytbnaFK9WWdgv5G9DXe7uGU4mEHrQzQe+plrXO5MF+Ipcyj+hUZ8Shg9
W7NNgaa3Hbmx1Nz+6Q60UfOg7HgWCQrjHyBKp0o7VbURKmIRm/4EXBtwN0k3WTV8
qUFEw207URqz0ZsiWo6G+B/2UJASR+UE/77TMFd7hq8p7CpMUNiTsvWlmoS3IEyD
logdbtl4HmB26+SBWsL3Yd9ABMaAkQqmSCLeVBTvfptBh5deqHDoWQxcWn/lsSNj
+6r6rxYi3rtesEfSOGKmN4bGlEGsOOttgHPs5XWYnsQfyqOmZ7cHtXKazTsgV9ek
h9RG4h72rzJgLImYn4EwL7RfyHSt8U1DaNqp8WooYpqA03nwHMDsZJLoQdzCNftt
DzaQSvduK75uDx/hEzASbClZR+dTfPOCsDzc9pKhR35EgGawNEUa0a0ZCWl8jeOj
iFRWoQUJRg5n1dtAfGK8FViInlzb15yqosjCHOi+7wg=
`protect END_PROTECTED
