`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmCx/LTkVWuKu2oYNT2WbStIrweV5f59KA9KkBzJIrXGKUMPG6Wli200kFcMKBcD
yzkrzZLrCvlZIKVosxOXaYKG3BgKF1xBShy9R/qadiU6PU8ej6BLT3ePtSo1S+bX
TDAVwoPkysgnvETc62pOCPVNu6OfpnRY/zlSivawLv8D+ur9gj4PBFAUP68Wc1BA
53064bI4Rmo0tN8oxajaEJHFBK/A4kNWUP9pnfuQZeNLq1dX04wwgP5FMrAe23BJ
poCq9wZZ8zHhJWX+2HOzz2C4L2EzpwLUoZ4Fwdul92iZtDSOslCkMb1hTsdLQA6c
P7DALmwIVzOTlKtBBnPVOqzSiG58cDyhQC7zBThJ6DwvMl8d/duy2YhDnITelchw
ZGiWgyu1mPtR/ZjYuhxEBE2ohSsAxSF41G82IDtngZ/y0EOgIdFRV/QnyXBtNed/
y3tk9WKwjHrXBw+d6tQaSfKbx0WsMLulHlzm8a7BOh7JVKbhNQr1KOD2ta/Xx1KX
sWpSuHo3ImdCRKeSvZcqDlOkKvWTCwpIkl7lN2KE/2F1zoIHIZNA5yWMyavZlOZb
S5/Qet3P//0J45g5U11E5pGHVGs5J4eS56+W9kjttIw4xu74lqDaheLHYk+gS22Q
N24yUhCDxGfdiktxG96IsbeXsnQPsgo0NhdXn4abwyY6DQJy7qUXr2apqidKDOSn
`protect END_PROTECTED
