`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hoqh7lbHjH47p1n/MhpMlHIHvqRp4etM4LhyN2MbL3k/C87zpQVg9THGYocJTPSW
sVzn2IjrrxtUbIJ97vzgjVJ6n0jynsxOUfLYLRzyKU0NBgNlMSStZQV8yfcB9qXP
oeYQPiZxHknUQ4P/XFYR0OJM4RVFdwE6izpXLd8bgtdUurGjxf01FIAXWGLl7xye
GR/H3Ag3t/bXW60fv3m8a7824ahMgi6IlHh107GKO9yAR9+A0iJhYazR1owfxJ66
nmmF6k2cWUTuJlsPtuc074AxWxfW58/HwEYRILjWQo2xDCxrA1f6jSJx1zc1kLeD
a5a0r2R/yO6RInPZl48P+eWZlUNmHZ1o8wA2etSZKmGxzzULtnLLfysKOyq8/aqT
`protect END_PROTECTED
