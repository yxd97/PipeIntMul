`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMEldyYf7vQkq3/xeyeD+MQojvq9r8mFvo3/hpdHtu0uaWMQUt9/Gi9HSKkahOwj
y0ITCtl19CQncInkOmgtEof6TxujQKe5Z7Vkq9ogk2rOlEp1Hb8pbGkYzFHUPtZw
VlpREMNEPi+AsyWHy7mToEhDuOnEhdNehYhkfHzCqEajf5/7ZdOw4K/9Wb8Cnw0t
0xcX0iKvjBtbfP9P7xPwMa6PqXdgTz0RMBPXnqyS7cBebC+wnd22E1zFA1rbmKzL
o7E641636jnRECmC4X1A4opKFWsqd8J6M8TQYNi0s97EBaz7kzImbrf1N+1dIyMA
iXLLpGZmc0s1zUgkGdXlmR2EI3SBwr9qVRlvi45JsXWkwS1OsjaL9C1mpLPQngF9
2Y34cqqZzD0QohJRbMiT2KVO9o4hZzVRLkNc4Pa2deAnn/1ZE9mO45rmmBH1hw3m
HkYs5uxgvnHhzunTxa7z3F+bi4v19YSLaZ07darIN9ynbFelIQPlsR5CSxOGhPSl
N3fbPNJV972Q2CjaOPo4dYqyJIAa0lsoa4zND4fUbnX63aHP4vIM9PeyKj9kFZJq
UqghlCuBKqrM8kC1AMA7luz5JzCU/8IQL9tdIlH2Xdlf9c3ijVWtvdN1JmC/k9bc
eoGFTSgiIeRn3/keIULFItNRftbP2ns0qt2aAe4fUkn/ZeCsBTJJXaa9hYeywZpJ
uHzzzHzcQWmFUq3Mq7dBZRSkO60vksFCz7w4M5xWjt5wlr3AX5Fg08XavvLhZkjN
HxXxefuSF/nnOr0hNj60MEy4P7P48qHlhReiQ+OCECz8QXRSd0uNHaYASpvQBJFx
UrU27V229ivwfrwe/6LQtAX5D3m/43r3jk9sF5EPVT+VVZX3WKyvXPnkqJJwsph1
Pgc8G3laThADEQv9IvbVqGTok5SKWZUiWhdPtkjZRplrZLJgJYwU/63BF71cfVtq
CTv7Dwj6McJft+3cTCBfDl+xNjRZgMDbll5aAP1jXHXQLSPOD8h5I53iJlg2TLqX
wPoESNZ4mwV8qpi/h3ZczAT7wdP/rbkR6MAKU+L6YbSWX/ojikhT9Ty7wQf5kuPx
Lp78V+4d/0Rlo1f5nr0LOE9JvtEHMiJIl9bWf6sn2b9h+7yoFyHN53TxT5VYAmN3
FQI/qimaQe+cmuPN/MEz4KftcWEGtr3AFyT2S4snuVwSbmDtQab6gXl8tXtsvhgF
QwPUjjft3U1EQqtfLQRGp531j/jT7Xi5jVZC1Shgk5o8De3m/paBOYMRJ2Nrx315
+mayLjJGTA+0oSWVY8fllIeDL93gb5FNxi21VsriwsouSzWsAnYvp/1636oNfjJ6
9i3RMc7SrvyeX8Q63YCz18e4LsAaA0a0iCI8gZwpyQt3VFY2lo87Bl0/e+tFQE4M
mTUJkszuLt5yhQXnV1dmBRSWkYOvICXSz0fz9WyVK/FSbORwtv0mFVl/QsBVtepc
r+4NTVRNIjqEux5WaNK2SVKoaFKA33CLtJBydOLSvzNE55jW17wEE7D7iE03fYR2
wVJXP7qwM1Id6PBZNF0LoJMT3V9yRE2KzU6LGk5+iv/7DU6OoeEMjGUrQFi24GQJ
XEiT08GgE3DWTM8yGDug+dHlMotTzgINT4xpHhgir3yNtY03RRaNKuqwDQVmbjmI
tOvYoWjeQDaxNSP3N1qUtSvZEwoBXZOA1HxPNIysrMV3p/vQpUQwKwbPy+Qc/3+3
DPZXnyU1uU8RFyxZ3FJbowldxmYG+iIlhtRSyLMgI8++ekkJaoziKf/tF6dJPoHG
BJXlAKON9D5Qb3flN/rg/yxbjUVjJAh2qH2Vm5xMH29IoiYbRt+m7Ynwe7PAVZsC
4+JcS0SZrenXkRo85vKJMWNX/ozmntSYc5qipQkK3lompVBMRNFemgJmXvExPuna
XYXOcpAKhrqDB/bR88UtlJZpLyapQRDQDYOszcgjBWxTOkJu/4+8XXVpy5/D9sr4
4MTfe0tdAIihSAsQc03ug4kVUTxYg8E5GsSzWy3O+cfGUiCA82QeDXsZyGVcYAgc
pSDs1FzAMKX3/1MEUPGj9UjaR1iRd2hTivrxNqPlb7v/s2tSj5R651CWIqH4GrDg
NkS91CkKOe1HsIC7vJIivxHCr0aOVvoBALwGq2e6rE/QtMqzWvSCDzbKw0+p50oX
`protect END_PROTECTED
