`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5+lbkN8ase4u3eyeaW1cLJZcmBz6xqgpaTfn5OSANO9mBpLymiCxXBZYszznKlL
41Jul8XFFzViQMroBW0upJTTmR9p2pFLnUc1OOBNeEl3vrr8Gl64h21cOX52u9rb
hOE0AmYZYMiGnUr7si+UML3pRDu4wIFQAnQigSdos0oW+oCk1F/5k+JLxnf9Y8J7
LXaYXg6uCqDpmZb9GFO1SmJfpzInLNWinwWxHXzrvfS09zMww/IeZj9oiGDlqPs2
TbmFY0Gy7nxi9RSbj/b6VWbReldhi/otzv2nRF18iF1gZHKy4Cn7b5/go9zWdzhu
f7qkwGPuCpC6EDFDFcSC+zbFKK2zu2o+U1qh4pCFywG4kxXWyZJBUl3KIbSOM3eH
tz3nwroAQskVya6quDIh7N4noVTS0rD8uNfym4nfG+ZfCzl0LHp8kYxEeK8Rhp00
aug8rLN0qghFYiLwrrkUl+x3IipYtc9ljwrklZQyV0xTT/tty3YR/R5kR+pJGIc1
`protect END_PROTECTED
