`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EXVBB8znA2hTQkybRlb58Ub3sQxiPCe7pjT0xc2E/BXZuG2zXaRWhMWcJKTyEh80
UwABevWHkHfh+793shGm2Mnw63toQ39e7wi95xoHG1uZWQczigRci86RyB+htN2k
C5aq9BbRM4x7RH6IoKsmSrcK/ptgbfXISDcdMTouoSxA6qzhv9INggUwQro3OaaL
kWz0wex8Lc2kS6oOukYDAU/p3md9upwGEIrx11XmhGAJMHXOmfuBhWN1gamYte7E
eZkLAVE9FzwX5JSr4937wws+tlYeJoHBZ+25ErE6QCuf4YFgnTexJmbbI87LvL7a
TdIROVMnOlNUc7mBXhC6rtudW9Z2CXbRzPMGbE9Vhe4xLO/yjl5MZQslM+c1jZtw
NIweNur6FkeMZbwNrTWgomxL2fZwrBaYFD3lXRNxL59JCwn5NoXURA8eZAEV9WSA
cc3o2aAT2Y184N1wDc+gG/pNaqR5F0txfRZPDAP4MSVa2NW64IoQFndjfgMCnSFs
4MH8/w2SvqFHiAdSOetorpDZsK4L9kyzKwQqsgnsp/t57MqhjvEM87p243NXT7Ul
yDAc60fkJ8ZtPSF6/VjCCXa2n1YGar35/vSIepRHNvVd0bfl5UZbFto8flLb335G
bhxYMfwaOEx0ReTjS8BHOVRyg+DEUoEpzSHfFKhG2XuHezrqh892q6iOcVOUVe/O
Pr8tx/4osVNWumbR/WSqHbaL95/LCZLsse7qznleQQRRjeQnAIqqi2DUAD/0KegL
`protect END_PROTECTED
