`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMJ0gadU+sGNJPA9rIEitsUdurSw/DYQG/o6xtE+MshUgJn13kb+VxAm0mfCc76d
TIpCgATG8nU3qzEz03A57PpQ7THPz4tRzn+tBjnkL/UvBIdEm9xB+k7EEoVRmfJC
xUsFstFjCN5K2M8tCxN+YbdIS/8edXkLV2qZXzKGsBHVciFcHEGwVk0Rd1znrHlM
AHGZ6Nn2N3S88vnjJeXuV+96J0Zh2LxX4IJ1qv83zwepGrZ6CMRMBsNWqMUySSEv
s0P/l7IQbV9TUPYujAoP76kn4bARryeilsGN7sM8jVwbVWoPydwFqlPUkGu4Jxfr
0pDdkC6aJqLgm1cxI+YrfAiF98uq+mzdYI+wyXOXOC4hkqH5W4XLRz5SkGQjPDyw
LQxLrfReulYiGklLXK9i2x6lVL7AtPrt4HBsFlpndL7cK22D7df3vpiVRfdRSWhx
db6KrWALJfH8OuIXVO9EOKavELRKeIpSCGPSvFlHx8xkYop2lgglPr+sxpYw4QDi
SFICL5K92hViprRW3hgoNalYxaXMwTAZNhSbvwep9xBHTWbEG4msQlydj6X0/t6q
iKnD0rbD8MAjO+wW+Rkz1YYZa1fzlSPuSAcNN7pCBPtDNRa5JoCpS5zbRIxrFCO0
4zNGaun6K9CY7k37Dd0jw7qxAZpH+sgaWJ2EA1ZdM8n7/BicPvExouM/Kn+NG5GS
s3tyJ7d5+6M82y1Ng0sp4kSsRBcculc69VzkrdwNY8Z7zT0AFLGjksRSVIZWAqm/
Rchk32wMw4ldT9y17kjglsxxkwK1IQBYfr+7ZlgK+UM66cHKKxQU4B+32v2TL9sS
eWFjK8ajKJdgsQ3kc8bcCkNMMB6RunuRz0niR6q3HhW8AmJcMGu7SHmgQUx47ynM
a+/Y1JOZ4j7/zcLIfCh50Q==
`protect END_PROTECTED
