`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGcBcFiwwphfPMqX0HkHRAso/IQUKer56+Ky1RjOeBEwNFOg6U4EylnvGXBMha+H
s70znBFlvnFPPm9R/ZcpnJVl/RnqFdwFztIKAhdXkci96Iq5sypdKmH9ULgBHLGD
Hax7DBnZkFVcl8eWTsqs1lcXnlo95RBtA0mDlGFGyGZPxbqc8clHl/y5WpB+JDGg
4F4lczioSygUiyRM6T1StPYu1SOBFXUQnJC5roJPMOM8HmTgrEo+zwpK1QWi55TX
XM4LCTxqYfm4OzkK/yPbyfeDDN5Bf8U2N1zBPsvMr5Qokwj9r4mv5GKIoEPykIW3
UA6++k1RyvaW6eypqxxCRNHH/FXCpeJ+JkMfZjf4J991OtWLiONGv9AomzZvbMAN
ChSYfundtdXJUYKOipiiCdUQzEOxqYtzYRDR8DxjFL7F6Ysmq8dHqKKw6BMVm6HX
s4TXg63mUOvbbNcuvHdYGzfieWzAjgoufk3dkSN+u0Nf1Kit1ONEXtn8KeYpRPEt
zLbB6M67dWAkDRvzfU9r2zsE+BzApNwirV9izR2CesOtTquCM7tS8BXyNzylzkrH
MOu4KNX+WkQjCleaz4dHMg==
`protect END_PROTECTED
