`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ceZ9HipkUl2NcEfJhQ0dTOYy9sJTMMKYKtmhOa5vXXXVuTk2lx/HFHBYITfBOgs+
J1/nzv2xvt02c7VDWVANxEM1IMipDyJqy7cjlhji9pJoUXLndCgB8S8E2RKdCpKD
SgduSdedmwDWx++GnjsR4p0E6ra9wU6BuDpAi9IlXBC/726R8Bxz7E4fUvCHQ76A
bHxD5XsmDxMT48a2eIHhW24m+F5XXY33ghZheXG2EhK7u65/lqOkIu3JQq7yECzl
kRTiQGTapXxDlCXx8ONoyW0YfErp680Y4PS6YqqWWliRQOzHUjDP8tvbVBfBzca1
Wk1rCaMWC5HA8tEK46WslbChfYVw1awOIKM+QdSWCuxkePkMTEq3/YPOGcJaOvtn
I2POUAOn96JQDGis2t+MHz+mUcf0sUavNWsYuPMZnUE=
`protect END_PROTECTED
