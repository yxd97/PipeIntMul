`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCsCPO364hW8krOXHUjpzkTU7vG2mKUR21Q5HB+1ypr7EmLHr2GneVdMbYuS8hMB
ukAnaF5uxOtowG8BpMaWhVj0p7GEBm5vFv7E3cmlTiK+PZd8bfVWdCehXIcfy+vL
DCgJc1WsbGxzp+dzESnHT8XMyMr9jGowVVRJv23jGvO8CHgb2EGRARbf7mMraTXq
0YVhIaVzngvPJQiSDB8zk4VAFNLmwwVO3+E5FuBHG1qn6zJ0PJyhYKFEx78MjmY6
sB9eGsnSvxENeGnXeiTukteLxcq5wfRxscDrJ/gIu8IzAV5YQMrx0cBQ5n5M5ybQ
yen2kb1oh9q4rbhAwHLU0NspaX8CqiKFyLBUZypjgZElJfGSjSyddc17bciv7kQi
uegj/UJJjlsM7sxy0Gzf5SPXLWMCs+/fzjDQx1PSTUO2GdajmuYZonH3X7iM+ZEC
cKxKNmTEkLAfPwSn8msxm/trN6lMtcW1VL8Ng9kWSMCUI2ImuQsNKAB66rU19N6y
/tNeFR0QaMLyDb8t+6oRxwTRIZzH9vjcG4EGC4nj8aqjBuj4PRJQcUGim07oZoOP
OFGSCRWjcbSHHrlEn202+k/McLbug9nB70g7cXA7jSMlevqe0mELInHMugjGTuA4
lSqnL+pe4r3H6HBqmDxGwdmbAFnD36k6EsY+3amDcsM=
`protect END_PROTECTED
