`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLIJ8QqkUheGBUJQdaVFHYzlZDnyAQ4A/wushEiAepg/SWVNoZh1ljoF9a1+V1sJ
zWE3dRcDnzIEpfbPlTSdWmsWAY9wn5qJ9nI3OuKYYk/3Id2X9tOdmYoY91fMG5pA
lSBwJ5zvHJLR645uxUe50S2ropUUZ1CTruM9FZlwoEID+JDspc2vK39+tJ1KIBma
eXUZT5u4+pa/CRjw3OTUT61LxXdQfPCATGJTQPqUuMQd4x+82roV/cpNEsT6CqJJ
CvU3TsbEA73iR+kY6JXt+Kj3sPg5VSG6Mbp6QLrnFmnM/AXHlqDgDSLwC/bsWzcZ
He1r3rWlor6/FYEFkoG3Twu6tIcei7uwbZUl3Ntk53DFRsM6cNH4lYYOul4/apS7
TpgUlYnTRFz4HIgcch75M3tZ4E6PLlMXzfVV6rfbBCcPNp9sbDquvv2DdfO6+efP
MKRTIeYYdVb0YNCveudBsM5GsSHeDJjMNPyggdezHvGWcSV3HIKGlz5ERP1u0aal
NHWZe4pI7uyBPvXrSKwVrGQxnAYHPhxSeU9770ni9d1o20rUDkpkRdaS7kGHcTyA
LKgj22Kb3Ye40tQr4JliLInOUf9M86+DcmUCdi9s03mQpbLdsFK+s2yO4MRR4b0i
alA7IYjLftutUTTl+KXVP4wqTIkxMZW9O5oTl0/XIrywAW8q/ufAJjeXm2M8mImG
xf78mrPj8IGWGRzJSTRsgLMiL8IvpEK8VB+7LY2GhPeAJLJ/IMBgOAwXIOxSqL0y
NCAztDvbWAF0TFbc21zQsHFiAevr2FKK4NRfIlFgoigBywTgttP18BGBhwOUDyYh
XXLdp4TX0WAbqYylZe7KFebW1w/xFvOsxN0KCBrdOYm2AJtfBZANe9xYMMmDhkku
2q1HVHar9udtPKMm+/TRow==
`protect END_PROTECTED
