`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gzlEra7DrEPSGjzBGuIFuKUKVisB55BXK5sX8v5kkEhrZtcFyam2+el5p6DW94mY
yK9QbVtD0qGSWr4Z3Ruzj4+p55xB0cDclxlR3vjRKVjVJv2XPaTai62pk48cB4ye
hDOJTlnw3MJPcTode6o0w0+7JCvEfPwvX3OWAhnJ3dE2goUlBpowY4Zim514Hxrv
vSaRwA+G25SelQ8cnpeLsx6WDvnB4CRlxMHvJPN8rqSx+gv9bzo6A5rJfWjEuYM3
1uhm3yX/p7JSEUYcfqZ3LcGLdyyWzxX+cOyZwkHIy0QxxpxadLpCIQE+MXwHhF4j
f7pbAGDscuiG92+ZRIpHJ47Bt95FGJDesO0IMBwJ0xL7xN35SOnNroEiVnnBl3g7
vUdZwY2HR5sN6OgAkucElw==
`protect END_PROTECTED
