`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1LvbQXjF0vixqRwxjhEYO+W9hrz4Qjs+7fjsNgXZ8BcxnEzpZxAYK34cikvqezKf
dYb+M5gsGO8X1eb6yysOrztHtyfz1eGsh1qDhNEqA2AvGtrutiW31x9KAW/Nfiep
usEelNBJ0wvw41SoXGedJSrp8cG43g/FtldXh3fVA49WZQ4b+5IamlQKXuQ2RLOg
KGvty2FQhoko61b0K6jShd6Yhe4Ykh55FKgql7vrKm1T+srm2HbusbC+5xesb/Wg
c8N0gDTQ2SU2Zuwa5WrDHc1/0KZvM1Knh/v5TzW7fPQdgbC83x8uMhhFl0OEQ8WW
xPMG2/9MZ0izCjy9WQC+N4g30gDYpA9sv1/fz18qahbE/7+zUk0M/ENWHkWRE+v8
udUwhR3p5XVEj36KYgh5Ye8nCYgIuzJLsKhvItIl4vDSpY8QmvPZyamCROBKWER5
1b1yNq5di9t3pNOtnD3cfjIFy/U1Sk6kcDDPEhlOdb15g8tu120aoX//PoJJRuT0
LXdsasxqBRaMqbGuJYe0joA0vBA/5ZouT7G0UTsA4CJsRC3OsY1GUvRk17CMSEFv
`protect END_PROTECTED
