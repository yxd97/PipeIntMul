`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
apMyTmH0WQC5esa+M5DzXsDfLIvZIzD+XUO1kJtdBfXMEPo9yyfMuJWs81S/nPdp
SFj9NiCtIlLS6cKRy4n6Hf1ru8BaJm6unaCXhUjrKci79Y6FBveV+WsE8xphSuPO
HikdPJ0hgqKEPkbI3/2N/G/99PYkjZUWNVD6/uNh3ZGY90I/qrLMJ7fbZP4zoeOl
tOzFjdcWucwpE/vszZDaKvcD07dwYkIq9v6boAx1c3XzFkftNw58JEijkE63u7B0
ywVM+er3PfWBRgsCfHbgkz4a+URuQ9gKbLv06GtUFBkOhAnl6qnYLszSXjkX3TjX
ACXwaGeTLz3aehMsWHdVRrSSzMvWEg1ZdDyJavs9YDAEnpH8GaVuhf8Yum0t0leW
+G7EopF7zhty5Sr0E8VoCmw70AXVstd4GXmabGydLBLRjLZnKwmMbakvgwFoI+Oe
a31oZBXqczROrwVvqrjy5dbPfshOWUXOmbEKZ4h0WR/77xtMbaQ+RykX9mxOtt5E
en5xjNo3Z09aLoXMQ37N8Wy5I4ZL/0RzybEWUGrKbZp4JMyVJAms2o8pHNrG5Ygc
zzmMt/Y17f5dPQMyt+MX6vRLdXnzE9+MlXU/XBOumiq+fvJQIJhPMzms+e3oXQU6
J23WiJXlS7/mNKOtQ4xTU/MkQW9RtEbVSN4tu1sm/iMsQZ63BvoTK25tRGitXKxI
0fRA2npgd7xBCkwYZk4q40FoIj/ObyBZacMg7cmzy01vxDrNFTwGEKtigP+40+hn
YeUvBAdkoDsLacCM7jgwZw==
`protect END_PROTECTED
