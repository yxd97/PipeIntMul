`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rIuOU91pUata+lvpNHvD6VA/U3myPP/kT2Y0JmL/yxFbEXGN2DhFpMW7qZD1Be8
YKpS1FMvX+Kf5Ll49M0k8aAC7vOttCAsaaloLSzOGOC5rzJxh0/tD2SeUTj7DcKx
mscIJOBFoAYhMaUKnPlovDx7F6kUZ78rthjlp9tHKcVMbC/ibY4uKoAg/pDrGUdP
G3cke2PGXpRoA84aIvXg2iPtP/tRVaDTgjlxjrqr2W0cmgIo7Ag72PBJ7zjRZZxi
A+hHIMGity0RYrFhnorUSxsRjHlwbPwau2+uUN9WyNGFPPxEK7iLD94PIk0AM/6y
FQt56IN/Ge3zCRxPbsterUPMdR/I6VFeaU6Q+yrYACN5eLAvXjYNj0wfhj2IKYI5
pvHwe2t7ALGseVFepm32dyrZvOrixZCiadSOG7RCROGz0BM7WgoiIyBhvbk9OisD
VOn+BNOW6fl7GDSUZj81M2QSe0SdRjNYb7e14Awm/Jn1b/7eoqT+MsR3kXTjHq4J
IzO0Vm3ejyqsoCj9tk8Rkwsp+xgjDB+xCxniHUFa73F09PhN/rqXXmn4wx6cxE0E
zRY9iQElyxW3BuqzkvVpJyr86xtCMpq0+1DZBI1rVT+D8K0M6VpmbUgGpYFIkEyD
Y3CtdG39Rh8zrDNlqOgFeAlrbEmbop6zzY4NpJMubMYjRm97pRylr9AvFBz0AdTj
FEYdb9vOdacc9ypb5IV+3g9AhDeNB1Uuak70PuDlczL0quWVJxq+RTF0set2f4pD
xaAITZVfhG0roS6PT7WSblOFfejkCWPBNm0izNVqamR+06tP/kNSA54GMj3mJ6KB
Lq/G2RmkDO3RUsPhbRc4M6g1jkTbTK9uUXVU34p2unmCHidGHjO33brmgFuOT5JI
9NQgCBB/vywA8vw332IWuH3QlPA+dNk58G0daEQvPAi8ZdQkyN3T9s7Y00dJV4p0
Xc8yWn5RJKONjVDfdFHC686GwT41PmNIOXJDXaEYPQ27b0IRn2Nk4NqgM4BT/LWV
pAWh5aofL+hc7MxbTa6VBfE4e05g+HsRbXB6R8H2dH3i/aXwMaPub9BSnCsjPnk6
aGml5+nEwUZJj9KC5csG3/OGq4IiBAm1QplvMMOWR17x8yiPGKn6ubS9ib7ZEYk1
8hDAHoR+XMi3gSxNgQvVqDMPcZV3Gtzqu4oGBFcZKcrl4lZZ5Th717T5vZk3fat7
WmG4Z96vE0PCJTj5Aueao5zihBDlem6ci/Nwr5ztGnyfFcrI8eGEq32/ZIcAxsba
/ekWHmGmEX/JIBrLsOS0NB2dAuukNiZ04zP9EIlf8smau1r6rvi+pYgb5gVC3pTK
7JxsMqV1JeQhf+qW/BqZSLe2Y8HMBhH2brkbl1yXlfzexTqy3gdsrbvHf8tXljDw
QX/TPL9PQNxq29CSyk1NqbW6BfL7NSO3mY4TGNxuAvjqBSYpxjZYHSc/flquOd5G
BrPD5vZ/RzjBJRwfLiwGlWiQXL/9nDTeFSNtep3YdVe9lN2cI3RPhnQsxSTaPrMa
WAbC93brP49cWF/+88sxRMHxFEC3SkoyySaohEetmZs/zNZ+kWu6BEHdm9u9j4yj
wpJPYsvIqMIf4FaY27UAnRhmGCC8QOdlPuWSkwADOw8jvLQHDIbnATJ7/fVzZTtP
pN0EO07bgA9Ygpz7ubKhiDDP/qqVvWWCULV0usJ8f8x68oTO6EBY37S8v6jBZPfe
wS7O5wkfPKosxH5IWL6A/lsKIG6DXnZokdwNqs449n04SqlJ1uyPbhjzjCsWwFxO
2xZRBjrPrQH8OPGmW0ufNgyXflY5IbK1q5DoXTQf52Xlhns7ZQbsgT2cppiSIAbS
MEvHFZ/k5uBhHkYjUaxqnBFjCgHnvLLcoHFvkf19lXtqDB9Q2Yo3LwfkH38OhH1A
rAQYPB5608NGpphabtJA0M7p7RZALXBC86StdGOGaJt3X2c9/t9Ct/RhW85j2SAb
1741Dt+vDktW1CrZFl4t2tleXun1Xl1rdQ6ptTkOssA7dRpqdymxroWNbQGIJGKe
R2QnCFEzK+Toc7wJVb0Mw3goS0pLOcIM619cGT3NGFtb7HI50VAgj4ACIgfY63SN
AupkyYhDIogEM65fM3AksCeVygvI07bSeMaNyl+rW9zKf9uObeWZayxnoX03VBdr
+hFIHj16i+idPX0lRMjWoy94hFwY8OQElqyvywhheVRPqCquiZ4xVS+3ZMfJNtiX
pQaWhiUs0343hafbt2VT1amt1RNZaRv1LVgQW6GGLbwaI6mWuI6X24qsbcC2oj6z
WEKdUghvM7AGA8+tY6jkUXe7ptZ5ltt6xuheRwrBBhWeR4GxCrw0YD6FWfNKue/V
B3pmqTrHWVGfvNpSG1fhm9lDvoA42jRc6Ct+OBWxCdIYYwAOVqgqRlOBAc3cnGyZ
uOAyucs2kagTDS1tddFRgHR2iULrXnSCHIt9uYdf9YxkBZyGE1yAL7fb4yvHfYll
qrmdnjKg6nWMiwPCJYKp5RvegUqzQvaAsyvfoivFmXC5PUgvTjd6OiiGB9VzUXYS
XqCcmXpZC3bXLlRMX5rxAm7lZUWLhgvcK3/xMbJjdoC9vaO1mKKWRk9EXs5DHYnb
Ffb2o+TtFgKBaUXXNuCj2ou6y0QbHNycgGR3E5ov0zGXjWhkPd5NXrNMl5ZXG0Md
B55zagHwfcFWF7mvSfMreYD+TkWF3cc2oKwJXsOzFd4BZP/R/CnUYK9xlILURSxV
L6bTkgpbAJcg2IST7xo6NCYadiT+9T3nzUGMSX3Ky78eItecnFE8EZKjv6fFWOoG
iOr0lDrBzGTe3dXEtN8KLs6mcK+y15TkZSzIasoZZwTLemOOTy4EQ/1Yc9X7WyT1
yn5OhAA3e0s0qnFS/urZWjHTvNPutEf/txKmyg/iJeM1P5BUbC1m5wv0u+L5l+9C
ImUsSv9aWY5QEOuBk7qhpcLY4FEFhbhMaXnVPnxqrLozuRr1x+YUE+P9lq3zObWU
/lQjaZBgxgrODfjbRhZl0Bd8+B77UUhHvfM0OCOnM+2AfhSMwu62hfKdY9w2KV3u
shaVygzkRFMXIhCKkmZHipJIiXIqyMIwPReXXBgZWUrcT+634P5rScmVtd8Qgy51
IaLqrhG9UTrWTDIeG9uZpAQCg3ntfG5cPFlKCqOK59JmmwWhzEFmLW0gND7hKYIL
ri9sr+BKnjK7x+6t5qkA+jsQFE0gMvpFitACHk52NHjDD1PyjO8so22G/GafAzIT
75aiCg+8zMtEtS/3/0fED2LrXcD5CAhiQ1poc4N/KpM2qpFwhH0EA+be8VERyHy9
vJA9em0RsWraliY84R7e5tV0DC/WrHNkKyuy7feZfIpz8ElRnebU198Zc0qhUxFP
mlGaW7iupj5LL6gEbzQdfuhDfX7RSvHBXPYZW1NTVvxqcmorS+VZwhkWVWkujH0C
wD9NjOcKfRomsJPh2qHLxjTSWhVfhrn6yVtmBox5yFDdc4XAmDw1kGjG566ixozy
GNu0A085u6E5i+SjXhnq+V2ItrLN+ELVO3TGjmj4pVOTaMSXXiNrlqsdKFGlRuOu
ppgHqUyv38PhbE0L9bpjn4F1UYbLxjuUi7l45KnwTh+txQ3waekykYaMdvGLfID8
xdBPef+WsBd7284uVqyT//pjlR/LAz0/rxvh40zSkiuEaHEdiVU6TlayXRGMfVWZ
KtqfJX5Iekqg7A/y7mo/N8zLZ5SD7+J3HBhCEeCzZuyMtm+5gCHqeaQd/hywkmtF
YJQZ/MWJsm0AzjTUotHcMhFrP/4BxSIx6DmUOBPG6u5oLc0kydCmf+cm7ZDLndPu
aebgIYVfbmFP7TnUkNaZz7T6rx1vIVvmc8J7i0XM0lm+yb/wwhZ6MiO71lK951KW
0qZjLLLO63WAYgfNljRVvsjXWs3N1/Ec2x3DxC14VlF0pYSr8zNAeRrvn8ubMWdT
fBOG5eKkflj3X4CpBTja+YbIWCg3gjz0arE3Lafm6ojHd84M/OHObDaDp0W1T7Ff
PjFiuGxfg9buNm9QmgU0IH16n3l4nOLWEmMQ2Bm3eFJjknLd/cEm5HK1I70HQo+B
CWR6IsTNeFNztyV48Fy/JdcHN1N6OyMnyCK7OrKb2g0CNo5ARrwUV3Z2ekA70MtV
p9Os+GOQfuKz8HyzrUc7ydHwU1L5H7rU/L+t8YlNyvwyQRyVJYk/f5BwM0HSskuw
T3PoknDpTpWij4fCbi3x8KdXgyo83Hsb1tPkjmLmMnUtQEBqiDLNi+092g2QmGSD
E0wOUzOmKeoPhNKszwoVe46yRi4bPnbjajZEVnqQEb9gXCO3X+cF6C6mx99LGIeF
VMiW0Zaj+Z71TnY6aF7bqNgcej6adYmSxbenDaYBfIArsLHEIygGCCinwxlbJp9v
mJkbjeCB4Rx3NgJkBwM54+OlSpn8lI1oVpzKZFGvNZpfBvZ75LzkCL6VUoa8sutU
QmBwu2KYrtqyX9lRvTYhFzEIZ1iFUWHWdTuGASfT0U6Zpi4Cj8IBH690FEaPIheh
UhYFHF0TeFUw/WxxwG7OkJRP+gNCV6hd2RTIVhHHWGr48DhaORR8xa5dxE0Gpo/y
MQwN+o14+7Is7MEcxVR2FZBiXd+zHGO5H7LovW33AtG/Zwarm6MVldG7mNsaOue4
9VQQSARbEuo5xceg9NLb7iLVPeKH+Mg6txtGthYIhZySi7UYA12OjDxj0B7XteUn
0e8FlIrdm14iIuJMLudWNUoEtAvUlwPwOgfmDiQsCPkTY39ppG7Hjz/JvAc8C7Wt
pgfe7hODwe/HJn4WgkeO2TWVNxzol1Kpij5EmCf8G5vskM5EvDbv9XhVk5shCqE1
GlSGWiGnEWLBOH9U9Z0nKohNODYkLuVnvD2IWhr1vR3mVTxtgIIIDv1D6itcNT5W
U1m7ljDaDxzDV+W27XIbE3SIpCbItacCzFzr7OMxoCxI318WQz12hnbV4vSrCT0Z
Nw+rQPGJQtj28SQmMopakKKB4eC9tFdbWnm+Q7A8jLk+z/C7xIqiVntLrFe9+H49
eAifq67V/W43R3DPCZt+/zFV3HofH0Bmk1TADZ6iWWiXl5orOYkpm8rK7unMLVdB
mhNhU/LROyRwY8NxF0YSfXuTabcN7By9P1F7EeyNei983CZaGPuVlSQUPnmqZIat
dEK3BDezi+dzPdvK4JnBy5HIfrvA3uftb8fyMtygVhRkQQ7Wmrgfk8LCLhU011WR
Wx9mI20gfJ/X52L3wkRyWFfo1DcLiXM6CB41eeRhbQP3yl7ckYnR8xfZIArsnRir
T9Xin3h53wBtvdHLHH4dmS5cZMJXvlQfFg5QlUtfeMNWrbfPnQesYBn/HNOxEVWI
YUG5fJDxElTl6EBobixd8hhG6Fa53XYQ1SQRJfgKQ+0pAPxD3EnAm52E3GYupPBa
UoTnGXLPtaJGmKsdzOna9bBpWLuhby8hjOc+dLz235awUjU9BteVSrgKV+18daMn
iNTE6stvP9DmACQvcs3iDtbJPJe5vILWhaS25c6r9zu+VfX29YQnoGNzp1XU5jrc
XdFb/wKd8Rwidk5GmGZqaOX3JHTE58K7vHFgByU+W3BV3zMjmxpvzq2bLg45APzr
t09zD4V4z+gtZnNHC1z+WZUHD2OKTfh1L5mZF4cz2wtDi9OyREW9B4PCFq6dniKP
D4LN56SbguDKTOq0mGB+NXnGcAXjtv3oSODXVimfZDPutqe8TJ7tDy1UyAHiV3tp
5a83nC2NqTyIOc4F9t79CPv2apqqVzkY2HgJ27B8UI1IDIlsB1V/JSljC7cl7EHD
ngn2WxG284URMWHik68Ioq0x0HtGdjB8Y8NKbYf6eVSmmskCQnmuHmtGDKukAgg1
rG4TLTevbsAOXynHml0SMCXdbmguV2K2iEiFB1rtKLf7158qtrTuvtOgaSKqIFgr
sFiPemFTwSPknbaqLkqEPW3TNT4Ys0sTDLZEQUibMsz1hX93Lcmn9VdrQRWUoC2L
MCOKY4dq9T2EF5elhadpzbcGarB3mITpp/g6INuppfs8rhG/chf38AUALPXMZwxc
drZzcvEhAotJWm8x40vsICH+ltDpabzf0vdtNKH5WPGuxGJmCyj8kRmGc1fP5nYb
O+JxASsrCAlcRoIdyG/3TkV/T7MdGHvJ2uUC4nqG/gdgy51G/GWDq2X2Hu5ioHGr
rdixJxxJZ8BZNLBI6Iltom9aZLumzNBnW/fwn+meP/GR2+G3vz+hq1jxTMT6JEaZ
xSy/Dg5vMyeDWpNvGwg6eLdkaJiC97K/IoU/GnTLq9V4DMk203vyU7AqnuOeZaWD
xq3A1IyJ8WraOr5FcfBmvkZ4UQLtcTelDugUYeGvAVSG5iHSNaLLtyur7WxkR8i6
i3K7f0voyZEifF296N1pgFAe0VfoHBywxF2EDHHVsC1ErjdsYpQXq1bUVEygq/IR
7QtD9b1ReakAG2RGDhkqq6IvTnYzBm3InVzTpDMSU7owgrgbNlCk+a3loZotj7yX
2b7Ig+m+BgQjaUm0fCrusR52A7z77Jb4M+ZsUVFXJPWhLhpEa7rJQNUUBpYREC7d
jLa/Oa//8EHguq2g0ufXs+Rkj6xQybQPfTxPpoab4a3dHUoSW+LbHHnX7p5f3AZY
II2eBnjqn0s8XVyhr+n2mhY8pN+bCOy43dfwxjJuLPsXuPfsJE118QxucXN5hCXd
39s+xYaa52CgR4POYuCztkUgi7SZxVAJzYFXDKUlNArQ5UbGwuiT+VZS1w1g4T/D
1AZUd3nYg1QUIaHHGCI2/kTUeD+NKP+uyDEZEblteQ5pCOELX+ZZsi6D2k0fiqsb
GR1ZFVRGiNOsRig3OUK668scB3S9Y2bTNPxYOd5RrGxeAqn7HuldxoUDcvITekXd
Ma4KRsUCCHLOjnnPFE3WF3+sgoSxouBl3LEXJaHJXPhkdM1JIRjeRMmZiD817AP9
TXWcf8iSgaNwhLkrJMfJrNRYX7d8S1LCTqOdgquwOXMJWnqrrjDiJ5SiD1o4gTx/
Da/7nyK/afJa5sDgby7djd+bEISUY89LxKubSD8VBpK2sjsf1D7UlRwa7san6hc3
e47eK897dPQQQz5EHPivXUKHN5nl82RcP1fbtGtMGGZ4fwzST6/zlOcP8Hl/t/G5
mgQt63JeSRRvqwWY3VBoYuKKqunBVyAgHFjExDgGnjENm6lajq/w5czhPjSb49Dw
SVacl3wZU79tsnXlfH72zrbnaSh1PprRg2QnVWBKY4JTm4xz0cePTvTAK6vvqfhE
6DhNTgZGBvjZifAcQIpLkcw7SY7kjgqkJOMIrORB/UioycTNuFTTCrIKEsYrv3HT
7r8jkow53n33gB7AOtx1SB9RZv3CfU2bRZUrJqtOJ4rbvfNa2Auh1DlBeCuMwz5J
JeOsob8PDGme5H1Wh6n9ADiPv4SJ1z1UX/ex212zP7sX2yyLYsBPZBWUQtdFG3zG
BkQ7BH/MW/kVCideEtqRGi41W0YQfQj2EjUTSN3jsi5HIV/9dXJwd/4z9spS4j6q
DfjfjLNnXB/vLOeZNB2d+gpls99RzE5r81F753s8QMIrTh8dY4tkdU+Rq1AGR7yS
5g0KGtQaj+ZMokFwHYwS06BBAuOfdOuhsIcnJ5mQ2mPdtA+egBMHTOppdDe4zgDh
c65iKimu2N5VbYTGjAGzZXS8oGQ1gjE8FGAf2t936TsL+eB5vC7eU8vf8067pxU+
ImDvsD61Np2NsyxSQBUMO1xrvMOJwU8L3eB63kEFF2gKUCOYSAY6nFuIOE7vNihL
hbbwE/DkITfnc6rJNr7387acza582NOrfTMiqFxJ7X8fAXDrMpILdERviQyXzpQ2
tqyhaEkc/1wijdbfULLCJtFQjYfToublcW1i0IxdIdZwlam15mcJMaak01gMTT+c
lJyY56MqeQO5yCCeEWJYz+DGBoIJEWdj34ewQn+NQLouuYULky0iMVZDbyPB4cd/
5MPE7MSKqool1pzP2dTuXimbp6KEIC3WeTV9De+TP2lVxYsCdW5mKBm5+kYOAQOx
cPXrcUmVAM64cX0x4Xb1SVFxOa9KBDFlN8eyQDZi5yxVKXovchaT9Lmuca69Pa4U
8u1lxysRVs9RCaFRuOnixvuvPwqLvOI1+Is533AmKOeXGmCfJuGUwiEhHIzgsJkO
1iYlRC6gwQ5X9mRTAubGaoc19O62ngjibEo9KdFYYUmdxsMjf2UZvjVOFQ34ZY2s
rHpKc8PsenhwcJsmHlaoAVNi1v8dfB5Y+pqfUVLYZzfS+5+BTklKHgdoR66H28/S
vKjuYH2x70Cz66Xae5E8ANvP8iemOLWs/GVCbYGPmbbjLTuc1Ccwnn4bltnShxA/
Okg/jsnoEQt9VWfYwsUm1PRUqVH9JSMFCYmilDcUzHIEvp2PaET/DvFaqvR0Yax5
3312cPVV8QwJ0ZqiPL5CXFf+t9PA14Oty6wnyQaS5Z+DLBCCkUawwagZhsu7HU+a
5alkf7ZLYZ7I8d5HaGeeGWw51jLD3Ab+KjlvMAcdcJ4sCnFSZCUiyA28osTyjYpA
tuRcoqQqEnCrV/HheKq13sRxDMJnhfNlcRdQA0VedIUZhcAWr6cdO8Ux9XQsxK9x
0oc53WdER3tN4cd8AHJLoS/RQwSqdGlfC0KgwpYwTafaf68oSIAWS15nZL1gWLmf
6rn2RJDTYh+mPD6KpWsk8oV1pqdKMUWnOTKREKCDffo9DCWhdp8qMOODskd5gRZz
i+VKblVNbKF70ZGRm4OMKD3Tb2ZiViNJNjNHKo5gN+BH8s7D9nbHj4P1jp8guyx3
9/bIZpXFIpU1LdFloyoGTPr5zNh8J5SnJkX6MqniWAGDB2EDQfCK6M1FP0IFfdPc
ZpARtdtO2oPLAUH6AdcrEWacOrUm4gPb4gJ7ZSmHGqi+/96sWdTKKrmGHJxjrBPe
WydF6KZITAbIvKkB3d6iirpO75jkCf4NSZulqFxLJEgqSCUMsUuMEG6DcMsCH/t5
/kh9S68+RbUH5ILghBXl2MAjvRKiG2rXtXdNHkODfK7MDvlhgV5uqXnzCvQ2SxYP
yZuifEYSzQHd+KI/oEZx34KwNxzLy36Y90MZQFejuAQoOGf96eM19ng50hQn6tKo
faIAxekP/gqBQebRKl5ymddzSbdUs6cyED2hN+MskJhQrvF+6Z8hiQnGDhyct0Z4
Gm0AWLvtt4f7suszwFUo//EZv4FEJW4ZkXJ9j5oowI5ZyBc0wQiL0u6ZkdU5Zkru
w2S+EqD3aK1lixDSAzPZf+V0ps57pXjiL2m0+a2CQuCpQoh8N8Hex/bQAVEZUFkw
FRgDy5SZ/pBoUk1eCVHRlxGEllCcfKrGSV0sSWHIVxHN1gszw/3YvfJaonpH8ekx
O5L/K87PVfcW3yhqCkXFWJVfXL4sfcIOTN31YXSiDOopGXF0DedCv2IxKX+OSqBi
4y/sPS/lGaKGlj4EnvFlKKn+esey9uQ4tP0/rX06flUGvljWLEZkbHYH1o8ZOtzm
LswmrA4o5q4QRYKRDdhEMNs50y7/oOr50IRzS2ZTpA/SZfZGUmNkE65JfNHLOHBX
P9iWRxLyjwbvVmzQ8/cU3idXA7KgpWeVs6srWQj0K6wi/lkze/19RKTiutgIgbYE
KwCEw5y0Hsr6xFwgDJIsq6JSRA/pK5Jr7R7/KbmuLshV0dOzTW/pxdt9AL/zawTZ
fUuqATmNkSdUjkhW2k7AqOoKM5Mi6JYOKQmViNj0cakFDDGTJDxiqHoRpcZPeYMn
/qTl3jzexA3AjFIrvIL49RyU8RLAlIlcA/MzO6T1zkKWcIXl7GFlFwKBOJHC7QJW
dLNyACOIIjUJO4APYsh1fm7AgxuSENOkI8qebBg6XYTA1UUE1JBiJvUi6ioybDCB
Jx5QEy23TX/P7SqzrH9LvNUSq5FS7uuWDQk8ukBTr9NCH4+Yk12wUkbCZxyNIAdd
QW2abKeIVovtwkZcpK8OvCv11hjnH22NPcqSyNSGduGuiitd5Oo2WIMHxvnZpMl+
qJONP6golDCSbz+mcF8YoCsaUHdeXJ2IkZ0NzHKSA8/u3SYsXQNXBZvXc7/XyEiI
433I4D2iiFf/cL5Jee8xnCkW+PoRB9jc3jc/GktjO0lbK1HyNwsYViOG/qeRQKhI
p2k2U8wUCVL9YfKbZBEDI9dImJlA7UnwqTbzMAONGAXvCLu1HxY7ReBScAmLPNss
Jt1Jjbt+x0cMQNspn2tfe4hqtdSaEfiQvB9HsXZYHvLy5cZVY2IsETYTPqfsQup0
2kl34ThNg2/+M78KhgQ8aU9mRd8k6Z6TGWQ9Ci+8A7V4qnmaoq2eURkfPU5Zwssk
VPUI5RpzFRvvmpwoGhg5fdo8YKfgc8bniG3+SEg0217RDv8aYd25Mq9frSY2Sapw
yvMUGeqzZsYKLFXH3RxRT0WPD4mIx/fzsl+ixdQcB5Ni2LunTR1cJo6ryQNzlx/p
2kXj0AJFHQqU9G1hrEWxK0ykg1zvqImKf3fEDrD81Fnkft6bBCtKpvJzthRIdkwC
ytKaZRZaUuVNSjXEWOaKlBNWaxOFPqsD9m6B/CSAOCiv2oqZWo6jXRxrLFIcf6Qf
kzT/WXrO3kG2kiDap59l26QjrTfI5vNnblWtH+10iLdgI9wzTOCfz9qX668gDuQa
CutsrpWqi18jbfL7FeOUrHiJmxPF1+3ydzZVmOf930MLwPRJHr3+rVWBDX8w+P96
wvVWCVVabOeIco/WAPFRNXT5/8llqr3IqJWDUhOzwYsx6EO34a0Jd1lW9AzmZeQS
baPZgnIO0nm8FHRFLmuxZiwhcVvZLI1Fx+spanp8MtmFCddwHIkrEyQzm4tUVByJ
hDpMtgYUUwhFkqkD1dNbL1dKCMImgtb/vafUBcUrkRU4GoSbCgYj/vKuwEo13iXA
PDzJiLJssJJnt+ub65ZsGPC1SqQDfQLtbdE+yODldbBYrgWEgyru9pRN0pyHb0nM
1rRJwSRljdZX1ELFKdyQwb44J9li4BcEuMCho2SFGsESesE9w+6XRZIdZ4qQ+X6r
Y/2JxlRrIdwrKf09vuq71nhvUzXDYedfRn9Eex/bmJzetAdO+gNeGEZtnDzXOqx1
rKbYR1m0IfL8ZAp1J7OXxib2zNhVM0fq8D6hV5V/zeRwNPj2x9NNZPQT1Yd3gaB4
UKOz5rL4i7w6csFZvts337R048Rmr4w3qSmQozpTEV62dVFkKaDsOc9LywwCRREs
ggA3Po8dGHfyifYNka13ByAibZ5VOwUsAMg2TGtceMsaSR30hdy5rG2Q04JMbQ+R
uBgNooh/uA98PoA4ZAxIIz7I9jp+vCiicWidvZKS0feNXH8mcHUurw1l3Wf5A9hI
hf0tNQUEZxKNwiIt48S+Bt5OUzomdNtW1VXDoO375rDxphWm0UGxmiz9wloOnloL
FHk6F/DGV3C2YQ2RPXNGUODU4zR1W0G8WSDHyO1o1FHUiu1o0USmRrpnf5droqx2
7/DzTHHQFC2ClM11av2eiovnBpF5iwXECnJbUKEBsvROHErqYDU7ICenBaD6BA8I
bVdNXYR2cYTajQAJC5n2GqPi1gYtqcwOq96ecvqNug/qWdO1bN5LfFYqb54eASpG
Eu5Do7IJ0IO7lKiIFSacDUg1M1TpDkeKymSi/y7wrmwVczH4kowjH/xHk2eY9GdD
Bzn577ZgiKRESfZeMlBpSuSmrf1lfTKyg7ZgvKhZoJAxygaImC7p8abMmNZWYbv2
cXU0fp3wNRnALvjtIGc6Uux8aLxDfVuH15EKOtOZyhVi67VBvuX/5tI9Qb9L9TUf
duz9t0TSapIh8M32tY5FPbLpZDR4Iecpllv2xz59RhSavV451NXXCbK+jhIE4Ifm
USi5pI4odq+UfZvxLTRlAuCkHPoO9eOyCGNDiGCrtvKYux6csioH1gyRu+KLhoDo
PZ2A7TYnqNXTKYpXWaeUbR6VKT4QRd9I4ANPWpaBGNLJ4MaGssvgbBvmwL5HdmKX
r5TuE0ohnIDhPqDXUVNhlkISw+dJRFXrtVAT3zjdgcsXoNWgrjW6xWs+swp7JYiS
Ojl8kQMGh4EJZ1zqX+puJokClZn7WyEvc9A/Gp87xO1v88GAafY8mLAKLC3Pgpig
WYvMHOPjedKA25/LJ0jeYBavcjG/Gnc6HB+A56urPKtaqzBY0EUqfy2qGSauPOUN
T1Of1FFEUnzetLsiHF4D0aGqg1RkvdN8X0253VCRfS2NOcRnlZKvdks2Bw67Feyh
nv467GbIQVxIiKfnrNtFy7eXUDVreUjLueqpRxQLvS9pJBSvOBDZF6/pckR4Gnle
HbodrPLlhu5cNYMCPdBM2bnZGLqbfKWyXLTmoJ3k4UVUj9WTtf7jx/K5+nzWRVug
Z0+D8z3+AHlyGtN4L3JApv6AJ9mS+6GL/QLdt/fgEyWEWsvw3XNNAGf+s9ga/SmZ
VXFl0HcSx0IMROGTaRj3whVVSWoKDd9raBvlQ4W+Atd3WFgO6Z26hZdDpMgGV3wi
5E4M+yMeb8/yfpi5g4qbNqrfEgxnBykaVnY2AOpYHR9nyB3zggL/YBA371fbHMza
SI5CIkxhq1OAkfBb9THbxzyLOE5k03V8wEpbuMkhDtVH/fqXMCtMuauRCVRTsByB
5Rs//UIgJinCGTtcjV43CxqzM2BhJa/GYf4+Sit7AOuuprOHo4ZoyjtkqtuFLkqu
4vaFy9dp4qZXBU+XmnHnMUlmrJgs5rv7fWXagaCzxLPUraqoQ+TajrOjjpjC04A+
7Ewgn2O+y7+gJfLmu+aIqD3u4PoXWmdQBrvZk+zadi//P+6RwceHl/7ITWY/UWu1
i5/JgJDd3WOAhDldJkds3ywnu7oKotUpa7ZH1FpbetlLL5mr7aGpsNXqDzjgZrCY
vE77bEYzeJVLzrHU0kJZlbulCSP0Z1YXsN0Apt/mAG5WiraDWR7o1uMX0jorLgV9
OAQWTz/hHIrqiSj4J29sgtcVAL6aNmHInuRDXCpyW1BFevFpIbh4YGF3sqshawNF
K1G49zz4Pnl6qbHyvNoyTCHk4QBfV8BtMoCey9Xj0aAMpORG8fxxr3UeUAcut9nn
Uz4bvjatglnJ+epuzwS0n3EN3i5E+rIWOG/SAxsyxzL+1ro3AK3GtScyUt0P5VzY
zjxztjHHHAl9PVAXvtqFSMsOp03vVb8jrEFGe7va281kct5xHhfVcGsH6EFeYrc7
wvgEx56evP2cONhFwH2qcFoD7xujD/AzzQBfmr/XU9JbMT9Aux3LgjZkG7tkM5yX
v0OE0UZC8t5jsvruqNvHSu0nPDrAsURygOIEeiE7oE7m3tuQbOe/ykqmtAzDfgbD
7lR9ssycq6BjuchjbmM0+xQKCGuf1dkFDyCEInhmSMV991gXZkCYz0ylGKhnD/vF
dN7yAwGDc3zR/DWtoiUABFMrBlYeol16fqCo3LiSTzVzNg6NVDDxR5Y7On4RGOL/
uaK+71wGtqrOiXbgZZTfioqYXGWJWFr8zI/iPMBxo3/2Z5enIZD7WmShGjeNuUgC
1IKqKA/sSA0Vr1S9Fk2eZf5aF3hLBn+BOOVoQWBKV38bjzHXhazJ3CBQ+0l1FR+6
1pZ4F26AX75mR7QJvjKYMGkq9tWhyyHcpDg/lok/+b9bKNXvkKiHv9OBGES1ThLB
xdPdJBWLeNuGNBo+B0keETJNO+nG7F0AhTykiPS1kHHRI0KkgVgF0R7B6OBRCp+f
XiaWRZZ6yjJCw5bHqjwhNxKixqx6HFB/aiAmA4bNrmou3ZVkPxX+J2C8+RihIRg1
3n/aa0QlNlDNN8dH0XtI3y2SXwCkcw9tfNzWvvIfOqTjRusKjU4QMnodMwmFrSj9
zwM3x3PdtyoJpqhX7jVQ+cQ89i4TJIOgLHxfgagNC7FHo3WbLe5/Hf4w6q9ENp/P
D7HXHu881fRBUUUO3hp1AWe6XrgAo3Os+59WlpxPLsdWCjcxkYXLbhPSNrVRT17C
eAmwkMt/6HE26KambjhvsZneksAUdYZMk9Y6Vnpl7kXmpAm6AvNtgYfe0zc254bk
SeLbIi4JwoQCPm+JU0wtHPJP582ZmF/V6HZgczVBiHOCvDLOCNU6FpW87DadzsnN
dpTRACzr1t0IGEvcwEFrz8vWk6TqYhZUMac3/AVNECMR9R8MQJvXIgp7Bj8ttNbh
FWy1jbD+6aSYjazPj3qbGl4byIgBC46hevfUQhleLuseAw6gYySDT+2C+i5QXjZc
tOSOO6xR0jTtY4EFJpa/LgVHPG624YBrygrudyInmSAbtOR9rAa6LGOUzfrEwO+g
xzvSCyBPyBoX41+gBKeexIHvSyy5Rpxe2gOIbdXcDqj3zn+RVsBubb3UZqPVoy+V
BfAaYVE1zcwrqUaVy6arH8d5duzF6ZFiuSUXOYnRsPuTKNDQ2Is4F4Y9lILBovnb
DA1Vsklq6gaKjaPXiaKo1te15Zo7xbJiPIGVnAY9t3S3RrTqzLcKWkWAMGptSuJO
QT/+DVcTsugXipqbezHyNuF+SL2b3pBKqZBn3J7W8pLqarUEPao77EXt9+OKgqQQ
wK5P+EWMAj2V6U2sld5iHv+zY8bSxB7HMYet4qXlSIXj7y5du2D1yuIj4Ixlv/BT
XBcRVgOYCFUyoNTU50yyO16AN//P35Jasip6bkrh4FMynVlN0ejKDFMu5LiKUNOl
qVBll9jPolLueQDZGN4AMMxe9akB6b+0ddCc5UE9rN/wDGX3k+NXr7HsxcW4TRWL
S+CxiIzR7BaLzpHlDChSlxQjPMr1z0FSSPK+Qva8BvPy/XjJLFcid5kJdomUiNor
IyerZ2hRgNwUr+bmYoYmCHVzPsgQolQwr5fLj+pHkN+uqwWlN8hRhR2H+UOSl9BV
kgPBr43JIDjsJ1jSFYq51LSb1nQGB49yqlo5xBQf1+GLnI75rD5Luy65t12Ph/yp
Fvfoxo2p1DwMAV8psJN0OKlLK+v5dzdgOvv1GpSZOJTSum2AEW2N73kBoRZAEHIT
/DuPVbBiW24rm/OafMysLkh3lRHCxEMkR1MXOnj9AISG+wffiNOPy9LDmXRc/5Vv
MisfNsM6Ujl3meX1eimg0zMdzMMu+TGS+D+0Dv/0bUGHFa07VZhlaP0UMPdd30wC
HcFq0DJolqeeXuXKE0KeeWc7xqA9vjxB1YAVTEorl+65ayFq7UIWafPyzrrSjs7M
DCxGtWq97jKZBGsWF7wzkoZQaV1SGh9XKEQRhCJcUd5jjFcbyYM48ilEz9sI6/7j
+2SDSAxJ/mFTbppGB/a4iemFTtM5l1ZlZZr5VxZhSSDzR9G/VfKnndds3i4Mq7lg
uEaz2LxOyA1TTEAsItoKMetjrgTKSSZsHqEoP2BxXsZE+XLclIWXd5TFWNSSHkOI
qwZfH+sIhNFzhtd0lnMtab3vse7/O4rNX1TdkzjUUfXqFbg9PgTbaexNNXprrzQn
gnSpmgdUqmmO1eAQVsvcMqwqYMW2BezjlIemWoS6T7w=
`protect END_PROTECTED
