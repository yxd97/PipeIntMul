`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iwz0beQMdhG9WTIBzW8Ftgkw510HPSs45f05AvuHbuXP0oJ3WWKDS7gjZTncS7Fq
d6P9EsSpqJeHQEyrlxMY6gS6eRzUwQoWGfaC38Ml6BKMKWAiBNSbsZzK58AgUICj
EFdf3s2/LAVeZlofygGv6NHcOeQkVBOOC5+w9nbHt9IHUolA92oEF6xhot0ZFafY
gKJnlhhTI1qpvAsEycFPD8WQxnnPhpAc9KldAkBweZF1EMOKEQOWv2ilqiIHCUWn
NfonQK5ZWTRC0AQatZ5skEAGTgt8L1KsbkEPamfHzld4oU46xZhCQbHm2OM5YjER
jk5hFaaaTw7NOHzMZ002D3QbS6Out511kPgwg+nqZuSdcWOygmiA+lwvZkitBiL9
6ZULQIsgkZkHtHxQUqUmCLPiGlY7Oxx8TFsjy47UrVIfbgf7eOMqA9JsVOpVa9Eg
+6w1TrAgiqLomfOisABbiRBwJoYDcR75n0bRKezNaAtWFu6l4OC6IMRp/p2WK+HL
8a12k2YhJ7kjzpqkVwKNEH8J08bOw2jc4ocILxEZgFkORA1hqaK4U5ZfyzjA2Q4Y
FxGIgmGp7GYDsC+4hppRDEADoSvvSlJU9wmOW+01YE3tVN/TEXbIKrqCCSmm+LH5
cpEerscJ3oAZAEi8g86TPlSOVgHl1qG/ZQqMrJpMUM59ma6FGq+/RIpayKDPYKdB
UblwTcogMR42icuvokkwiOHDCrYJAK1+oSb+vkQcmej8NVLeTPEjmVdg/CTAMVqx
3zTiklJRQx9T57vTwlrIyDlHyBJxotSUbm6j/9Aka/kwR2xxoHvdjmpvlMSfsaKe
0xAiQrZBW0OGHuX01uhi+ppFtyH7rPpV/w2OoElpa4mnYDGlzT0+dkjvJlC78HE7
jGRNaQzxfFq+3NpbAu0wWwb+w+p6Xx6v3M5qNVrFax8y1AOvl8Urfrg/XsEHWI2f
tYw36Mrm1g+sXeHHY3jFuBnV3U66OeFOFZaij9SFfSAuZy9CLd9bu3gy0VF3BELB
MMTNPwtBdqfMn7zWdeQyu6M5NOOVMP0zordckIM28+nuEJUA5XJTM5pFR0Op0zL1
Rzs5fS+9uXfv0edta437DLminKVWfWXVhq6l6ayDkevLmDfbahrYaMea7XXjhkNN
0JgKi0T/PndSl5RYhFiwmPGxwnDVCdmambmql4NfMRY=
`protect END_PROTECTED
