`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fDTqaIuGcSt8lyTRqrtyFYL4iJ3efcw3aCokmnqQFfSBwj3KVoljiIxgnD8aQEB
KuBdKj0uVSp/pjohKvslkzGwcq+eOeiferLh4UJzOwyGE1ubAElXTpf2+j5ia5rb
1/fsWOj7saN7DU2ZimKBj6zQOgJmtzquli+CT11I5aT2b28hntXaKPGO/AjA8LTB
Ru/AxO0X7/NpeOq3uvrLxW7wNnbv7UVLxe8hecdfHtmquT3iTMA2GB9hSgw5XUXa
xJVyv0svcNE4fhFOG2YHuEFbRiYvjzCxPdNIHXyuO3HUlolrWl4MVbqY0tnGOwx+
kfiIbcIm8JlrtTMEIsWGiQ==
`protect END_PROTECTED
