`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zzghvXw5/AW6hxQaklw/24+pmP+gZjyTfP+YkfmEWRxHYczPxL/igWJYRokMDrn
Ym/9kZq/PMpSVULUaDUcHDmPU8WAz1OHjNtpkj56oggZmxikEUVrxSWwO/7eqavp
U5Q9zf99IkPVkOSPoyX7PTz9Mt1r8NFF+ASDp27gQRUQ0nmsyWxHyFCutUW3nD3C
YsISfjAh/i36nOy+WTY6jZ7V/MEzkBOkNXcAJOzqlganuHbhUFqAx6hK47PxeHx8
Hv0k69V9sdahZn2dOIUXtUIXzuuQBvctzykNzyQ6n7ST4hYrlWRvIYDtXOSXN2GH
/1AUfHwrhRuZvwyClv0pQUGXmXvalCXZQZRPzTnhSnuFCsDAdJz2whQ4oJ+mjFts
77zxdiJqSd1sD3Z7p5Py9juS+MXB6Uz6sL8KCqfl6Ws=
`protect END_PROTECTED
