`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SRy4GzIydvCU9bwTlGHnn26nEMvvHFdw47LouhFEMCC2lHSjlyqnmY7PoVEhne4l
cP+mRc6qCbPqbeV0HrIuALJkDWuqYcHT4osO6WnF8YVRR0OeBWg4TFGpWxIc4FF+
cUSXY8BnFCNQ4bghdANJXDP9yuBKbciFcOFdcRte7XTpPuNlvFy8JtEd7dZE0n60
4adHGVFCMJPDKW+Ulqsh0iUCdCA2wah0Z5+vgRnZM9FyNeXY+cOofR94rjKQbmQm
VShSVtAhQOPbzDA8fJRrGxHUHABc6PzKW4Av8Zc+MgAVAGAoGGrSlnVIjWu/IHF+
flMIUm87+i7jb77nCGo3CeI2+tgS92oz626NFTWJtG3aLaauK1yRbXYXQZco1FAk
Yy78WZg9YW0UlKq1E3PziEIG1l97Tu9clbX81pJrZ3kz0PLfYqXw0CISdUfZin7q
GGFCs8G8iSsVavEDf2Tumr1+64sTZ8QITAC+8BHLksFUEDwNHLKoKd8OTd71XeKR
M+KK2F34yf5Qp/dO8Lk7fIUaCQcfm4SULsCwgzfmuL8YdBgXYqEAQg37RTBSf1z8
TAn7+1w0SE/LBsbgUbEOkXVMfUcv8Evwk2etH/gxUw4jvQyzfWfJWtHB7Gk96YRm
xSY1sY4AK4pP2WbL6uLlOQ==
`protect END_PROTECTED
