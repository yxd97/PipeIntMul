`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xX+oeFdEdwR7YKGlK3vNyJdhAl61Us5aB5uVlDO2q6m0bKXVJPJSapbU6yhOVoyk
y10kudmtUhX+TT+Ib798FrhDYZGAwAGfzhI4OT/OQuUFLczh5bAn2wHug6Cz2u8N
zNDVQewKfSwkQw3WsDRtKfIhPRue/eWumnRqgenV+YJHrowNKF8SmhcsU9YZ4I0P
dB8VL0uXe74GU5If714cEAMP1fJ5T/uMQIgxT2M4d8l7keV0AxNpPpxiMt6e9tXP
omHrReMBIg8Tg6Rn47mEzKD1OmyDt66Y4tDBefl0JskddK1UjgAil+938oCq8ve6
BlCLiYYC2JD9RDLmHcjDC2NOZy+muOkwiW5uEiqVc5Y30hCJ4hZujLelnazK+Wbb
6q3TIsuusSSsNdr4veCn3Qe2KnnwY7YpJvxRR23PUEU/VYXA1wIrLOK/eeeRLaNR
F1boHvvPk4NNMpkLaaMMLEW/ae+JXEMw9uTpFDvsBTqyfgrqfleGyVQY9cD9Tja/
ubOoPV3/Em7CboGF/n0qnPG3t01DWipF62plWjmvKnGmlxthkGYuMAYN9ILgkCCW
EwyM5Ao+QxixVoRVnyy/a/TNh1iBt7Gmgto64Pofwzbz99v5ZHRquhbp1BA59A2Z
lA+K/LBJvsQu3jzCdXFCX2gEHn+ti7nluitypALlsGdzBKTMuVqWOW0Vqhx/vdOV
CCtmwrJZvcYm9C4CHjfToj+UKCAZ3PkQi93f0cBhYOJ715/dP0tmbcN05VrVvOvW
kD/jp7ryR64/mn10bJl6W4FkurJMtYpbAs3g4EVmhlBgqBbx/4YV4X7WvF5VcMMc
ufJoix5ilYx/rOfAoaHOH0EoYaMV0nIxmYrIiExL1sFE/B/8pAfcdnBrmspqNx5P
4gR5hrt5Fi0Nev7e4LgSiWe8embRDyvjqcR7rJFqawAd+P4HMYYxhRlImX9f3ayE
sZ1oAzDQjKabBD0J6dwrHC5km6tGNN/l3dwuiHhSfW6tv7E+pWKcFV6iSPyGBr0M
X/HBQvhfdApaGdspjRd+DVKUDwRfYVaBb+bU3At25qOGINkeuWT4EJ64LA634ip0
qoEB+N5hMArieo137Uv3cWtmsc62vCR3CFuxfyGVL/DUxB6qDAUOJpM3AxEiM0ak
/8HdkQP0KOzbq00t44KnkEQxZBsej4mduL2JsLnm427xM/rviFLOFW7lxk4/5HH+
XOLc8XHeVYWWoVWcMHK8sNY5BzNMe4DyafrI3pHSXI/B1/qGwYf2lglStyY1gHhN
HSMVyU5mmBPCD+Lerbex/yniU2s010pNRsQDt5V211H6uBZSgkyd8eNgduEtSC3A
Lbuv8fEVxbmEJB00mF3Gle3UEy98e8AWemVxa8mGi2Jgq4BjIc3wZ6UJHOlwIQ94
g6aS7dm9Zwl9VxWZVV3J1Xh8Z1lbPkEYF05Lk/syg/YsNDsbnvOpkQf7xH+PiUZA
AXpqC/szdAPOX7NX6lEaA7hDGcX9vzdcWfjpjI+b1qE=
`protect END_PROTECTED
