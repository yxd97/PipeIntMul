`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SSOd2z/hH16Sh03rlj1XnzUI2+xnaXOprFLg+k4ouDmgtyKtOTwdnxXNq8/MBi8C
vqFr5Z7NTEId7g4zpjGdV5zHKUsxgisb+xDz+sRTS2aDNt9ZEsBXm78E21OqUaSx
+6zbt9gP/b6l5Pi4SQYFpMMESTTllzNFo8yZEjRVioUH4eXWKmnCtSxPkPqr9gJB
hQXFcuJo9HNE5Pq3JyffxjA2VD5Yd0JxHAiI3BbYrW+Nz0nC9u3tDrMwH1QBI4Rq
9TbtoU7BiUkwPnCZvkiWGhEhT+k7fEHLFSIGBfVLV3yY37Gm97QrHhT0aO5aFyJu
wRtPBnXp8UAYIU47qRgKhO5mFLMa4FYzbTNE90bNnBSxfuj8aRa+rijtHJH63f0+
CW1gAdKKERTpC+MBGsfl3fnkjBhc17kp8XFR+CsMJNHwY/Db48KNOjuXj8Zc2PYF
3WINHRsKuEdot8TR4Jii4pZwfmuRn84VQLsxmer2wr0WOhZ2nmLD6gBVcQU7f1qM
DA15HrkIPWybo636IQSqbIYX8n4NGm8arJz1aGTjrUGZ6Sg/5LHgOdFZ0iZzoWhr
sIQtTMiPk5xauDnyTGySB6+QTnWLEmdlZCu4KpZPJ1loWuDN54DIhUa1XQlwyYmG
Oabxdv2RaI4Hs90eTLTzMqwdADI9Efdyddu0k1tN/sl87uHTQjx2NDgu++UaeRMt
mrGQbyOSQ7beS/8RxD2wymDoiWkca4iDLnWoZz/dwXJ3iPIMlXX3q/J8DpmEqclq
5a+TIXSSJJYUNYzkHPDwHd57nXfF1SdlVEOb3BOiOn3ukmhVFxJxO3eVUj22jLyt
t+8PJiAYzYASiPeOVBE4GCEZ9E05Jrgz8kMwP6smaMdLPnaVEQ/YR1kxtRD7pP+V
Gv5k/DHfkBZps+Qk8yxHsuR7kAIHlMsHvsf8R5Uut7ZCzeUwyX78GEX/VmFSWIty
NsYHuyPUcq1tLdiMdLzxWMJsPP46esffkrjF8ZOfLHbjYLKiG7CYzv6q+D8RMt/d
CQU1ji8T9jmXqtU2v0rTPA==
`protect END_PROTECTED
