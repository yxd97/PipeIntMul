`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJPc8D7uXALeQAHguRbWhjKmnJghd9NFBflIPBD4FttcPt5+rWRQEbi2tkZlxMvs
vpm/sqvv9kGza4RkEEpEcnCHHchiUpwO+SlehCqbVpjtziGfTmu9bTy6FOt66qmu
Uaafrlx9t+GtmnmAQ5d50jXmR5UpKhP4f4O9R2c72xVc3HXcAmAe+opUNOOkSZj/
D4Nh0oPHIhJPIm79SnWB3J0JY/F5V6nPWmuk/w9OdKhYN4pGL6VtMgJRjacXyZ/s
dyk9IQRhEZS738L126EPnk/WtY3zMfDQ7EapvVUnC9KmxIFoVEI7GjOGMQ/BCZwG
s+IvUdTMeLjNSutbQQ8J8A==
`protect END_PROTECTED
