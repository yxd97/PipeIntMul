`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xq/ehO1g9k4NQHk3G5jOtEjia79S/lh8gZOHRc6rcs5xec/1DocN1xPD9D21fOeZ
dQxBwZrz0553s8iWjboFI7aP2dbwnTta5zpfEoQ2va7UqQoBeFYn7+I97CpCPoTn
BiQPL2ggGz5+Z2ZsSuUZqet3q4NO8RGKO+e4VlIoK3XMY4DY7H10LAADLbWUB5zy
ZozrlRHsg4R3eXo3Y7KfJ0Iz+gLMrKtlHgiZJ3ZypzAXgVUkjRUGXI4pk1eRPtWw
FPZaiVNA0w32p0W1plP8yhg8/u8aNvg2SILBK5QfBAqW5SdXWOpAWwwLjqx9Jlum
p1cgA7CdY/JkFIzMimDifgX0OiNF5KIdN53vkqjsj6AyVEqICcWlfWkZy9YmBDDv
hiZtbww6UTSprRNDggtp4+skYIxvCuT4Gi9R9wOZcYhBI1DcBL/4IfUx6/9o8Jit
xhJalonZ/SZC7+9FLQF0fDk24Pe4CfSm/auiaBmQhJyvPnjj1sGeKGU0nEEaE7Ix
`protect END_PROTECTED
