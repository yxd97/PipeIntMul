`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwhK1L1xvcGV0qLv5C4pL+CWQ5AEThn318t0DdU60JFMEZJ/53FDYzj8HoH6xdir
FqQjy5e1kQvgpqxKMiH6BNTbc6wjJMB8ViAbikJamHlF04C78AbovQQPnI1vLOlj
m+KSLrQNF6rPjyLfqsGfR1W6qsOG0u5jp5ssb3rE+qRB+1TsCk59Dj1l0z+LjWjt
obzpYScTHYN/ckpg8pYObvsEL8ZlfAbt9SGLuhCKmu1PoUo9DP5w+cTTgzTxqwad
ABIFNqOeVRiaDS8qoyqp5igrrMtDjOlVsxGm2dp6YitRUIzgujp9NVoDjbFgltGg
zVRlv6TsuETa2I0q6KRhR0H22vtMcdyiXHwp4YNSGhDieRpvAgPq2Otmyoy9firT
Ed0DJ0tREzazfPLP1413ii96WZh5MF0f1Fv15L2Q8OUUkZL+1p/qJRXrYN5JdWl9
QPOwEVmC68XeI7aCZnKJOVdlup5lyV1r/5KSukXdRRGH9OJSVzMfDCscmVrcDgOG
MX2b4NxrEF6jcSYaKtCtNm54aHwyJ2VeOaxGXvmaULqgUUzjuTq8N+8xqnW2Q1qj
Rcyo2jfesybTzsiRtNQHCSBG2vPdMQrm5cAFaprrWvI=
`protect END_PROTECTED
