`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYU/oZ2V+Pm8jPks3G/lVcfUFXkrG08K0kDEa7c2j8aihGlPDhIUUB65RpMQVq+V
2aIxW95TpPJDpqXyOWiQCM0dMRsqcN7RFvnbl4HFxzivShdb+KBBN1HzVt07Qn6V
BM3DkvE7RsbH5oxZ5Wyas5TaAqdrwyfJy5ghoSHvnPmioX8PYxaneKxzg8T52xVP
FhrFL2ZuPi8D4qeHrwC+VyMsjA//qtsO/42uw4CeDtUs/NJM4ZEgA0Uj18xqYgR8
Sbg9WZVbFlw24LXnl06yk2hLOu9S8X8eYQ91CIStO0q9q5nVl5K2Sn5SMH+bcDRW
jp7u9v1Hv/R/q4IHOjWdqsYCv174IP+7MpS3Xx5hKbdkmTgUB7qc3JQ8dhmkuZKV
Z83dooPH32QegLNZJTgvPTrMQrDTcMsEZmFRDQjqz8Qx+Pd/24QVT9KZT2O4uxys
CORNRqPe5OPXVhy1/Tf7D3C7Zh5sjNdQNsXICoIv0gpt09EPpV3dXCnO7ekFfkDb
`protect END_PROTECTED
