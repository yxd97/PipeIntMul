`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkk8duJ6Yo6/a1s6hObHktwekwpG2AzZlWs77KnDzYcWMYJVmFBMi7jgxJ0hm+Sc
oed9g3GaOQIa13w8X0YHi31Im4QIUJRtDr/7gN4WvN1rLSldArEDE0Vs6rjY0ykD
dkHIAdkhO+2n7AW2gpjnNSSLpoqbj1as5uRw2urd5q9VD1Vwaz1uOU3G6jBdZZ9Z
+mfA0fdoIIQdCVQ2Hv4xi3UqjGBGFOtVPpl010KQrWp9xHJN/mqwGnslNp/Lwjpn
co8UMJVAvhB4gYv32Uei2BTa7HGRgEZXt7Z4pet/dsJHMZFD4bsQwbJ2kjNg/kJ6
ESGvnjgrVgVOsHivAOYBg0csZTM7Z6Nbtjx6e324gijF7rbueVuqIbQ8kEw3ipdN
vYlkhxCC6e2t6F3AUF7JiCWfjm/pY7LUmvSPOCUQpl7N5tBp/utv36XSzc71VCHR
4YbKRjDhaUKzX1iccQa25A==
`protect END_PROTECTED
