`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zywc2IWtL3z1R+Ld7FHH1tNrB/gn9cr4CyeoDHnboP1dUahsQK7Wy9ll3BGLP/Ed
hdFB5wXk0RseP2yZaCsVgg5B92acbTvgrWMAShEKfNC2X6O90m4nV06bZiyXziMl
O5crszDCTBMPrTTeDorL8bXL1MD/2Riz/ugzD4VVDZFfr4Xr1h8HJjj1TsgPw1u7
Xlv74CCufHHx0P3Vg3fdDv/CFFMdG6kfqhQatjFBd9BwxfGmPpT6xYRVvHS3Lrch
mA+CYhVl0voPQyZz7jiUNalWRR7UJ+yJi9J3Wx3oY8rhZR1S3lhH3cP3Uq7oHpxX
lT1D6DZeAWflJmmLE7EW0HITDY55lJC+u1FdMBeVzz/Ffp2mOLofwT0rFLMI6lm4
MPs8wdk1iLYThGCX9szlUnZPqJ0sNw6i3VTWBZpqJMFfViSDJvQk4Q0rMZYOrrrf
e8vpov8YjW8GUVupjr9Kxn0vDQANEMQQ1J6SnEMDalrAf5FonAgTHX+nFAjI1ndj
0pAiTdJovbu0GyK5++kc2PKH/QmFZZVtFqlypF8JBZv+hLXvS9zhf7C3WRYEdPta
5eOoN9tY+4IxsOeIf9JX6Ie3vvop6Ni9A5h3jdbC7wnIfDYA0IiHhQ4IkkBpq/rk
`protect END_PROTECTED
