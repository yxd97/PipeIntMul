`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uu/uBLDqjmqawllAU0SZn190NWCeghH3AEFGbbCtm9po8C/m3eB2qH+6wn0ZHRaY
a11eFnqAvTEp57UnN0vqW2kzhyLVFD1JyNpWU64jHDp9RspgpzjA+KfyGSbmzxk8
hjLM6j2yGtl4UCDRJObJA78IyGopoOFZdeNtXSx1XgrtPsnFaio9VQWE+wTYZ/Lx
AQvsdGCUDlNn43N4IyT2/H7V90wnN99qGcciMwjz6AOrmuasjiwPT8UhE3BZyzPs
3qSQdJwIGfC91jlCaEUpZ3YV0UOR0zp+r91IfctTR3V0WQNZeSiczWeV6vDi0Hyl
I1nlBq9JCDESliaPvuVhJZW3ZZE4HMGl7M9u5d5DxXRv8jOew89sqFX0TACu3v5M
3SbYMoRNQacj1+JAewKozvop8pVYe5gF6z7DDraegyvKOehWDnBA5wjyPAOpF0iJ
AqrAav21SHXsBNQtlfmrtqUDv6XZ0GBx2jTeL39kbGrFNEq4zavz2096XRzwSJ3a
9JrBPMY6PKRU2LqtAWP3MnFSAEfLjd/cEOy4Qk8g/jaWyM1MbFbWt/qfEnWvzivN
`protect END_PROTECTED
