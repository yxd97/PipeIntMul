`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B36wEXERPlpmOU98yGmg+p1SJ3baIOCGWRt6ofjh1k2l+1jQtv9px49LjI0V4iDA
4XQJNBqRWdtD6WDtEGE77BAlyIqa6qyT09vTSLf6CQkb234anBcbaqDx5KXKWy3v
xjezDJZLpUv3l8BvJAT8NQ==
`protect END_PROTECTED
