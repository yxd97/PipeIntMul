`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ip3Ii5xogtW3LfsS8eljBnN+3bmMr82nWFrmJJPdS4V42LyrCZiPO9gznDlRQ/g
WgPCNeSZBNM5BDEwszxdIp1eGgaMxVuxA4OE8QTzV90dj6XuLC3SVIzRGRcfJtep
doR0seGcJdYJcuVx7G/Xl/HbW5Wi/jdXjmO2Hb2Y9pu2oo3MbUCWFS26Py62yMs0
vMUrvI5um/6ZX+cy05shGy+EwxdlrwDsetP39KKBjH0Tb5CeHRDzfIspXgi2k8RT
sVo/SoOsxooduWdPoThe1xJYrUmMW+Z1JwyV3FmPxAkukPOr8NjCRoB2aXGAQGcN
jwzun5PbOMBn/ksBlVN53rjnF5+r8F4/bWcaHih9qsKw32+eqrNtM1gMZyd4ZO4r
gaMiRRWC2edY2LBYsw8L/Tz0enH0ayXBcW/AnHSu2G9T8CdCH0M1K3ghWlYr/aR5
PKfUp7N/asPru4C6z2YBhxrmIuXcCWBkp5+xg6P7cyeG45iIc5dlg+n2Daconzb8
6SIjAn7ix3EVTa5MkDUGFY2jjKLn0B0EknZGx8pIVE8=
`protect END_PROTECTED
