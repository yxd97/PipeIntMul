`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D3bHDhJn7xRSPvIGhxKxMXq5po+/Gtmyls7ay1yp8zoaTkaIV8JsOlgEuAGWm32n
dqom7pmv5TK7hbwz4ZTifNhMFZV/RZdPZ4zEQzK7ZlJIoDPxg7m9wl9lOCkuYbRM
SCq3B7Pyonb/leVWKKtIaDkTaWZRmaSJNe4K/kgR3q41Q/1IDAA1mKo1/0gaphIc
2ZQttfhTTe2GMjOTWQu/QiRt6sXeWs2MGiH4ABQyo/12oTnNZpZ/HyjHwRliRenb
myiBdiavCHFoOdSB+rU9QVFjuw2xxk/pfnvsQQiY6qhmbuE3nsqNOq79QFMesLyp
F+H07hymfVu1N6avMV9gnMA71GE67biNJLmPr4ltf78ia/JsLChWlFn9xSC8ChUk
FHZTDuvUQKf8eE/YA1qCgoYcpjsfjqWvxog5edxc2VUWSIIQnRm68BrDbaFO5sPx
t09MvZJG9MJw4bf9aZdCknuWZnmldCpmxzpYUtEUeDn2CW4Lalo1r+hQHrop5i3+
HAAqRUWrQVQgh4uV/PRLV8rDHc+ntLnFZcRPgOtSA7o23BWjMeH/BUP5Q3H8p8vj
hEj8CsmPF45gurzbgmAgQwgtIYTciO6bNHWU/KL42KZobBhvrC2nTKLf7/WjWKP8
aOPSEUl5CcAfZC3/KshiAg==
`protect END_PROTECTED
