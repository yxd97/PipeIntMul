`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTtljQm3PcgxNgqM+eYjMIyE97XgSKKvK5N58Ehb/h9+awk0mXqIaDxE0KmmN4G3
OHX7VTLbb4vWNgSriJnagaAAKxM5hoxfKJ4JvCxKNhqv5gCNqb3GsAjaKcDwJ7d2
6ABy1KDR+Ko+xPN42QI5ZpPSLFrbBhyKiE9+HhFYUEefbK/OLAhArM0xHMM3bzf2
oNzidkxvYNsPDvB0XS/ZKZpGXdNnI39uaWxH4SwkHbEX2Tne7ZpGA0qRYBTBskZ1
TXcXI2qyBaaYVWP91oTHIbQ+GL7J96Ual4iOvVibshbUDOJLpy4k4lEXDFU9f0B2
`protect END_PROTECTED
