`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pfrx+4ssfkjL40mw0AoVPE2lEaJSAwebnIWT4l1OAoauySjVohX82aYqi2RiTnWQ
fetvZpNCU7PWNwftNQTPWlaoHk23XzX9Ih+cQCNe0I7Y+viNzcvjlP6dKxqD3Lat
qhVHMslJRdot6QECd3Sw7hexRYBCRNkBqVXP1I1CPKFlblcb19uj4E2PEM87+W20
0bVe9DpfMqHGUbKr1fqaiAApbgZkJZULkvpbnglKfCnWDSCrr+dEr1pxbXbhVEOJ
TH1sEzremAryOm6gHU+ZA3T47xhNtd7yYxSSBOVnN/kLUEene0bjeigScN1SQWix
9Zb4ciTi6T2iofvO9bVRf0YY+2PGz3mpe8MrhytVOWL4BYvTrlKAzfOpn8+ECKCz
Gl4i0tKa9xcU8BbxHAnRYJKpqJWdqqrtKYTissMzj+miubevnLcXYN3+QK9ncLbc
IrWmSGzsbczz6nt/QEJFJeyWnQ7UmUGf4h1ngq+yis9xHiCeT511k8qUz9fO58X/
J25Vdv2RtcB5KAjEL9eyN+jhpE4HXdwAnF5TTwn3idh1e5wKTSTf2ZKnK1lirUQy
UjHQZo5PfsXRnF2xixh90GMzrpuJUgTU2O7idIH8/3EudhMkYBLHS7GClqWP68zk
CCT5XCeLgvidzwLCiWWvul7+dRBTLyiXHGVllYHqqBFfyniClSWjVrY12kbypd8M
uwjpcEZ/ZMmSWWhoRd/mBa/nfrn7Tnh3VVNLqQQ9BU5wXpDtkcYkkLJNnUicklrB
B2V4onkg3t5ApHf5o3/OpB9nMCCwwHOKy6R4oAEZwyQrmj+JcLSDijJvTQ0LFGKa
HIAqBmV9fR7RGSUgR7/VYR36B1aRAb865vWXlud3Iv5IsmNAUi3AgqEnSrlWJjmS
YApCg2oKLLOLNq2F6YT3Bi+XcdvD8FYgFfHHa06wydqn1z1LqRc3MIL/Mp8qPzW7
B9PDRdFi525vlCF3LKDO4J9O5Lu6WQAyMQbQcZbgXFSpOhkPXU2rCOjjZTdVMP2G
nJeTyTFt5WFGH6Q1ACm90rZ3Ab1WvXMan/TRvSkyEz97j43aCMTQ/HGQYHWJ30K7
gI9S8/z5RCV4Yt/XOhISbuwAxdtmmytxho98SwK092/NnK3QDa3cxpjdoiqTtIch
N1Q+A6iVd0Q/FbuVslubVP6LDXOi4Fd4I3+QUF3chObRPee5BoaZiSK38lkVurrO
9z43XyQkvPuMFEKsWkxkBXYC5KG/XyjL4IjxXCfil4G4nVBzq6lOd2GZsEXiO4c2
PKfiqzMfdmGJ+sBOWPk686I7HW6M8D4IXm3RZyGRtwXedLsSf1QF3UNcmh/rcM/l
jAdTKJjvSjwPW/Ke9BZU8A7Vb+2pQlyc8GxpjlW7oxckaWFHbKDKQJwlir+wuivf
qETwN7lKR49wxRsgr33qdvDaRSzaYW+hIYR9W+NYT5Wz6nhsmqjA4c0q6ZNVEm1j
YX36AFJ4rNujxwugAQ500MtUn1m3Ud1QRK91L+4Hhjc91Hf0JpoJSoxWBCywWyEj
wqhI+VP18PeHt3JDxHJ6WZciNcyNDjcufVBiukNQ9LjWNDWe6wTSfJt6NHtZCxTP
Pyyke5WTdakTWceB3AgMuvelonMBO5hZGtnFXR7lX+8eGb5NPrco0bqw+8jsMfO4
+H2cyj76bpQNkcNbFdoUXjNGZFz9taaHAyJJ0mz6ED9GVmzv7x1OJclraTZbMqlq
dWgG1LxNp9s/nqnKYUsgskNXkJDDWTlGex0AI5vuODYmi1PGTCE5HnMQL2KpU9Ow
pYZmTSTamavT76/hMo9pWWtstKmKlbEY/ODglYw3ifUXKbRQpU/5HPpXCblsRjrl
CExYYdn1A80af+H/8UcMLPtT0d8o3VnIMVXV2HLfcHSDBryyvE849OQbr9lo49V5
E6MYiwXk0OBFSrf8DmBsQsG2Paq7+GwK2HckYpHy+oHKaXE2G1oksk3Y1BmDuyEk
5zGQcUmaO9XfsG+a6EIvHn6xrXuBZaKVcV5OYcLv3iGoQwd2dpcdQFvvGWAv91is
xR+BDDk+whlD1KwHBcR+cUXpvCjTcuWUOizS5fQP7G99xf0xtyVlcoNiK2quTOnZ
PBz+BRLrdhQ2PlpkxKNyLyGN1KeA4+4wCJPtI7CYlJpWj4JcKUU6X1yOHJEGEJsp
lNLMf3djPlGEAfLBlN9pyls9oJaeDf99GycgHyGghiWIfpOk7G9pDRm2+L3hxJeD
gqK/jKAKN0M9eR6jr8ormaTLGTKRhjLh2zxXs3jH1HKZA6ClK/+HpPqq9caPIKS4
gTxyXzFqWLfQ3MwBEFdAxbkh75bD8edz3C2+Jlq63g4ckcQseb7PMLmJ9nWI1my+
3nckMCKugKSN9oRw08YnkGQ9meNEAoX77SRh2m+So51MuYp0jBzW2QYKj4gx1kHj
Qcq3VjVeWXPr+NLP5YhXCgq2yOZf6s7FnG7gkV8QQPt3ij0nfk3oY9meB4VgmRxo
7UVoOxPPZTCl+EHSzo/akhAyqWzXLkC1ikl1p+wipx03+QocC7tXUkq3RGDGXQ1X
yUrwh3dG9F/wVNRcxcDD91Z09a4JLvs1N9mz7qFgo3jgu4yIHNCyz8HbMjXf2Ir+
lPAJbfA4AgSy5/78X1McAEj7Y0m8UMAWXRGox4XyA8IGV73pWQZdoHhuxsQmKIGP
eddwThyHxEMLnp+McYU1RQubRqO7NXLFNiE4fFoREulvgy/JJJwaihOqdDzTXJn0
YM7cvTz0VxrVY3Sou3IyWUYpXjyNkOipinIknI79iI2fRnk47Ut5HpUFM0MH7xac
ZGzXOcXz1Icb2YfTiB6+ECIHV4KdCqiWgONgtU1O/KemtuJoaNSp5QP/QXjRkUZW
rneTf5Nxwtn5MXkfOl4BqstndOiPOWRIqgNynnQRluPwKVeClMhkjvSNClGrOyFD
n805VaSCFbxGDgibvR9nbojvYJu7L8U1ccR0EGWNafkCtC+Qhl7hsS6pdrYUuoZR
UV2xWVxMLCVRSOuxcyVg3RtDLAySUjNU6odXVhiEHhKRVE3V4lq62HRGoCMWSvAQ
ocBpG3+GG3oYa0qi0ANe89fgPgob1PJRlZN0Y8KiFECVyWShbj8gax42Vt15HQ0T
Qy+3A1SOnCcj9VgIB5VFmoLiGM8VymV2wvyNZ8zhCII47m6Xa3VfcecJ8dlwhfNk
qXONJmvWiS4TFwu4siizlt6S4ziIXVKp9CJ+kXttlHzg1L8IOVvVlTszlywa+wfE
j5e8Nt33xAspH05JRb0sNPHlaVKpUvOVLv4+ikxidaQDGS98FGOy6NnfbfkB1q5/
8NDS8BknTkbCx/zAClA4cakKChvO5QQLuFktqxzbBrc+CtSDD1WjLwcI+Nzr9Li3
24rSIrvsnWi+lljiOos9kW+9S9F+aj9nLhKG5kiA17+rRH8x7RJ6yn/Z9hTy7Msc
ETtnD2TCpY1A2lKDDEe7s9dlUHwjpyIR0OM1jqbq6dPFaXrC3qzap4PP3GxFG+7K
ep5DpUvOggNDqaWW2HjuiCpIdQ22c5HHZFKSuVXwqW9l9jS3A8fs0pc7mVyKXISc
AClOtUYsZphShs+5RzMTNyrT7PBSqQ2mlt5VSRyhtNUKPtA4KG0k+h/S1w2WHP1Y
axVVVJ1PVUqvqUpQDb5amkI+87AizzFYmN2GU983d/9A9La2ka/e7ZqIy5lt8hjM
8Wtf7rv+WFcYbMd2Z1j9cXQHw5FvyturW1Aprcrv1s4bE64vPfNi1AVUfdddWOKw
zgVocsiH4Q/IMkyhPYKGT1i5DShfihq/rOwJ9Ktp4dIQrV6suzZlAEdaxfbIxkT4
k84nLWJ3+bUoVE9EdJxTDObGjASgCqTxcVw/YGtQ9PT6ZmnhbTCvyyLCMwsYMdCJ
GDv/30T2iSgY8UwhCELueb5T49rlNBER1N4xxErPt96IqFDMdA6qp1flDbFKbY1+
wqFDihoXy2ewujNxbrTcOM6JDzZGbODOeT2kM3OCujOwnCLpdlu2EDX2koy/jxDL
wVf2gUMx6eWXjScksCilErJn0tO0EhXdUagyVFZf1AvVJ4oGAhaaghl+5XZDom53
jEvm17M4Tt52NEABeVGKSVXK/rl5YRrT8SD7cABo4g7FC/U3B2jBkJRkriZWCXdi
/aY5V8UVGuJ0D8U95gu7puOin1l5DCcYdVpACDwJrEVUGHzldlWEXDFQx1IX0EGr
IRDVAbIYvDcx8+bT9v5zu00I1X31TKJnILobuJIGnXeTbcze7WH+IecVWNAPa2/i
I3H5Hf4sI8ClYAtgwpU78Gz/gWGXN5NaQrVMYgoVZiD6LCWY1L9KOeaq9Zss8dCf
jV5rsUGuEXk0NLV8FqPj8omqq1Ewq52PfWuBx+N28lbdRC9sSBD+9ZvBinpjnGqO
I5PFUqE2LdhAtHymyLR0nHa7l2rduFdc4LxE/rZIGwFar1tUNpIO6DqUToLzzts7
QkbKZArL7My5J7Ao+nQHq+b58K1zq8fVQKa3lVzfWvtWGpnTT5FgGq/k/D9t1uAj
wq6/0NXFbCmEPkDQ5zfPXxlJvl4JV1VGKBXWT1IlVJsylmEoO/9XfaG79Xvvp2XS
usXU1Z/zuxo+yKPaEIeaLdqEUurrkdVPJi5bxVBx72Jng3lh6CfvrymOOim+Mg0B
0BM1GJqKbfOujfEVAEj+oH8/b8Bh8gPYc785neoyUSkhWFb/RbKJB6Jz3YDBWrJM
4WV/8ZjenXA+ErXDsu/acoJfXPxPYjAZzMZIYWDDFlznGSiFsRUqAxggcrDZm98d
da2T6zUe/DDb0mqEAUCnXdYUHjbV8+C3iBLvujjBWVOA4bHr4+Zsr/T83XQgkpNT
DmYqLK/jsi349Fborc9kL14apmptp6sv5b9s54OKWM3iLxqi1a20ocn3AOt1nx0E
ZFFlhyigGf4UY/LmB40yYS7iWIscLH7LAnScNv1Hy6UdDednHWgOdavqckZfoO4y
mAE8SGjf97qy8QWPwkNdMl7soddwp+oeXnspK40+zHIgMtYK26qdIqEJtJe5hp1j
kbX5hz033Q5xvV4VXd+MVAk6gMiq2VHlsOhuA7VuB/ii/G/1zY0Blp2cDrc0VYpF
YXTcff3brSIIOC+VaTaJpRMv/Luj+KnuHazKzrIxQ3U6BhG44MBDTFXxOk8GajN7
RDAXme/hp1GQxxbvM7AHV9qmcYHY7iy9v6UjNRXhPv86ESeO6Y832+EvmHxzCD2R
vz4MtCIndrrE9pRcF+xZ5UZD/ZcTqqXU9qqvgXrPt3Viv7TX6MWZ8tVh+1vNYQOh
iAJw60X/DIn01eNy0wW/0UED8oszTYAdjGiWUj1l5Fvj2773zTsqIjq4QZPAop0i
lN3X6e059ILp2Htek0Oda7IDmw0jSeea7eUuNL/i1nLFZNIdGICLlOwioWxIj81P
8xH8bWIBd8t2I6RkbY/d/LgUHO6g8f+VqUdRofD8BWFvOao/8kqiNvOEdbZCxAdK
TkM5wFHgpv1rG9quN4zbXryW2RwIfFHGCIasoD7EXgnJ6LrPcyrhI3CQpqx/AUv9
cNZqzf1kpK/C+9BEUX2ijZLYrY48xOP9whGsFvqwNbIKnIlDq8gp0XD90QHbiyXM
yEvSTL2GWfaXVEoJ4OY0y1cOMBJmhUguvHoNLpUcZAoZV2kO5NYrJF/5dA6JYJmk
/RJJlmWxnFyggvnaIVgVar5HeIpPb6mLLJjsPBnBt6xXlSstnHvaBimKAvlz0kKF
K7TznN8VnukitfG/GzLUFVepliQCGl1MXpp7pgoHLQawrmYgoZCzSf8pH5EbMCyQ
zqZQ85QfNw5PgBx7brWyatEavZn6ML0TtVbRyw4coeU2zhqtAguwCrVpDnjc3ALj
CaxA2OTKL6xx24ljqOiNvm9sIV7VzE7RlxlRsO0gkjGYehyYRTeKuY/+Z2I8u/cK
LarupkdUtZBufT0glSPT4kD0rgHIDg4R558qPodEbrFM5m/YgIfmcH+xZ3XGpyZ+
OJ7ewc9ZKm/QShmCSQuyLuf0nbhW5OtrZGLnHhJAWSq9jJKVI8XQyH9Qmc+hPmZG
NxE3B1/Yz5uhMSQ0lSFg2qCTKzdng+dTKIBt25MC8Asr/XDvJ7kFMGf+QyQlSAqs
XrBGU8Vpq+AvxLA12sNiAcOZDoEwGfIvVSy3niebbDEhyNJ4UQ25+2qR01T1uURX
byxXZrDUqiHeIu1nczlJqTaD83Wr3gd/Lxxo0zLZ4ExZAwJoHk0TY1/7uofqvv6A
cu979tLXJhjPZpM8EpwRjewrPC8KALgXGrxHv6H/iYRKpMfYKHR8Vfoau2xeQrkc
csMspFSNgygsfmKcMmVlt9vDlX787ywx8Ayt5IUNdXaDkwEXvh9wt+vtfKk8rGed
FkD5iav5k1TtN+vqyv2tKfIztK43r8QMCKoiABUZxNQjn4kCbmlXNS0AgW/ahw8M
Uxbm6G8eNYIFVmLcZKC5GYyl87GlQgn3VyUxEMxtARkUZ5ZpIzZIj6xSBbWfQvw2
Ac/Bowpa8eJrS8jOgo5zqLucLNWirYnjUM9SJ+tzBzXWzooyxq94QMYORT7JRmZp
VJmQIB/r2sJO1OSYw8LivnIb3kBb58FgtHWIMBK8CwyEW5RTQOkJukbUyfkt/hFv
q8TWBu5LOPjdPDumJPWZIzuBXdg+c2E8WUQrBFD+gULqu9fVHL9qOpE2mKMI3H/b
eYM62cUjnnMv/yBNuuEVAuIbokGfuKqTByphPMmEDSGWHgaDVaGRAevKAC4jBqIL
WDm2sgCjS4dUBg0CurvNMIVKQB00UH9rPF/CqgfYQDzycLxgddgr0ld1Ys8nWqK8
Hruh8r0DmbZ0AISVU9TqToKfnOsGK6x6DuM/6GEnxbDqpLMs2XEoGDWZM4P2kByE
auFsktcooD3epYRSb0ODeKRA7iK623wUB45/01acFzS/7vQ8LExWffqg7KrUJib2
V54SkXh7WwxhcaKwGm94oHVAUcttkrT+Nai3+l+Oz1PkVApwcTEvMBEWfLxkhafh
9t8vd25oaUrJvr0Yge9TTYx63/mYYeKcoqt/OvioOfwUe11hWoLajhqeR2CBsKyh
l8PQph5+Wo/s8HIq9CHUC8tvF9Z0mpe6d7YjH/I7wgDk/Sin1tal7+IXOONKQAIQ
gvNqUf7BF4jCXhdpizrH+pYoW2q5f0HbSKpVjt/Qop3jIJzO4K1Z7e7exfhHT+9J
Fzkuuii6X0br8NvIVRNgRWsxMugKBVXwoNWoDr4sfhLGYHGEC0dkuzhzYJXn17bR
07VPGG7+ULye6xyJOe+j029q8qjA5vzXc0oPnIG3nNWvmilgjHdKXu6dhN5FFY1W
tGapanV31C5yCa6NYAQvA2U1UY/h7i37wGcdvaLT3BQlr2UGYeCgkQzFnsF1KLOx
AVOzopT/POiweIJkyzZtmnONWNbc7wJ5pRf6somd29F/paqluNuJaKW9yL7V7y7a
guwNXfzWotx/nnuX6T9aQzOSvMfFOQBm3rhxIsJL+qMit+7dTYM2AstN9OLmDFGl
tfWqMAnbwv8QaIpwicsUueDtZ4FjQl6dlLjPS4G5aXazjo4MdWe2JOm8/GsK3xlw
RPPvOJOjSPllfVZ8zw7fZAsqb752jstdIoUWh4ZfcdqCJc5NC+b/VuSvAqWdF9i4
UmbErzMa2dUnCP0EHHVwrlfJv2cP32dlvJAw53If4GAnxhdKQv5Z+W/dB76lDPhZ
0hBrjfRUS1uUKggO+hH31aybh2X2N0I7BeTQ+9shQm0+6TQ52g2HDAtqWAImYsOg
tQWA8UUGTwnslncTnx2K5bFzqw1hLFBwZve7N05we+VMHx1/HC+r9/DOJ+ppFtXy
0tnc2gWDaP0D7CHKTCL4RiGYivmMVR7se3UOUK7lXLr3K+xiev6omZOtfklrZ+o2
7mE8TxSM7pi9xdZRm7ZAv1oNLHq+yC2tiOdvORnTWF2LKMLKta1qMDIxMdG701cH
c5oQPjOWCSvmf90sN0LmdAmRruaZJePkonMQpZ3UvA1pIr7ZsvP6CwnifLRNfDmU
qaQfU9GA0YE7A7hucPoMKoSQZ5Q9HNP0ywbKygGkaKnf8z76/QdItDv/S5CZ8fd+
eVF6Hzv4+YWKD9IMBM9DZTtYSqS2VmzyboFndGkFHbUz5G5Db2vz1wuecee0RD+/
wRgi0bWc9PSzcFON0xyJKskUitPX755bspPOFP+nD8ctwEaZy3DC5+TBUOrq31kS
WdEs97LJj6vP2pRFWEh99E8ecrTz3WeliAfXN/nadu4=
`protect END_PROTECTED
