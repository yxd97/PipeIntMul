`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ym7Zq4ARUMUie/8NTqN3XrYsLssQGs9IrtlsTlLMdeABKO0UDxIlOaeu8XFaHXXY
OVVg/BT+sMGKizhR10sKNq+qXxLOpArGEuakS6/w7V26b3kTw4suEwLfP4TOAUeG
wWpb8tMxMHUhQsA4YGJydTD1zP96dHBQpDcBerprbSCaRKlbnfbDBN66dzKFito6
k6pjlqr19PROwZIPn9DRDhC4keWOrkxEIq7Z+Si8ljkfnXupwrD02OnJnv1NJNaj
os4rwCK/FiX/LDZ+nOvcLgP7o63ZKsEFt73kKZlTvUD2lZB2O7tCEQIubFEawFK2
qGfQFSE6YaiZEczqXKemesnW4kJJAo3Cw35HqTeTanGxHyjBXXghxg2eyyFnfkAm
Q4K1L7PZxXGV1ngo5Kx4eS7BSaFIGc7hGUCSz53AfViocxMFfhiW4h4fV6yYykOq
y7EtGX8NDqrZcSPdInR6NgsSDHwn0RdA/DsV5BrXvXM/ZL+APH72pYRFS/CxhgBa
7qS6ud1A9Vf93oGRapNuEmJFkhIBWU2pCE9jsp1LzCy89E1elw6CnrgOYurKlvXs
MYnFbTAEwU08xy8m+xoas8y9Zcdo9nhZ5t/W/m6HkxDRPjIE5jFI+wjW63Pax2C+
`protect END_PROTECTED
