`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
upV2bxnAKC71+uwU/w1ZOpGcNcJsVGhfV0TnxcFmDXZwpP+LYYHhcK6NfYlR2IZe
wQdSz8IJFkdPCzY4P5ZhyxBTiovcfBohxD6N3T9uzEc4qFwhzHHXruSc+QgPJbi1
W03pATPSgXs+XHe6ZrnUqruJ5dR2DPtc6B5bB5YbCY+kggNhT4TIWqE6KGzHR49F
90zSZAEGFHE9gazC6WRRPM5gg4gveDR34hEGZ8iHiPIiWWv0HU6noLsIrXXkoTgb
4LRtDfHOTsjzkZ1Kdpawcv5LhhwD4e6/PH36VHG3lruvTbYMfujDuyn7A8XJxt4T
sJwbjtVRIEUBATNQ/Y3fd3KCssoiKvSSNeuViOzrFgpnZ6BOfQNlX+R+O6snj6iH
ylchqUUemkMjMkwAS+ypx7SUr1Kb7DR3GEZMDWmg0XA=
`protect END_PROTECTED
