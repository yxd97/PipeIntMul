`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/8ltbuD8SJeZqGekBhlgU+O2ApmtIhGKWar0pel97Cd6AnsNLZzOoZqr9gvf1fq
EOCiZJ/LZyY5JoNmWmXLOy6BJE6GSIjQOWKmNtGNDObECVHxLPlwrFNPaBZX8+n3
KWPLuVlrP1L8LPvFbtr7qbc1ZOdn+4uwqUvbzUNy71BCHbWJqWJwU18sB65a84hv
dIBahvubAz28ZTEUHYc/3l+1hnjOIJO8bR4VETOrmg+W7afY27BOtdfFPQl69rlf
OtAP7p80g8y+gpI6fojaLApzOyHDOpjKyg2QdhB/RgpqXT7HefG7ajSZi72NY8IT
CGR9SNksEm8abewgslwkb2YGgNSwZnQ06TI81QW9CgwwTQLB0g2kDopyb0J6raEF
eSrZhqL4vZYFSwp1CPURZ2wt5JpSYBbhBh9NQrzzvXEv3HvDxakKcpWtaBYYa62o
nrCH5gTSIkpAbqqJ5KKZpNR9zc1nMYRsqWQkAR/h59bKvd0MbD/GdWAqtLDB1KjM
Ru6nXvDqLxJdcvmvY5dlvHkzBto7ofoUMoYpS6U8tJXno7aoEbrekJ1aKQwerQVp
hc1VqiZIOBnwB66m02VaiHQ0wRvastLdYU4QUty0RSqgkUv0qvOqyCnV8JwLQIWE
woveTWBc63xcM3FeouH/vAzoCRAinogZ0iOpTD3HLAja1PeAiXJHwSGP3CT/0VkN
ECML7Nv79y17O4/TF6PlhlS4sbB8m/MRpoPE2pRKmTWTBZTXbRyxAeGTp3Kx38Db
8KitmkU/OJr3mF374dwmP172qjYLbLlkOYudLKvxnK0sxDFzNZ+Kb7POCigpHUcV
Jd1dJEnEHagcLEm+n+OqK+psuV/cIrgVlvBGa2LkElGflieeNIHHARaYFs9UGsHm
hXolo79ZIaAJq2pTW46Y2CVO9rtdGZklWBH/IL26jlLXsU9UJsWNrdZ5zwyuavUK
Vp+BzRt1cv3qtUXN0nZja0ZWvc8FxMrh0isjc0LVGvS+y5LK6ecvoBR0JVYYpNBi
`protect END_PROTECTED
