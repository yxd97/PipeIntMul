`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KallPuDd8b/O7cefIim1NVjz+60rcfB8EHX3K6h9eJxfpFSJh/tcQj144C3Uj6CQ
3FYR7R4PCitiFh/KvjtZbbUgD+wc1FzKehB9gnq4qgbK9uJWCRY2/iJ1oNK1k/Dp
IOpDrDBT8hiU5jLjFngnisoNY9OMGUtkkAwswVUYjF1OPGdnq9pD+QUfsGQbtpHI
74vmE97NdvX8eEoSnaBPzfDDPLTP752ZX9KpPhoZ5ZFQ+WBxZjwbkwY6CkB7jOoB
m1WSyyFRpXeu/M1n6C7Acce9rGxpkXnIGyOWSdGta0Ii6lHdoZmkp44aYzDoJrmb
VaACk3/hQAGuksUrYvxn8EK6fPVttR9oH0CVFduCNSGRN6yseA8H52ePxLSJme52
L/WmjHmd5i31cLIxTF0/dQnHnSqwW4XBRyKFLrvWncjofw0+16HpgNFiPAOZdhjW
JhmEFZxRhYKbu/+46wahYTR7NaKsq9GhyoZGwGgbBEE51ajzQDZ8vTc3vqYmNHrZ
TR4VRqXcEXXVo8Wq2hz1LGWTdaDQ12CSy9pDUpRb5p4U+MILnPvpnf2d/m8csa1A
yj9R9viZduTPepMGWpu3+c002zJ88Wo5Z+ngykooNBOzrfBPiVCF2/4CEhZ8Qebh
veZwRWOh6Kk33MEe6b3IiPhJ25oRgWfHfWCbmEh/BdQFtz7QR75kSyWut2nOfXm2
mUKpgP2pJJw8BYGiKxiS8+ipkVsCTFEcL97Wz8hRHYnPOjoYH0OkLrp6w/AMMIWY
BW9i/x1rT0JY43uboMwnRudCkgB5e00xx5AwJXOfcgHCNEXxx5y3eLF4nM58cNGG
EzRTJkFSk8idukTjOYGlZYvLZZesWmRqzmomNfs8/jASa2+HTAfGMmUzpLhfPxT/
EQXUZn6I8QXJodcP8SswPV/hgyoHppX6YgXRAXzwsvtWtnJFKQdrODPocqAi9Tmt
3WlOqIHpQwY99ICdoQBPkKJt2SCLo+WkRAKFuodqKBW03Y1Fbk62iJBBwlJvQbz+
noRJKdiPb6nslP30MaXsX9jUJ7WRZci/YynqRzdiLYnw5j/BJKkENmEJs5hV6Pzj
+jUCDqMM1fKS6r21uMQk4swBrO+pDNFvD0DioUyo3vPJ/KNQ22krVjx1idIsMsdl
zo0+Bim62oDqJsnaJIaf5Qguy2iQlsdzzc8vnkoGLmRxFZGb4QK2BPvbkogPIg8k
HFhfvXKyl6YRqGwT2QGltkysTJbhprAjC7DhxQ/HzbU1LVf/S+nC0V5UpC9Yx1Bg
2EGMVfRh4xS2i4BA50k25Po9V89EHa49BKYw04sp2tyXiDa0HAYkzc/waNno/Kyn
cU9KTD1kiED5jW+S4+MZg/OlYVOZL/sWpA6aS1EeshBsaK0+zdhuTI+CH9SpC71j
VnJnFoUKqQ8OeHEbRGR8i5Vac9tIOYDkvFAIad23FHI=
`protect END_PROTECTED
