`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODiZnmCT6ImT3DIrqthoQfslt7X0HUfsZ79RLlRqazl8ZreFlZypUC0PZ7eLAlHI
0FCFBj9tAXaVRprGm7ZmDcIU6eB6Z9lFz1YreOZVZ/tyGVS3ET2vVirZmD9dbp1S
8lELfW/8saqz2cNK+kHytOhTO272fA2XaNtAXsMy7mXE3uokqA/3fkJwzJkkaVPw
MNv6uxiYlEcMU1Du8fREboi2KC/FrYSJnZT5nsyb7XM+kdkJIDxd6u+SxyGOFjYY
Y9Xo28m2FAMn8sxAxSdKS2YVmyC6yS7vm+5PwDiEf1yfQrBmtarR0Eb7kXXVuruE
AsYcLM3W5RkmmbpzlCGW5qlKv3E9CDJUdmnsXiqEnRsuHSIgS/QU8eQbKGZZAUAr
enVSh+2Hl4VQucDVxeQvyLOBDlTSW2J7B/E7PJj47oLd80hndYtJZUSHRT/jRK3q
kxh2IkTmCZq4zMnL8zYYx6Oils0UUXTygR2TBIoq9rQrTFKUC8AF7PJHPA5uE4lk
xKatl88e2kt0+iRrSvGqcOFMqoeBE7zbEGs2O2AuO9L3zrq6zXZ9BGZzNk+cQkqT
zCG+lkC8AZTZjT0euaSW5E1HeFN2Ud9bDfNWqYrZQ5/KhaiR77PvrIQUmX6OY8Av
5P7qi9M3EYsR19T8hDtqCsv9UWEW/UNs2b09DlCwam0mC8wBdvY5rihVEDlUimc5
jR8W1VGp9i6LGQJEYjo3u6tKEFAavZ6ltEHxEkId3RdfWoWChhmyU44hlxy8cUjX
MBJqeHepzhGhedodqiqUwHO2O5hfVgW/jDi7qM/EXo+X8j35e2LraBYeuX31sx3N
GXSUa/Ai27pM5tc+qjmRnoz75SkT1jAcUkhEE7Aic0TiX7ZgOdBKUrE+/ZuBGi9H
lBPrGcHVXLEw0+6uuU5vUDxKByjjVhWlvT/zbHmOJ+PBxKFWjtzSGMETuGUSD8sd
`protect END_PROTECTED
