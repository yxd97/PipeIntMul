`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P7QOFLbYKGolIytV5z9/hqX0SDapmAnlFLi8zSMLhLDHExawVp5uCDFFSDroKo8Y
0BVnedPThn2ataCZp+Ax+0zoY+ppnpCBve3RTFnVzYCMzK/93hUPqZB2EGC1YjTh
uT+v/jCFozFRbeA3dGqKrb9WUVKAOgaBzl790LYMjSRxL2MlOrpo4/FdZvFzvrTQ
icIx7oAV0KBWsZp+rNPiRWuXv58KDuonNhstobs1xg8KzubFaVVBlQJe0giwXhf4
sk4TuwzcS/qhcUni6xOh7er3iQE+DNj77BqnNDi6yBz28/GDh64zmfsM5w18g3HU
h45x1Tw6iryg+dhlLrs8VONBTm4/J3O4VzzTVc3EvqzC9iMU6+Fj7e0MLOTUeASq
ZRTeDgtB0CkxsJYjss9fpxS0SHF7X/MeAB1huweWe+Nk7YK153r4jdoA/Aw0Jcrk
WgBs5FVECdhQOc97wiLOlYKc70Ym0ZKpJYS4vV+KBbLEqDFA7LUJj+qAjDp6pKn6
2Ncb1kpYRDBgfJT9sAigzWh7EPQo7SRhwsuXyyePK8agYvtxq67+4FbF1NJW7NY8
15jjJJjNEw84qFnIMF3kqMKIhfNLdixTM0iM3x284yYCjLNMDdAsh3OVsraAjyBk
pguXvqqZi19fNjZvrhTn4w==
`protect END_PROTECTED
