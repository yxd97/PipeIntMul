`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ed8BgIm0vMJL7Wz3OfpJaoWZbqfCkZMhQvcqYERdcxJ8i7HkVomQCaUOLe5ajL6q
DCOZXWAKgSB6t90jHCjEV7AS301ZxZqHJwd2ACuX2v5b0ZprTgvhWTbr2w1gFad0
u65kYkFK0nMU6QIzUNAFQffGqydBLnkAoNRKRkw3ak+rmSQyJe5dgMqVbqXtNLvK
2TtJ7MXOFRz1QCH/EWXHXv7JlDkZtPKuxN2AMmf19GnS3Wq4iotOQzHzJmNnwGwz
pa+DhSp2N+t3yAQVd6jgXpGlBbnh4ijPCuOa1NBUEQ/m7OOIwsf3NGzeQIF65TH8
xYXCR7mWcwRzbA6U25WK31IEGA6yN6ZKp4amPwgshahvvF4s6drt61MpwLvdVgkC
GGuARfTM8xpWuWV0YVFY4XAOB9BPcx4nAbnqcZ9wOTDQ7qKNGQFmEvE7qeNrd61I
B44k9hnKUitGdcYJnIoLwR3OTvNc2eVhv1N+wW6aj47T9b0fPalD+ZZRJOI9lJrb
d2QvMdVddyXUe9wxdvp2YpH0J46aOtu+MVorxLGX7FDj0RQgQb37uNjqgg8xrG2k
8fjFY39fO3EmA7d7EUQYwise8XpBlD8NxDnkHnqDWA6tbxuNZoJVCon025+VST3K
NPefshbjEgFyFt+Bd+nnYosoyc7ZgZPM/kxmWGoPucBY8/E9C2DPBN9lLebeSxNf
zzK+D1J3JY/oMWAUT92Yq++rGkc57XlKoBwC+uutA5dsDiLjlRAhEnl1fG+4Nr3T
zjUgJRjexBeA1liIWroWxYdfaagt71P9zF/2s6GHRMfZPwxRU2MdCWFlPP7V824L
RmBaWibxtu5wGe0EPL0n+dSCFUQ6hY2RPl6OTRTNsOcOYOZdVuflUI1sXfZvrMJU
SDlmvolMAjGzFQJolXsZSEJTxc6Txv686DoEcIn3M2ZtvGrQ6dR3Gz4NaWSIHHjW
EakrvBpNw6bCCNQLwvi/KA/Fylga+onIPgwvcFJWrmPzZXQczgQOeb7KnSTJ1u+y
+cT2A+UWCZ14Qk8iQ6+HyD9pqYdM4dW7JiV5loWqhFBW7EaV21UcmxdXNCx4QG4I
PQhHbhK2By1IbBi7HybZtGb1peXbFYuTGFXXQ+oGti68QXl5eh9Ysbv0ZdOvsihs
Kxe3EhqQm2uJRT8dvesl1Sn5XjRWMk+3H1u3/8l8Si8Du48dZp/uNTRgKqUhDF1z
GnS43kboKe8YaVcSFr7kHZP8xsLSBAhGmHk9Gjti77KA/LYT5CWl43nWUv+EUhPL
5nqcnt8W60I33kE+9nm7E0paGp/Y70IB4lQEl/O/nS9kdeUEETRTFhCUf26a95FE
PtD44h1Ul0b4741LlDHV6bt2mLEOa/VZxQaFtwOnwVhrcntMR/p469z5QCuN3Zws
dadraJza+9aTpuFD90Wb+KZHI1rC4/wsYKKcFcl+sNVnRc6OqSQVWDB+G8bzwL0+
saW874FJqI0fTNoA/ulTNGhH2f7RFsI3PMAHek2KUa/WaF6I2Srs2mZdADoiwpHW
Ehcbbyqiz74t+9UoDMize3CMZLR51eua38Y8XJBI0hY3mTP2Ccs3DcoOQlbYdP/E
eTtarTAoxM5ulO6QCT95KjopEnIkvsi6e/G+1txrHW1kwpVq/U/6WxrRsmxP26Tk
Kok8SFSTtl8nsq1XT6gqIzIHWg/bz1ex4PVo3fXQtp4w8UzrKO82S2AwJtNQvjlR
Yh2Ofj8X4vMaNQcLqt9iSQxpWzwy6J41OXQLMUQ8DbIlTMGqFjp8zsWSVpLFLpMV
MusFScWwIe+ksHAEyyOA1AFv2KtyEPEmE2Jo+WN0sUC/atv9rXufXk9VXhj97Vbu
x/9ubD8gdELywJgbBOVlgrgT3X0tkTjxwZ4CWUVj1mfzAZ+aG5PIjI6LCQtn5QYp
UWOVcA4M8ZoJHdtiO0HCjV9tUTV0nwErspnDSXyIMeW4D0+a0g54OQa4SLwGm8l5
pS3Mt1fs22t16LN98zQ0F6EtY5+v8N67Ai/hLMG+WSYYhcT8l1Sj9qEiq+QMJse4
mrsBmTcYH67vgN7rQAHkSITMqCXd6i4G/29XedVfxMxpuU3ZFmvnAv5mUkRCWSPL
UMJnCPxwn1VnJHypNcUn5vtPPXk6nYtso5YVISI1CTLUu7K7G82UN4LbU1J28FHx
isni2xV/jzlcrIijTt1I+EJII+X4wGE2J3jNqAq2LgD9Dxa2EjQOloads/Fkkyip
em9OpFbocf5fMrjisT+QKo+/jisWzVhGVgSNBPKO0pEN9TJKvBzHIqTfYxKokkti
+1bfOUR2ydy/TwkjLSwevzJ/uqNvD4TxoRFYsaJoQaOuZo2Ft3FTqP0FFVsZCw9y
j4RHt2xlXuUEhPeZebdW5urj6zSwqiYFRONaWjU2K0XRKS3VMK0b/VRRTYlaGBe/
Z9IRAGtDx2MqzE8z6s7h+clh5sZxzI+mc1n2wFPOZPcfsY52ypIZlAHpcCB9ub+w
MFSj2PS4iEbWYxRCcJGRd/6kntWqY4Jz2EKxQ9+1QjyJ84+Eq5S7xy+k5wC2LL5x
KKJfP0ISDtnc2COXxYCfqga6FN/EhqBDLtfQpyqbjoT2vdFQiTWqIGa61WDcCYa9
jU0f1qc1fWphyuuxWYj5XJCpRxAPm4PuorXcZv/O0pNqQxd6bbD6joWGWQBRJffP
+ESLuF7kEQ4pvh8hbp0Lznggzl8rFa132ocDx+7u9tvyvHndgB8fle/Ky/F9ZgLY
D8HpR/zLI8aLGl6NeE83uc/vY59QOOlqGQfu/4ZmPuKF7nJzz83J6XIFxTt4nEEq
lXWi3Xwa/AHnWaYtbKgoV+SciPX8woVeydyjuoc8A5+b6K2VwcTLTPsYTCBJmpJ4
bFd0ZmD/0TJ5NvMxDwHGTuUE9KSCltWRMLH2OrD/JOGbolbJua/gFBgcZwwoEhIV
TsIPoS+Ty3I5srsYdyP6aeljKRzFaYfBQdg6SP+I91chIpaGRBCr/bVam7ThKz3v
PoOS/17+wGiYDr6e3NDhJTFdboZCUSftJjRur4xhNQQY7M1K+nd3I7qocQZomoAo
I7lCkYRaDXvo1f5F7Z0gBxj79AkH1W61QxG31KtvMT+ij7r0FGHWN+xnvtypy+qo
+wZa5nE754IzvpdbJr+XXi3L+BblQ7cq9lZDu0fKnYsLiRCX75ax64gQGS2o5eo8
LAZ7BU0rm7QHokWLQETYdzkb9tyKulexqV7WPbg0XEgrARGtxSfuNAu9Dmhykuvz
9JO+a02SeLlGHcMARdm35w/yBE8vm+sQIbH/srazOQtRZRY3oJf/DcM6BXGF1bcE
EMek8CXqGiFzRuZs1SQtZS4yC6IjKf7ZpxHVGvTYdTgnpt5iWgoM4TaMZScGcfog
xCy/olSQbHC7kVQxttOP8vbQc+mRmSTlyeBRl/ach/U=
`protect END_PROTECTED
