`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JQK5BjHd9QpZ0BPtvjVGb4hWP7ZEAABQxeOUdMmic6FskAINQQGzD30aK1S66tg
d34ArFEp4IRwEhJzzR1CCjMA8WNXpOXkoXqw0fzNfqQEby/AOnEhRmQYpzUWx7+H
7FIOqzb6tB8Bfarax8bsOJtaQad+79hw7TA0RR83bOlpzY4ONuZZnoqC/babchOv
Hi2Or9NJKt+BzUtda44SuvMQa1tyAqfybW5MWkT7oSmyTVq0TjzkkfmwAHkASiMH
RJCYwGl6xjh3U5Of/PYHxdB+BxoX8qseYqSepmAI5XSDs1GL7/bXDOR4ysnaA//+
9vjqlFqH/x0Xtt69YCnt5830szL3o41JHW7p7SKzdfPqiHNa9+08ZVCw76eJRx51
uqjQomTL65oum7KjaTAOFQ==
`protect END_PROTECTED
