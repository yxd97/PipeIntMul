`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2sAFkCcRnekTtMLeav8weY5X708wN1GyAOo1uJ0HRMGIFCXOKTCkhmp7XBeD/HFV
/OaWjGtYJ7N9MlpGj6ktNwKJ3B0yupOBj/CkSnRXsitjUfMmA/wY+3G8k+zg0OA4
krpIzpOTB2c2yP0rHX99wtDKcfmLV2+Wqh3dADYmzKZMrKyxjZIPKGa+VV330ZBj
EH99Da9bf68XXdmrRazekFiqkXvtED8su+3ZtVH54Vjkwd1C+s7unUrsCsDKsRgn
oEimaOcb4P+qZ9XUO5dosmkhUZ2vL8X8R0wAeeHZX2HXuGwM3zHVrjaGSJiWJJZS
+vrHU8RH+y4rqvsRq09f7O24qd+jbEeXbc2NmfHHyB/pldPpOIMkiymxDZdOjpb/
bW2rZdXqBKMxsH0DSBWUFW75GooR55xq/UKa8WxXkAlI9lSw9IGRmuacf15qrw4d
dw/FTmv43j9BP3JhwjyXBlkJOkKp3jxCv6km4w/bcOCtLFQQNwQX+s6JmTGpVVTr
VBi5Wor5Pcvz8kuQilGudxgDBwsi5rqdxrxdNEDVYbCjzU5NYzQD8E0NuYwikVRj
BjLU2YobXWG2h6WLvUxO7frlC+rvVAtCvhNH9RZjMPJyftAop8vNsUTzJsF7x4sU
ZrzmU0AuSVTdaMsOmClGUoTWn+4e4SXgpf2KJtfJbaCHkTf9qE4PAGS8KLRdwU+c
uzNTBkXCG4bYwAEQVxQtKDmS2p9RAIfivDWzuekq9LZf88YZkEQ3uK5j76p5FSJ+
rJvcqjd+MpVToHk/ic5JnBIFF6hIzGENZxMVn9VgqvvTnmNZH1gWMgs11zm0ORr3
bGRwVThhed8vSadeTWeNbq0gFf4nYw0/BizynWgLwrwkIOldqFm1HoYRCw3Xa6Wo
Ozo9c6mv4BGggjOUXGoQuZ92fqJniJnsTLp79h+ffZJb4TSA2aRYaCaGp2Zf7/Uu
tE81SjY9Z4PbLuw4sg5jC7PiypGK+OP0yl7e+wvuiiplkc4xPrQl6xDlKfsxrCQk
MSxGCEeQ4W0oV+2gxj9xZAQruG9R3WvyhJ4EdI4w4cIuhOF925vzqfPNtMoWTm3z
Ccj2GSz5HgIrcHd7KAJBy/Kzx2HB6yOXb73vtExA1OOHVb9xTMCNXpAFOS2FTSn/
W8tZ/3axA5UlSQwVtqepObKaaFXyJiM7DfKUTEhWsbfkU6v9VsrV5sH0INnI/d7L
P2aF5g+WKtybM+Ph/FAthuDxlUA2+bdg9xvKpMQH+safrYUgCVn6rR2SehWtyPp7
SyiPBauk+cGrm58DddH/EUbMNHFwW5LGrc1H3BcQ6QDZVHATj30JIar+hmm9Xt5e
UhRsKJHvuVbOiKBolQbaoFTSF2pqq+rCE58XlSQfKd0p0TsVCyYhQUCuCJrdQaj+
pNtDrqSFRT96AWx/6f+4Bq6dt8L9D6ywytX+AOh+NAGPAZyYKcaJzIb6jzCZO+2X
VpcuPmAvZjhYTVatbQFN70r8luygQIn0wFB0E+q+zFzsHnuSxYkDAmUoqOouTFAD
va7uvO0tLSw5jvA3ncwCvnQRjD9PRy4wmUGqO0IR0MR1HgOc39GQkBt/W2gM6UXt
9VVH40kPLc5/xEvN7+iQrTKUoTh50e8R76VhpAPM9cbm/fgwLWKqkkWiLj4Wj9dW
fnhq7lbDNANw1Z4cGTvr3435u9qTedCIzlYAfuMsZwUZRCvwgdY3vMlOvubetkvd
1LOYUPLr//x+l5Bl+7wgoGivLF7oiIHV3d6FsCpmEVZvEQ0j07kl5uXpXGhMgCwv
cgVjYL+PB8xE86ReV2pveLVeQxcXg39kt05eYJgYxasFGQ0x10oRVIyYdP4J2+mM
/Sri09zspLu7cI930ExrPKk92t7kj+OoXIJKsChUGbcsufaUMqvml6+eLFMR7VS1
+M+j6kPcwKUU92j6F+TmwXkJa3KihQGDuNC5WyNcHhmyGaWJG/MfZsN5CBfSCBYx
OgImy4DWDsNYeQTkzRchvhHKxKxgclW6NstN2yLeYHr/N0EZhDb8eNRNLc59tyEE
KImRwgiQAZ+7hMwGPkIYhT9+EEbw1LVFVO9WMeKzn/h1TrtbM98bRwSfQWr2TyRI
0+OMXYS7heRJRpKiS4HDU3hZAfj8U4nfxSYoFuAoBo4lIXOqbnloJcp90AAoqCUL
20gdTQKI46v/UHj41N/9bNdjio4j9wKQSizNokoxXE8kLvECwt2OTvjUQt6hkenA
Ou8k1CaZwsmvBYv8sAHnCmBp8yqqup7YUslcscD2LjMIQIXcNMt2tTIuI/C4/dZW
WB75bDJhKgJQIeeHRL/rtdF/d0m038UJKUBJudA5s47N0vFK5BZTn8FWCwO6jnhj
qdLJOYcbL2aLmDP9VwrgcBIYgsHXKfeGLSA9i5Mv3kvfBNyqV8V5zjrkKlKbaSQu
sHizNlER9eElT4L1JJWFOQPzAJoOjgu5c9PaGSmIjaPHlLewoTLvXYbofjq4DoiE
NfGqUsZAPineRtG7mQqYSjs01usHbHixdDLz59S5oNwaCqZtF0+vXgiUbe8zYJnE
zTNJfO87Hqz9ZR0bfMd0rJ9DyyStjWW0LrC4OulrXOGoBDnnl6jqTndjRzbC2c5+
KM+KAHmluDzgTjm50HwiZhEGEQH9zQ4x2aF1659VXYImTa9dhcvz1kVta2WF4uPd
2PWJjbjOdmuuguxS5jfSNKm4cGobzt5NKtoGiOal1D4=
`protect END_PROTECTED
