`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jejF+z9faIOM1PARBLOMZiV5X1scXC+m3aCVn2xw9/MNitEd+PYD5JW/PshV1jPh
zab9CGX20tJJx3Souqt4wjZSizrzAUhX4RYNO4g0op5J7QHjPqQ35G+mNNjE6jEx
6mm/PPhsnMD61pG6wqQQ0K6Vxj0av6jl6dP94Ik8MDVSYINXtttn6bMyMqfdPYj/
6C1VfJbogZXEdC9RVOpGDUow2Rp6KnJQDcjIDf8MOByESlLAulKRV6jhbZWP7vwu
rZ5By7GTUUBNgEXRBiNO2qGTUD8g7ANrzuVa8pYypxOwsiugDYCYuxMWMBt46zTS
7ssuJrS6bHLAJhbm8XwDNAiEXX+3tgAR2QpYk0PkjBvZJq7hbGEGeInPLP1WTGXw
3aaifKOA/WqVIA7lgYzr6n/KwjcbSDV8WVr3Y2ZGF2hvJ+W+QKQUtj6iv9uybwmo
70jEehGwa98kfQwHqKgMSc/auqq0TGYXOZRzOHew2+TeXMTay8ir548/xcGdTkMJ
boGEAQxONW8c3z90EWNrmP68+8cPdIFSr2I4UKp1bblMGTSWnw0qmOVg/Xgt5Kb/
xnGfzA/glOWpnXh+mA3aAhVAoDpkJvUSLsD3e63f8ht+LJZ+zkG2ApuIJ7OPJDDa
6rC6l9j8DENlxa41jNeEst3ge7aDWkvUtdE1HWdgdbw9UH1nd5iEhaKwlHjHO4P0
+uGDFQ92Y4vFPOsn7OT9UdhFCkc6Zt+GpUZDhJbOR76NjlUkfAHf5uGf1TQbRkYy
PFHAO5d2KaPoOAI94u7Hifi8GCj+8XN+y7NtamH0VJbtRhWDIq1B1F6Gr38TipDa
XmZU995HKmWyVpjSOeOW/SVlxImApykCph/TBgcg8haA4Lcfim8IwjHce5G93ufP
U7E3gZ/UgmEuvnc7aaG8BkUYz/cF/8PlCk6+kc0A+6S1x7+r0X25kKD7Cb7eX1Sq
uVT7Dos4BZarQAKL7i4q81LEAUaTxu6kyD3Zt66hb2xCch7rCJf+UzZygZM366eP
PFqLpUYaKhib6sdySaA/geii8cmj1tQKU82PO0gQqiSBGYJSbo7adBQTZ1mvRJNb
5qMjQQp+D8LsjGOGs5/IPqIgz0rAqueEXfv1yhyZiGd1VaurT+HZTIChwQjXOLnE
M4Dg9OittUYIbJWlmniG4S3XnW3b3qlqXnX3BZ5PZeZTQKHwRpdp9XV7NAZ0RPi2
BYaJL9B6ewvJGYoCGoHesARORnvxt7/LptKuVv2/CGJ6rbZSVXkPd1LMgHOnSeUU
2Qv8TJQB0D0fN8waLW3FwesE+kXjdp0kjg/t86AiqnMv168AbdkcvvHXAAq8pNV1
9kfFvTp33Uj39D0/EHbFqls6renXiFGeTnWKU4qAYeG/eDW7PZY72Y4mpKZB1brA
Gptw7Pb4qxUJqnReou2qFJK2lr2QGhsf0Ihlm6j9LXni56RZwN4z7yeMm2jeYmL+
tgwYCTvbxk38xc9IaLmzLCTNZqwwS7tjeaMsfuo/hmiUqoOFkF7cUu7E1b/wwkuO
FfWzND/9kjxykXwZ7qSjq0lKohWXhzpQvTT3/mgJfQifLS9pVUqFw/g7rfwQIaxH
cskPkIBTTHGuCiewLAjGvQaGqHtJNaOSwtPFCKu05Au4JuIwh227qicEratOU3iv
h9kKhcq1WJl3CZ0AM1QFIiehYMqu+FGPh5HNFHIUS2N4FXLd1oIWqOiifkZAcSbk
hkU35TX9cjWeuAJUrwtFBo7zLFS9/vIqX70he0ZgIE3k7QByDAZMkWTBMGpIYrQF
RX6STxKMpSGX0PkgZdd3JGlcLrNbVy9YfYCfbONs3gZhCL7bEW9sUXjZ+2TOLrFY
lNIdNXRQGyCVKZSIoMN50GA2n3XsaYCJ0/9LIbIdo0Vx1oIoSnlsToDK4CQFVpQz
F/aGeO+YsvE9DaNC+D5m4yxoRZzoKdT2Gl1xQHmFZ8nwrtzhSOvo2EWH8gNsvUsE
xXuuxEGeYCwKsXOlvssPFJW5451AOkYiCzq7Xum4sqmG1jN5gtHzd0SDZ9pVseIe
AWqLVEdRHnoYjfJvpdcJ572hPfgw08ZAyKtQr0hZzrIk6FvqU6MEroBi2Y9oYugU
W3HvA7M+sFKaSJYGmkGrdv4IOuXIk9amAGMtj8Qr15WOF2lOSarfywb/7n51VoRz
bFnHLkOdGc5NQIHj5LGJSh6va6Wz+42N4lU/xoHse9Cwi65X7V7AP3zxjdzBPLjL
IwfxshKj+45ByYmn5bGvevQ5ZPYVZGJ09dl58zHf4fj1LdCj/r7b/n9rhV7+EK7c
GARSlVvr0bAYRi10uaP1SVnWkZOOq7Oy1BNnVEYHryrYGg6Oyv0HUrTmItyYHAtI
iZcX1sO6Rk/Bo+ptGeymOFVa/+1hyZTfFf0C2TTcsizROs4fgcPCRTgeqZrCs0xz
RmuF+ffTAJYHfxu8vQlIAEV7DDiOSwmnZPhiZGmQ7gP+r2cDU3X9V0f72m03aKS4
LF+IFj1yNYeFzzBz6mzcxbj2s0ukoF9WYGwNDuiB9N5pHQad4oZKKnRs9Bs7NUr0
tfpHIti1b8jcHGbCZQBFO5N1hn5t2DU0MQUK+yi1su16U/JczR5w8VPIWjR4V56I
FJXzft8FJwBrGSV4zCipz6yUAg7UPZ8DYXuuS+9hL/dT3UcTjfKrdl42QHpkD9Wn
gq+Ocboet9aP1pI0ufTXYaf+Z7JnGesZqbRcLdwOZ3Q030ZYX8H8UWKmFwePSAI2
OTvpZSu6RHFYf25c6mO/hhQnw7cg7qMYpM3/QYu2wyRHAkLxe4CXRa8j6oiKJbHT
BEkxTAZFymjox8srB+BSCPvXxUtKk96gVKz96bspmgmzgntA4k866WzXUzc2Nujy
H6UqtffaKLiT4C8blTyNQWIQX8tnz1pU3I0dHI7QvEvpykqVJd7R/9uGSzpPQ7k3
FeUDG0qj6a6NP1WTCaXrqTAgY4ZMn9GNGfxDnZyYOzgRlRKGpo/fKT8fbnyPiwz2
2JbSUL/o7TyZ35Lm/dPew8TEscXl2pR0nRCyHE/46A5PshBpIBqahFvdyUBAK2XT
RewdvYEq+w2R5HDEyx6hVNMh7Do43tQyjLyNqHlEBqPFWDQk4sgB+p1qkqiCepoY
ckTZD0A8MRBMX8cCMK+wYiSOea42TNPzY1aP5eAHVPDzKXqK+7W9inNMwJVNZWcQ
hEYn24pm7zj3+vUk59c7tZTlmB3bmmHSGqEqeIZRdBUIPJyVH3ndwx0jfWP15wGc
+/Tbi3oNlJiSeziKjX06Ym0SyShIS9BbvQycKf8dHPCYH9uRWfkCwsWOx4TH9NWY
EVu9mke8FyVDdV7ip6nHB/85pXB7fILRKHvqH7N1ye0H4sjedbli//eGbT5dTKWs
01PAnchQXPaQxp9LlW13+epLpo27+y4cXIBv5AST1wc7mOybvd5PG0Ji8/gTufh+
Uv0X5Ssbe8sjHh6vDlAfNtIonVAOGWChYHtVCaVyieYY8SyY2q7DZif/zHpt6/hN
vhPrZN1vrDBzTOUBYD0L8I7CsqXnGPQC+/mEChOBAIQvpFC5ukv0dZqxddEEd+1s
tUapQs+cNWmuajknvU7wUczQqDP6v7K6T3zQrMoGguP7Hj2u8aWqochCOKNnvAMN
K4I5u0u3jsIYLs1RO1et21ivzuLy8PRz4UfWqCFkWuDqcw2npd6vs941Hdv7vpEo
fXdbDv/8O3NC872LIzk8jQ1ieuPMBPsNVokmDZKFtMLgQdxmF6ElNgdR0oRZdc19
sxHZUGm6xatKEWhMnEEyYGS8uQk+fLDVTsKT4T1PSS+kDgvEEJVbPvCsS0yCx3Q0
2tUQs+RSyt02ekm96f6PeBsV2k1nzuEWZEQq5C7oZPVS9H4+dYKIuZq01410LODL
SQHeNSb9ex25G0Wqcj1SyAytfzloSMLawApPwL9US2fiCzDHO6anZ8s43tLcPe9d
+4VZgQsbhA8v0WCQb+hBqJMKST7wh7MZ2V9kB8Q41GYCwsqlKreD3O/GDB2RGIe3
ckNFRXFwhNu2yz5A/zH7MqzhEhdBdHISvqDcHzDmlIFCdMFp+jv0pccmyYC6ISwE
Wj2kP/OSITTPmbIbvZeel8Pelwte1zXHqvRw0ZJ2CxtOZLmW7Dql/c1SPSdFiYbD
EvFBO+YGuCgUZ3sUZt1+qSYtCqNXXxOpFQGqp0DsRRnjEPSzrJYCmSRhEfFhqnQ6
4vU4AoNnp3mtEfr8o0atjE/W8yXrfhQRxrI0aaUPTVcSMP4IFQAZ+5JJWBBqJDqZ
/ek2B7VM7XaOkipjsxoFG89caber6lpj6jPgAjpx5I6aZDmvRDnRbayPUALQKCyQ
NoFKtfzWbKI9cqjFDPFLwrTJTePHOM/77AcsEpTOW8yXJYwOmIgB1OkPBo0DXdml
buC6OXmM9ESeBAUfgLNSVbILI9o9jVxWKh3BQU/4WkhwScx3UHwVwLlR7sveZe6x
yfX/o5FIhGOBX0ihbRKzyutsK7C+kWAJsDaGiNC2enZwu3w8SmFe7Y90DOM28qBz
afsC9VqpU10zHE66HcBuCqAcb8iDBL5AyWH+ZrihPqG2MCviqJR/8g0747d/g3Bb
j+5JiwurVlSwQqwk2XFUurkAAtHDXAN/JS9Pqgp28e42y+PNaZaJBXyY+JkXG5qq
GiK54Gmf6ZYpquv8y7dV8Rz6Ls/D+c0BWWKEUFKY0gYOyYaZ1Bpz8LPQ9ohlDevE
9Qpxr6NNvysdXAz/EfPuGteFzUO8310CXGMIzvDgleLk01ZsJOGeBa+DtepwuDm1
1BN1hrrvcYPm+HqbqKCIp8YV8tKifV9B/u/SENMvR9kzfwbkv/LP1zhuj4TqMZBF
sUdTn/jYD9t8UvJBefdv7KUekHDEHZn9q1hdTW2WLDarGalnzwdSMbtcuXjwZ0Os
Cg34kOsK7HUPFuSwcXd658ft5luyQEx8ZaK0pfJcBK3DdSP+mKfTdcLz5wbYlTGr
aM6J9lultb6TVsN3SX2c68BBGYAOArREfqNIIyltnt1FGkYGBeQFXxDLwiNslutz
7fPq1eoOx2ploSJxx6n76LBE7thW4rm6vUBZn2/nlVxEr7UxmI1CpmxKSBgOfeE+
ZG3u/eGcuacmpCQUnXkIXKs6dywOhXw+mRhoNuG8pfptNQv0KP/xwFoanTUyokgK
mZCT5SwRoNUuE83OZ+WUylD95WvgVKCX43kqX5WRo/DJspGUoDOxh2j689xBBEHl
cd4VKLvYXmrAPcu+m76QoQ0D635YFR4tHUkX89uOhudWvxYJ+rKmxdGVE67jRd0g
aSl/LwXIH//340PlbT8yfOFtGoNdZCVtsdxSihq4Gl5CSbA67yDF5aoMQ7FfdHbg
r6B8pHFPjaU8IzGP9srX4skGQrLa1OccQ7ai2cAJ7AEvHJeNJjsyzSjfjPyIEyFB
63TxWaJVCc7f0iu0EzNuRKthWAMs7v9oWGiLvPvhbx0bYT1y1s4gf0iLoBHjb6Bm
grWwlSx5UDvHep3a+3l2k9/UdLSqeeiAO/rCq/BNmyfqBJGWvVS48We7LF6RTbRm
Jyoo0mtyWPYvfTB5cE0QVhM4wcbYQpTPENEBe/2kSTCq/kFSJwe/cmxx1cL3H+0x
pK2PxVk2IdF+fRLk807jIQIEAreYpzul96RtKvYSy7UHpPujB2kRGotGIAY5SSAC
//9J46T8MRrJCeLqW7CKafvMcDA89PBC10flO85TLqZ19VPk2pG/HFZAdVfKDTji
LONjD3N/toJbISf8Cb1E8pICgGUfnoIS1NwsUUdqLv3G1nB3bGLA+dvCW4Z9nAQT
NaxXZxoWqWvmxVmeSyvz5NJERR4ZbyOXP+2/ZZhW92+r+Xv2XFAALtBaGxrHZegm
f6Yfch3WRa2TFAg4vfBWk2eFKZGCuETf9cV/rcOCatPDxsXS6/7oZCD5a5spFybX
TLpoX9w1mQ5kFTfyKj9VYPpAJ0x2oFOWzpGUHZvYdJIvk/g9nVQrvQSZ30ICktw6
wyWMGdTo7Zt6l12fHpSvHzAybn2qUXcXbwkn83AhIXUBf19k1zD0jo9tXKWDjX9I
HvlIsZZcD8CESBv2zuLz+4MoTwaVrxPpOH/bapGUjX+IJNvXvyeAES5LGopOgn/p
akEYeZSFKZ0lVVFWmYaljLT6mnPr+X7V81IocEWlgv9Z5e7469K6fhr1bQR55Gaw
deDQqgxnanOKuWhx20JwS7eEpK8jpvotCNEs+UCE3S4IDE1jUzkDzdnb7TfKIJYX
5rS4aBgnxtDDtn8+lfstbA9mktEWkwvc822LCK+JhcNS3pVPwTijt0NI78MtF66Y
xLAg3p1GsImOsgy7FD8K1JGAt85RFTWub3NMzG9tCBXNqju2QY76oDKD5szx4bvW
Ip9YpEOKzmPqVTiBJy9cUlpWyC1j6TpN6z/j1YfALMz3volb8LTYtUFIzooCK8I1
OzY61v+ebhYmMZAijq1F7zT0FK7Jlduju/KOeeXR+E4DBXnXNv/DF3CNjik/qSbv
8sp+TOsvHABYFd4/0WP4NTXYX9sKs2e1LSNYIL2hQIBcAVl4dov0Il5jrqGdEGWf
p3yqzEP7VHKgAXGkKa7PhlQmO8JpruvUwEYfMWUyTZ43g0o3YeSi7+d894fAzMDt
erGMboJpCUptQhfQLplEbMIyTAxgruPULARAsKidztRVxKuWP1gg8SCBbr70ISzE
lwW4CVeMfZFQnWtB683oFghjn6keKKyCJUiqcVRm/ChvRdaqI24f6lx/0WKylGze
R9RN5pwSGlUyMNkm2BMpTl79vnV8wMdlrgZg4YmEbqitV7SS0QWpH9A5zsulJ5xl
MxfHGuIabniCrwta6ndJsxQ86ZknzjoY1TRAxyFk6fmMlgg9rA27I+P7TfnpBBtu
fOWiQPTHFfJAhr/qvsuE80Ua5cN18eDku0rcfr+5gv7fAbE+0VqvDCNL4CTByT+q
V2ARwDf2iAZH+Bq9V4HLdiKsIXThZipXfFoVVX9c4fZlrQD6Q29Lu8NNZV//w511
3gcAfvnGnlMJPZ4AzyHfv8ilN+D2CfewLFfC63p8bcSwReinNyIvV0T/Z+fo5+e9
rBVr8ZMQq458Fvx4PgzYcPw0cQQ3Ul5MBNAm/DegIUma855R1pdZvsJDE7AmsbQV
hdq5+uwzM3tARMp1BmcshPxBHBtUBB2petZAfoo04XUYbNdIMYDENEPcqxQqbOnD
rJIuj5GUNs2SGNPxk1EWcgG7iXs+bhTgvi9LVkEfNoibDzZPXMWOeKeH2Q+wq7SD
Qm88Geog+4crBr+aSLkfVoskSr+Rc2jQtZ7FRQZgP31RDoJHMnMXFuz7KNyFiPVW
S2q8vaG2MDCiRHhkFIhbgHop8iR82Us67nr0ejkIJpJ0lZp4cShrSvZsR0dMircr
9nFaNN1IRC0nSDwf7LQhi4lIPx9qewrV34sV2y6i/M//LHaZXk0MLqUDzEZMGa9e
VOR4Bwps7WIYEqwhqJjSqx4Wh5vP1sqLFt8Nas/CTiuULX3HVscN9R+34y7szVCq
FYCc46Z3en3sT1NSnv/T7RFPKNR6liD0YW9jhg9Zhtc3XXdPaB6uELJibCJYLNyI
3ZD1RK6AyLxPUBlN6vj4veDZs69Re5FNbau1xXqo1Ezi/JHMzsnACh9TnLUQgrjQ
dNsTlgUpFhk1B5LaOyTU+8iGzj7CuVkQuQr07sPAjbS8hyZ0UGKu0HHVcrZaF1LM
2yfo27I9whfMiQ/PE/4Phw3tL/L+hn9nylDnW0huiNFD1TTotqhBPYf0AfPgZetn
EMjOCIdkv9oMZ/SM6Kmi2+V1XqUF/bz8NAekU4VbDgG+lc1sbbi8sBbxf/mlq6Xr
xAaBKl+Wmo8SNpJsVFN46Df4YA8bzw2SgcLt0STnudABPuCqEtycDlEvUy/hVDo0
Hwr/zVWNC3rp7oQc3vzfUcEkCRpdDG9q7kX4CSiyaJU8MzrlWLoWBiBpZzPTul/p
BFKAh+i7aAgGFHOlsKcL01YCyrjpRtm7to22Rg9K1hW9UtU1SljPKjfYO/E3qKQT
4VDZmbVWU6qI/ii/MXgiGDEHpMtT9rbk+xl671JFuZevEuG5b7/UTxLYxD0DHVum
vVHMiilbbuHsj+sZs3HAKzBfReD7ZESxTwUN2EPKVlhMVN6hJk/cYXeLQOABN/Hc
kJCLSn81ZfQNMZidD+fj0uBExUXNojW90bSxZtzhAauxF4iuojRBQm8+FhXwOCfP
+OL1bKn9rjMiRVMahHWH9qjTmOzWpKdwl2Xu6ZafUudsLg3D9t86AYXk4bzNWStR
x/Z60ZP7t0bB32U6LiWaezV+fV8QdikdnTpRllGGlqki5tdwd1PGWsZ99ga/DcNA
hXaRZq2UfeCgcETk4I6hJTvKQnBvvBhjjdbLZ+IOuvM6zQhk3EXRWEhMC8vE7+1z
pjM46ZWXW3g0E52DUAqoupfktQHWG8lgjNIPWRI81TvIhPnKkcr5WdaUwe4ZnRYq
3fS+85W64hxCH+4GEe5qNzCUq6d5D59eenrPsY/xKum0To9E5Wf8YibbSIren1X1
+HuP80NoTiN/jMZBbGpkI3zmIYLPkUx0MgtCDQ+pDUCZg/cBII7TQC10fT/jYTJD
TaQmUUG9NclFqWR3jCTEt7R7TpYFKXsS7T2BWoPj5hOe0e99ykIYDnfmjQnSwJfb
P7H9C/VQUbMcrpQ1BLVtM46MGGt5SymNBgg/0VbvacHTvOsfyh4ceo6+VASiypkX
Uo7oN/wEWI4pAVPL924brF9d/U59Qp8NPiqe2LHT+AYnUZaG/CKCZiU/cwLg3nf7
SaYgeHMVCEU8vH5A1a8YcEVWdy2Q9eCS3Grq9/iSLIzknVt9VBVsTpmD/25AZZeG
P1gtdAOedptsqfUcI/qDEgBGHBWlRz/FcygZCJ4P4Fepi8TexUNs+LeReA8QjHD3
pR53RKp9QNaax9U+iJ6H0mAvuUO24eYO805KpV884QeI1waTfXW5YCeUwbGSCNFY
To5y25MDtZW3kFHdXmtYzXITPPWTPbeEeaujFIW87gp3YDsffbdeZHoLpyD09hFI
V2PuEL9PdxG8CwDv1aQbug7aiybLyanVkwEakGT0VHHvae2WuBd1VitPyAph9Gd2
lMNq/CjOKTZCeGROrR0rfNC66V3guAoLd6lgbrotMUpp3SDz2oWhuVTel2FWzYES
NqhDYcWDT2tHowuTO6qatvipeGlhtor50NHvfdK71JkzK2yzxwm5kAI0qId4h1BC
Ac9BEwnN59EJLjx0qsxttC10CNXMDfUESLxyv2pq6F/0HUhR9os/klhNSdjpXnQy
0atQrxJ1AgFuBYbFBnVgySF5ilnofGoa1kKolEKlPV+ui7L8nXlPsyiHjqFzOEfr
V3GKFhbdOHOeRAe6oSHFynCNYCuWPnNfS3HUJ/z/3ykCoFGQ5CAAmf9yh3/KlSFU
A+OF07gSubxvs9ny8B2DrZprMeyobnJ4rQmZo40YIvwBmjSSoU9qM6ObVSDwAfb3
3e+lJE1sFBYmQ2WlqZCe2c9JLuK6uU56MJ9lyGpFhHiiqzJG+l79Y3MQ20U+/mY1
tPFlmNvnfeucbrLxRyH02PNoLaL85WGfxUjXB8alE0xpAtK+aXPELbjjfzeCKa2g
Z02vxXTwl68Uq9TtF62+/rLglX9Tmfkee0Pb5Cm5gsnkEfPouuOlNqxoBpQ6oVB/
LRDyo1CV46aQpp2iUI6E7gXxDILE90jhsQyeJF7HiDriuNdS4nDtPST4R7qY1taV
OH+2AhdzJN6LhjeVfwgcE1cRneLLPv09BKJc+6hhZlsT0gY7nA8ilDUPNxHNyo0B
4qj/sinKTVY07IV7bQTF+2+sAWznwwhwrm1gwXfuQhF0zyJXP6yzaUN9p2nSX6np
k0euSnC737u4tbgV8VnceXxtQwFDx8wChW9B/bmR7EmB/b9ZAPnP2Ssdt5iF+Ohz
7miRk121F/1E0hY6RzTm4WeOgsWcIFpEwlb9XKBPTcaIBegMNPLsCr+nIPgGj1PZ
/UZupcSh+BbFYz32GdU30Ou2qRp4ect0/8ZwMaSLIlnFqMwisZ/2pSEtEiL7Sbs4
2+dA7C32wYw3leQke8Cnvql1RQV3lck0Mu1pCiyDJLW51Txkb7hmTnYlRY+56mA3
NA3uWAEQ1a/vuQ8S1Zc0LaqddfHt82hYT94Xy8utI+ltaK2eEvN2NXLFVkFS0Zph
3GZ45Y7pykVnYDqhjIayewHBDPby0M1R6SLR/RosaCdJ4P+7nxN1l3MMn99gTniC
42MpH+7mIFpH6BT1eR6FcJvCERTrHdCqd3FsN9/vGct/Ks2yLnAD0wJu53eP3izv
Z8MUlNFovlmMOP5cjarB9t4H5k+wQs7hRzQCNwzyeSyebdZxNhlePXFWHjh929OL
btAcQOF8qmb5TJqBcayIQVGgIJ0O6pDEgm2PeAFA/Y5CkVAqmRYoczv6TMSA8ekx
yQwgl+7C8pCF8stTkpaBD14g34vwzJqEaxYbatjVQlu6J532h+NUZDrb2MI6pOeF
0Vyf55Ps3Rak+9WeK0COlJqCmlsZ+1JJtmOSUDlsDEz3EcB5ARoWZrMcxcWntOd+
64jcbLk1PlJhtlkGdZF5tFnt04R7cqYguOtYAMaD5ZnxcozzFpe3fzDG/ECr0fMc
9CwvjBv48yMgUutK1oM5RbL2YqAM4Jm3sCRz7p6/ruWygI33Ux4uNEj6TzmihqHg
3YHl/zZJhh91BCPOBkxFDUqj0E5f0l96jjpgu6BAzx+DTyezPMhZEeQOeg/KfZEV
L8nZIu/8cpfpuYpSa33pP8nkY2TMMgs0/eOYkYzt14Kt98GLK9T9uL+LlkG7ehO9
MWwg6i7KNow/5bZ+kp1s39NKShDKdkn44EmYgF68l0gotk/zbrAm/fXLQtMDU2I6
LRqmzsgjIcnls3mnRBOTTW6n38tgXmlpLJG+YKQPjenb8ENKIrfFPtV1zUkXzLQ2
iEPM3cgekd3hZlOeDOns5Bb8Pu6t8HUC010yLCRIf2kl401u4sBsBwr8sg3ZHu9d
50qDk+fjevwHCRAb8MkgVNXWfHG34qQpgk9e3BbGaRu+PsqKS7YlNf19xPYpCNh6
alsBhG8lu952/SAa2HQDem1T78h4+lKe85Zz691o4h9LHkS4Go5k2Zw81GtZLx1W
/xli9qt58KQNxNRUmjZXQBvbGHs0wQBHNcC9YZzBHxBIf1MUlTTrCpoRqNLXH8H+
2PzxRO1HmIP+7V/bJ2ghHcVzwMiX3XyxdSoG7ZAmZPzBnflb6RMmmckJTnbCGEgU
twfQ+25fg7OCtJflhAHnlvMPjcHFf19ojFoRgcM/guJXDKXdVN7WAAsRwMn+yTQX
ta8NRYBUyg+Y5RRVtZxEgmhRl2uIFAQ0u8vTY5Z9R4ULrNvv479BaLq8ylYf+t6W
CoELhjy7ZawIlu2HBeelVuefM7F2AvnjnzeW0YiHYqFZjm88+015On2I6lMH43hz
+3kwUWkUwwOOprLjiwPJ4aD/r5Z4eAxb8N2FMbSiWP+hW+KnsAFhsLtW5ZcBUCAa
/oX1ZeRgTB0BGURnclIswC2ApSAuZhyU1C7I5XVtzIAzALu4VFwVuG+xvph8XzO5
M6i0e6XewkKAex8MeDFwNbICCV+yaEW5wKZmKOEbRvBHiP643YsztoYw/4xM5xBp
+JET3bsB/x+TCVuUZJCn/3xHO+5qcVPpsDr79RSN6h+PD9qqOn2LhushaH8nL3Sw
mVdoLzetEZ4q33zQq4hLVEeFQWvvqvc8SZLdYZMUReA0ocnOZOZd1UX93b5E1sHg
WLJkprFiDo8+i3rIYLBDwuuerbae+pYGG+pIhUnPFD1w6HxdyFWuzTbsg+m2K6i6
RUiGVIq53S4eFm2sEa3da8ILbd5ydByojvbHW5Tlmjp6iF7E0gkVvNnccVngeXr/
Y8j/oDfmado+0gs5C3Eym3nvaWNhYR0eYu5/HpcMnudoXDL0lnw81j3KIYLAZ87d
Gfj4H+SOwE1KbcCCjJ705ggxFBh+Qj4oUK8cxuLEW06JePeqW3aYv3S2FSopKcp8
hgSmMB5hAey9nOqN0T4b8AhvCw2qSsAbWMhK6FMISDqp0wySPSd4RpLUg731mCXj
dCCvGN0fvVG9yVj3CxHXgEUsQxbqZ71d/DaN+eMj7zfe87f7jr2UX7GEjIQpkXc/
J09oewzRLQRo0RE4tFyeOBrNq1tGOJ0tbi+VwlB3EobOIpkTLpL9rjQUDzzBGDBm
jlD7/nAunP/UJajk9jjsO71djmUhWh/4WAjkQ8ycyTxxd1nxqrxeqh9zuK2dOva2
lAFOtNOjY9MzqpV1wVjheagM+eszx4uO7yF+5Zc4/AnqscGRi5zCfWvX7SbRaMlU
82ZVLP/FwxlsghehZpFARaTOd/0/VfxPFP/JTHrW8vPNn0IPdwR71SZS9BZee3Oq
wGBxf02/zd/flaJ8tj3F20ijz9NIrFuvTfIEwj0B//+YEZGQzIhRA3E3CAq5jqYp
Rwsy4XIq2+rN73lLIp1vPjSLlsUcGRuGnJoxGsUmHNVjMJuDj3lr1cJl65AzF338
/yTGHk1lnh6elA/T8bYNcwIbqpTpMyiwHs2+e51HRVVnNciIhlj/1/U9YUdTOekE
Gsds9Sw7pBG7lu483JY9koOBHjUrY4e1u2D8GUukTS/FElN49FtWbuOpEe8RRfEu
CO8c4nMh9uei09u6RbsasHAdMWRhIUrxi4QJF8WqoFNOsZWQLg+Z4htayPu15IOv
ER16bKbq7AAcFrhvcD4ep1Tft+nwX/H/U1U7N8KVRLr0vSoUeBQfdHdJ2raswEs7
+T5qKfaatPAWKMThEccLP4xIfgxh+bHC3N/zDXi6nQbX3WZqTpoEr715qxFoMwC/
pPSXmERWKsgTnZBDAp3jgXmOJaR+7HgBPLbXIU9BbMJOLoSoKqr4vovFpPwPdzFz
KlsXmokzExxptEW8y6xQOBEIcKK/7mq6IN+eUEDcTYS+xfcmQODHAlzjZaqJ46kd
UXd9LfXo/Ux1TRjOoxlAuIPdqlXhbnjBtD294ntbeB+JonWhNsaf/7qUIWM2efDS
qcVG0vG5jpMSSk4UBiboVjR4E0TJumE8WEz3yyfmpxDUZV8q0KaLrhXk8RIbcfGB
3Cb9MjBnRreWlRmJmqG3N7wppZhMhOj0TOBdZVWfGFC5nqxpDxrS2XXZUPOBQZkt
oFlx8WAo2/bhuubetse+3TEo6B3iCQ+hjwu0scCZmaOKUXYRsSzwiyd0HYiRt/cf
qgQ0w9U/WXLwMVw67I0otOw5b5tsM8gacZTx+AEaBhnydFHkln0V7eLNPyRAudj/
sV1CEmPZfL/RVXV2WnIN/GTlbd9aIPDt+vLwcpXDdVU+1Y1jzTty5geVbnZivcHV
iowpP/KFNY0H5yQhOtVpUryAFm8PKfpV/tADNDmhVlWKs0lt32v/1/ZZXd7TntjF
JzusDLcoN5bRoCUpDbCaIRrQ3ofJEL5I/52rcNmCc+Sig/r6OaxcfyUEHCMII4YW
Xk7XofCWZHOS+2ZZ+ntCgm9MjW0UQmL0h5RB5xy/W/nF9NXWJUzczr2Xm5EW+Fye
4LXnbbvEYuBlZmUAGg2+yql83EzlcLfpZ6m/fkYmiQxTgKtSMs8czjAoxkcVJNsJ
dE8FmvP3AT3hqK5RcyOsvucFjBc2xuDjfv8/zGWLbmwK0a/6FRSEObq0o9xod8WY
clT1JLv1CUWHk+O3qN/z5hC/li1w5FdcOC7zXWqF/MqXtUB7GxJZ1rodaYmGKOOw
HDIPQeP8wI3ZA1KEggaO1rNJO5EG3QXgmjf3xUmDhwPm2dKSeLrt5PJwXPy8w9DV
/AjIwQBjNAi5jEc7VXZ3WV3xc9XYv+drTketijUEKURDdishDwugBbfGizx0+uyl
d7s9mLuEuuBj5CXPvd/4M8+td+p/EPckwx5nVbHN35rZf68Hhh9xtWPSaq+R9IMj
928qMejjJDXPd/rgYsbdGUsYzSKuijygjVkFOX0og4U3Hd21Oi99ttfp7g+1jcVo
36yXLMYOeEoGcSZm8A8QmlVHdz7QSPSWwI3pljCq5He6xg8/y/dcCQwTnbvKd+3y
tIXcMqVfHT+mrk92/cDLDgzUbpSTAroj3lghCCheD5B8FYKtM4jKWY2MgW5JkMoU
XHKqo/6DRVOdBVqln19wqC7Hh0kgv1Iuf0F0msmUGntbzj/To4IVkuXiJ3p1+ARR
QgavGK04TtP+S5jrLgeyiOHil5tSzYyEDKYfzEeQ2dV88I8caP4h6RZWzN8dDY1X
xFl1vdfftrb4C97+Cg3oBIr7TZeeoPeoKthacp2E7qFKjp8tERGExG379Llzs58X
2x3X2vDRN/w7nvdGYYm+Kcr38EuP9IHLeWUFHYCmwc1WZkqQv5m4yWvM+3uTDSkQ
GuJBX7LBdXsfT9ESGgr//NeW3rJmPZB8tXzTDMNJI6W2z0w08bko1MjXU6GOGs0b
KWylFRiTGfxzon5qe3JF5LcNlaEug284Oa7xirb7pN4+1nzzWkXeCKBe0907QOL8
J8v/TDNpgzgsS1n4zm6tRIPAh4/2yIBNNhvwRX0mptmb1qHF6xbwwY94x3mIVJfQ
BxWwXpMoU31N2VNoJp2av3uzzhhrIcRHyZIi5fcw0o5edB8xuaNXlXC3mtQtc/Qy
Pcc6fwACBxeLdwWi4Pk32JRE89Ttk+40hqsNpL6LaM6ymw5oDdDy+4CuV3vZsYBG
C0yvpqdesgETxBAwOFO0sPIa1nz99l50sYvJgL73d66Rq8EQB+9q84ZPOlsQrqMU
ldM1Z9/0neixVqnwF6iYqW9QX/No5slfwT4OikPtlR9ZXIOdqan4WLn5tDfTwV3C
2coABf4tw8qXFzm+J2YsYf6FJpwsiHvd6rLii2sjToA/dk9tU6JfwbD6cgbhG/9L
SS0OhD64IyIq27XAK2oym4n25LMh8L4XWE1QFN8926iAtoZ1mNfvAOcg3GDOFfII
zR/ZEc2vAKB+HL3GMhoj/fxJUrMQYYw3mexQx5q2KOpkfm907624CAiUV7OnLBc3
9X3hzfrKt+LuInWZkftn0tXaW9R/gifxC2oWvAEpbe8Imr9bARbrRKLe4TKmvReD
LvtAyUlmVEaR776O1SMLeeN4GBPV+YLfceE2fSLCHzpLbU8nrnYpIwMzRt6Q5uN6
ypozbaDKsvKi7Uu9d0RZnrqzPWwuYey0jqShKMmVYt4DGb9LOP/TuDsWPIM9kzm4
FzfF1Y1tSg9lLAUblBYJz7yVCzzOzs48PnRfzdYCpkvn06OgN28VA/0cP3SItgIs
OT0oQhM1Arlyb77z7IEN/wnb1ESRxf49PYY5R78BWI3t1gRP2EuMWF5QFb2HumYL
GJjsbCRAAQi5uzRsVWI32Ofw17M/FnJEf1j11EnJh0SJnqG8JsytvQR6gHTqhWf2
qgaV0kJe7SqzmsfgoP3tVnDQuv3evIqQUoYjjqpdF+A1itKHf5i70RLfbshsfk/n
rdT+ZtDVLXYgKTWf8aQSKlzGmreBQEhzhak2dZCPQ7HwSsBA32Y4D2zkTy885rsf
Jm5BnQ535J+8ogpPrf6BGsRCsL226Z3Kwp9zWfkQMxFmAN5V0K9EayDI9ze+2tiW
T+4RbrOQ83TMJfq/5Agog2cG7N7x/GGF2e4CfzNpak2gcGfkquiudznvX56RAGZI
j/xnGIS7lBi9X42/rsugX54Cbnoe1H89RgP/rEM1+KJVVgLOJB6eVTb7gOud9C5K
q9XH/5L6zKt9sIAfFNIQQ7/v9RGd6TZT1lXMvMrN9vGrMIMnQ6QK8Tw1tI1zzxyC
k+qRQLCGqG864JL/g3xJHiwsazQQRx7mzKVwyONzPV29SateBIf0sYIf1GKaLoOM
I2xQokyjASiMuF0M5Ywdp4C2L6utIjZlYeDRiX1Umexg3dDUp/WqhywIkdf4Hv6F
eZyyxGZ1DO9Om2PgFKDZG0bhToaxx3euEyXrWJQ7oUaBB3BbZ7W2pNI4Ca5OPSDY
nOTw/3VssZw2PtDy02iuURUxIiuI3WzNHH3iCNBzQBp+UUKXSliGhyqJ29aHPATl
+/TewPcqMdXf+OVtp5CAvPt9WKhYxs56E6RT7Od8RIJ2hRpvnRqDaatybusxR8CC
4KlTexoVCjdUKPNoPywJ0f6gn8e8KslCp3j2MlD6UkzN1ac1Rb5i63dggxMnqQ8k
WmCSyssLPMJjN3o9TD5KO4A1tpN5B0G1OWTvIuaCAhDzdB1d9/TW9PsEp9Rh8vCb
KHgwMbwOHcqNhg/3xn/bneGfa3CBfsHulsQsafGZc4/vvyp+L+TNEoGePkwhCP+c
xPl4Q/1kOLRp6cSt6GYRzXGtvLXJweugUvrlkzETG1OEwZgEdNCzkzxaHd602MBr
sWzMIUAT6mlGRXaa/b/tOBrllRHQIZMd+C2srEaqm4jPAOQ5S3rHShLEe9MmqiTW
Tn3x+GI3uJVtuH5Xu9tphuAvoqfNGS2WN1P7DiNdFGrjOxI18Nl4b8oxJyrGI8V1
8dXvWd3uoS5e/ahOztxfjFHCrgifc/KeXEw6SaC9qKSpKjTQJiaA8cWEDxT6w0lF
ph+VQVe7JfzDSIJdVEbxKOgIezoiQ0wFKk/l1frCqdDsKvErXlxs+sk4h+10EOMK
COOi2wbKA+0qxxvObWt7Paum06l04wJTsMpjd/X3Hl8or3yjeXB8X3wSwa9Tso6Y
Vh0jsbhbLSn7kMvWo3vNbIk4zwtvW0+xn9/jyOfkEF8UQTQ3Bal4eDDEusb5jrFO
WoObacGcEQVK+X0w54QK+bvqFzQ2tUoqZz/9rbgdnOsYwtmf9vWOroDDixLrCnbh
0oa+gEwi7EPP1W1JPosXzHuEkr08BTuNXcMTYM/P9ZAtDBUO5n5f9/JORH8OIQ+d
4ddJPTq1fKU8Otm7bjNuS4tm7R3Z+jewC9A0ONi6AwCo87zjb7fk37KAu0qThKIy
KDB4Th14dO4Dw2RH/Ze5ClevEpWEtbxiU772RhrrQ6v/AX00tQ2u2PE6SaKjctXw
gN9Ow69MM5mGC6h+f4DCzewOs1v1AegIpj4Imver2agF+eCzUvZtDOdPi2b5XRnu
kT2CYL/9mosGAnhJRaD0BC4CvDwwF7NW1sJVDqRXKw06IYu3fN8xW1dPfCCQLOZO
fRR4uKYhxKZiIuhFigQzYo/N3xwQhPqJhhjgfu6/XNsXh26W+H2rAViNASttcOZI
I99j1ecNTmlTChAmFR2rc1EEFHMnUBsWsiDUfJkUEqpTvIrJZ6MrxRpwJ0tQu1A/
VpPL3BZySs85/TdEblw8BnS3No9hyaUNFbUedZCxawzaFiiFx5YkoPxZky2F2k7N
QbOGGqFAYvyko8rOuvPL5Zsf2CtevHs/SvGNVGZPIFq5I44GyV/r7YwAA+BCEJYp
IboQxLc9DoCSuoT043FvfromoagJCBNQ+62JHHvcqTfena1u10ba4CptxNIjKrWg
sph50/XWV4ewtqgkc2bcutvF9pJNad+HryC3kubrcrGdP/4XIjIuyqeVphs81+wG
qy4uh1FotokNXEPehCBe+zy4/m9ueePNV0RzyfUjM2PgHaA8/CuDyXCkI4ve2li4
334ER3VfiYoXS9bnflxzFURXz2dhbPz0CQNWYkJd3avM+OZZFUYoYezmcMUqGCvw
eTF0hyam+Du+ozEv4GJ7NQc+rpljKyxAUFbD13HUz635Do9TyaqbLlrCKtDpHQ17
6xP25wQLSyDHphqS4GwCwMP9vRc4JLH/qcTAaAozagu3izAHkYNEeUbAtQG3ybZj
CEX6xejlWa0AAvtN+mCaXovXOgZ348c65Hj9g90ZJdLgxMbgFeejk6nCJFigloDq
yjKF8umI7h2frBO5MwDXpt7OzeEjSKEEdn/5hzVrqVSxmm5M/weBSAtV1RJSd4Ea
mHcvZHs3q30hKblrjQAOI72ER+yTbFFTX88rwf6qI8eBJ5k4yfr/Op9Asio/WBVA
x2Nq+lt1Qjx4WxPf5hp6Bi4atdlVf4nEB8OzgAlPIzIO8D2SCMRhNrvNEu6Ixngu
RzlZGGLzoMWcJqrFoHEpN8PKwHhrzmzHZoabxn+gEK3tvSviy4cjWfGdd6dmbNhR
ax98FAOhIU8qiXL98qf3tMVD4WvvMa5/b6M1OBcffUdDfmlPwbUlKgoCWncgJEof
iqXzzZFYqJNJO4bQiBaweXXQwCWHR+JR40Q53L5rjDPr2M0Xa4LvYnEiSihV99AR
+ztO1xzopIX807WKHYRndbVfSaD6XQ3CnSwAK2eHkXAfHs7sbIxMTuzBaC/vZbQb
nEPva4sVtBf0ggyjAAJ+uqqv0UhxIzpxlBUMi0kpOLcl/5P1a0jsQ2apARP2vqKJ
O4kKdvcR06MHTesq/72LT7cNPpgr0GY5HWbKy80mLylS351sfCTTuk1p+Y/D49wR
nGLrrb+foYb44Kls98juP+pQr7PfhIvtS1igYlB3X4CgIbGDmiM4dB1QQQLXDzub
EtDzbDnWtqZ5upQrJ8W3YvuY2uw5MmGpzzRwJMoE4soZoskPNA4F0xyvhBmnyRq2
JJwXaG3LyaDnCHKwYbuq1YZRbsba3qHNKLGJOFy6HHaTkxn5DjVFvvRJGPmBZsK3
0YS2gSTwuMbSLMYkB4Yif3MTErToLc/LATNgfpk+4vDQRYnX0e6h7E621JLfY1G+
pzi1oGrPMn32n4Bds4gniLpdgKQu/YxBJD+hf7dqY/exhom9Nl9o9rjk+lJKNXHh
Du3NfSb46JDq6r2Qolkek2J9J+LGF2yoDe1qbP0Z3XuTfufYsKH33I8ikbiUEim3
DcoQ2PFOPFl1+6G7pVVK9P4OQOGdBhcJ/oazLRxaIHGPATxlDSypF4NlFhr2KVi+
BVVssPjKKtKxI+Jm0KseeeW6yQ6eNFspR85vQ3C6INgh7t3Bb8EMiVPyWmNPyZLg
HtbM9xicRpYZYjkcdqSYVg7FiMspKzDvwM96KBLqRdYjz6GucxPoFQQflWdkfv0Z
cCeXWqI0aGlYnEkFZeUoiR0IBzHe0AqqDbXBcDrsFR9zcHPqZjz8r/Hbj12kh/Bl
W6HYcGjCXrfaK4YdvOkZohVof5l3We2TTDm+2fJBPwMR3YH7U9SDHavEnpkqXFwv
pMRIh/6ou9HaHrn6TLekq1F7FU/MGY37CFY9xp7wYwcbJUJfNXKrPZWz2W8onVy0
UwrKqPKzdhO53ori9gkVCN237AK54Y8PiQaMzm2gux7iC9DbfOsL4etv0KZFYJnw
GW7zhZfxjisE+dyS/DPFnx1f/ckWzBb7jUSEAb2pR+zdtumgko/GXM1ob1Y+L6Jn
hkKgRmBXQ8KD/4tkW2OFkyueqz2jyGd479JPmMPa8tZSVdAgJMjGPX+S549wAWbt
2QZF+YK54XHz/7KH/zoqUxhHKDdMDNidLSZnG/TIJs7+MT3bHrdxEbcK/0oo6cqf
+L2ukkOd47pRz7NNM1FsMeNFZqpOmiyD+ywj0p+sqy3AC1Wm0eiy/PfabGqWEK04
AdGQMiJJ8tGEIvdrth00d9SzhlK2QhqDurAGVhM0GIThNe0KzOB6HnegvAD7YJsT
duO9yKVGvVLLLYxOnoeFgjHg8J+qJiedsq16Pmr7HAGi0rTd1SCC5kzlGWtMzVnl
9Ro3E6UII3AEf1GsXAOVK9TDD0HkBNvhwqseMd6MyruUc8k2Ma1Zl48u621QPj03
+uZ+MURw08TMgKwnnNZP0tNah7h7QMwEeilCLV3m7AZsu6gdqIQp03b3gsdoTrea
B5xc9/djvoKEviaudLVM2uMmt5IJGElxY2p4zAiPlegszrS+iOcI4v0pwzD5PpQL
9TGQhhx3K48F9tXgDN7YPzV/HQ74hW1Hr+38wpBgLzyUTjPKanWWWvBB4tG6XoDt
KkuiY9NR1kn1SZ/UI4dSjDNMuXBFn8A4JP5QqXkiUBt81UeZY36naMevndxdHW1C
meajj7/6Zpk0jZ482uy6YzW9e5SuUD3viJwGiAmNat62gFLvn7iuy5HUIEFzejcV
BAfP6SHIutL8GK7I3JnTeqgTZ7WHf8k9YtmTEXpy8M5qCoTECYsubkFx87y0ZcfC
Q2ckhjXu0Cnu8KGhv+b1xLs9BBMhxaQxCbnAoKUJZ35aNSX9w+b6Vhfr5CyH75UY
9Iav95Rek7MgALGVupQKM3EJAKO4+0ppcQsLewAMj+SVjGlhiubF/1GR+fbzr3Wl
yVhwPQrutGehFJRzwGxOH9NpI8Tv/e/dUAFd53HddNqvN+b+Jajlauw8OY8rbeR+
qnL7wnXA06f2j52luFJh1U62h0i30c7+VIGxcblDDhZY3068qYZahQAdiq4TNVT5
CR77w8ne8sUa2GiLAv/7QGC4R36xMx/YCJgTcuM0FfXLxQOP/W8EJWByOcqFkMny
xVfMKG6dVrABfgJFmpYp2XHs1tp4uvlKTfEPpq/5NIsBk23aWjOdjswooJ/RffVS
SR94dGmSudHiwrqhMO/JTR6iZkESofrXUcTSXlHOrTZflTGWMuZEFFxJYOf8+4RN
BQmFhRvkRUmY+1WTZcjSx0YJsidgmoUdXheP9fRPt4A5hdf3b8me9xhzr40ts/LV
ZErLznaXIHEsUdMbx/d8xD+tcz9wKvtFshZmWddYuRF+GZczLxhhjsMB2dWk2G3w
Nj/giOjvVhVhBQxsYA/lJ6pAJsMN0AZ9ZolusW7PUQaGMXu5/nwPRty6rGUWyt6O
z515uop7jCKHL4IHgOH6g/ClXrNRmvhSrIhSNasP0DaMJd/HpZu+Aco1SarGdYYA
ihAAXxi+765r8lei1BjZCeV7BnzlbMdXSyYlJRDVpp8Dz9x0whpFIGKb4BDk/+LX
ylnZo/yB05v7tRpplQhuMy9fWxpJj9USQz8TV6qmVNNKbk0s+96QTyPp9pCsZneR
IoCi6BhDDP+Lywum/u01QhtYFYdy3kKQ45h+bdc4uzcQup8YAfoIatyfQSaEzP/b
zkRlp13Xykt+i8ZBrAa9EY6U2uZ+wQgEVBsorWMx10Bk1MTozDUJJ0hUpKD06qrt
qDnfjRVFN46pfhpTrjtjq+FCioyANixKjlKLgFNIbColw4I6s2Gkd+Ktos9U5Lrw
LXeSSFTGskyl1ik4emNIgPjzTWj9F7rt8PSa7lSAcukKuW3wC/g9YnEXVEqH8FSu
b6NIfeXG85AYxz3cgduTtX/r4mKZAk/jgClv5hwhdZFXl+RR6TrZ2PWhip4l9Zrb
3TzrJPdk2QvT0xfehRhUICWMyslfU8ykZclwZG4OfZWTRR/Hz0P400TwktaXC52S
xNNxvqccT11FU6b//0qRyX2zsjRg4mzJZJhRShePVnl7ql+BCuzPNNOkmDteroCs
ZmZil1Un8Rzb1YdUw9Ye87YinF/EElTlnO10Vw20rJX7Xh1m0VkaYdlo64D4XAo1
4FWBVuEVmd1ruxRNlxqbJCm5eUAfytXx2056Hs8sJTCpHcWxjePue6+eZWjIf8Hh
i056q887xSscmVuVF5Bt2J1i+sTg7q6Mj7ahSyQJcMw+pw1EJUTom7TX1YKEGzmY
uVbK38jbmjbuRM554qqQyegnVAZXN5ztP/oUjtV5EvEAHDcHlRRraP3fpyOinIVX
ujX6NdCkOWihbqwjF5sg2DI/SxPKi/r/sZPLwoZKewacEaza8qQTwFvpWwBZ9y06
tjjWxLezAu3ZokVAnUJ4J2BTDZ9G0iZIz56PKCPYswp3QEekr/T8QCutsgD1jEmA
u8USRwl4VfCKwkBpxnogBK3yMVvNBIUHyZnilGKxujDrC5VXZeArosF9DbLcgDp5
Ox+7J31eJnQu3A+I8V6LYga+T2WUq1PMD4gIZvtL6KozTYgEAvqCy5rdGINHnGdy
HIv/+nD5czeYyPVtX0MjyLQu1Tw3Lg9XyLy4+aH9twr+1NF/VG6aXmd4cYEx9C5v
s9QgX2y0eAV8RrjdaWFQM9k/PvVAUtjhoMzMuII0UvM4/jhEdDRvwGFwjc62s1pJ
UKt65Kr+pCOREpH0g5QrIUfxwTvvOLo1XZQbCUrzDpuZouf8UMyAk2WaY0rLGzSf
FEBBZJcEds6lb9Tg8ALlx6bZ5meBvnA1YoLQ5mSE6Wqx78tQ5m79+LKHwFEfCX/a
IJdScY3hJr827IVOxc/spp02bfKsLxzQNmyOOMGCsrUojXtF7x8n2y3WFDZhphPt
EANw6hqG2JBQ0z0OGlHrBHeyLfWPMB9XO7aVIWUInEQXIK8KuOSsm0TwN/0x5hUd
5yNTqR4WF6KvO9I2Mh+8T7GTrTrZ1susXEKMCQm8IbR4EyDNEoR6HIpQVn5TVTLV
Lf7YrAUUb/AmxyV+l5/HgTLbphkEm1/P8xQy9iMumTs3wgwDlKylQpqMvU9D3XQD
xaB6gw612mIH2/GEl+lnFagBLqLpY8xAckqF9KDlMnUQtVTJiKL+0CskoP8Sx3/V
4YbrTo/Zkk+Zvb4aYwsOMJe88RD9kcuJiuSWOyfu7IXttY2cjD3cu8EDAOH4bVF9
c9ddoh3gZ2etFDZ52Gsc4sjGe6EfpFQZYekXLwvPLpXwLorRqPCqO4GWFqkPRu/c
ww3luMJ1XJn8dLlACkPsxaBf100FBHCmq2lTvbKD6q06RI78oYfw6pqm/Ag3wsBo
IR3hfyfAsxR9K+GeIca96BegLykjMvCaxXnp+YD02GSQkIh+cD2YwFk6TwxCN0XO
0D2yaRXSLv9R8AZGgp+R1EzYC8jhlGpksagLnyxuZZ6LxIxklb7jdxo263zYo5zQ
e8CteHM3J6VhppNVeqStvaKhY4V+ORY5r2gNWZ403lPNNimqewNSLQOh7emMs6a4
/6NAL/QNyzhOr/3FtQWkfjYGhlkrJzG92ZGh4THdj6DikVecsux+1qJTK0WxQDC/
Jdh08qRYfY6tbT7FUGlzHM98wHKM4/J6TOAycGQUW1Qk8TUClPrKHe+wjDNj9Jbv
FOwsxY5dzrxkN2iI8XdhYhidQ1G+5ipO/sXo77YWbWAEY6Wv2dP2g7WGzg2jzRxh
oSmiywNLwLWVrSXwEu/kCjqGLPasPjsqsvEVDymEvUONJUSFa0AM7PvoTNgOm0Yc
ZA50xqwMsKEY6KxPBgri9RXMlpzkyCnrZ9u1SoRbgjFjDsGVfdZ5HUv7qts/ic4m
4PCJT0a2vFCfFpMwTRTZp3wbcnLnDhYOu+IT1RSGReJLMDCiYzrrSpBNOdMHfCQ6
v6GzoJVXdgwgHaKsMiuVXmUv2jkbGl72H9OGAFO/l1m0iE3Bhr/00g3cf/ZV5kTM
vedjs+PwzbSi3kcNnf2jYb6LzcWsob2hVtv+BPClGyrw0lbgNx431/3OBJd/Ql8W
/1HlTvN/NrOOpwz2Tt6AUblWdZibapsKV28RVWiqFSE4w5t2jDNzFUCfgcN7XBJT
ncDicwpi1kC52TYZdYHQ0mJuWeWeSNZGCuj9/QnU/q/TTvX4ourM8LjhQLtpMCD0
uPAkcfojAuQW2RIs0Uf+g25lxGZ7EUmeCxSI2Pqd1NHrwjF6AZh9/U6p5YvIKe7G
KybrpsOXua1Xtv+Y68x95RXJNDcvJ1gN1rHDxVFC8EV2VNbeGMhtwvGMueSzlLPX
AyAKZHzAr6bkhHaboiHrG+fmWWEUy8CaKK9i7tDPxUcPszx3cpblHt8F2olqowfd
6YuhJnQyCGXiD6SPHXNfQxl7gDSTvyJxNzltqQNMwdewSHrDrlJrw5UdHdcUJnA0
ph6q4chHUU6MFKdpV4MuuG3MUINA4wc7sbS0PJQ24lxJuZvOkEERUdD0bUKDqk8s
yx3aNc5WAsm7IW4yURpm53mzNl3V+VJMv+O79NLpvGYgGwusMcxR7pyJssGs7i9M
c8Kz1JVYREtX6EE6+wQqlZnPBGpgH1zB5Yjr4epxxn2Ok8RUB3gjJou5eN64nI1y
YF6Rc6qUiJuHK6mh2VZflSDiWRV8k/NTh7DdXPNmZDU2pwLfWECBRwoIyUrNG8EM
FIAJtD1qpp4jR2ElCb0HbQeRRvmiWoEAVtWqdNp1X68qMUK/Hsquyj3rgutBn7YI
LIL7Adu+awXFJfteruwSIC2X0l3po4zDOzYiGFGdudjiDhBYw6pXw0A5iHOuaRgY
PJJ8Kp1qQOIPAYhnLvwA7+IoQE0H6VodlltlLnR/LZhtckJb+z7TTFfF2HPeTTcF
LB0aOTb/Qi813/W837yvwyVKJuFI1h1pI2HK/6YLwmPfd8pJLbj+Xd99frWD2/L0
2EWupk2ZhyVNAvWz8klJeV6XF9l7ijL57scGR5GtzFHUlAsRGjOLteMFOanMmm/K
u276zMTxeQ5qpkU5BantqmsmVe9H0280b60FW+E7kqCgTIPLCvx/Tiw8JjmCwmkD
AbcmKoKRfn8nfa3T/tq3oEOpqlVDg+8pG8RTMZst0MsGXqIAkRIJGe+Ofy253HEO
28lUhtUjGFhp6vwb1GC9PeRcrmt1pNtmRoKdTE6xO+R0BJYb5Ta8nLVSyY6HPpk9
nMIhV4O+jaGkAiJTaQx781zAUuIb5MkSXQUhkzvvAvJAZjY84zvEG+oQq0Cu8obT
/rbPaNiOX91xyUsNWh6NDcAq80uuF/xri43XIINF3bwWE/eXgdIAvy3SZtUyd39P
flht0DFig36LS49QCkePxcYz0sC+80r90Y2sg1Vno9wJ3dkEtVPPSMlKYgB208rv
vFWkSp1DvFR7jas8Ve1sdFy3TY6fuay6rC7UFneSBKkFKDAKSV0aa4M3W1hArOXb
fAgOhdEd+gSA3/DLpZarFMiSVuFSDEBwzG4shqg/aOySB9KuCslDTnWKamZH1nOW
MJu3iDXhypSYWgc+PtBI/DX46r1G1Gl6sbyX0CnZwB7sJCHEIaMVpoYjsjYFjSI2
XZvJ+AzIyqV5RIwK51JJccN550A/qzdWyktQ1FurN8RAFS1ehOFUYp2RDrSeHoxF
b7GakQQNk9Ug3XHE2h3bqzkB7ZkQJNDWbC+enNREq87jVRoaeF7MVppSaMDMczbz
eQvmwPFAbocchMeTldINl3GZWNNvu9zFOh3DO4AgZrqn/7Y5zRAxb/8POSoNxe2G
iCqg4R8WXUfJgKH4LWepemdHn5zDkB/jG1E8RtPW3BgN4A3Or/rt/22e/fQSLugF
RgdCyJouq71knJlkXLg0nSn/D/V/FW3AxtjVG+H0/WlFuhxxXMy+Bt5cAvy37NvM
7YfW2pojYNmvy4dXyiImzNJqhBfrUHQ3OgJgNCGpFfwL2on3ep4NJ1vTeSLobFeA
lOInPAWsGYARRYBKdoY05/qbVQKHcFU/q1yW0Cgg+SnI3hq5ou2K+IKQKceHFTdm
lBcGNx7IevbuC0vZz9Cq8TpTs6ps7uVDMwOoJd7iIEzN1Xgn0UKuW4kvHL6bQeG4
buILcxlkPT1GbD2OlNUbf+WFHpatcJFlLHzPM3botOYeKg+xQW5aoAOquGn0KWT3
18XttpynJ0v96wsiKDeEmwxuN9/YMTNBXAjimZOyOA+5OrXIl5C5TaJlB20oCrlN
FHdI7OrJln3aGwijJoV3C4I1iJq/P7hkJuwMe+zfmK1qkCLkjnsLpsfbcwMru2st
78YaefgrJQ1Idg6T0qi5vK79gHqSjGZefnzJtPONhqaMRC2SXyTM82Ybo1ZjMdIu
kyOD3LGY8sCXNdRq832TXeWkXi4fE50/s7eh45vFDB076sPiwQOXPcwqpX39L9ra
Vg++W/SIXPwfHL+p8Pga/XB8HIT1HmiDZyYaQaSn7Gcg6wjJaBETZDMSd1I+3n54
Z4ahBDUMpRQO8Qpx0JftToGYgG9ACf8+liVtbgeQ9ZQ8illk0SFO6p0MJBePzz21
gev+8wC2sIfrNmxxB0C9dqG/XQLxsXgGSfteXLrOKfVXeGSmshRByxOEmWlO+jqY
1uud07u8iRyIZ/8d9Rfw5FTddnw5mFbkzZAoROXVy1rncjvvVadkW8YdQslRD26C
+TKQEqqIlk0PrvnO8MCaliNcIgfRQDgy8OVZWXOtgPEQQTT4fNLtfz0bLHAkFvZA
pg4IIQyNpkMNb9qIiKswEuUvLbi/Ctlk19pt57q5M3JjKurRceWFy4eG7aIGw1P3
WC9Sp5fupOWONV6T24QDgfImJgxhskfPWyTr5DiIlUeQxM7Sz2FuUQCNx5wgoSVb
heioMUbtaBd4mlbEUCUFsY/h6xqcWLNuI8JEhzI/ucWlXWre8+FKYBiOR355Fn/1
9F14/L/hXnMVGAdURpaPnditZLQyiBhPWrC3+XjnMGRBhXAMsnoFiEVem1NU5ycS
SXUawiC/p3Lr4e0LQPXSqlHjg1K/ebLQCaurVaZ1x+DDZE14EQalHzCRq1SpyszQ
HzAZyfxOl+Lk9+w9tTZUwB53bJSRDnYHu7RYP3a7MYBM+P2dz1QB81OcSKcl7ciG
7cWpPlylI3P/PbOrtEkw8SIR9abO+duJbtJ+en5TvdLO8u8CaCbPPJHBHDNXMuJV
UrC+2i4KfYWezTUx5abAA/DhItkXzyxm38emOCCtid6o61dMqEMB+7FkDBxv0rwh
a3ZsdwuRwxyRYJ5EL/J60WZ4ACWvIM03uD4iKl3bW5WPGsKO3tj9CsbhmZdwnXBa
5Ii/vkkAfkIozmEX9OL/6VSIR/7q1nUDzg8tvjuNP79Fl2eVwcb6f1IOfZS4oc84
KV1MhUcR+x2BQIQtz4E3Ys4sWL+5rK+Hui6orv7tqCBIKCkDqgwh+fV9qp8LrjL9
C4w+HMC8y4OyuWoVZ8Oa8fbhanEPmOQGHtEyxx49S9dKXpaxBPDgdcJDYku4smXt
RnRddGVWJEpYDuIBRsnkbumzRadHxjfa7FIzZRdo1HMmF2a8ef7762oYPOcnnVYM
s8zXSu3yOJbDDZK17+xq9T/LCj66vReg+CZjiVbjErXKwPEvk0DNIqtlquhZ283g
XUqsW9DLnYBD/E4kXcE/JRMpCjOEiOnM1b2WmNSDht26UC8mbtkw/O+sikpkSZLN
Mh6+i5thw7k/xDLS2HlMe/48M5/Rm+EgwGZ/s5B4hVjV5ORfpvfBaKoSZJvPgxGO
wpaULd9KrOatVNwJpvuaB41M80Tv+heggm83+ueR0c8subQkwftJzR0eC3h838P/
BZvv9IU0aADMKEQhbzLVTEiFO1vcLzgNeY0ASZ1KK+R/QPXCiGtQ9QedraL4YO6C
ul54ZvLosm4aoyfDT186hnER4orxfS3oZGymMvgIWU0L1c9NCP52nfR6Z82m/Pm7
r6iMVKKpgUvN1X9siNNz12n+fJWZoLXkmxOc222mnAkJeJEQBdzz0wE3Y36PDHJQ
npmBOm7xtE+67bWxZ/wiDor/g8Ap25JVlmRVUeuLz/np66QXmNLMdzdCNbdFU8fq
gghpW3eJzJZMa/4b29xy0rO7hkHyJcakNayZx8ebvgcKfC+geQ41XYH0U/oB0y0f
Jenh8n9qao88BkDSssfEJzpO6jaBfqamF5Ms9ube9ztXrt+vnrNu8DWFUdq17Awi
cauEdDl2buY+Is3I1fxOTaOrX69uTXl/wXUYBvyEgFXYLzlVC1Q3ozYDTiZgtzFX
RXabRUz+ucDawP2fjkVO3cDRL8G3yuIN1N5AL0d2Y0aJRRipjWwxX/A/Myofn5F9
+vKBOC1cbjHfts1rASC0I9POOLk35S3X1TjeIwSE1dFbUzu8x5ibmDuyxBgKC9Ok
n86ZfQqj6xmmq+xvuIBLZGyJ7LuTZ2jCqy2Z8DW9pTXp3AgcGIBZ3Jgbp89rShMY
f314cWbPbVipcfvoMKQeNsiQpjI6DVHKe9GljoyvIuqDW+M0N1RHnIDrMXUhyyGL
3ychlimo9rNI6Pdrdu2o0TuK7FvsABi6xxrh5QQxYfYN7lkWKFvDZOmks63QuW/9
uvnG5R9kT/dp7JtBH70xCYLFzhLyxd+avrfu8qhfo+3uGun18gVbJPBgkX/dNqMF
qtaaUd8u7PyYqVLYgukKK30IWlnOnc0JyTDX1xhWShWrgVCWFVdFURCh+1O7tgJ3
w5ydS4B4IVcHwpc5SqP83sr5coKT9KKRe1p0QS7dtR5nBhPIaaSHFmrH9Naws5Sp
o/fGoZZW+DgQLkXpMopFcTjnb+oRYIkie0IqFczOCNcCXKBj0ceproth/tm5w8d4
c0XjBV3DsUZjPK8vtBLF+TACbLm40KNCX9tYU1QcSzsdxD/IgcTnwKDKrPtHmTXT
DG0bpzhhbsZi706xOvKOe26f22BlEJxhX4Vow9kTqFxd/IHEkexwVXLHZ293PkJU
tVEZ5ScWfRYkDy0lYmzoZqFijWddP+VYO2CE879Q2ohr/w2z1QNfngYQOfuj/3Cg
cxjdHuN7dA8wDiLQ86xIgFLzZ3fDoncoayCasGjZKPo6UdKJNmlTmGbL99A0KNmK
t650HDvQSkGpmS8oxmWJeOYW0KYF8NmqgFu85Kju9qovTGqe4S92eaB/ZtVDvzf9
xS0nOf5MHgUyKOPSf/YvyqOTgI0/3vy4E//SfIHsdkLWypyny9Ixvk1MB4OHoV0f
BHzaW6jzsvWi9P358iUE2W5L4KIi+wucCHuCa4UgwpV44+tCYFvxgaRFIqsiAkOo
zcVFUEjDtxquD/XTD/p2EQxma9RzrA6aF1oGCB48u4PgJtmkCl66t8Nfpq1QI9FQ
EUqqVYTc3aeTfM5zGOUaUW3OHK5BwQYGRSTTPJ6tlG/1zO3Fmc5R/XyxYTM5B0Qj
Gp4HgMl7wiR72w7G8xheXNCkIBF3DZUAaeu2pO/9Wv6GrmfdGJEhR5iTYqKGEP1n
VWNFLZTBkfkq60Yzv/jzi3xr8wcvnMPoI9IseqYayf/G/wNtKaj5cJMjt+s8/rn4
QlfgU2oZYoOOCt01/n5OeAhW+FmmOpmgch9KDVbeqw9wB8NKnigobjEJYx7IvY0M
TbpBkYtJ2bXYIEhLO1ABPW3Yl0j3qGhhku5B47GUuBq1OZUBZdbOXU7nxclULqZA
WYG4sJhGehglzuqt6XijVXiVQHMCSN73u+9q4Fb0tVzt0d9eiiS+gdt4KjWJHA9y
fYY7I510KgMezEn0GD52GJEOQWdwsLYBt9ohoiHaJl2cxfZ4QpniQXrY2lR4V93l
ORpdFONVOi0OP11fYCsWRGhMcJ2x76wu1OtQCYwUqQalFS0E6BbP+wEFGkNGrOCl
ti5K9vSnXXoWjEgu6cAuCLk4xPb6OeG2Z3mVoVfJ5IybbKa9x35SFdvL38/eH5Cy
32dKiy5UIHkPh2LUXnlWs5PVmIyNnjPezyzk/rYRJkUWAOMobkVx+TUujXRc5QKd
lrjeNkjBLsqDISoSzgk1Wq+QpB+UQ88HL8nhJax+nigsjB/vywLjLYp8Z2vufM5K
BCgI7eLatnhKpEkBjgWnM3VK/BxHDunCzCPB1quPUhf546AOJQlKtoU9pLQAVpnh
G7WsIswCkoDAZ5HxtOOKupykc5/1ZD7Y2C2kSD+zBtmsOfynuaPDUeHmKOMxMDM+
FDoTvcnm9AYfSZyupke0VGpwHtiWoU3blqQfOdOYsvYd6Zt+RGHmzkqFRA+Kjr8o
zELJPeaFqmY7MEIjptPSzfiW6jLBWn5Uabz2wa+VO78L59mKkUR7maIETOERPabn
mGo/tTCIcQ6jMjP33vhyv5sfEM/2zyILkyoy8WInahd3nS2b7Dr/qfMFcoYGfTqK
ee95cc1dnLPTjGC/F2TfVNJGa08Ttk9q6z/HJ+LOEITzA/e342vX9PVFBoweuQ/Y
odvsJddcVgeghdfmWYHFfb9kBUfgIsCO21vTgR7Y6CORbqykPGJtk0hnnVgbxdb+
sHAgkiHG574zpx/2Gc4snehGXX/sHAlnLOMKyxkLO75Yy2+KlQAs7RTB08b6g7EY
N+H1YhKLqi7/owcQdaqB9y1S3GmNyG/gzMCtnGdDwR88/gHBRA8De0w5C5Yi0+DF
g8kugXblZkpxouVegc/nLbkdZ6wI00ZiM7B8eAVwHEraqo3X1yLxE0JpEdPfgsNx
wpUlYT9SIJLKuqWoPbyDXuY1PbyrxSJIcIlx9UbO7Ez8HMKTPhIyqjz3UWld9iH6
PlrWFkMaZ75sQ0LDbbaOPZ+V42HvM2+wKkD7wogZy0LlJZtpucL7IFY+5kYAe1Ug
zA/MYS826T5fXvhp+rxoSwgWSbruelEI0gC+oOpdfp6Zkn+g1x1FlnxK/GlZ1/MU
+ZUmuZBsEXeQUpuNkT2Ig6C1MUPm7DzsOzeoNtqBi6E0ZB38yY+x0/vXtkIg6P5u
+B2hkZ8mIrNP5PpBulZWiojsUGlNSGrKQoyLsBppNs/8lqwOnv9wdQ0yPeFeU7rm
rvEFDKoysxjwpZWZGX8ZWSpAEIYsLTD72GJ/18K3SfVFrxs4UKtOdD4+yj6M/25k
HO18AD6GPdMVsL1LKrmrGUI47sJJpa06zqsI1jcPOsE3KH9lF91ljU3t2fyS3Si+
h5IZxYftZRBypow1hIHAd5IymqhSjY5/0JPS9IbmEZ9+gPCjpOx3P0g7YW1tS6DM
KPjeSZETE8GdeWYULOle+8zxJF8+Fizsvj4156ai4IySFlzCiYJw0Abr31uvHoME
XOIC4ud+buuLAIe7OHymiRz/MKDN8FR0RsZ4CxCLoBTcGb84wWNXl4aa8AT0YAHw
5g1xg1Eyyw4QAxpFLtjteDVYgqct7iygcv/f/kkqy/LGIPzrc+D+hdVdxqAA0Vb/
CCU2XGr0DdkQv2326UCW88dP1NXjJuPf27693rQ6oVIXDGV289gYDzDm6I3hli0D
7ftEENOiJKz9TRFu+Lgb8Fd3KE4dtkou9B6Ta4AfZahcCoVeA5WlSusUuDQAA950
nZsTrm/a9RLklbLBnc+GQiYLziJYssprpjtOnxHHekDgfBSRWxkeA5oRQGcaJywR
KL4SbvLzWjAGUioEhkZx8QmdbnsQ8ZYlwruYHcn9EqXmFAer0aEOnDvVKjCorM+5
0D35zJHJG88eopcUYfYl/mgBUpYOjuiPi1owlCdfJbIl9GxnUe0UfndFPyXoLF42
zd7c95HHbLuCsSVx9wBcMKgOAbiRHFm/+ujTUmGP2j68AQu7IZLl9+o3ciY92dcr
L5m8A2ojIVkZUV3neXMwug4bPHIeUQdJF9oERvEQ3cKhgQrZiii0C785RCR7Kvmp
dQzh35SfsWFFZ5NQ9WO+OxpVQholQ97NAR0I2Vst/neUKNjcadXzAZEUBNP/niu9
o64pp4spOUEr03SN3K0oPMpQf4NjTYp1uuM4yFyGGGznv0tvTwJZY6GsfkEGBJDM
IcnzCt8UNhOK/kSUMp+U425pmqXZqosTSTQooUsXO+jNgStixegwtpEzff/d4IGf
Wb1O5vOTSLrLxUeKqyQTa3i9AVZzl0dgapWlLObX0h9LMZuH2Yoaqg4rvIOVRs+g
sjQtaSstWk3cpESspCC4VMcOx0lk71USe3Ry5SseR9xuTbRzyqu6t2AqYqP9lF8/
soamWCL2mnGrhdtRj0Gs8Y06UQN84Y4OY6B4bVRvN6GqpF7oTqQY7UtBd2WXNstZ
DwzmyfBSRancWpCS9f8snTQa9FC0C2MCMVg32vu198lvLvjQ7jHVdEwVuHZC8ACX
ZxpnEz1DtKtbyUyzuWcUmmsoBhtLWJKiVF7zlXn7G7zSxglV+qgaKzDXqWJL4+KT
DLqrwPTLZWonLpWsaJLqRtjY6v2B/jnd4HXV0DbgDV4XVlESlEWuUPhCn4gYsjlv
CiUtaw6pI7dxz6rE6KYfqFoDAtGC6Ru/trU37aw2uQSU8LdAmcS5G0TEsRGWM9Ko
Ixt9GA7O4pfAD08hpjaYZ6IbWP5MwXwGwfc2g4YMRYe0op3b0IOe9KlbcBN20Ldj
e77VpXBnhpLBTaFysjJhtgcmyGtHsFY7AiUjkdlDKAq1m5oXXS6YUYrk3dzXFneq
1f8UTlHFjnx77NmCmSF1HXdHU4zjVlMxHGxHPDFDUiNrVdFoc6bLUmHwLVXj6hgf
3eyfZXUVbwn8JMnXxVRNCpY4wxd0ow57vPOhOdnqD1mXEDgRxlpLDArz1nOSXFuB
N30k4dZ0VgLQFix0EFEx19yflz5X9tOQhtOJdHcdX8c+ra6hF9UNVdqKQdVtJ3r1
pQn7iyFowbL0CeDLMK76+cMqxL9C3JOBeeHThilrciaZUKFEg15Dk6wNWLidoxJf
VnCZJbaj+WNSKl+xoMmyGMQBZyJToFFXjoPctBk8zqw0a2S8xOBUJvFAXPIRZreW
HIkL6kI1kHvOSgRywWKomzNOrxK6l4XqT7+QHb2VX1rXft7PZUYSDPZirKMU42yf
XTsn5bDxC3pnb3tatM/0R/WjLd2t3HbI+gdgBTTEJFVPWoeSKnOV6TiqVQoYX4np
acburOQb4klnJ7d+zgN7EO28HxDNRg5oBxi2Q0l1xzprFwIK1ibwJp2bcuoYe8Q5
yy04uAD3J0NILn+DLLzdvYuOqLeWdr06DjNqFPF2QQ3mt4AYeIIbIs5jOxPogNX0
fYuRJspijfAHpSanBgaXwUqLXiZEiNlGuVvAKVqA4ZXoQcKGEMTdJ9lTVVKzgtWo
bf20nNCfWnxSoMEHTUxEHYdp3o86AQggPb+ZZGb/OvsrgrmanoQpVVWBMjhf5Jq+
zLrhmaKvj24+Espk2d++9/VnYDl4LZkHpigIIhxjT5zmrhJTeh3KO3a6MlxQgdhW
EseZis998jEpBsc5dTBXZaQu4ALDpRfoKHLEWZYMd04u73/Jwc5eOt+lbmexQgNX
fUWNwvK4Y52R9WZL7TKTYtuNz9lxWgy0dYUhQfCPpI8ZRZyjjAgn5gL/FMoQUR8k
X2igNOYp8r0+HHwBweSc6Mn/QI3odZ7q5bkA00gtNaPg6Hqn3wNIb2FtRWfAmosu
KM67lA/Nbqbp93fKIQ4uqJz9Ylklf3qg96HFxV0cDIX/RcHeEbNNOB4x5v8Lan/d
sfKOblD116oFk3GSDKGA1NfIgjplXsBmR/rHbdr5RfECBxOGlu2U07mPfXHpHnJw
sej30dXExZ8h8UM80wOsOG1GHCw6z9vSqaOcQvuVV7qGO8cMBORUQr4y3kHAnSwn
MYqkfVEP3vvS1V17c+300BLzEqYrsRSfvw8x9E22YZVf1KtBocFsUre8NXZxhBZK
E1BcDRL7CkBoXfUgG6HNt34tJbNHUm3wPFzaJKWjE/mTbTnQhEriB/SI0t9BLYbX
y40NuMNmG2u5225R7X/TKW137sqfkylQSasmiXo8+lAIepsgEcSCjTc/whv6WQN8
YZyovhl3599CbRIFojeTHggWX3jfAeScBZBsVwinlzBtQXR959y5cqng6abbapbq
tgY24edaczeqxOTOevxhSTwbnFMb4aVGJmr038AkvjDBu1s6AsV0LRJGc4inr4H8
Mne29jV60qmfo6IsCg093hfeYYVts+Jcocq9eyxSv8CDxNX6DCcUQW9QqnarV7YD
0CBstt7RyBqSlxHj0KbM8hUmC8MPloOW9didq+506cxGFzRS6yLg/fIahXbE0v3y
p1/Qblc3GEB5+EEGIp8P2/oL4KqqzjEEkeQxnA23TUshoLlL/8Eb6hRYfWoWqOvJ
ysUA+F6OqX7/+6Bx6ZDpxWfz3rAKwR0+usxJIG3JvjYTG2W2uBeSjG6uaRrIrwH0
eyJdKxLOgPHXDZ2hi1mG3jgGrWcZehGt+8VkvABU/q7SlYeWJ6v0RdOcQwvV8qTg
kgLzhXbq3by418/PMabpgnxEm+191Px+CmpGPzutsQAK1t7NyKeXhRRcDItQdpe0
ngBqcyFrqMI5dNG4bqHfsDYcStAs3trAfpPh2oaSswofZilziKhuce3yg0ZrYSIV
ydVOFUOA8dh5k++NIVVl8LWUYHkLofsoHDArkpO0Uc7ICNCxNXSlIO5PwtYQdL3s
ZpL9fDA9cyPl2M3vacL6a55iXbZ9MnNTweyNaW4dVKR+sd15S+H3A3v7jdHhps5a
1s3KNSbT+hJe6oizqCg3XI31L5Vf5yqlSh7mGHChvdw12nUs0/hFGDnZb4rqmVTj
6x7iySaicbnjoYGJNHzFFzrOgnWtL/Xyg6rOx2QRGpAiCtPyDXyamR8FKb910U7t
gEigq0Ok4sRlTWHpW4Klce19akC0qSheCm6sN1tzJho+mwf0jzQZStt8sRttN16P
xnmgu2SjQSiTpoaF0JSzKE1T0m1i96naDDLSmNrbpZY2woNLcKYWyhdSMRJi95Pi
UTSa3IDr3HIYo3lD2lXt+m536ZcS2UZwSjRosNUExNX+kHzk2FMsnJ1KOz8D/u4b
1bTkI7KJDC7RNwlGvkWUDbeq742dfyoz4D6BRQXB11t2TiExoxAukmOl5UuulRKw
O3tu5tdAZ3V6fr+QmU0HiyW0his4au5JCf9tNK7JytFByXKhmknn2/KIQ6rxgAL0
quGQJ+jkkJh9mokE9PcNooGgVrVeIXjqayrJcS5AoMqKV6UEDP8ZVnvRsZ9a7160
rWSbF2pM6LhYt7R9u9CIvxl1VwJylxity8TzAv9pO75ZodLPkt+HTBwa0flCejBf
FFh6+t0jZwawJpS+NTf8sLusWShsZj34z3zJ+wHGz7rt+By0e5MTp+bQzO/AOcj7
qVVuhlxkHh/taCoMYj2qcrmx4i9DkumjYHDfLWTYshtShtymx34EPLMdTxk12qv7
FXt6/FOQc0LMMPLKGPawEGM240PluNtINlXEysFfqD1rrHnrMnx42swRVqgsCXSk
/gbu0Vt/FhKExusNVFey3CkPAXhC3GQ+e8GiskNyX4lRTVlcjF4svDgWUy1KwGAz
0KLNfqRFA7wo5av1wIDX/EWUxxAvU4OCfs2x/i6PCb0cCsoy56DiD8kl8W6TwWvD
i7485cQfnpH6GFFIUEw+lpFK134Tq+ZICXbs24Fv6fCXJL6PbG4KAK2GHnntncf6
kIhTxu4W9DQRV3GkKBd6JH2uH3r/BFkj/C5wccTO7BTiJbA4RXJojsEfx3bbhFWU
fcVw6Lmx/P1NvOseCoMmY6Fp2ia5L4RZfP8MMhJhizi7Xx0hJTRSf5LIm2eDCnWk
UdEAcxSN/moUSPVhF/xGrNOHZrGTkbudkw1ugK6dqro=
`protect END_PROTECTED
