`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwzs4pyWo5cfcL/CHbV3vGrTwg85SiiI30jPsSh3/aOUGNmajUWyfuPFy1dj/jtm
xtecvPDKJ1HULueOUr7v464wM/6wHBVpPG8DTEM7V3AkikRaVXME0/76+4sFzHxm
Fowxd9TlTkj6Y7rNhrZEVxAxlRwvxzpcKk8S9ChDnr5vzKKfjvc7pWYxig72yvug
qhmNrEIutnm0P/DrGwWCWZIAWREsSSKSHAFMLtAo+MUZnYJb/pASB602b20m4AqG
LmMDYTyafJPoLPYZggvTv1CdqtiP+6GKTIB9C4/M4MtitCJDeMXaelyYJ6Dh1F17
xPLGKsvNbDh54bT0/J/zViYsZRfwea6bcW7hrulRHwrSERJ2oTADKa5b78fezvKg
nv/N98hyO+VMigI6KAqqfw==
`protect END_PROTECTED
