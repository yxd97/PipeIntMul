`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Q10/GdSk4Ho9LkZh99ExbB8ApnvsCMjNoyrfFXAl+XxK2BnrkB4Vs1Dc+O+KtZI
YZAc5La97d6vQmKxRYMRqIVZevOR+n9xwZsnxkAywKtpRIcyX7mJKsFXXFXk0xEn
05DSizMXPAKU27pkSRsaj0E73eog3cXvKdxi3NDanrDvNlSVVbI62FEFqFEq6qha
7+EMsfHkj8VJfaK5dOL48ylX9v2UR1O9DRst9j2OjtR47Ap0f9H9BsRH+AiDRKh7
NMRv4+9Jjysl8Nf2S9fnrIAOr2Tyz+v1tC3jN3N/hfoaaDL6VgLtzKnM4oMbs6mi
nz2a0xopxhg2HNGE4OK0TsgGtwMwN27yLejZcEExjPoSisCFI/YgAUqXgZhNCipZ
8hO1KusIMuysMunmV/4QUrH6amDpA4zSPdt+p8yXn3SLL3GmIxOSrYVsf7g0j5cS
5TGkkARahLU5V0OGx5elPmIccE0u+jqiD9h1+3hosLgBih2PFwFx0ies53dAzBYO
97Mdn/zhyV8sVv7OmCzKZDmoSNTpCvOU45zO+hp0e659h3WRcuSFl0AFSL/r3C8f
r8NjAbTniBDe2Asen2cQY/N1JgyVIKfKyxMQFJmyDUN/HKn4PUtivRzsSyrm1T8s
e7pvTHL2j/Zp5kJHbdJL7sRACHJ6wscGq7SsSTW65FRm/IiGDWNrMH2cedSVYxS+
a3Ow8Z9qDc4GpIsd11Ut8DBdlx8lQUzzPUaB3zZppis=
`protect END_PROTECTED
