`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zr7hOj9ey+F9qJ2hFg1R3ePKS5wfq5LZOblz9wLaS0WY1wXihqOrV5/r+XjbJvqf
AY7OMMFRVDXHBXrsl2AS8oQ+WQK95a9z+jnHJ3Q63JPg8R2aV9XESFAvxoLgF/MW
GjmaQA17YEKHOhVgh/fhjegqSWpAby3TkpJzt9l/YuCIL2mrZaYxZuyTzZmEznTT
d31dIStIdfHNKqb1+22wtXpaDSbx2A9VQVQQO9KWCArQzNqdwSxV8ked7JVe8AR7
537A6cBF8ELIqVcXFlYO2NwQHa8+hdziu3WKp+9G8ecfqLiZjp7UuHAOTIzMZKki
RLe+zVHfLjxY+8Hkx87zegLe765wT+FLktdkREUkn4MrHebtfnXOCFqbNKcoGhTX
DOiPC/MoYhvAITjLYLhiZTopGILivBqzZ6dyFpB8Xk28YndnMNIUaFy7ND6LEpLK
KgldI8dMgdya5rgpRg7rfk86JHTr0ZN4nx+gFNcW0N8OxiY7BviVbdrKBP+My5Lh
+bMuZ4tQLvwSpjRNinkEIC+uO4zpWtb3RF/Cr/arf9mBqNgh90DJ0AaVGYJyWPQh
9nmIwegUVez84ytCCkolfbY0/sVsigmM/gVrQsiNyEFouHLx5ayIqSP1i+Ath98j
GDMKx23dWt9FgYERxrSyH9Q6hB6+szXsLI3I4j8AAtaVDX28pUx4iCZFHjNDcyPM
TO88ipavo8PFRNsQbgUraWPNNGGVCVRlQTHmGCOGOBLRWlisDmd8iTi4vXT/aUuO
LZ82y9Y/9Kml3YuYDIk9rVkZucvn4ZxdTuKpnfr3vpZ0TRGDFfb8VCyF3PrUsJ3E
OUw6/wnX0VBRCDkw2kjbuFNqirjOM2vfDXdFJyeV6+p94CkOHKriIjfVA5t34IXD
LDJ79HuPv9oaTWp4Ml4Am4WtWzfFq4VD5BREDGBxrdNKxEEz+Jt6pLtumiGuklh5
t4IKwSOxy3Ob+IEGmEHE6A==
`protect END_PROTECTED
