`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbD6aoqGXHGr9cYMtkqfDp0F1/GVpn84Ig4a9ZFk3y7721UYcCR1NlPbpIqBOutu
soQZ4vyj4Mt+YOFTmK4P5xLLKmK7GBMHRnPDneDGRFHQZx3FHuKBCOaJ6BgVB3Sh
DUsmNFGpoq0SK+F6RR9ey/nuqCN2QZT0SHHE/KEOXjjv0CVd2ejwdhi/i45pQ9It
nweHDSmnlDRbI1T+DnTBO1Mo53GZYCJ0cdnIYeO4QLrBO+nGCIi9GzdpEw6XkDVe
dyT79/2nMk2+fK+eO5ZGxCu0v8OwiBrAvgQJP4PvxTIqYsk9TrqWt6pORLAOycFI
wfEHc5/hSWZD4NQZQD3gKU5akZwVfOeNVy0U78qtZWV8oXrezyd4jTQRo+OXwaOn
lrxdmvGDHq54EJkCJB3AeT3jymM+q6UTQkWEKoJfcKCMMYkD5JybPH+u4rW7ooxU
j5RxjFwYbXwY2uXVMvqNepS5Lqz9hSSuQMvC7cI9MAtPhBGNWOrOmOSAhsl3qegm
bbyo2A13JlvwDUxoU6XcsQ+xvGk8p3w3/KocXzfOYfbzQi7JLZX1Cs99NVq5mMfB
`protect END_PROTECTED
