`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xsbGdnQizF2XkvgJthc5v1LSgEsaxj+drEFNhWM6YLEP0pbZuizHMldiHOqjE29R
7ixKzwirc1LEeXtjwak3yqvcG2JCem1cYiC2HIU5Mq3eNzq/Z2+RSHmTXfKRoU4k
T3o4OHAXJ+9iMiCQxjilcSzheXJ9aTrW4cczIIMDp7pxKVYTFZOfOsLfWK5BcyK4
UD0jB/JXMkh2eVTRkNmIZYNctOIN7oVtcpN+7GLTkWivmwL/+eXcpovuYxqeA+Y2
Z9ObQO4/lSi9z+TFTj2CvnljRRgZbqDyXqM6hbBCxT3AkgBldzvvaQZccrbY/ruW
kIkbugoOtew2+gUVcgR3qZYiPMVfUYUMM9ggyHey5kdRAt62aenH6TFG8lZo6JKB
eKzq6SWkSZHU6UX4+qs0EV6boVelWqhGf3U2/5/Zh4ZWOkvVNzO9aHPAoYoVUhTH
JP6arosQD/V46pWMcgMiStj5c82ZkhldjOauflpcS0K3dhS1WvqtTj4+H61C4ywG
endsAH+GZLCnSpY2ILSz3x8QwqNvv2Dl5+PYVRIGaedhWC5AH0r9F+Nc8pIHSHSP
iu3VnQbe7ZdEn+j1hEIQ5EWZfTDaScVyyeTg/bB4cvTOAxgUEJBkJnf9JZj6lle0
ZdpuyjPkNEXTUUf66yeRxA==
`protect END_PROTECTED
