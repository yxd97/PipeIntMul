`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pHNgq3txfnKXCE7g0Q5ITVmbFpqBviNwpDGSLC663/L2a13v+XE++DX8pjaoZKeT
3A5gviME/7J+EgU+qr7FAMF7cWoSNmEI0Vso6Qg8NdQH+kdh1462Z5qTFqqiCbMb
WaS7EILGYB8Hvl3A7lE9oahRZWXxHG5xhfvvMewWYlxChZ/vUm1thqs4rfFQ7oSm
/wANVWm+mZMqh+77R7Nkyoi8tZGnEh1wZ6REZNiRUqUTRfyK09QkVH0iEaIqmtmp
kAvTXuQL9x++IFRSRGfl/8kp9j9rqJRRdyNJX4kGkhEuFPSCtHRcTG5UwMW6y03u
GDFfcrsgMbyvVT43d40AGIwJsHjua24DB3fbZ0ghel8zZkZLkKY2fYtnjng41gOY
kuq3jBCPVkXnmDKBqGzIOGx3/7cuzB3o5rUryNk+bRWFDtTN6ExYuOgdT+VbdfeP
83TlJURETMF3qWsPl4yfMYnUoz5i2tIcAfKFSO16VwvtNVOp1HS3e2xMPHgw6tTi
vcmUaOCxCNC99C2/rDeYchvzrBYEx4E3lFMdVZKi+rEjYZ2yzERlWJSHcoYaRbhF
q7ZGDf9XQZC5rg0suALkib9rOQyqMmtZ/jeMFCqlgSmDNhiKe/BC4oll8at5ZkBv
qDyd43V9el9i0mBmaQrc3g==
`protect END_PROTECTED
