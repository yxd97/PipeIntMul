`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgmEJpZ/+FG51W0fyINthgIGToGPVUxUl3agJzGqB3zVkOP6N5ZO+yCA3wIyDh9O
A2yjNMLuGtmbt/W4vE75BHtB9MNi3nbYDAz0KdambXEr9Opes5E/jV7lTOvF6/a7
jssi2Rt+nJFSshMUp5r6w9GbZJSxD2+MOUn6bj2z2b90/4hGhGfcJllrdr/bj+ZU
EXdp2g1nT91OWg59JAy1zoPwS7sh0sYVU0SPAZFKmStM83j2GNWFzuxd1NYrSvXH
4uepF8QqG2qVw5HKgAHjnbMwWYdtdX8VV21nTHS1Dqz+qx1iSkn5N+utKJaWwBt9
VHtw+dY1Pl0hTUihxdyMMlR90J7OSXa7SHQCLAcOgm4P5WItSy9g3WUe146Z9fC2
U1GXPwUUe58542W/MMajh1npqj58JVKOUoQOA/9CtMPI1a1MxLTXi+jfn1rcn3n/
hL5vAsOAxYBLn7g0APUduYhHbQ3YUCmPbufdFVBw9G0QoZfKMMp06TgkYLJY68zG
3qIqrDGfXRVlOF3kwms2rDnwMf1k8gyUEmtT1aV0S12vfmefiWbV6P1oAdYEYUdM
7wiQX8TojWP4J0XrsmA6gq15es4UVth6FOph2ybN+C5ZYa0VTCGiRFsudE1mJofk
dRFx1XVqi27EuQd/4h5/qVFiH+KoVh6USRiP5fwBTcS6XV5eE53rraz21N1c2lMh
5rnZAFRklYy+jWa9CFsmQXR0quc0BaNZ0G4A2LQRMMeLTdpiQWQkFeP2vJ2mIeve
NTI7YyHDfKN8L0GegTF6iZYyQHPyO9ZUmty+IjH7kdGMyxg/soqnuAF7hwnv/7/A
H+/RXvSBsXJM3cogR8TO0jfMHkCxjNQlbDhMtjWT6vbnPtPyQBmFoMKSlrg8364s
dHPlt+NwFshNqSLqGS/SG+IGxOOTahwYt15zE0XqFBHM0yMiinL+d4gwVKkweMDm
Pzy2ILdaq3d+SMIpcDi1u3/SI2rTSOaQ4oNyFU8E8zO3VMSvkguS270PyTGZI7AU
DVmT3C+NHpDkk7mh0S8TZu4jcF4D38YqkhVk/8yauEwwkFHusU2nBuo+jwgBJCo+
qytbbPmO2K/XEX8jL7kCAYE1bcPbwjovHyue371N9ViUET0hZRAQkAM1s/K/Z1td
HL5ZxNQMNzFDqtk0G28wZgIea1Ie+AGglU+n93A0XK16yqKdoXnM8hjOt+8dITs7
rNWINLv1jp8aoF6cspV7guEfC7/TzAVAbs7qKx+/q8reXQubru7a/uufxm771DQd
zmCv6oXYgmIzjMtvNf+vCeNzgvr4pa6UI1t+55vGX/HtiPgWML43mq1VR7PCoYv5
9cgJM/fuuBByW68hCN0YfuUf3jV1pWuyirb7kyeAXqjh7LCZBBSosrzU1GXBc3T3
6oNh4ypwTSjGaoJKRBLXK8mV9NAps63l6ue2j38fzMmYX4wH1C1XuhwmnJX/wOsA
NJrCQrhV1vvsLPlgbLejNcjA4K1ka6MLpusAZiMpxQW4iJ2yzwuijQ7L5GDfh7Zg
R9isYRyvQwpxDIGYc40Q3oJ0aTQVTkXyBsb7Z1hq8gocLsWHKRAmtmQfS1zS9FRK
R+s+MesX/ZgIMBwt226elvVa/KOXjMQyxsLln9Wq6pkYFdy9+GZ9e5mQxtVjqL5w
z2LuxRQ5mouh5+R/xzuPgdUL2hjP5MkVd7JTNvsh5Ko4Lax60Ci14GmN00g3rvSr
yTJarqq2mIoOiYnMfJKJTZcHigAU/91SIcU8NkSvIqMrDzD4TszJ2N8xPA3qSRNi
lpFcxcxrlH8/GQzWAXLS+d0QCoNzhWY+V9pYnVbCkpqeM7HmuJRsRy80XUsq9SI2
ucEPWSaqzJqz+72T4Din2sK1HCFOt2AWqhr+JNATfytN64yjiF3pakAAIlYwCazm
9u4bSLr6REqrjwSZt48faxjBgorbSW7BAqzpM0z2wQ8w5wflc6Uqlv9I3VfkD+RZ
YCUpWw+vCveXAEgd1+wgR+zpJXnuiT3SJ6NoPfkKWyjL1AvHtbYntcihDv2R8Rd0
WkMcZqT9vlX88VHf89jLZ3+yrcvpzaHWJT5/mgHlKyEF+Lct/uRc8xj984u44i4V
LZE0djyVeM8zD2oQtsK55RJjbbwc59+r0zhqwWpC6uXNXfrq58nwFIcYDTe5C53X
9VCT5j9vAEb1uDQza2ePlsEg8OzCfveaQKHchJ86AGGTo0Q8qRLEfbIu9l1b0CCj
+fc7TmXfOJ3KhZ3TwLSuw81mS3OLLAp7PUq9iNp5UzvTLP2p+/O4NFXO0n3NbMr5
jwUDqbhD6RODvYjrTXzHJN1eUrRVSxXbhNnWQH6A7YUrWlpe5C2Ry5WtA0VZElmk
1qGSKdfrDq2rnofcm57n8fWYw4e4NK2WNyQvEIaU8uAzXoJJanI18BuOpPJJ9jEh
U/yCb8MJlk15zd131deKyP8HhXHX1O8OPWywF9VniHdy8Zdyyf2B3+8FMQz2TMOb
JswR89CgmMFmSp3eusHL+e/gafRde54DFubRjbVIauM0TSyDV06X3gJHjbJCsEIl
IZNaD/hyCNTfk/qAZr3qJbdL8uNJisnCpNhm0ewrmNjAYd7Sjjg4R+OFxeercon3
uAHvKPZ7gvFFsZPhBgM52x22AIXVTiD01Qxf+0y5+LpPKRMuJlRn4keoryampH1T
er3qSR1j+7MQR/mGahApgcpW6uPy5GIxuxiBgNA2CJwKOTABkated3PkrS4xyBtr
Kbzsw5gzFNHx2q5nBwGRIZDwqINHxe0McVfC6h64zG9JvF5ptJIIVqOK6a7UV8Qu
Gl0wVm+jBdqaBGd71kHxgdXegCXinpF37+XBoXBgzbU0t49phUD8lbersyMsa8ei
xtJW4BLS8y9MhgAgIEyvZlvIufc2SNz5WTUuJp5N0Xm2TYK1uleGB8FgWNHCK7Bd
3k2CdG/XtNF66x7wRW8jrTP7tKfGZ8h8EhkuYvb8EGBEEQ0gdOEg3UcY26+yrJcM
kaUyx9g/xCpJ2kAWZvIqZWpkN8CdjDS2FFgeTqd79BRmcqjIIEfvE7p1b/LSHnqH
Ss6RbW15I+ZAUtGydFY69u59yIc+RMIfAyvQosP+7Q6EB9Nkjw480hBXTsoTTOe8
E79LxezpESY7KmKZFL111VF8TqN10bdMFGqlgSOudntcRnN68k8GsiofnQO9Q12u
6V5DFlFV6ANWk06uVoJAMXY3tkQmVeh+fqxjgwPFU3YWv6fCjGUd/SbdNyDITbzH
181HX2BQm608fLovJnClJNiMsUqESZQ5Q/v9P7fZIJveMgdsGUjdPzTuOnMt8I6y
Znxxx7hM9Z1jtLXFtaguc1kRwnw5jOL2GnX7zJHrAzyPxbRHqIF9vZZm7Xberv6q
DQxX8N0U9WGh45kl/eH9N3NF7bmR90KZkMJQisi5p+/G9o8kPqj19DU0sBRsxIz+
U5NiXk9DP92nWJ4C6famt3ziYtykmUbjgWIN4cueIohM1xYNnCDSfmkZ9gduBC/u
Q9aigBrzoJuZYIfBXSWEdMXdTduGcy0a1r9qwGZiBbw93HyQqnSP34KjuJrHm+0Z
dliIw+t2Fy6Yezvyy1jgXRJ2dN+kA3NlVR35DjZJozShVY/PIcOEu7BQR/yFAQak
YqJFbLH8D7PrMXi2ygx8LCJoKF2KIpcBPzOuO06dh/jrdS95pdyQC5VOGUp3k1HR
ymoxTDdx347Ij8n3R6oLLB1fxw4yE22t+zY/z0+tNHMapdK509a8lHVa1/Xu44mo
luPVqAf7Mt46EzMOz+u363uHmVsuIZjC3AxtOFQcRE6q2u/ZkEeJ5CKYHMtEgOLE
jBWSgYO0o7k4hTZLuG3HIZxc4ZRNIkrJ49Cc/L7tDmIuNuI6OFH4GIG9Pp4eBtjv
I3BVQ/aNPM+edbie0K/N14fotY8KONkNmKqVmAQBpideFLSfLGo2t0wo0eRgRkwK
XQmpcFmT3QsWKPRgkE5FWxaB6oYaqm6WgsOpBYnIUGbE5xH1RdCb4empa4bdwBBS
EUiQPItfyHrgq1jj2LyjDqmoyPPB8Ta1uebhN3UYIDXWNhMHC762rswC4wQS++Eo
QVqMC9C0MFM8yEF/rSefo65uQD5eQVXHXdAp6wkFjwKwY5dukatqn1LDfcPla7wZ
herhhAi1w0duNu4iiveG2ATJFiruCtDwBwDpXAq6ZiBC+n5FDkPQbBtP0IIrf6a5
q1btC1olmF363Mdf3ybX2Nug1NkR4adjEy5AtKKb0oE1o0LFgpBGzDO/712/uK1A
r3FWP/fJ6foOURLqGXJItI1gFIXftpA+HLqqAEC8nAyghwF4j9vA1D6YEvA1eJqa
5LMY9v0XSE/XU7W2VnMLBM8AST+2slZhmc/YCshEtlpSz+6+CXyRSjoD9zthpojy
OCPgsyPga4rJWZBGIMe6WDa3vy6YXs+yNdtYLw10aek83OMDWBPAq9KWDlQHeglT
2R9HJdoizIZ5ruenUEuLlzLuZ6GpVRRA0KZ491KaE9J4bYmRpsyPF3wnZe3YxQQQ
FeMvIzEcw824dYW5z6LqVIK8i94S6XQITHmF3gvcM5UUncu6WsDRR4AjGPpv6yzI
tgKa2ONNdDmNaixkYxRbeeqen7T5l5sZWvPPhFBKCI7Axwr8FN0W5A/OPVKM9TG0
tUOSDWWMC2eXpDA1RBQMjYJnUsZ0G+W56N6sThXj/zePpb3mPY79V+C6NL/4JA3q
Q+9lkMHnzPTMBVdl7meJUevVBXMnZIm6kg0NWqVchLbipvgdIgbs9DtugiSAkjTT
0+Lugn86zlEtb9K8xo6yTi5BaUUILvJNu5VBPKqJ5KPccZIxTG9BDLuejA+hBvHS
/qxgFDDt7DD73cCJNyrKYNWByXx6S+JKbLhImMPImnQVF52LoGuFXG2HJfz731Bu
8EvSOlcV6zlXqdYN6V7HTM7ySFOnBUt48GkH8u5hFKt4NXEcQoIIckdWmo5cObQi
TaCm/Y6e8zsve8+1Am90GutFHhRpBsxknEf58wbnsGJ2fnhKBWex1Vv5UVcOrIK0
mofI8FYuT5hEqCGS6hFW4Zpxzx+U0hZoNzMGbmUzvTQNsVQwkpgchrcEPvXiHkYo
ph2zbHffcx+VrZNm/LqSbYZ0NTiEby0Nr9SYQfVbPBHzbLsy30Xf8F7KAy8qrWX0
JGFNwkv1Yxw84wjYisG227AEEV53Ab8Ek1Pmip1lYHWAJ0blaVZZsQN28x3vBEvS
dQe9W8nPCiFQuTztsMGaA6PrAHW4Cn0rPTdqabfXanp5sRjB2VLzY2A01ejTA7Cz
K99g8CJejfyrCwOTSW/PzRvIfol9GMUaGLdD7bmkM7CP6ZLUH/smZe8SKX27Qt4k
UxC0UwzrIRMzwCS5ho1ZxR+UhACIZtLWXBd58A0alkClGrjgdtN3PfLZo7cmXMa3
aarjh7EIVsrnrfBU11xZ0XeawSiAkZiVIYsH2CCItslQgmnoWGKs19IIypMvvdUF
Jo9Bj8qE2P6vIETgitbm/3XGvvWdV9QUlH2JnWH+HJY=
`protect END_PROTECTED
