`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqZ5m0ab7linARw+KyR9htOagV6BecQT+1Af4syPkDLtJ+59pEhd8u+OEGJHQayh
gZw5coOygMlZoVVKKw8Z/NqRjdYd6Pg9fGBEQYS0cndF9CslN9uV89/EPSP5OquQ
E8l6ZMe38vA4hjEgT8m/H5QZQIDmEIqh2ZBj//bfAdBonaTmsQLJCKOSISqqVl9j
Z0zx4JPmSR6gSpXZRXIW43ZcXWOhDTqcmdMfSMp+ajYMwcWGkcfWOj8adaVwRkIr
KqnES6hswJQFCWow9iAySA5hT77d1cHkw060noLp2i9lE3LUIMnvQnl3KY+RXlc3
KJdjm2zqp6R9rUxKNR/uuFDy8lub0sPFRyWV5XY9vIbKLZt5x41cE8aHzH6UN6LF
4/w7lcrnRp/MK0OrR6NxOPfWWeQnIvzmxhZcYfbp0UyKiULEsZ45u4yvtrS7j31w
hL0mHXctmbCKOWSpi3WdH3I1+VBGG6gDx6Omp/HOq+I+T7URCzRGABkqGqJyLKOn
`protect END_PROTECTED
