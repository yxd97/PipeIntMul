`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RebSpDEoVHk55r7dEcddlAo+HcAFpq8xIfQHZC4H/cXIjm4cQGyY068xPKVU1Xm4
YBui2o8OLNd3Oa0rxXwOkMHPDa1Qn0wF9KGwLE+tkBwft9EpdPUlNhT3wB2G44/x
eA6OBtjLE9ry9zD8N5fQXzXTAkJxPj9qckuIPpd1O59j1ahmyquwXb4utbv1xmLM
ZjMaxUFZ81cXtvf6FAM/Pce4/IWo5K0Ci5T4aXUJsBVWyutD2o97bARQuO3AUPPs
Z0a67JVySvSkUTELzk8GQmD/Qcyxs4dMTMDlVmZjtiLHygeoQactmGDVdFkA9B4d
f+ZMBBsl41hQWPGkVsvH+jLPQjnfciPJQCgDTYt8CUKsVKjm3loy7Cz+hOKuUPkB
T9/nxiRAN5GQFjkeI9oEI9dtR7bEeDLBmJkTsQR7ldB2x2Q5h2BAzhbuuZOIoG+r
NctcS+sfnrsoCyw0eCA/igeVHlp5ELJidgpC5XGpemgA7A9zTzsobpVK8EYO6Xdm
jvZRop3SCu5dHs6J5fGRUGll1BJYdbujHDXtTvJ7GK2xpShoc6Pam78ApfUAKQ49
B6pZUxfA4c8ZaCK1+WT6AWI5LMF2lbtHvy5/Elj2lJjppajTZQ9smoGZbuNXZ/bx
A4c1Joq47wJ+vSadGMwMvVx8cbSGnEDFlNOUnC5TNPrvaP4iHZUcvYL7m1b2c77B
hEl8irD8O5GKPTIDiOdw3LUSvwzVWtIMnk7qjAZKdeXM6s+kAjvP+LtHcceqhE0B
dgeryY2ZAMMKudj9L1jFMnKePbEK9zWq9fli8CIjcdudA67hEK4dA7NT844wuAh3
nNFsOBIp0WbggcptzzxoOVHQSa/J1IWvam3FB3zDxnhxdj1oJ0GIH2moOYgtFLsn
vnh7o0pu0dLh0sTBhGMfk5NunMBSLd8TQDwfohHe7ep5c0rD56psv0ccIccUFtWU
I7JJOik4IU7p6EUKC9yuJ/5V/xz0o3Jiyu9pjFqgam6Xv5j0KOhvdHlT36LC37j9
Sdyvyd76RDCVlQRQM+l0yrduQyFMzX96kPR2ZXotljeq5d8IcTtVHAzcgmgGYDMz
oCXLvT0oO9EABGxbUfwtiaUPenzv0yIjBdPtp1RV81+kuA0JnG/ifdmZouGZjVuA
Jqt33YU+F2ODeZ18bpACbjLVJjsmKKMc+lDXZjZR75Y1lsq6wsDHk9z9sLM5nRKN
elzeogrtQork6SooCbAD8zk5yOrBnBTrKuFS8GDl3iSZMCj+jVScv0TF6YWnCNsV
nSjiKuEUGH6JaXxhRtD029G4rF5skaAGPeZJ8v/luEQbwGeT5rgPMj0TaOLN1qZE
cJuZM8A4QLVLSEwYKBtsF9zFKyNnc/Dpb/JDHwvME/dK+j6xnvBU+rZ/bXTVN/Bu
3XefZNs2NLNUlYsIn7Qz6Sd8EEoArO79TNr4d/JlPHqTN8zdfaia/wIxPQ3zypNm
oWg7W70aMndQx+XZ3vROxl+jYybxtk2onqUXe9RbQw5G7pHVG7pGMEz+Bq6zu4Ub
XEKHDOB99KQXVIcz9+/Lse6rDh/DLUk3jAHNRbjANW/hCco+VCi3/E9DnfxA7kM2
Mc0D6dP8atYZJDW+5qU4utqi5CqzUPYaA/gWvfZ6C4yPzzCG1DDqbhbr04D2wLF9
w6w7S2HcmjoKavFiMiUOwSv4g6pWOFXAvQU3Yrq/cLxzJW14TPRxUAcF+HNG4LpX
wpE5MwAOGUUF6Uq/QbNn0foYwuzzxim5Ib8fGqX0kKJvdS9tVoAmuhVmzht09u1Q
yQ6zmZ1it8g2MSNX4ys9b+nVDE/RwOTILJ1DdGuu8pkjpoggeokTSN2MneHS+wVq
V01MAf6niaN9Oa+lwQLAG3NyPA7ptr84iRM3oIZkRXg9K75MS2uSk9xkbrYD/zzn
iOmps7xlL1KlTroI8sqRSNS/7jMxFDPYkAf4vjWad9ITA0UVkTyUkEuQNND63jMF
4l6QSL0VJfyhXaxjAP6hLTTEy4dHzeyFSpE/ago/nWLdFbaZytay6n5k1XdwdAmC
oqTF2GsgzElFUOCQZpKnAsty4dChaSi5NmFGrb+m2KNN0f7wDPl7jf4BMAd7c30Y
bj2JAXgrATuktNnH+SQWH7RWdZ9YZNQJP+zuRdneaGmYCxh05/5HXZpWpt/08A+p
9GxtVbKWOHFXYpm4E6fQZnYIKawTxDuCNh32ME0InoqjdWhFP7sZFzxIAZfjkLST
zbfWjKg8LGCRyHV1g/JX9ceP9pAqHwl045an6jRy5b4lk34a6AfGJo3W4aLvXxwj
dlZ2GTXNJhhnxzcbA281pyVolWqxmuPYMfCg/jkp0aEOV18+Xw6ego7R2mHGRJM0
H6OcxrdwuPIqwjujtdr+RTowM5qa283bzgaW6L0vQmzBO3+xv0QWbGzv7cYkwro6
pL33tTIQUl6CZEPb0wKdKOI8Rt2G4yQD93MYvZKLlaA33koJgnXTUqayBF9/Q4Zg
5ZSQZemdsvfer+e8CiTJ2d3EE5mq+ghAOfQYAsQcmFiFEai3XUpl05nOCmkBFQy6
1yl+4GxPtmQvEN7QNEmQT+kHZbDUOw/ldeTKoo5wtzq6vfGOW2gvGboQ9t7x7AFq
x5UE01m89nvuRuJl7YAakz3dCFZf9jqQNARy93uYtdfMCpSOrMPCU+WUwcfNqSgn
COqhEol6t5HASsb53C0EF2c3XtNl1kOFsR/5o4QjR4SNPnvwloBSbTtnleu/YpA5
HJmEPpiyNVGtGshziYjYOg6rlioWb1qgTRJF96SUWsTa3Y/Ce3QN4WwwzzXzwySn
f6Xc6ng47TaZwO29YSmwjZm0fLJJH7hA+fP3umjf2zb/18pJjIBzIbRlhnPoasz3
a2vspC9VoIadgRpTm6es7ui+23j17aoINzw69r4cIIYGfNqm5yFmomhH1U0qC4j3
xWUAy34bPWjaAa5klFoLZ+XVpMfp/K6mFX1MZ74odmseJw0B9CwidhzynzmqsASD
cbnDjPvIM0jjyTdbc85R4uM2BlMdOfhgCgpTF/1rTPqLACCL44eFaMdUR+wpkO4Q
NuABl/uSi/UwyaW2KvtOVsoYBJjIuMSlgPtNUgKaEIzMv8CvFBhYDZZJvg5bc+K4
Lj9I3NOgwiJs3+Ean9Xk5tV+wHtkWAaBeRzQeg2Fm0EZsDkVbloLknzH5t1m7bc0
ip2Ot50onubpRt99YOWmxiqYJqae5MRBIH1v9ubZD8k7s4ufEK6YozDYERoYrrIU
8uySMnB1Abu/JYhyhxJkaQ+IoXa21t3nTfTd32E7ndGweCwEYOh5OnWA9MBVHKWx
5Vm9aE7ZOwIjgly3L7OrR3BEX9y+9pXIxK1wuiVEbpV30DmhQoOgRfCBVbxF6MD4
0xAQnjpfUvVcncGp3PlmmRwM7bBBzelAyOeiHboRUDAKpK92DM/h/+WvVZMy5uOE
lo/rXPWBqgozLatADR2yyZtB4OQj47j5B6i42/xcOTfMlSO1nrOFbayxTUpd6sQ0
wuJMr+i2FReX/2LqwTRgwe14fH92PCAjRJZq2qDACUucM7/Du58qQnoa/KPJENjA
pxqd32p0NKa0xmk9GMHX2kdFHVDKcCa4baE/tgZ/3Lpf4ijAZvyS9uCnAHtYtzXo
V/kVGA7TkAdPoXzVfh3fCCJfas918nUWpLKpuNxKJ4NZ5ZokIrs1uZjm+SNZh/W5
yDwMFq+tTDTc1QfBH1jxNkzo2rDRncO8GXrxk7mOFI6len3somVXPDLV2Ts7pGdF
cYKgqxryIvHYlZEVqVHPuWMHt7/Ysgnnn5+6e0JC3NKdJ+c9G0grsN6E8E5n4648
VA8yb4nUXPxz4jIqPYa7SBxhI6AtdBZ0bL/L9jchmjhXOGv+2jL0Y82iGmmrZU5p
2bJtarwP/oySrDewQWPl7x8+Ch19JSn1mxP0/jN/F0IV5L0GWt2oSAugGq6sefm6
DdT8sD1+0Nf2+2V+ftuPDMdYIg1Ne6oA3ZbSyJLANN6W1q914J7q2HJbQyasTQg6
A/6JdzxdXUk/DdxsOhB5CqrFypSyjHsHQjohjWdCmHPODMYGyFxsgY40sc7bDTm6
52Uawjwifi4bK74jXltkY6Xwuqrx+HBembfuOKRW3+aBomHOm/4F+bc6DULmpKOy
u/ujC9MbhgtCNB8mlkbCpa5PPt7xpgfgLwv9gs44mlkUGL4uhs43S3Rm0oNKkLq5
MymqafAB6Q81p14wedskd1Q2xsQPQC2mqZo1B+1r0rKbeC4o1R6ue2QY843o0daa
UxJZmfjqQx1koIDm/rvtNmX0VDbRiEXag1lWqnGtnFkQUZpACWUhYkd5k0e0PJ7k
B+KnTlgXR49DYoeyOdG0AOm0YRPiZgbDb0ROzYjX1VOBcHlb1wu0eCyMDQtBqhq3
hMcxO9fyx+X4Qi9NdvxaO0mJqpmYt92VFU7kM918u6l4/3zduQPWYDAVQBGHnYCg
BlmKw5gsP8ccjSXLJ91XARqTvOBa4BpIwKTXl6a5aYT675ARJmGTCksFu24IHcXr
nBHs0j0prfcYi/RIyyLtdlesq240MDP8nHWiPumAP9/rF6PvMSB2QYmJHEnPcRce
LEuxUbe34//CURjckTxV61jHGnRFDjv9ZoWA/tt0oS7SJG69uhmJjEe53EkPYDce
wH37GrkJblfd7Bc2pUlSmg1Qh4/SkGH5DEZTUJhaDyV8Ta61CEixfmFm/TlCuqg8
fS+3FUkKkhnYJTup9zuysVmW1MYgYN3DTWZTpJMn0zknRxyseeOUEEBobcSsQLSm
iWNX8talPQs1V9IeZ9NNnP1gYJGCn+myvRhZXOGuMtS4fPV5Pn+LhIvfbNVcInvq
L+RCZKF40U5Y2x2ZMuLEWQ+ZWJnavGQJBKsNBJZZ3iDOlrhHxY4PqPsM9e4Cl826
Hj107STVhPqVVX1/FQu1XhCioDJOI3z8z52nal6FzxZfBJTkoHLU+pPfMoz90fPq
pxAX5OAbys7iPBcVd0m6ZBy2jrNYSUfT/F/x+qwVwzYj5ylIEAjX4llkmAK32qgb
uLhR38qj9QbeMZDPhBvs+ZRkervsaFi8zGt8KYaveoY9QYUBQ4/tqkQCsu985cl7
Ad7rTF7TodvveZ1FlqRFrb0jCTDaY1j83XytvResUDdqL/h5oy4fjYE/cEBHpC5U
LLHofpet1aJJKyYyJN1rmrNRGhf8638fCk0+EXIQkj6tg8SLJYYtsrxdLOx/id+g
LlRVluJTpLu2yMDG0U3LJvAC+XpboHeYyaIewAV5bJVyPbuL2p64VOEcYGb4iepp
EQtB3CtiI78nTO01fa318OkTI6zQoudUmtD2Ct5oogNor5T2i0wnyfWjeLWcV9oy
NubM6VyeQLdlQSk7k1v3eGkJWRMEbgGy20L5mKg3GGTJDnn7Jy50xAbvAsI4rJbK
J7shRNpmlRvZ7Jv2RygBWK02IG55tRtogTJdNpNmTibJRyrKc4i6h/1Wmjv9Fy+o
/ujRY/tJYpCMWsEOMuBhW7i3NZUtVZXp1icCzeiE7/wfeR8LZIVJfQzuhIfZ88ky
hsyNGSWeWWiGcWOdIOHzKt3cx+CH8oU/vCfJV4b0g1xQdbENWLr+i9w1XPp9tKVP
poMNZGUVQtvP9OiI6KXFW8hTfhWJroEKtFInBBMeYn3o4f+DZQ1hSpN2zmZxccGu
o/anwTUIrgK714p/lFnXaUYGRQZkYZCmT03wIudhmEwvFgFUBRuiGiFy6pmmLJdV
YWdn85EX9j+xRcGkdaECltADr2MjRlpaeSFuNinu1b1yfYb9WX7Y5N8PDePYTC1o
vPJM8YIw2cm4UiYz2SLgH60CJzF8/hB/Xfa5hQChEVDGyarBkgZySzxY4CxgJ1mw
vxscMLCG3jQSzSZcPwt0K+ZjiAaodOnORsansbDzZbvSZJwmEmYEzxQkNu44yAaH
DrcEMLQfw0aayGhkkCFBtcxMq6oDr5nGBOp0Gr/qHm4rCigKnc/sKwyYRyy2hpLD
HqEbHFqq6ljn490AAlDVcHLhuweSMvRwrIqJUD91Nxuy+OElcqmnoSvH5W9I9Ph/
SmfqazIiL/B7iKaXFZel4c6a/bjwat4Dt5UIMqX1brcNhai0qsPdhhFPK7XN9TGK
YJWvFNj4S+Rame6aGTOif32mlD7f8i8uIN9CUezo3bdntEpMwabgxQzixQeGIvic
h+e55NbPm5sbxAvE01VikF+iQII2rDtVmixIwkezloiCUUYGxKXcF3QkRRc94G5U
vbanQi1NFkfoNILRIKupRI6NhaGWAX7143THleNptDd2eXrl2XZRJ955xgdLx2ba
6O2KvNa/M7PQTFPS0OCv/loB2RMZcA8uV/kntGvmyUl6xaYm6+Zq8UcbSSrKBxwk
AQojXoYgeqWZUDi7AQ7M8EFc1byKdLi2q8hy2FVX+9SAvG7zZQTAkT+P4oOSyaNk
9gdIkkamoRx1p3bDI1iFIB6nj1NJ1ZOU6Fc/SEHIdsJ6ySuXa8DVLL1j+Eq1Z8Xo
K4kiJcCNE3YywpDCM8SATKYSCFUTyWrlAEhUAKWKzcKXFGFZA1z9xF1kqa3amiCT
LIgankiOSwbUpstQ5z9ddcXvrE+qs1dM0aLWvqnyDwi3JNJnEfNTdij3gp2uuTwK
2wdkJ6c5/UcS5s+pNBAi7KlOsS910XhEIA+STLsqHfA=
`protect END_PROTECTED
