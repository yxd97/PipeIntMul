`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0zTICNZA/A5kpk8ABr8tSbzcUvebQJwpGaCZIemJeAHMpr1kZ46eDu7pNerIdqU2
55LavwhuejGDSlzPY8eACwqwQe59Gd8+m4KhKW0njNy4TmiI2XkkrI8m/rJdcvL4
DZvkEy3/gLr2a70S92c8GyJo5NJcnxvVSPF3KkCVcmWfQx0kRJ+/5t7yPrSF/TD2
aaf6H4S3mYQtLNtCe1GeS5wpYZSVwSzf1tA+EL+ex20fn+CIpZ/HKgHGnesfUJb0
26A/of4FVdC2kX15E5lAyi8t3um0k4s4FkCtaC0fQBCzb0izNUeTt6f/s57wofaY
yIW/FT9vkmbzK9ddVIudWeYwepUsNmI5tmENScMqykNstCwbgcjw3MaJ8MeeO036
Vv5Ruqqi9jKPAmUasUJHDf4HYyjprItUkcEAWvojYYe9AuGLXtbE2sUh0dLo2XFt
hs+bzUDkup1aAeDaTBYUIaR9KG6FAaSUoMRj5B57ZwDS/8WBfReuNoFaAa2CD0Ut
UyWt5FxMG7xAt7UXa0baQwxsGG/eR/hFA1ZBM2YXy3ttcfSXbufD5o96SvEMRtv1
mCkGbtNG8JrCG4YQG4h/mgcVXBp5tlBu5Ca3gtGRsm76HwGr/I4onycrRW5QXn/L
bWV1+4o/U/ydz4uO94qxXxhwXsBqdF/Thg63AYjHOsWVdLGbDESo8+CTK4OKJYIy
oGtlxoER4lZOv3/ibk4PbKEi6wSHcm05SFHndr1L3Xacb9eGcZX6k88g+o/AH9RT
n+5OL8CwGPlOLyHJ2RNkBA+yd687FBwe8fuT7j3nYL+xMN6nAQO4pK1xN9i1jW/z
R+CPZ+/ixrmLpu+3HDmFPlXuo5xbTStftWJtFhQMpnbPtKHNP0heD3O4OBoP2Xi4
E+p8zLEoiRMr8jZNHmr5PgX6GP1h0gEL4AuSYlHKtb2dFdbUzGOjuoF/+x8CyunI
Fki7zHFL9ZRpKsW25IN51rFRpnceuk7uBfcwuQ3gEdLrjqN04uD3Du8po60vjbct
Qus5869uVOvbUcoLTrSsk7vpVasnsU6Jq0/it3cynIJHJ6YUVp8PmPDmp6MsaVpU
l9IoKa04jv3aocD6lKVaicuLMFwjD5itF0cRZ1vvWT3qQF/JO0kSRBZsGs3c6kgk
06+WHtn4fsp5jZbxWKG2KW4SHswLWloECQGsEKn3did6o7OSVybBcj7NLkwWOS6d
kIaGh5mN6iEoKeJrQrjMO1U56El20o3syQUxZ5wtOANUgknNnafx1x5pCyK8ouVw
AjEd4HIjCZ0XtsDT02pmyea0YkIxO6UP/IMshML/aKuOMWZtEtpGMJ2aoiJFEbe+
KlrzANutO3vD2XVWTjJ+PaJMxaZqZBTN3jtaMnqNNHU+czuvA4UC0qsAEa0ja/+m
uRz7N5CVbheVRvxj/uamgTVKWWrToXLZpqg2bb2xZUwd4BodQDtWljLXoJbYc4pi
1cGsDM22IdUc8egAXLtIzZgQWhFWBn+bh3er4DZudqFlqBVT0gPKrMK4+z1MvGaa
z9MsXcijsrTBL5pM/yaukpxbHjd7TvJap1179zzCCjnIqsz+Q7iA8N1mQZyIra1v
9Jjy00ypSQEtUJzaw5GU/UBVnflhGZWfVeUh7uYqBmx61BFmnmeuhAQ8WcA/cM6V
lKY43pOdzK6LmAnQo6N5B8UYnTfb6ZfEAz9HrqnAdgotV0rhsqNoQXNtIHkczeQs
z8Rl5zI8pKm35Fnd+tu8oFnsOBkA057eluHO83d30t3zGLz+f8sltcHrW8K6+/Yu
tdbxd5A1k48dv413KYx63zW1U+ajP2eHA5MOQkcOD9YxtH/idspstBCkwe9xnr9G
+Wr9dFz7SbSpVwmyc6+DvdVN9XQvzgGezclDRLc9tGHWfI/gu8C3/4yqRhod22k2
4evXQAI/tiaKfJAsE4K/mnKw7st+6EVW7Te1VmYx9kjLGM0p+jTz1q8gUdBk6jox
JwreS97xn8r4mf8aNyyZJhS9RyFKQ1babxSCdNO5ClfYiE5GIIE0qslt5ZlwR1s8
L/skBXAmaD7Ov70fssgDdUUdMOIyxX12YYQsCchYy0HvnfvJ9FMXWfdc47nZhs08
Z90aGIaD9nd1zkmaTSWscYESQ6Fpkd/VilZwaxtDcUGSpb6QMI8xJxH12DTJ/DOf
tdmtevhw1QI3vQ/4zgAnKDiKv0oGWILVAECPAt5JuWRpnr/6vFn6khA9TkZtIjdR
OctB3CRwxuCS5TmrRD6b1oJgLq1fLQdUHgXUTh7CLKpWMqWpmUhdrhVJPvpNn4Ms
ZniCZOzG5iFJlgHCKYjGUiEXdd3dyRWuNdoYX2qALmN8guUayZ/wjFf5t8ZYQ93Z
rw9sisUBZ2yJow8qIX4SdLXK0I2pOaz8ZdGMXYDW4RjUDK+f1gZopC4MiW/xQ7Pr
tpS3YUz0XfVVN92wPX+g4iwbGBFmliaz15l+fEwDxadJNvWFvLeNYuAuHCdQEzgY
BpjzSEhJ7Df8dktymX2PONrOEDvmLrbKucYpYXzpDJnvJY3Dfr6KOBkgOUD7ZqEW
xnYW06nvJeTd7y81fbZpQazWtTMnv4Slxb9Gv3sd3njiG0wHacE2fec08StCD1jN
0/3b74zWDy1Ne2Zmj3p8oNUnjmYbluzDR49c+xq2Ujjx63J7g+otdh6JkuFkbdu2
/JfpEx3mv0B+ParpYbEkH6NLIK47Oc0Zi18NtbzwfsXUoC6GZaVNVWrhmYb7lEVf
OdTzU0sinlmVzOwLoznXU+vllqI2AfJlVBUtCVqNzOVwq1094quggWTZim/WaWFH
i11zkaSyAmVR+y0yj1RTb5KgJq0vIsCWPNjJIW9j2iQdPw4nFcDRxpIQPgeqWMFo
aBfwAeMfKcAt3XX49CFogy+l02QrYAY/xZzILGd1AD8g2pm4Livp6tFCuJ8xp8f0
xncdBN7LabsBimIJmzIHObHF7a9o0uz6QPBqtdq2ZQeKmDyCqNKZRY6JkFnkpw9D
6IRUa9NYCrNaGZhW/ZVBCpEuc8kD3bqb7wLwUakp54udzDdz5ROVr0wZnL27DAQC
jGyGGdYdPuVULEK3Y7CapQUB8zDbSM1jxaweAuMLSRemH/E+Bcd0fp+GsFBQ/+VN
/2SZRbupvPXXU+bGAu1NBMdtXtLLBkhBhfYNWSZP7Zq6BmTevNf6UwaVD9tQ57hY
wYhFlC+lZnOq9jiukre/jQJutYhLBKLFinZN+4a/mm3Q9MRZgCAyCtPd0i1YxVYN
8h9eKwZJ4q/QMTX5tGZOY9tZxz0oL6wYLyzVmuskKhbb5wKfGpw3fN6AHnKniX7u
H1kQRdSIrqh5k+9D/yJfQT1zJF6g/338RdAMoBIWx4FWK5qxaW/5Kd20rpWmLOak
3dqEYR4mrQDKZwJqgKwPZKXqKKoG2tmAgPxyPBk1OSVXriD4oGAJuPxo7yPxiui/
XjVK4BEQOikvs8TiVSdovrM5mGk2Nf6S5AFufuf3ON/vcCKKadZ+o+W4dRYiEZn3
fZ4ujIr9Su+7xh8h1AhBlip6ygIYRUTvU1HxST69HZmf1hCrkuUFYWS6+PXc8Nvo
GZf1NJidIle8XvjTvTvg0/5Ja6st0NyfI0Uu27tZmTxECvPSY5r0So/YhZrCkgZj
iBvR37POsW6b2VzYKzufGNuCvMklwFB0bJlu8qoI7Rt59IPPEFZm651BQHpTuoip
PIBN27ogAh3hoFIu965PpwOQBSkDp416+opg4356AkzWP0R0LIxC4batxGZsC2bb
MlAhbW9M/GQsEWoJjE2YgNnygBLz7pw6YXdlNwuUQycH5lRVwcFmCN9ZQkUmsbLR
w9KNsHZbkLe2IlJAk7sbKs0qFAQhO4OL6DMFURZGYWbnkSBc4iFY6PuKVzIk3mPs
WeBdujujia5cPb4MHkWgSLdYk46Zr9vdjqR8/W1t1R4mP8b80HusSgg8OsAeNLFZ
XKW5B9Ss3kbebgdd16CVS3DeklqGrzJ/Ui1CSx5cZfjQ2OjuQM7/cupyeQD5z0uU
D3pe5gtLNpo+1TEUrmvfRZDX6d5DsSR9w5b/y5HxCqCWQwE1h4CTJHINTrnTVaJr
eXkncOAXmzuQhijCBRqqZtasabKrBgELP6GYbCh4Iaj3qMBPKeljPfd6/O54JMPu
exbYvWVs04LxqfC2pMiLYlWPNDh0l4qCveSBj3OqMDTVptk5yahXgA6zxptyYOUv
4tsekRucZlhOnqJZ98s9IqQnuIcf2uWFoQT4W8AD6v15voLkG8Uv4Vo01ZNCfYtn
KI8UGMrvJlt8qLT5IFBWA2nGPyeP7823aV+WZTnBEmsp2XvYgRyzytZ0zoipcGha
jpKogA0MbaiilyUCaiZnYZam3a+XJ3oOM/hCoyKRNuqr5AJ4HWgSeyeNZplTbqpd
VVhv8YgNWLzlGDCDwupVAjSEePWwYyvcurCcevnwncBKzDPkpTTMwDhruIGT5q6+
wM4GpAedB7nXQ7snxCvvGf7KV2VkoplxiY0AxLqPaQahrcP+xhbWs5UuAPT22hPS
08KJzLuzFhsdC3uzwb15qXtRFepVKE8DlVwiTTqKVzsc6AUZ5CdkKoLBqs7DBgg1
0NDdlcG8YRo/HCOQph8IvbF/N0MuRcHsEpgwAgJlVjrZtfu5V82A2n3I1IwM8dST
oKdMTahhpYkZG52bAZJPXwC4+mVo+iT2WtXasQewVtAOVZwGsRSS3vTQ1Sty8jZR
CdKWVzlVzq/X2LN+o5WYYgYpZyyDkZvHnPmn3s/sBzIUwOrW0EQy4ilNxgX5UBN4
peFGYHjpUVKMgRsjUIxi7o7eHkQahH8pJIjjuhLaRhBQATIT/Fv9baBaKTmBvRUx
Sa4ZWcvqlWpMGWFNAZOBfd0MsVitg58yvtAcRA+gMbGN7v7xDeD++6l7BuWjmcKQ
6ekiXaBHBEfAtq8U0sMovARoIJ3KwAllrOnHpZH5/9OjNJstdJ1yzKDg7KjCLwCd
wI+lzRSoOTHP+sVUUFs/sOhhpCrQMdKWZnaE+RCIGFfwcc+/eDGNonQu2FYBQC5m
LSNpsw6FgGHM9RKwmCShXeDzIOpPEg7y6P+4fuRdW65VT8eBmVs/dA78F24YpYX4
MlBU2sb7vIHofuK48dRAf878zmgIBqFK3gEXIZms2cwH2shdR3AacC9egZKTzfBA
DZi+3EcqzmAGZZvzG8SYnvqNpP9F8JUmflBtP2O/SsPsz8SokQgbQ6YzVONF+q5U
PH5YGqHWEEErWCAL/5jK/EX8q2QnM9Nj1J1MXVGcVZOSsa43uxL3wA3zTSq5qdOF
AOKy42hhIE10R+kGrefw5wfV90QF06OEEAhdlARRgExyB20fGp4O5Hf5qSiuIeae
RRnYgshZWO0rJmN5vnHhDFOUcx0S76bjLIGKFNE+4DClyRD2r5U1haBMJYJPQmm5
BcgrDU3p18bi5cUETA/HOim3q72wIjxhHnb5fDWb5AyvyJqHESFrwO4Pi4r/3wyQ
I5BXIuvggXTkiUFrZkpZID75qAfDzj/vlqits6DwMpRJWgY4BZMdRF/qWTM0aNRI
vMKq+C3ojzy+3TOYVV081VrZ2INxEnRMcgL8s7bMNvZ93mD3Y8EHkiqucx1Z7mvn
hyt6xddJ5eQ1Vy45iV+7npAhPJaBTJK1mOMWs4wdjJ/sCWnqUBpaNbYKrPNaxtim
SkC3ZFeFPK4Iq81H0IrBApJX+GTYrAGBhRcjJ7tGWCk8OWAllJ3pTF0+V4rxmymr
VGkN1uz5JXaJ7IHxPdCQu2mdL4znzdgjjUxpBi5bQPp/jAnIVfBLPm5QlWMtyeD3
eV243g6oZYQbgmjqNYa+RmnDfnaZBlQSiNdpTRNDAb6IXH/6o22bCYgrjuGa/yFa
I5alAo1FixVwV7KP9jhcQychTum9IpIcpk/aWUENQbUSkOfbOoTEJLsAPEkUqsqi
pZqaEqJ2m3H2TeABCTDUtL0AYu2ntifGHZ4qRA0/0/Lp9ihPwbC5+V4uqDWHeMIy
FqCPUU94M01McqDGPSRqPquIqeagubJs8oIlpZ+QTuyQDXS5eoewz6HjqgNKLwPi
wwRAx2OEqdcVPHoccVjd3qlxVxd12sQYvmqNC/uKseNq9eiDWb9MTf1JfDlmUp3i
S/3BLpxw3vhP8Dgn1h9d7h/mi+lJmWsmEuqblih1evh2ojAoJIuPZCvOtsZiz156
XlZ/TE62qWJwX0mo+rBFDJDOmjwQW8Tla3cT7dMFzGompO5TuWFupVBs7HONocV2
GDrP/kOcJpkt7/yab6I1F9BS2fVfCKtIEO3uMYiqcsAnNy9l7KU1JDMA0IOb58Kj
IgKKIAC7pZno8BqLxz1RP52XoOfy7x+oSVIYETP8EeFQwKA1wKWiZ5Jfw0xJ+v/T
zDP8fTH3LO4xxWpCbpgKlvqGK+TH8/a7hF4FB3TCJKYrPDKDnelSdvBmfB0RV8TZ
Nm/kNaTnNfC+R3oJy5S3CByUxOd4Xc4GN1nV+82v3kETzUMEkSD+u1ll8zYXE8Ze
GzlUDz5EvDbSy1lNo74QwSXtAlyYZnJhOnd2I8vpPzT1Nc+KyK/fUwIK0aPZEDde
MiGZ+fG5xnd7V+/7XtPYBXzJzoSMaaUcqudQP6EmyVpT2Q+/djxoKY9w2cBsyHGe
UMaB28xRl7flVr0l/XaqYheRGOSjhUmIlWf7AGMMm4dmX+dTdDZKaLpTuL/m4Oe8
pVelQAhx44BS/Po8fkGvVyJk8MAF4cMWDcUo2JX3VHgj4P3KV7cHD/3/oXSjD9rQ
+N0DHe+EqdRMP9O8txGjpMZTF4VKX2g5sStpUkDah5WbMyr7bBJodxSgjXTzCtSf
r8DJs68IQuFVZA37TzbjzMHHHsuj6DbD4kNb5OD4P0mNWDXVKmhoCtI3PBHjkL6Y
bCgEgaLO1Lsp4cwl9BhmK4qnMTVaaM38rc2zfVNMjlWgaabl1QCdvR55YGt8AQhu
fQFQ0Oqde8CPdI3cwBWEM15dVana8TXV6LIqEfsvofM1O3aIHHiX3aByAwPuqqc6
L/ZxquotBw1/LW6BIU7iXGBESe7nt0YrZHY19tnKm4jzjoh8TrjWDpVdvuLGXJ42
jTzhWZ9dkvYJFStgkWMnc442v5q8xVeBi64+6H3AfQz4E5k2uFHoblV5HLIHAOEj
Sko+rWdltYlOOTjZxxz+ak8T1LFsMyejmVw+XxVisCfe42ZtLJcB2PKjjhlycwT5
8E/OfPaBwuOqrC0bhNcvVYTPyWdZzPuk7b5wOUIXLl+KNY2+pyBfzUttVnou1uPu
222F/uwPSRt+zm9HyT8cVen5YEAaMZAkwifgEv9ZvqIxlUnJJ7/2XQDDQ0N9o+mm
UZRCqAJuXK29+hFfT6AX4HDnc0KmNr5MBubSke9FA5CW9k7dsoCF/0j9FCMfR+ND
T7HBoVgwlbNOWkT0KmYN4xSjSV/wSmezlAWOIbY3H+GqejuXpZE4d50lJq0rgHyI
TcVllflJklxRf1LixWTyUU/OODqmI+tlNcxBv2uTjVgQhPxWuZkkpodfgdYX80Yb
/pdXoILbYiytUR7nY5Kiq21jwPahfq8CjfC+2J+GtDustCibjWetvRJu6Y20mrPs
PY2rnCwqtQ2wcPOzCqoNRVPgmCz845cIl3cKQ0je0jL1TOGXri1oh/zlcKuQWwg8
MJ7C3VRmpcAcBkWnjsb4ejjds+MGziq2C/oU1dcJo+8uwnvLcK9cLiQ1FuoRFeMv
jhU41eXIovKpPrrofbEficejLK7SneDBoa6uwNmrR1/Dc710fa0yjNviLKWB9FKp
avbUYpyUcKHh9eOrL24ebF6SKUPkiqgRHGq6rah00kcoAnXhO6Uqu/4bbLaAeloQ
h5fH7UU1Sn07TCSf4k1OFA4lmjb31H3nzR0nfyj/sog7WYaTuN64icMDNjMm5Pag
QpaIKoeN27tVm0rvFeTNJPs7kobCk2o/7R0Z6BNCjeqnyYbFFDngChYwHSAGnb4R
ufv7BiLQGQJk5XA43sdL0wofnPbT+nPCEBdmQ5pKa95KqjW+z66S4s6/SQaDX0Bd
6deOPpTtj5lEWBAM+Kh0+oibwxbIAdweG/Uu2Pc24EPA0rfyWDZk4sPXUzBw9yES
0HWadv7Thhn16XcWHhYcxE2p2gSddMxmaLPX7smmo/0WsJ5SBtnQ6KTj14Zd1Txi
gewDUIzfgBRnWXoU3gbgaRXKlEPvF2xU7kSMekSRgp7XeB57yvtl3LGuUvbaaANO
Y+eTqtLrajjaE1br7zwecqTd/z9G/uftmNMN4D/65vkVfEsP0ctz4NPfiwzfNZr/
kjDfNTpLnGyW1z6++pGkjHVM6WxUXNhrGHojg4oemaLu+lKxkreWzfiIJD05nbqs
Yv18qu7oA8dVfJQ1Zy7vUrQPwYXGJd5ehOnHQY5NSlLy1406EButuL74Mzf8vEUM
PLhycrz3CpCv7FEEtG1dYI8jmUDHyODIeFZIhzoRo6ckag21d5urZN8AVTtsaD5Q
ckjBIBEv/OhFB0+feOh2nQDeT2xJZ7Cw2vIwGDTeHkjAwUUy/852Wm6ae0KnWmZm
lf98V1I2IQCocNlhVh1xBf8JYEZ0DXzTLihijVjlqT6M85jJ8I3pn4S4e/285igZ
tyhluBn9bGW6eN7Si7Eqpy92S12mCYQJNQydEoiCh0Jg1qpPt1Vpyh1tzSZZvrU8
0w2HYOfhsb8xNtvIOdx73mr+nOB2Gk+eRrI+qvkOJwifLaXeyXZJ5xtgwjYeHZO9
H+/hnEA/Jc3LlHzym28/VlvmBvQsxQzqAuf/51V9RLcdiLxsOukuhba6OiJpW7nx
jz9VtJYNkvOM0qoHGsPmFA==
`protect END_PROTECTED
