`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
04ioIiaa6Sn79sMqlFUxlmsBg9Gq7oI1IGz6SZcqMRXrnvBHen08JltBsXuUg19x
vEcRCWFYGb3MVAB+RaApTf1Igr+5i7MC78n1UZ2wMryWy8jmcpsIX/Z1gLqoR3wB
BDFTW8ynwNQYxUIFVw+575Z5aFg19QZHH9v1ubu+neeBN++c1j6GqusP+p35mw61
O2KL2j9dK44fU1H0gCQlLkLlEnjofZZsabToC3zVHwjpDU24/Fl63aQ5eXfMPNS/
ZchV0cb/P6CLGawOkHEFBAjI1qjMTa+NwgNQc2F23SQ0vQF04NmRiWk0PW5TzNhk
+z70qWL5DuKAmt68Ix6Xaw==
`protect END_PROTECTED
