`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Touh+09HtvfBoGM8/iB6W3hU6UlFFgyAO9ZdYmSZsvqt6PBR0dDh2KTU7dGeVCPz
8wWMwd7ZPdyZuN48PV4bXWYkzfDcfv+bTY24NECgWuHXTUcUHbG1fauBANbiCDjk
tmc/ypfMvUyXp2fGEmv4/iBgNbXAopN/lfCPQ4pfXa0SOqGg3lbl7I5VY9t8TTeB
CnT8FABwACugOQn0U1BnzwhJAs5nuLTVREVJHCMXZNmWO7s7SMmU1mCirFN7THh+
ItkQdZt/vtljzJbnGTWiwvF356MgGMfttplYuyKvzP0YhSLCwxlMQlOvytPrUNM4
1HE4onu2aFjuUranZHzLlw==
`protect END_PROTECTED
