`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HnwmvgTGmX5LLDvddoh4gpMZHJIN+XHWaipATj7ZgrEhQc54TxZSidc8CAEj03i/
85ZKOsv4PtB+jHHgVbiA+ur7HMfTEzUQk4Cvkh7/iGi2zQCzI+YbtZIiZFj6fN6Q
hOO4pwG96g99pZPfsDoDD19yDWhUW5YlM77de8Z9/zS+49XOnxYgJ3xaMeprLvmP
A8Azve4r7iX5hkTaqM42iIjMdEFwBy61ImWRM/q9OPhGrSVl2LHF4/3iE/W/OS43
qTV6CtyljMfbv50rp/sEG0f2jRuipufXyGz71S9I8+d+bZ1ZOfFgh6XI6UQrOd4n
Iw7U8utgGkOEHALsFoc/7Q==
`protect END_PROTECTED
