`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhebQD9p4vEhYX+ZnT2ZUk2IDcXjKfA7YqoEhAMKlGqwyvJ4edBIvTqaxYiH9/LX
AKQ3jQUf10gA3fCrHQcRqyAKy6TqZIXbORW+96szbsP78EbLKhyAYF9bfQiGj10B
Kwuq1DBLkaRkswPFF08YmQ8VjYof8wEpxG/lA3yaVcRJ1ODTQAqaXBkfzTJGN+Kf
RWFSxnYx21OJPC9fnQESv+X//QvPw5CBhkaoo8o81dLAXNRTya7S2utIO4gXvgCl
ZuKNqVnF/75Eo/2pYcZ8dmKDt+sNdFuHv9DvdiAlV4qGrCyYzUgCTk9VGVvDtBxQ
ixPCc5aJ8VVE7AjFBAhDP8RPseGxeZmMk7qNgfk47UebLg4Akbzwb3AWhWAYBrp3
McLBd9T/FNhjufkFOCLPx96FPh7KXCO2rZPgEloQbUGCeCQ7Vab2yKqtW+bwpDSH
V8+emm4XYvc0fgBXEKvicxWHI5PAYI2ai/6MW90OrxmlQY+uM7R+8pvs5LKCyq5a
`protect END_PROTECTED
