`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZzNWsCK89LiDvH6Ee+jZZRI/c4nEoKV059b86dpsg/cadwhlO9Y2IyQOrJ0g1EYh
fjO9FuFMernVy8OTA+7ig+Q6QIgSHKHm/QnWQnQEtnF47weYSSi7TEOU/42lCs2y
fI777C0Jw15OnU7r/EeWC6FY9upO6/8ZjSHqkpQzovSGUztZz3bsIoew8kd306Vy
KO9RRPcBlNiLY2HF2hfqOTJ9XmVuDo7roidtO7DuTGQ3CF9DpEjeU0cKznwVDFqC
olC8JsBP0nxZ6JknV2jibeTkKZnI7336PZ0ZiA5zEGBAaMTMUUzUNoSkKhzZP3Cl
I0MGEhj4w7wEPV/Gw2Kat49mQX64ukBj9c8k/FfQUvQH7bjoTOXD/DP7VzU5m7rq
YbqrUoo7snWMMpoPqGABkT4pSjOQbLcsqHz7D9Wk14L1PW9ahylkFJWboUiJ/YvH
MyWCCiLC4swojB1Y7tJPsSPuma6OyxC8n1j7M5825zxV9gS8bgd0lq56LtD4Z+vb
X21BQWzcwZw4sOFwunDXRduOYXWW7J/MCMLHIfnlNdXfWPI6CwTTp/mw8CerHRQK
P4mAdeaZGOTwvWcQpxFfi8Z+HfFXFI4Jx5tCkfXBC9nECuHWh5b5SqfZUASMtKQb
cLuPE2VwlPW2K8UAG/GDMqIKwnqSEr8aGXfMxm8tIgH+nVxdcldH3aT7w9MrMutc
cmCSGwJGNLWE6CEmmJ74FHEwaFfqKvINCWnr6kaMXs25TSbsvB8XKW1q0pLQqase
irj748zdmcP5/f61tzbxrSbqDwUdr0jnNcKe2RJlFjrtkofoG+5ANIVq/aKHg/Qe
DSqhTaVep7nxWPYIdlLZdurVLOdz4tifjAYziTY8zf/doBQWvjI+x20KtqHCByxz
2mq/svNAYNHU4YcLtEgdBo6gaWUEGTFYul3gZqgualv9PfsLZjy5ltOZJENK9yw7
iyZDxZgeHCqjt3Wzs7yPBC8PekjeOaZqarWqVypAR5HpKtEfr9GlIrqCOCGViSfp
dVlefl1HxJBwpbWEISOh7r39Hoz70nphTLhyB7MrW4cbbFKqyO3W/+f3BNOg/IbL
8EBCPcIHQo3UQZHEVGZH5sJC7UR//qZBGAX/9pp7VDdx/iwVHohbf3qKKQkM2dmY
5qLua2eu86o1ayhXK6vbr/I5W0frHRirtXxHa1v6OcaA4gudS15L+aoQ5YKQCqzT
a06q6RnoGuJwf6dpv7vCqd2Od6/Jl9VtNfgwZbq0isn8gkv5ixoItD09sGsnea3/
Pe9bzRam/+AaNiZaxU6NyKdJ1OUD5yAQu1i9+eye/FRTylCHFdkzy25IA6y1A2oG
3fz23YlVpwcUG5HiH0L3Q7egB5p1Q2MaLSJojxCRfPUVGNwtkczf+injiKpo3VW8
YzdCdmfBBXnRcGDgGMhpbX620oG8UKgyahacDKTOy6lskam6jqan29SrGOsqbT4D
FN/y5OC5C2+l+MpCUtcKrYLa/aq7EWOnG/qhs6SSzJZduqS7UWMo757FLrRpjfME
cbtpYw2iEzFJyFReuy6h/Y7Cai2kNg3Mq3AKzh+lHGhdT7tJSCeq0wEWeA3tD0QD
u/Mvu4FOM+OlbbjTgOELyqVdHda+6mSY9N9LnawDkfFc9aga9pRfmpNLJ8brQvuN
qVApDTr3fIxSljDED/s4qUr0hQefl/E7aOtKvrAH6tk3GifX0nVp7dBsm5Of0XWn
74dzAecQNMFMT5ZxBgSfRxDWi7G1d0T/4XQTe7iLkzGysLifahMpOGHDJHR6Jr2q
cVpo9ARBGv4gPX7+C8KQelLVR1TFNBXGG91WvhYHzjmIURfmcxVb0BXe996UBR0w
263i0JXoBboYMU4N/Je7+bG7UiqYhLZvzNAD5A5eMvT5rcLe6tnU6xlY2wr/yYmm
QI/KRx2oyzMAR9scYwV3YzZ2A9O3DN3u9exS8FAdrE5E7af8G2azT7TQANBTxXcU
LPb9hEbHzzhufi5FEPTPj3bR5sy6yTgs+NjkkrbcabfCX19Qgtm+LYAjtIn/U8fF
11fbQf3kQ7XAUdVIOvfwOomyjDPnqAsUe8sVrTMQMwC9itOggx1IA8aFKDH2CjQ6
Xm8snp5nRqZap/B/BlI7MEQf9fPAdOKaDcxdxfpo1ZXpSyu5kwCT3TvQi5z+9RZT
YrdetskOfDJh5XeURnmQMyMDZKgeVG8NbwkPfmE94Z/D9nshLkbRPqzI0dkxVBQZ
y1UO5hEh4kYniT77FwQE6oBVYiCYtQpTsZxuDbeH37Lwy4rY6EiDDWh6TIN94RJz
R4ZpDviToGiSuTLooxsc4odAZme/ToSNZbirvxni4LQX0oKNCua6Xk0n2g4nK7Dr
sNVY8nMaBX+6xeCh/hC2t4RUkI2i/HFdlLHDEt8xtrVYnIrppKQf9Lz17C2U5yoj
anMenrtOquWcVV3ACJQwaPmSgVGYr1oVzW+yxsiJGEFVxJo5kEcdZ/FNfB6E2hy3
7WqwidPh6cSVp+jSNzsvDctReVzR7r+9tPkpy+QVGxJQS+yIgr8xwPad1MlD7BC7
yJqeWI8BQHMW6ZtJZMN55xw+buex6TWX5Eo9QHq1B37cOAK57zsrVEPr8wIx9bF2
TMUTe4mqzv1sYppRdYXPQN14qz7YoX+wSk9LPrRkiRj0FdJT4KXj6SoXg20O9XU6
FlQNTr3PlaoxVAYZ0k9Oz/nVdXqjU6SbaW+m7fwkq46IxOAOgbHiIXXTgj4aI+tZ
jgd8L5DIcpx0fPZIqMorVHs14RIIbFNTicXVGj5rqZbTdtYQws1t/CgET5gDJMmD
fnevbIJXEM9K6iggFLabkNO8gIq9DAlHVNB9KSR4w/1hdITkX/KokLGhIC5UokG7
a+yYX+JsLlRQQnotcPFTa3C3DX0MRVJh/UeAj+G2wSrrRbYnv2P1pMc6MZW3W7p7
n/+KwkEtaJdr4SgwnvHU2625Tv6RVvI13wUg3boKrSKXmTZa2KG/T8ZJafHZf75E
uk478TzNQArXJKtmvlHxY+IV0q/CDQvzvYj17sM7ucnP5yJrlm5w/++hjuFKNM/8
1Qbsuv9xs5Ihp4tICjF3pkrRcIxTuUXivyJoJi3lBaUqJjLA2tymeQcj60ZjQ3cy
IbhAKjRwInRLbVtiTnM3d2odEG6/zLTtYJ7rRSSdjcdyuxhn2FTZOKADn5dBrZOO
madK/9vuvyFHUCia6ExoEMBhFTQScQWXf1NVCtLFBuRlsZc9ZCEVcjwi7aZOjmtb
sOuhgQ3QFaWjVXK0ZxeuXz42SeJHAZHIjyKIxbldW4IVvfmHvHKYQR+ISt8o80i+
ZVe/WEScJ2Od2oXABtwgSDCbS5C8vqcE1K8+DqbHRmhq1vQhbU8VtjCXAEZezlzZ
DjzL5I7W/j4RBBPsl5+KdeVfmmr7U92iQqoLC0w15nnoGDGr9DKOd5iQkxLZF+Rk
Po1yGETtLqWBPRmnH/vSjIuPtviinYf0iMdZfgBaO1jRbtBWJ5aUv+OdLOJvpds3
cpjrZWKdcJmtKTT8qlheEEZJbUhkun8Z0PDRkOft7LxifbZxuECHKybqOzTeE7Sz
xE+O4NTPuMigmwXdjjCIq+WPjCPPErqqDRvRYh57JkaDkc8oEad/YUWPNXFK2r0e
OWiUOxJOg+sRYSUmpNip8OVWhg1AkB10+OxuIxC+ds/OnaXq97F27+/yZ07f6alh
bUIgQ3hbMzKtYbgXUJAStZkWPgFOxezGyzXz0r6ygM12AlOsrdg6+ckO3tawPEIt
`protect END_PROTECTED
