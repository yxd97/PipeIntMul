`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tRzqaRvZfQXlITSKxD9GlfHHyVR9FAMaTkDKRQtJpgsycOAJu9phsUqJabxj2Q5q
FUBHsgbcfSOP4ozdg5NopojZU8ykXGWLndh856pqfKmjj8M0Idj3wzmIbskLUjtC
hI/yHMg/IyXj9S8NMDbMcYMUDm4dkH3FAEqoDaP31ROBoPII8Zf6NkyJinmNJiSb
4jpSByt3I4sm91lCt/OoMzi079s+CrsUED4aQUofSZstuD8q3fhyVUcVUmoexuLg
T7Ry8ywMWrlbhWXNwmpE3+/T1VtrIgI8hW1jHEr1mL7xs/UIfLh9V5AjrWKfsiBr
VJDjwyix6f9O4/ng92GMksN7jfI2l4GBT4Cu1cVHggHIglWJ6wHYoW/cMd15PQdq
G5YA8Ha5OdaSDuwbYkSC27i85czOfLOzqNpQ/MfcMy78ucuMcYxAiO8VO5D70WpY
mQbetZ3GDhe0ujs7gZeIaQTeA0gzky+t2xzGSK9X2+G1+Lg8XLQbCwPr9pZ5c2A4
j02oiBEFW9nCUMRRQSNgdaHK+cCgFHrB9I9F6WO8r9U=
`protect END_PROTECTED
