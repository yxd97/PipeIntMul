`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Kr3mWuymGN7IFJKs4BpXi5QmpgnAb1zSC6aXk850D8z8ZTkUlIPScVeTKy0SexP
NcR1j0Xa6aOQ0GAI3LqkUsHpajN4CxHugtReFBj2FOxM1FacYccIH9pWorLYlB8B
t0PULNnuCe5Ti+R1s4bfW5QHhkLtoR16W9dFm6i6NBXQUSQXhiZbAmGzwxXDXz+O
IkZ2R50VUqGg1suBA7+AIg==
`protect END_PROTECTED
