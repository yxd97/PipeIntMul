`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pt4lHPHsm6IuCImsF/mL5Kqrj2V84cp2W/WXOhn944M3xfvfhn8cyEOr4HiNUaFd
VGfRPihxDeFoAkpubKXQKbD8nFRNf39pbR/0MBzbkc6uwHdmvILiVtrPe+pUtM3S
bEIH7lxx3XQXLKHppST5gCnw3IMHnSj3GbqRqMrSLNVs8WfWyOVOZERxCVhBgfv4
7/TqkFat2YYvmo1NHilcoypvN3cQJrvW5goXrxvvsNaZdr0FipxQGIsgvJNEzEJw
F7FcRAkW4HUQEUDKJyMq/wFxecWXhAyR+3It/aogfYcgkq7i4SWYCrGWJJ93l1g+
HcjJ6cpI40vvLtUVL09yGBRg5uSAtnKh4k4AvtohYMP3aNj7gZrqXHx0V3TLDESg
TeQWO2MDjH9dxqE5BVz7IKfNP3/hLkJEe36HpVVUYKz3/BRHsYHI36sAfms8sMlT
RUynwUko7mGY2UaZtv2hJ9S1hWM9E2STMvjC/Bh+mRf671w8DitvqJTLPzPXS18p
so0x1EChfZHbswpuJBpn0aHIsU85J3eOuYhtqSNvzHMBpbUfblynqf61VhOGF8m+
nbYi6C/Q723rI13Vh+r66Q==
`protect END_PROTECTED
