`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85lm6lctHiFCTV01R6PShoV5E5LbYGp6rycIVhFeOWL28hdq/lOlmsE5dpG15ADa
sNVkaL9LevPgFsG5apgqgxMrT2dPiUHg3wDkFqBEscxy6v+q3z22Sq0Nj3Lqo5a4
4vyq/pdkaX08Ad1RnUHtPwBY+EffJL238FVq6ZCDS0qj6M7u4BaWGHLR0VsienZd
NOilgxeEZKgOlWyfLG0NJk5LVwf/WZ+sEAQlvIQ4oVLTPhYCKsagy2X8MA+1zoEx
MG6glW7o6JnqVNuCCTuGmMAoqw+Qw3Nek0oMrM5E+upZ8Q1UHgqwk/YV57djv6dc
ZdvbP8w9xxodPXwGVy6MEIs3rphf6osQA76dyiyYGANtw8ah6HdNix3njawg7iL6
nUqfyCfqnKfjJIPeliBhzWw7JthJH7PvCqzF2rXo77UomHEqwTg0NcXwBQllYPwo
RDMaFl9Tiff0Gf4s7m9cs7JObpzJlvNnFI2rifz+1vfrK/3wsjTAOL2nutkoUkhR
JgKBHgd72dXBc7/7ZAg5NR/jO630n1QwmhreFqAkry+L+EkcZC4ys3vNomu0mbRD
zzR1ZWFtOnD9GNzOrH7dHTDypPitsJ7Uw6pN2hwuCn1BTtrpOE/IANskrp9ye7wr
pO8jG2EFCtgN82vnTemXufOb5YKY9gEPkGwVvx9PGjyMLjOQLH/EyhlTtzdXLeZ9
1R57vTd+3XsI63I7TnZ+84eXlA2o5+jUUH800iLVKi2rXIYIQyvng14Xr0Af7P+o
0oed0QOWyT8kV6WljCoSjE1XsawVJryUaeSKSFWAH0ebjDjy7otlWLZ6FRRTXIO2
433uyo2YOAIOL0PWhvNusZeXSlxOc2DtMIZ5i1MhMlA=
`protect END_PROTECTED
