`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zc929Y+LCihPSbPy2EaGEtvPLj2pEqqF0+1Mg36OOgMQNQVPEBHAxp28jKVoOYXk
r59LAVYFo0Vacq3KRnUqMmDtBDwIynrex2rqSvRLmnKOVB18uRiQALEJYj8Ysn0c
fZXUY6G7hMXLSVsXd98uZKMaDW+CTYIGaEC5E24JqLiN1/zpV+15KO/838Uw+75j
odygfm7D2p6O0CGFtiYwT4PMiR96SeQ8y1acTFvH3acyKqEKni6SsJhs24KrtuHL
09MA2LaTpTJ8yugWk4nXYk1SRXbokk8F9vSD2O6mQObrx0on8vTGDkJhuZC6pJu/
ahqt/GAhbs0VR0rnPcDrdlnuOoszo5ffEdPgKxl3XX9l+8rpHh3Ql0aglqgFkLMt
qyhf0RmTdp69oiud2nCs3Oc2Da9hNnlM03W9fhESaSbNL5SxF1mvr2vZx8Cn47eD
aBe2YpW1Vh1Wf3bEUT2S7fgL+7fssjbrjFXAM8e3YOoTQas1rc0jdIzQ48VgDBfA
NWl75zgJ+3y4xeKzc7mA1+W0pZfxSoVKNcULb92Ke5egqH2rEPNiTMqu9r1znGne
/p84560SqtE8QXYa2AviSZEWkTB4laV88IhZj62KKnHULjZLFxFpwd6I85QomV7D
/6rgU8MJIC4DwuckWIUG7XnO+4Q9YP6Fb1khSi/aRcRQdOAfIMrTbbgmelSm/wwU
5DyswPGbsgHMEumhtEctjgUzHmlhEthSJlCZRJ6HLNrW0QVXSFI4U+8jim4mZZaO
6Gy1aQWWSTnNbwCxkBTkjxniRAu/jsZktVVNExNWQgwKVJmujtx9ZnXr7NskIT2a
q2tw8Ldukt4dn3CVPDxi7Y+Zoxw2A/0fQa9anu6tMuIz3VUZR6FqVTuLrqh48MRI
N7aOmHXFoj1O4E8TicIrMsT4s5OH7LPpwG/DQFEsJyf1QyLtK6mP31v0AGzyEyIi
0FaRv2OZped4oeHRdEwJzCoXTNsK/Aa6t+IUHPgyiCE9EPq4q7p+dlR9FmbvEIoe
NiIHNW0/UVPl7XDwwLD3R0kHLSWWVmepU02OVtvMDKnWFHvTT7TMXgvpE1Jz1ooa
5RfqVXwbSNFFGNMC0Mvelg==
`protect END_PROTECTED
