`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vi0EUWJVu1IlvpWtMxJokT1kv/5XR9WnEO/NiTJRmoRR4X4agBRqKWgvIxQg4QBq
s5bZxmQOYiTi8TzeZso6VTqtiMSGfeLRPSsrMQtkXfc04oDu/uSeeLzJSKSOrutA
++E2GdQ3d6U7lmIoIkWiqgDWvwGAAUe5RPMxQyUvpav5OpWBAumNdkcwV1KXRlv0
0n1GXOSkX1dS8f2j8j40v6PFW7UmjZyuThu8aIa3WzFGYUm6c/+V1Dk6ygy3XLgP
F4lZJeZpGbvqXtsScheaLhiaQ1kMJ/zVEFOIgMLkZyh4rPgRR+kQUAEwqtfEpIVJ
cHklb1AKgTrMCcrcUfUDmcRETjjdAJ9375NSn7Mw29iFxVUagoJTd0H/j4LASMfD
c6kymlb5fsSFkVbsJLE29g==
`protect END_PROTECTED
