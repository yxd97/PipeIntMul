`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDzrJVNiGaI70abIb93RcxmGrMUOvV9z0LPyCXiiTXYINXVzp5e5HryqO8vRkYmu
vehgzu+6I1hXh4Jum2xwN2rDEXzDhE64rE2v+krnJUKHSKYbJt5ycJYU/l2Fb0QT
unBtKZfzqICYJ63ESRchiGorX6OZ3wvn/yp4xUI8mvoDke5mxhCyXzt24fNYMwhO
I8ntbotyEoXltnuH+4QwJYNdnmHMRyBXDdK8KT9YayhX7DUIX2a7mhGaRUKkogcv
C6U99CKPLZw0ujhitpiiDTVG36QOXzoX1lnhhhj6v6jMIV9YNOwJoOncpCzrufjL
E0A64+dyRBSklT1JA3hpL34HDtVdu5e8l1j+2XG8J4EQ+sh2ZEuTX07rD42z/boN
dM/KENOxmotMLYs296IFoOSJVy0UwUKXV2Sd9ecUFXSbr3AZ0xnZXCi81S2z6nLd
3+0xFd8uwGfEKpa7UK0Wu2K7VcZTpRu9416G/Q0D/i9OYJWFi13CgKUXxrHVRMTc
jrS9itEDgKt24Znbzu1evCOytYtqmDgbEyilmz/QaUts7X2ttNDwLI7URGNV1AVo
9H6IjAe1cEeTCGiAJtHyUgEnjKdZOvv3AR/RRERZxZBO75f0Sn4N25kbQNnCoEMo
plNOCVL2PzC7io6HyaGAeeYDeq2WF+RPE+rbYKT/iRlo0VmUxeOe7br6HbNTXIZ8
`protect END_PROTECTED
