`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txf0Tho1eRENYgs7MLDj9MGlNU4TRfwBOG3Yrbt5WKNcYc/CQ7p+PhZMQ2yj/ebt
/gDQM9CtjSDW3uFLdwr5Tk8JiPUIMO+d5/brw1rMCF8D7wI8PXx8jysopoKsaM55
yNfm2gwM1FL7aXYOjvHdkVnNC8s2BdTtLCf2t4SDvmGcNNqKjCKpVvqn01AHxUtL
psg6Hb4ykxPPfhPhfJBeoWRMFBJhI8RHkFlnRyYuxHphrVMjvr3gw2M4UuH1i9GD
xi86l+8tKr8lEekgH1wHtt+ryeIXmgyJ2KmXGagH8RZzF1SJHIBjuWDzXfhf2e8O
+AFk+0LNglq6bcq//t5wnq7lvpQvnKKnFA9eWby0EMdVYIQiZMdqns7/Sh3VEwM+
EcxG8YbPMWBDNjccnVlQGu3Yp5eLaZgTErHcTjTBsryRgvCHdvW7dhqZ7lAyC/VV
0+3hHY1JWVwo/HLbPi6yavPeJj956xVdsAXLRHEJGdcaExobzNiseLbbLYSjZRSR
UFtgFfN7E5NGTzyyHZID/JLuGMu8D7QnYoGt1kzqTOwZebmChH8mFW2ZZV8pojLh
hDiyep20TiHtPOFOnMHM4oERl/mLOz3d4Hd8AyvIJ1Y=
`protect END_PROTECTED
