`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9GLfFBiz8cA+s/XIAtqAluA9joZvUvEJQPUCGGSjKvX9OxFhyMjPCsGo4Qm0S5M
bDzdjw7qFUVo8SVvvHd14eUkf7XL26L9LZgKKvtR0ALUTBwm8wbJEjO3PSMqM4bu
YWve5KsSPCOgGTADk5d3BqZvTbarIrnH6sSk9GxXwcuRhaSNB1eIW8yBxhdXCNez
bv3RLz+G/j82xZnfMs1WQRKvi3Bfjmvl1duuOAUw/hRzUph4S5rV8r65Sb28Pca7
Ybsp6p+k3PyCMkkPK4uYBcuUQrOCnNkigjxIgEP+Eo596n89oIbpur4TbGMtadma
dzOaNUCMI62chtIuhLHodEF+N+3Bkt12udKwP335wTPPRFW0i6msz9RTgGwcDAr1
l2dFI9+DaHtSVAx99AfNO6ugZgp/sP9WkSQtJdCTeqjgJDQunUfSqTJKsRYa/KuD
0pIizhfS3+WIFMGhe5FgVU0k3lDHR7RnNOAJnIdXtd29O6MlnXqKdxfGhlJplwDC
gE6Ix/StZod6R9znjGPgum7NiaOwOdRUrDN8mtF3EdTNZV9xEnFoDqnKxwyWVaPX
TTKEg4549eIJovMv7MgSB1Q+0IAHBNSCfS4OHqRDLZKMpFXKzE5vXLLFQG6nZqql
yX3I+u7vORL8rSjf+8fgKsSr/mUXs3ZTKn0Q3dJgzs92UQq4Gq/DdXRXN8FF6gSl
vYqtbufVjXwLISc8GuF1E5JypzSDYeeSsJdXRm6IzmdPESgAUyhRb5v5NsuQzMK1
kk2QNSLFxC6wBuz0DxZSU0v5D3PyesH1yKFVr7VIb+qqItgOuiojfn4iwhbJFpVZ
EHzI+Fcy2yqSCK6gKVGmIw==
`protect END_PROTECTED
