`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mDfFWW9BDg6w/NOqeI9KWlqwSw6w7n6vxvNvfKP0bfazyBJTpYDabPdjViAvFgr
KnURsq9yqLue1+LxoDAcoy7ggdWBXW6H1aTvye0DVpplokyzbejpUGVhHBa1+nCk
j9v5J5+zkp+XO9VH3CovBErtoh01W/X7un5sH7Jslsb0tMHqxd5L0SWWHs9rjpsz
xSjcTco1F5fLO3IP/6k1MudJ/VydOSCnb+6pd8PVtEfwol8qjLeWJ2u4mWQQ5bQc
NSDDus3pZAaCs1rNo8MmSoCGpD0ZlFX8WPfyaNzOxpt/4SkA+p9M3vlNr8cgH4xP
1QwgQYRWCTW9xICWD4c3WliUdpeUnMrgCnXDmUtRIaYEdYrHSNL4kyG6t73qxPDN
/M0KrgJQm8hDVXZgLjCotX1yrO+QBGvSEtzmr9scWiRMpo85XFZIV8IdmF9P5rzJ
1IJomYmiQWOOKCK7Cd16aejcPJckzMru3jOi7Hkjk9aIhJ0nqESv+CZ9r4Exe+WI
RLOx29HVApOlAQjXcan8vHIGIkA7HKBBp0PsNgl3c9PMRxX+WY62qtkEVdNWCPuC
L+DffoqPbp2G80DuxQUoqRhbxdcd8bSyXeumCkccQRY8CTaVbBudWDy5kBqd331f
TZCd/fQDAYc0uB1XwploB9XSeshEtIRMrGHScA+H8uaV0uJ0ofJZCCF/cJz/+1uq
DAf9ZeQJrxqhfmN2EkxytUBkKZslO8sE8dEcH8U0+LKzTuw4dVDb+fJ+hv7OnOLL
m3KZkvJZox8t7e2Kt4gW7W92Gh9wE0OA4sQKjS/1dH/wvwcUKr5IYdWnbHlSoRD2
FJ2AKucljD+k21HzQe5FnEL6SI3bBWsqTv1S1pozMK15IdRSf0cLTlB1HR1CCdTa
vA4MrriCyC6gGyrxOMTfb4mYn+B63zrX0hYp5ObsqxzdPMv2Ou8mXiyjHXLC1d5E
I2QnXIiQbULCS7s8K5Y27L8hfoeOxF22KZvSYtf3QY7Uxu53fjFEAdVn9HBmDfCA
ultJOjny/2mxTeCTetyfEDDrUSbEUABY2xvcxAEQWdZQuzPDf8qJbdVV3V701H86
bRUq98VBr1IAV+VMJacp94DxbdKqrdCqiIdfyNAjLRGW2NMq7tU7TzUvbEeSc1DD
eDUjLYX55FiBjFwkNoqi2wAYN3X3P9RrKfyEX6yCTlxAvjsuPyyHKLvREeryk53+
7rCvq5T/B5EznLFrdj7MtMsNvay8w59QlD9tWdW6cnx6cj19YOAf0Kbfw5fTif1M
OPgakZZjBGVtiW3vuI/uE+c2k8FCvP+BblgQlBmeSfMSIw7n3f8rGBPALoZPUwJ/
TtLxbt6sk0upLNR9eryk7kfKTNNwWhWLgy+QVI/LQ1WYlvFt7rLFj7FtFs2KDCHM
S2FHYO8okshJLaMABPPC6dU9hqmbSl2xEFRHFq/u1PYuc96L6IlEtbgpW2Zn+4tI
76eZS0zFX4AyL5sA+FfOqIDHqTCGa4bMn6NmkNoL9pzo1U+jU6c1HXCPAcpmJtdi
ZdwONZbQHuoCgbKaZV6i7fHVKq7r0bbZGgDJJx6PBY2MAIV9wU75Zf6HY7Q5o4w3
rpHbSuDfHDYOVbsKvYq/onsyQdacsQHE7jp928DzoqD5C7EBVV4WuEVhjFKL6ZHU
cCmBMXHR1P9T0s/6l3vZjj1Sthqfei79/AUM8r9DR83hMqLeDGVzev85yqcjJrSh
S6TZm+M3e1J2beUJEoJJ1nml4I32qCejUxUkyKCEOAAoTocqFrxQmDV7eb1xsmat
wdFSXPluBwSPocQ/QMwIQ8Gno6nzBYNwQb/4UB+TpXteL8964pAH5fxffHpjth6+
YGhUOs/MsqYRAJRNi3F0GZzbnSs1onbykxNtxKJqoQEV5ULfF+s797/ZT4Q1Vf0q
y0Q15p3HlBlK0aFUKeccOzd8LV6rkyZX+Kt0E6OiatXX95bxUjg+UQNoRdY7XHBH
20tEIZ5wCMm5pOmZoEamNdd/rZUxsDT8QBI1Q1XC8ZcYQOKXay3iz8ab1scUv+tX
WZFiHXsynUWgMr8qyY6OwjPteCuUNGq/DqIq6zoUsS+f2UkJ0/ADvOxzTd6XRJjr
sF+qJYeLfV50GTQdPXKZactfdlbDWVIggRpgHcMLFklG+WbeVHQCwyC0zqRDed3q
EXHzkvOVSwnbwvX1We1JnXloKNZXbEnqWxm2lxs50BVF1toboc78K9Gsu2TJSjIZ
E8Q7inK8I6p7F//nsJi9372clly/S03ksRZjp4KNr8k69YUf1nmQDvYf/eDd9F6e
d5HnASGQPlb4sgtY+FynO/a9aLh05wmDOg8azUbsCCnLAvKssG+aKOGlMWk6dCwH
Str1fX1qJX/nmN5EmYcCn03hKkchhmAWNp5qQlS6laUeR67/+WKcKK3zvu9ImrK5
7/3Cq3VxZkxQLQHZ68n1qsOgthZr0xwfInYNNN6hi/ANkDzmt3wziziGM78jUuQx
AAlcf6KdvnC95vYaLeJFYYsCMRzg442VQn2/0jgRcY+9I7zmE7prYvzwvH1HXfTO
syJbrpdY7Ohbt+rJC4pChhTqbHaaYlJ/ZeiEpHvYyUbv8pVCI5Q03tO5wk1ZkZSn
ERh54eBzrP9GdeeWviiHGK/E5FWw+Rf6wLtulsfRALPSMA0dEiVSvulkuW29ZDZH
XSy0RI6JoxbWfJkm+qYDKr3fm4HHcx4X3P0qDNH44PBYFi96iIcsLKJcebEBZN9e
oSQOm0SMBwZOww6R0GrkO/fk64YGVFpuNdOINYx3/XaR6E8sjwAXBLIoJM6p6hnV
2kYhNiI6sfmIiuL+CoWzP6W+vVRUrQ0h9UXe9OxEVKUIkIYwcOhqMvhqMriyH8v2
QMYkKxRczpLD2phUi7HdkqzAYpQZA1cEQZRX8HKnS8JZJ3sHdAZtOiHAbaI4Ex8y
FuxeUdAmZ13c6p1DQo4Ej4N4qBbylmgA/sJq5D7pJvUc/IglXZf+4r9TkQQriMxU
rdl1jR2FIsnp6t9rq8vatadSIdUK3INvw8wNv7QTToNLsUdCCSIbdRd9P0FLK10G
MCTL2Rwz6DibD/c5hL82QEiplNUeG9CxE+0C9bx1aRR4WR+8ewfnswIP8sqn6Ote
I+5mqLPbIiuYKvCE4q7kkSuIThFlFGB0gtfevFGNPEliX52Gu29zBlrQ0XuyU3v/
lgvaZAqcy+aQsaK3afaHbsyhqlTTECdJhSZVoWGndRVAxMGCqFRHfnl1j05HE/cW
XBTsTrMi8BzdjMq6JagfP18t3GbJib4XLv4laSYkmwXIjXNuM8QO1+44ybdruumZ
iSg03Fe1JkL/pG4qksoxmVM02p2UuIkotHTmKaCEPiiHDocojdoWoV4ygH55WUyi
HUhfvpYAUZo5CCGggMAlNJVHnw+r9eXVyKLTbzgktY2TusQTNFuDvC5FQFgCmSpx
Dzv7WP1I6mao6wh9WkocQe28Pv60meebipkolG9b6guPrz/6fNN5/UABNBwY1YuV
NyqsW1s/fTS4wOdQkmE7lWrqN9qJCoMPhXzkans+ORdQ5FAVXqOX3mEX3bhWKJUf
dh7MgYsLn856qWudqZ0aTJoc6obU6lAOTE3ui7o/MoIOOBzUOgXpwx0od3EB1j7Q
9kDbRCd0BbdnG34xLULqU8HbHJg1uXxgYzDWDHlOV1yp/vKEwvO2Oz4ZltkFIeSr
ygwWmfGs9lCDqPu/PhxrJt/80MCX+Tm4rkIkv2SP4YrnxU57nVTyAEXSryorDB9R
oa/g24UdVl8C9I2JHR9t1aAwPBOGqwZhv3BZ26U3Jcmb9W//PBNWifi9NOzpkenH
ST84LP1NhNyegchwzWEdaTNBkSuEqKgn9jtAdQsR4GCM6Fym57OAhT/Inin1X+p3
`protect END_PROTECTED
