`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IrHkP+uIfuKky5s8so7HLq01BAiYo3Y620W3TesAqBTXYf4k4BqSYLUk4A5F+W6N
Hx+ARqF2zjSV97Ub2HMeIpyqPW/p5iyoqexzWK+I6utYzXzxXZhZSC3chkF8Z5Dz
uVjGrLWDwVGZG5QkvBSoapSwyTjqAjo8zlYWM5qAFNyLfLR3JKN2z5eylXAOXVML
D3Ri87RkYMGqWJ/q0xggM5A/unNqFqHdrdRULXVdk1VwKozm06cKH3tJoQcMuro5
eDf02Gt+5t7JfUgGWao92qQWkqMbGSeifvUm86nHoDJTZx1zpDMZA6YRcpK5Pwbq
+JBZ/5mOtL/OkbuCNqIOBNWwQl/vb3Y0m8NvhhrEjULIc91+qlgvbuxzSyZOiAtt
0JBqIRCScrXZfnv+Y9axiRB5N/f2/jNJjFwYWEkjels=
`protect END_PROTECTED
