`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VvtcTwcVapAWuwnq7z9naCwI5KRaXdPvOiL5HKx9MiseSuOEFu0ak75PzIq/SE6j
TpxLyLamnUCHVWf2glAIg9YaiTZAn7s39AcAHXZvwmZmvUJXwv5wcsA0kMVLzocU
HjQgecThBKytyslI8PQTCMbwTHYcah8Abmb7heI63WKqi4/NOZOmw7LUuWth8NgL
a00NMSI3h+lPPbesTgwfGVdz1OV9X8lC5YnMjqTWBEEZ76zDg+XQ0n2esUPmoVlS
5+W4hKnF5phxcHkNHnnzpcn739j+SiGkkmcsE50WZRY+SB9+MxJNsAz7ICrk8t6l
DKlYbne1jIMgwb4/qotNn639fjkKAlZlmCl11bM4thqcjYHj9/LVMo+B81vF6QPH
1SEooTB/Ld6Lh5jm5VwiazKCMSOyl975Nt1MLf/jMCU=
`protect END_PROTECTED
