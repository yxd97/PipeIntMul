`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R1ASjYfVq7x9FbdlzMKa6SLanvHN2ujZX22ahtcwJPo6njKrmLbab6O3WJzFKyTf
cDi09RHFgl5t9r5wKmZV+uWTKc8IKsKycyqGvJjnfTJp/MK3XtzxTSNTxsbT5evq
IbsWE5h5X5muBNlGs5L3x/Vw+LUOUCdgnQskz+uwpTaTVF5uXaeHwlueX3xwVQRK
+0aU5R8rliaRu1V4xqrslPUpmZuJrQVsnsDcq2EDJ6JxtHKjNITEkRIlx9OhHasC
j9AuBwVCXzKuJnsekC3zVheCrKPwJEG9VQEuyH4MiMYmPPiwe3bfqc7vvrgnyGnj
QIs5NnaITVYAVgBMjrAZAMQ1D6FEOD1folvT83H6KrGKBaMwzPU2FRqIicui4I/k
PzLsWi90+tJOVo3MgivOIw==
`protect END_PROTECTED
