`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfj09kiBmo56Rvrj6VZ6VfzlCFifVTklYPvD6v44MT1eiQ4E8Ko7ytdfCRlJFUP6
LG1BuzKpHPcOjbdfkOIfnRPPYWnb8sWIMDobTc77CJ8PtvkQvEwEd9bqIrlZT4wc
9vCkAphGklr9tv9Spyfy0CHAOVouMlhMMK101zuawrxrNIfpJeHrHnMVwxlQ8HrS
fYEK4FxpTF8vFUouGd7p2EMO1HL7RQ0Zt3kThPsn2IeL4vLjHybByG0jSncEoYUr
nsTtsTv7K6l+YPsZzXeAtIG1opsa0dH1ADWlqrcvi7Ird76AY09pLP5BV7/MGiTM
AvHp1uDWnMQDt+VFm9MWkIKry63ppDS3ESlmadqC22jQtngaN2IL0bEorF9Je+cr
AxwXednVLySFssgtC76ACJMGjvDJKE6TloqgmJTW5EeT1uPb1i/tqY5glY4A05/A
xqneEKPgRsTQZgcBpE3NCuQ8YheVLZKPD18LF5O/wr6MjCOLYJ8qR8+aB4SmY4cN
tqJqb0MGQDA+r50R11kI6Myy8c4sxbeZ+mmgm5iD0uUjY8gDFkYKomzKvL0JBBij
BYzQQrO8wwQ6ttu5qXZxEQ==
`protect END_PROTECTED
