`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/BIVVnD3MON/YBNGgjfIjGkc41GJpa5yx04tATRhc/pKn3cWEUqsqxJyixBxSZcr
s+AAa3PaxhWvsSzx11P5khOYtAW7KltGLk4TVf5DZeNeRZF/mNp4nzTph5YX7Dye
pJji5/WZ0Kxru4nmER6tIh3Z4oLqgyPvWSn16ce2AJFpTde/sG3TDOeuTRhx+5Hx
W/ESDnNGVAtOmDaVUUyXTBAYzJHlt2LysROWcrQZ/3TuE7SbTBGGxfYUy7DNmBR0
IFukhShIDvqXvo2jzmLlIEJbA50q6N2VpUDyAZhz62rBNXpMm1gnC9KrwhuHaluf
m4WTkuMzvmBUdNxtULDbd60+yYFdzQvbpArDtwjHLGCZZa0SEcNWsKeSSY3a4SoV
gkY/mWOF15ONq8Dd6i/QCZISKn8uUDBNFj9lpLpjE0sx8rmD0ojQVa/EWWkRleqN
MbTryoyv7cnciCBgOfeKQmG8UcNBL3La+o3JMzvhFy6IbnWNRbHd3SLLXrUvZdQc
ihT7xkOoNktuC6SUZU5+X9+Q/SU4qCI+vhVXRmGaappGIDxlP6eEiyyfuaa7PdPB
jpVop337pyqSBc8U9kVKjLDHiSvE/BAALEEbGr76jCFyXNlRWPOTwlisCin2nqJh
ZcUxcoJCcN6QbAk2j+dpheD2ZLTyptKOiWj87bjTBB8riZP1qAPOrdocjxnP6YtK
jiy3ezzqe85JEcj2EkaZMhKgsgVCp/5mHRHeNXY9vPQjwgJNYFNkXxrALlCugxYU
zHolEsFZmAgduryTk+84pOsz9/2jie0p0G+zr62pulI+Jq/5DNIhI0NEyHCTn15u
HozcqjSdcYpkw469MBFGLYMqUbquBZt8fizJivex8aguNx31PQFwFrdlYLrrXhtf
+YSe1qTT7Hg5tO98dcCsqcL4AzA3FSVS0zaQh0JFI7AsawhsI0sVIJkDZmh1u4lN
cIetcc84YSTbLKY3ODqKGoU21FcFO1x9tBTBsF2YoJeejkQxkilp3BrAZgXSNrh6
VXip6hPWiou2ImsvptjIqGCRZN1nmBrt6VjwS9jfQjfmKtEEbQ2/59RilbAXa7M4
z7I55iLEbEfXqIjTjOi8z0t7zgK5pzhfSfoiMb3L7IKjl55Nvwmz0MoBS0j6yKuU
AUe+il7WCk79MYjPN1fUWaIKFL/p+kLlbflaTgdT8eaubIeudAnPFRnUsQUFxcxx
EhQ8oDbZAw2lar6mdIbhLxjL2NoEHX5pfoUOKEr3iOpgk7gZve9dGmmrUhs+J2Nq
Mn/jzwePTO9wZjSuIfmgJAYCYVBqEIY+WrOInX/UGgapcrkIzyzFTW/YLMBPIRB+
tu6Yzun3Dk9i0H3Mqe2IJ4/O7f29/TEq4vGWklh7SzZaCIMplRfah3jd1qE1/myh
am4oH7ge+E909xud2m7ALqv0rmfD9x0gzgHupsVYokYi+AJUuA9cWopRy/OA+iM6
OKNXW/lgtaZ2oAAmjnZcn6Z7MSBfaLVYX8ZFeBh560WhXlJJe7YluOdq4T6uGPzU
pEcPn4KQ748WIJRxh+LLHA==
`protect END_PROTECTED
