`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxGlRvAXcH3L6qa6e67TzRkpYIjQbUtx1mRdwugOp5prxJYiu+O6hlnjyNgZAl31
Pt/8sQ4qDHVEr+q9uzhkZRhTHx4a09DrOPpfbXIgR9J8wzSLCT2poluOHse+WG9n
3k5nD31oZcRaS9h0Fs4yOAI+eOI03O3bbGPbL6Ju/rwfJchHDQZc1jdEX22hpLp9
GElkBn2/VAMRldvEnbYJV3hPqfYwOqfWWJYjqiAvzeHXxFRmEx4YhqV8lp+rFJH6
lpg/J8qAdETKN829akdtOw==
`protect END_PROTECTED
