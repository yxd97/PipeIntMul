`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YyPVht+SU5exqH8Ud32/wqUgmyBccS38p54QhKS6Wf9L4MP8suOgZaq79EHtXil
V2zhjfzwRyTIS5/a3L5UCSJnfACAgLNb8pOVkUZUBuXrl05kgPFvu50BVrItrDgi
FuKg5gDtwKvRRnSJsbxjlK98eP6Ea3tMjWoZ8sYk4ttPIk8/QFll2zeuaV/Fa85F
nflbLvgO/OOk9lh4jk8DND5ijzulKlpYHSczPSrbvQrfa42BiZal97qlq1vEU6CV
IubxycYUophSAc3LoMO+2dD99UOAMYwXbsm4Ba4DAs59iJJNTFyi6+o7kdkIgPAA
QnZMEo54WJ2okHWJ9ilvSA==
`protect END_PROTECTED
