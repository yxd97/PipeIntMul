`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ionq4JleqtGPKL5Zz40fvc52qygQ3V6D/0WLf85lG+9a5kpbEOuhQDOi0nysAhq0
v4sbGSeIoxS/kz01jSHB7Zp4ri2z8Ddi7oLJryIdvMvLgIiCbHrmlph4UF7YoBt/
iz6JVpA0BhNVZU864NmPdGIqgUHd7aM6SLL1PaP2p862NJDh21RrNswIVxhwrMn6
bFY7WjugyiY2oDIZ3bRIcTRsxvnvEIRaG/brrpyFz5Lf085RsXPPZlEdqmVGhmZz
A1vdju/u1gUYMuPhl4xNq+pyhjlXq6SfDcj1gv1GyjN1U5PZqwS0PON/Ou4AAUYc
fSSxOeonXcapHr9r+GIeMKae55cx5jG1CnHVQnB4sqhTLKmAMRVdBFco2v2fGYj8
Prwcb+58u2y53kc2OMaheDD7DyAZKjeRxFtdLONFFrjuGDAghlY2o7w6Zt+5S6AW
IG+QbCLyZMzCjcyDpBFt/qYv0ikB+chGG8QOxlZp8X17AZbftip8irdIo/0BSSn7
kYKCBHHf//HrK327aQI1uGicggB7IixW4PKRKXMoqHKeyPT1UbjjKsSLtgwC20dB
XnAfDL2g8qp9d3Ob6MCroBKnhLQkR6SKJZQkwKW9gOP1DAOsBjTaj8NsiAzF4qVE
AYM80amBOpAaVzXsHXmMp6/p3maP4pRaYYSrH+TvxeUwiyodpW1NWuwG0CHYwCGm
S2HJebbfDcgU3H0k9IcLjknvl6hVI2sJ60Y4f970gG8=
`protect END_PROTECTED
