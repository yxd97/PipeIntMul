`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qo4reoo15uMz39hksW3HJBjdRckk4R/ukOqaKUg2hmV7LTl/vYu7/V0yXRguCYtj
HwENntOzarwywI1/7+Dx6Dz9gcTstCQTKqrjTz6jglOrOV3sF0J2yIqcYjxbUx3E
CJV9k4O0MKXK7o3unsf6RfnXM3oRwi8A8tGWfN3EtHxZwtOKn2ugrq6TNmGQ9Zve
X9bPmc5CdvBFxvKT1XMRaWhYqjQXnfALGWN7rRHdR4O9vHO6UCpjhWhBMaqEeyE/
YEFhH6puqyiyW6M+yCOR9/HjBj/6DbG260LnTCe0TzassJ+pcFGaVGGemxcxTaKq
XlTavoys2SyDKtijbx4ZdA==
`protect END_PROTECTED
