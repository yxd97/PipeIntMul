`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jw+uZz/sUUsmU0DHDMSfFgvjQ0JT5jLikWMKlweCmrJEE04UdqMT90ahdK6bchT8
zVFYaw0Ag5bTMd+7E3y4g1K/siRtv4I7YnpXMEM+rZg8B+5dlFmsqrpHQ+nQpFar
bOozkFFL9dUv7dtM/blAXrFmDTuDlsQKeyRypojOYzS/3mmLTqLzfjw6kyAoJQXx
9LV0ge/nnYKdzOBzLP9SAChY0NwXq/mZnAmT9PF6WEzAkXhaIT7oDq64BEa4a2I1
FpSqA2vyuoj4qExoeZl2rAm9INNqVGqsnAIs4E3eRdEU2RNHzCH5th9ZVARPukww
5noqAuUNQgrOoAWk95sve0svnPwb8SoBRFv7LxHtxT5X4+I+Yhb36SrMDFkVFok3
JcfS9Q+depiNHl+dP8CQQJQq4YQLD4D7l39h9rU6ufBg7EotJbzuwJ8g0EwPvMfP
7VI1gTZkHOv7dlNO2axUTT+pJvJriy5c9u8Vi2F/DCUQpeLnDiNVqOGfPDJXYsgu
qAYCXhoZWazAs5BAfG51K2bzKcF89N4fyU6TkiHaUgJCaC87lYi6jjBqIBxMB2e4
hretDcd5XYWWnRG95PxQhsIFzLqyYo9IPaJNmXRINORynOHbGp4qNepuJdryve1x
blT71uADD2KMsLyI6XOyptu6zFbdT0zVzFKis4/sry1/11usNXBbhTAOankJcft7
Jrhi7bYo188TbGXwlcJy9iDYefmtF30g7z5hHS9q9xnSVtmE06qKU5Kwh2NiNcZ8
AqDiKQnMdYwKlVIgLG5bNuaQRca+KAgVQQ6/E9wrYCU7MumCI+S410DPfDzxtReR
TE5LmSEb3MAC051IWluEMkP5d6uscwdEtpgt3Rt8JSgfLL1bjHOu42jXm0nDIm3A
sNSpFK56Aa2agH76KSTAeMU66XhGtr4S2ugM496D9ehsML1tTmKmEGpIPY39ez2M
85trxQg0NWLN5x+CVupqVtD/bdStCaRZAMMaIPi0zIBu25798Z5xKwj6hK5W0Sa5
tzOFwlvrFbFifpFRvS7ASg==
`protect END_PROTECTED
