`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ABQ3/G+UX3LIUfsJFH/JHfvR68WPXTKOL7ceOvt4s9nWFOx9CoE7tyld7EDUT9FZ
h5VnK6zYe91OlsHZ4Tjej0lsJJDHZd6fyVSEoL62Jo2lDyXUgWdrp0Q0GpNHCwE7
vdZkeec2RqNqpsloKm2/2dlnl46YGrq5+LPdxn584w8MSjr4y9KoxMmN5e9IwZuc
fkgYPObbzoXsZtvKoFJT4w3WyGes4wGmIl50S2wOmv+QeUulSRnjsPekxmHf1Shp
zIkIMyz2eR8hA2g+jb9wC9b/STOzBYKHgTtkxNUgHsSWKMfY0+vdFcQLoBpYOIdF
AgWFuiMB6FxjxZC1CEyi2Pb8fQylQRsboaJGVzF9WBOOF+KsWKUYaz/K/xUteM2E
H1mKQUwxHZN73m56rkFQ330xf/0axSdvXkHeg+MsgWHun7uXuo6lrXjaQ7akdIcZ
2hg9Gi5fCw1LtwGEdLsUZQ==
`protect END_PROTECTED
