`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6SuXqVwRgLD04tijw8aggkxbWhnWR04fNa+4m9HwjXamhDhPjhaImUSAlWtSAOyF
F6GqvTekTMczQs9zNDJmQYFTX1iYLgofcvpu31XYagW59xp4DAok5XBZk7g31KIN
HUnF/+5PdnxK/qWMwQMaitB7NEMNVxD52esMbfojx+uqiHXawoRnaYzNgKRLJhIq
G64OF/yneYFqL0jzFRu7g9TLxdv5c2yICJgJNKoISwYCTln9w8UG1TozQlhqUWSQ
WvFExexut5RNTMVj9oOghPLx2NPAVGAb59blARHjOauH1P3f2WZzv/SDJPIFESp2
GEap6ZTDv6fXyN9fUTLSlgH7HbDNtySE1kyNlPbBW7/LnMKZ9usT8hbGWQOfC70G
TqY4dSk+xqlm0JWYNDr4K8DiI0YFtrt+sjqacUtuG8Jx3KxjIdmAZOlUlwz5lSs2
VsqnQVeiO1HS4scZCE0ULs+q+KdJG11RAtp1pHKNgpuLNsboqz5wkMTfr0SuWR1z
aLrC2GbPq+5I+uWRSCHZsoH4cf9FN+v2Q4jTRuRZ/jycOZMNizN+FewGrQ5+ouaM
xwoZ5kehEC6mLJv4fTyYw4jMWbgdnbobKqyzcjM4U7hBaWHdPzRSw24/Qgv8g9Bx
DHBlZrRunVDNE/BJuT5PWToXq31jW1ltTr/Dk8JB9NWLc7Xwz43fngbwdmLD3M3R
fP8ms5+npvc4h+YVGLG67z1QPD1kFdmxPY6+xqtQeXU/xZ6mKZrY6hEEtaYlWgjX
IMUiai1Bg1zwNBzfqSFtauXv1m6pzs4X31eTyWn8S3c=
`protect END_PROTECTED
