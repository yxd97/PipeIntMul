`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctmdV8FoL7FtpV0XWSALg4IHgndxNfN2rZ6XiVpqn9z1DzM6dGAbA0pDC2X/xNIJ
bPzFj3D5kCqat1b7h919iRhXKSGKzYPn4wiCXaiiMLDNK+YH6pvi2eCTFigEk7ED
ahrkv6sMDA4pMn0v7Pf1VNfqAOyD6924rlKsukYqL+ulNMPxdAVrzlnyQvuVOj4H
e4ckUnzHD4KL4nmDyL5ZuBEILSvTOvxnsK/ou5AOq4e1VXwRcNLmA+pJY3EiHCYu
8SQDlcwnTb3AkI9NmYWTV1Cii5doVoHzlXeEX8BG0rDizULTC3r8888FmB3h98PD
vMrOi5CRVNYWv5FRI+ta1BubE/ZSvO0md70jI083PHrveVAm2fv4OG3AmoLNjRHP
jxzRSUyfgpLHzyTLTcqd+Oocdm+LKtK7F+Bh49kPv9FqF15vxiKRvlyi6+uEA729
ihJikg8pExCcAZ3yNJHdkeSl/+kU2fS3pOqtRzSD39UgxCnrWHzDq89S8aPxqvkD
NyyrsjOghu5B7SykHY55NBWeE1TDtLC4m8crXnFI4s5hu4/cESA0ErDx+YYRWQ5W
UI/oWqh5Uo+ydRVsgmNMpBi1MBigpfzawSl+Chb9AzUib2K+uY3if5UlhkVGNQ81
JoiB2fEljh4PE7zOOSeEHOfBrROgp3S8yJbnlsAIvhlg3cQoD5XD1iUAOmZvGIbF
ilkBBP2xCXmR2WOS+OtXSGlj8RLbDGQ4HO5FNdbHi4zL6WBKX5flxdRUmAtOzQT6
zmVnG/EgAg7Ey3RcT9vbBVtR6woKwNKx4wz8ulmkhwNpM0ytJkIc4ToVrUbWr4c9
0l/19AMhcuJZX629BW7XHAXXQHJBmSQRvcRAp7osH1zeXYAW4MNlKiid+zsuFPCT
2fIEWqVFtQN66ohB1O6HXRRNRfywhyBdFy+UaERY8V++MdNo5yakgvZAYohA9BzK
lZyhUkVhQLexSlSESe+VjzorWwU4jRUPev++3nZUDtshZOH6UKBtr/Ab6iI487mp
G4e8VG8XaiKNX9458rCE9Bj0MOaTkypkZD8yZmyxBtVjuaGB2uKF9a2fJvVFGSDC
UtcgleGqDIpjymmbmcwIyXTtOCrRdGgzwJiQdnklJOyg40+k2EaLDhNvOesluhpU
HorWKFZqJ7sTrC4gKI+t6M8vI8bV/SonoZ+zB2Qnw8xPozMg5vtAj7n6irJ4Pusc
qGpkdfIsc2Y7cHq6eW4SNlbUzV39CSkkFxPzoDEIY1uM2R0c0k01Wt/IGT60XypX
JcBkjDakrlhbnpMNGYHhy2ixgIZbvZIrNu+FH5slDNI2db3jhMmUhB2TfwR1mGs/
+1FF1ak6lFFAl+lxJY67KauDlW0IfNQNVRQ1lp6ht3hJ0kD4bvGO8kBpTJiwnBkG
jQKSFIg6k1ALAQDmOiWcplWi1w3ZboukKQGE4UZuv+5EvNxDZNXvoOwdm4a45Y1j
I2X6c9M6BZYWFRORbnjZnXD2zUPNyTjORp6J2uosE+ehbOo4zKnoz+IPvad+X2zP
NLGQHIX8x4s4rUAxCsbkL65bS7sQeVXGNmx48IAnUPlNECBEz75QRdg/CiZxCtt0
0pfsB2oeJJBf0Mwz0nqZtaZVpGEtu9zXPC8anaPWIQzA955BlaZEGBYrhdUuA5Ak
qXKjVbmvTxYKC19iwq7XZqW7mG5+xFTiNqSiljlkObFw29eVhexFMKub8dVrixat
tZF2+ljopapYfhNk6k6/wKLpPwxZzziGGFVfWKvuuaZorvkO0bElfAzYO4F/QOV2
`protect END_PROTECTED
