`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rnv6oWSovhr7do1wPGhUUndiALConVdBXcTtlw1XZtwyh2TierrtkIt8ohHzNNNw
XUYUoY37Sswvi14i0sutXL6ONIKg0kBP7OmS1TpzECnNm/bPhx1Ez1fDmgjUzmKe
EJ4cD6YAAAGZLXWOAKPDHaehVtW1Kc0vsyLbCHJK40yZZvs1FErYnz82g3OzpkvA
Tv3BA5OYb2bfER8fBU/iXPIOvoB9AsBUq6tmzCcDwU384+nPqBA7XmO0T7qY1gCr
R4n7oDhyVFH/O5z7psu78WsIrnomqVij+HZxueEZa34EgO1ZH4y9dyRJJ5vL9ol3
H/oF+5vxd7JLbVB6FmRI/V+D78ryqgF99FNK4nkK3zLhuUpBJoz5lp3z4e9W5hAT
1+kEo/Lh07ibGU9QMQrR4A==
`protect END_PROTECTED
