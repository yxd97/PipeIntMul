`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGB+FNgwaii+bH2FkJ91zohCFLa1//5sIkGUseVqT/z05IkQ1lYwX4o5W1cml4zi
hw/nCx9T4bemFRDERorTIkvZBFBTniepHBkn+ub3YB0OeuFWetxv+E8FlUGhDZK8
56funokCjfiYozFRVixr+JX4v/ovC2BoMP/MW2vTIfE3/B8S2YuHx0nEZjetXV3y
argZrK33FJdRSjyOm7r0pIOkZ1Q9ICEC3LDZkzgJrRfbytcY26k7K38xJ40NpMDj
c7Wu+Bc40WB9E19DYS1++qMrImZaUpzi5egnXQRttW1lBm3bPAxgosqa7ZI/KwKL
OufwOB5THdUGfsIyUA6C56QJNjukc1rZKjrD4hlWizOA0/KNZagMjerOnxFAG3Sj
BlyHqReXGWkjoRGX6x7wcVSNdNpwFhzHWPhGCh/AtFTaJkRZVoyxVlYTiks4oVBG
MFJ0ppvqnTdn5BGPAwlyxpUxJSBLur8rArcaegyazRVC8iTpfnW0mISbPKSn/iVr
nAEqBveyeMK2W7rJqmMIkxt202+yLNmZ1D/YLsA5LBREE6LGAfDoDsKlB2eiH9fg
8rCF7SebdpQ3uLqy/J1C+9YzpAn3A7IM39kjUggw7HIg0HcOYyTq3xZHsA87O3h+
bxouSjuS+GcdQSQ6uI5RJw==
`protect END_PROTECTED
