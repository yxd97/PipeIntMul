`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWWUPG9m5WjlErn9xRmg5obFixr2m0Ve4xAFJYRxvFVjYSOqHGLrCn+hTcCSHhH5
s1ADjD8JhatJlT3iTMXrCWzG8EzhGgTvvjMpAh7L1q8DVLj139ghuBZnWt8Qw+Sf
uXzQ5usz98rD2CdAOC+wxmEysHJbmQRZJDvj5zMjrq5o1P8g6o7fT5Dg9qB+XgkR
rMjOpwQgi7dOPJjzd0T2bnxRsy7fgOxQXcg7VTKt0Qq4+aRKyhCyYE91c7p666FH
TPXWpvMZfec/GSHLYVjO3RbXCXq9JtQ+IbvPfH7FgozWPy0X1KyyYOYlPscunzbX
kHgK+ENh5X6/YK/oP7+TiJ9B8FiwlH73xgEhPcr+f8D6rfCgs6IJtfCcUMCDXXTQ
hXndT4gftUKWYlKSj6rrPRZGWqQVSbnytxzXv9Ir52T+rSFtmG//pP/A/BbBZ1Y3
tZ3jd1gGl82h7qWjnUnqbysWZfOtGN3PC17H9EoFYbQNuuHMWnf7KDKLPT0f5va8
`protect END_PROTECTED
