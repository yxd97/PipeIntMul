`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OwLyW4alEbKn88r8g6oPXmI7ZFMxiX9JdAbK2MrdrMntXmFr3K+T0Wylx/auNbZl
7YZh2sf97cGEJSF7OJR9N4+Dq1u55VQIqF/nDtwhGGtvcPoW8ftohOeTxGTNp/zw
3qWOzbJohYxrjBC2U5FT0KwFNEJJ+u7El6zLvJQQWWkbTV4Cv9hR5wtEXnSjVNe/
sL1mDj57EiGlh9iMmT1BAdUCncRSAdR7n6zyFoQmD4AsYDwRu+lj9BkJzPRZMC61
evEe6RBHusTHsIvLcyRQS99adqiXREAOqOXy2Xoq84w4M0uzAT2Pr3cl5/ObI4wK
2q5+Icm+ZJd/6R1CJyLOZgZz2sa+RC2jr6GPYNLcg4msYLk3z5SkbHoDVWwcfyy7
hcr8f3sfmdySLrIclJph92AL5XlQys/0qTXsEUYUjIYwlGztRD3S2XmKdDctH7rQ
Sd/MtdttTd+nz4fZQNn9QYc6zl1hxyHmJvFx6gWM6nt7N0tMIoJHF3+R6UFy4xS/
ZzyQXYB5EDBusC8pIbW3/dthSn8/qn/VIqDNJjfpPuJPw3GG60fCxT6QFhje3kgY
SUAwjOnc9llcBFZKqXNthLQZTbb+/6gpwrR6Rv2bHtiNFa1YbstvFhPtHitDklYc
WIqoI7dsnTA9EzHjjXogMnKGns+mzKArIMuRoVf4UoZ0h8HUxnEyUFb6wWDYOfqV
0/TS5xoT/zz4y7t/rLJLcciy5SPgn2plRHJ0ZkDHoGSOfl7HPtgm2TYujpLguR8E
PXZ5zxdFol/0PhN8+3H/WpmuXYq4wmvEPM/k4HPry+kCgUDttKd83Eybj+DbUm3T
0SFzK9mcP0hM5u1i3h0ekILBUU7VlBanjgdoWB789Wb+gZKEUat1MYEZNfQu1zWZ
sUktG4g9pms6v7+1WUiSJkK8vheapL1aUy4nes+eVAElLrUrdJjETtTgBc4Qi7rt
Wb8EETeU938HD0ebnlkVop4tr2IigCRatwzM0Ll0toOpRygGk1RuLmGP2A8Q89Fv
aAhhi9MQZFgN4PQejrAhLP7ValT2slus1gKofY12C4bXAq8h8etz1+wTe5ye3e4a
geSp+nmmbdZnOQ/iP3CZjzJ54eVobP9vw9X+a+vH8lVn9jr1HZ6XevTUN7qfOyZl
Nat5i3rjOBpP9UnSq0i4nv6ItU4kOZ/L+L691bmL9lnnh+AvsJbQia83FmKP9K6Q
x2U+2rGd2EQIYwVXR79tKAfjcYXbrKS31JbtbTH7je5CNlZLNlc8L3on8VZhUY6t
1AnSIOJESC4nftw760SWMGt9QQ5VkSgswFZJzJTpkfLIiHy492scdS0aD4ks1rbM
cnsAUbjtHoEKOaowgQMgfKswV4vy11eFJeheW8SOG3AzUJKgwaecKhx4DLrzGSLv
Qm5Or8W5iXSgUKBuW0eFqjHpUY97KkJRza448DX3Pxs7ryeGDqnZKlrzs91kV66j
Y+vVWPYcRLITSVfyqUxglRJBqg0lQe5z6dXpARgCzATS0sZtSSeyB6zSSZXDOKDF
oPTsuMu2NbCsEJQ/327klrfus6MLcwbWlS3GRj7BfeaFCWILUddsoldBA38GNxiA
0k02IFnnqgnLUbU5GEl8lqTynCXbKyIqR+ipNPoYtnbPpzTsvrUZanhP9Kw/Izrn
OD2TW82cnrS79aujbnV17X0lQsRDZM3B2AkMhtk9hKGrDyGugOrFnuJdYY5VmxW6
AkIwpZtAOVxE8M98jEIu8HsyKj3Jsb0RhIn4vPzE1mPW2Sa0PyEbYdHLfEHgxQqY
Ij4CRSQrXjVxJQDsMBHPGicmsu7A8c+/BIRrfIHhUqasE/jGlDzUDp8DsB8+BDc1
zFILR9C9c09G+Iz4zG0IHqtjfgoahs17euOzgjlYlYsackKHjrLJTLfFvaIyi3vL
orhISi/g0M3XTrqqXQAtiWdpLu6mZuIAIjKsZ/B43JT7T1GcPrTMQATXH7tmT+v/
qgrCUDOuMPuQWBdknGiMPItLD73+Qz+4Ki2yLbP1xLWrieTuUqrfjIQTRefrYyGR
bQ4tRzSTec8MqjTEtrvdHrAhrEk2XajIEqa7RsKB9yiW6awof9iKpj9cIuW70Ybg
uvS/8aYaXJc2Yb5vXyzTAGIki6SWsuG3Tk5jNU0YX1Fr0LL3Htu02L/8qqq9Rfgd
0X9LK7p/4G8eiEfHP38yokW7OJEYua4v/+vgzenwO8W79om0Ccex6vE+r6iXuU8+
mQUT4tryFMhSD/xDOXYnCTKMr1moLGwPxukRCJQt/ZXl5WfFoi+c5QjImkTOD2c9
TBxY/8K33Ew2fJbTbwxGupSdIG0xae2nrDTifSyhQUKc9I6aUZiHpc/59G0E0UGM
yNb2qvUnmG9QijfVxAeYzjxMeKOGg4C84z5NZmf8g/UYNeP+RP8HEc8GEHAT7iLJ
Rn4Guf0QmYH6Z1+tEXE9jpxzKxffnstZPux7TrEXC6tMwTpsk+SzksNqYwwIHINK
LJ9A6t+QeeJVt9wU2gWA5xOUTX5il8Xxwlc8LoNDPS9nuXVqoq8XjySncj8gKOF4
SUEOlf7aMy6Kmt8G1WbvsTaBrAdbB0Zmwp5IwTY5i4vvj0izQBDVF2jBkuqXioLk
X71vlL68uFqZWNuZoVJlHlaZMB5Slvrmwmp6C9snvUWEviCYrdmNoanRoZ9MHGeU
987LgGpaVmTqcvJUcGPvnr1hJq1N3bxX2sFSoAfNIaARJAda7PyOCBj7QRdjAyy0
vwSDM0uBSrMoSLGiLL95PxXNtuvD4jlfjUF6zFzs7vDmFIU1Vl3TYmY/gF9mOyDJ
x5JgeUKQTt5QGRfHZbx6D0AnHRCNSd7CcXou/vmEd1R/ZcwHp6tTDHmvXWF8E09z
kMuxrlxlzao6aU0ZzN7Oe29Sarn36pQir3QTivDEeXfxZ7jmUXIv2rbZ5tg6qe+3
/h798dliry8juxP9Cy3DCfz4v8uqMNT2yC3/cPh24R0XNZXrOxptQaBERpXPaCnw
Ate71A3ltTdC16Eq3HtTH4hMjCNMPIlw/kvVdDq49yYzy1CCcy85Xn/ny9pqRbzl
Pc1KLKzT63FThW04nQiNf5r1SpAxQc3rZht+3kJel0OZvVtBFnJVz4Pnsyjr5zyO
Hc1i2zAN/vAIumlFadoDRZazUROzvMybWjrKdggmdLtv/1bB4eCXaG6hJPFkJejn
VHPjxS39yx83M1igj+x9DEU+SALq3J/bXrcjto9x18v+FVFmQdDDW2p+0ZLVZTzb
bmNvkNFpBsG9eist/WcsvfQVaJI4jDVKHp29jGb8JeHeyuz2Kc1NN0HgP7cUxaVR
E9Hni8lVlXUPvk6WMk6ZTISKlvrlJ/kRlzXOcUAyJaUs77guM+qpe45aKqVFdUBk
mVFeXUHQ34Mg3aRMrNqVU6p336ZpICWS6DOaZsT0fyfBHdNgMARlw5knlum/OVu3
u09KFcEAMEB6pdW5hS7PivFSrPWw/q69tCIYCtR+pqh8UV6TFIE8+SzlLJvnja8e
R+1SCFnuF8TiG0RcN/D2X9wjbBRbu5Udl3/kQqfNmixLxi0+wdcLfVP/gT6p4kvC
j4TV8mzuBaUQoF2KwX0i+FyKim97QFlG5Hss6DwEW666PFOtD23QTzb8jXHTtyZ1
D6Hmz/+h1X86bnQBEBiAenqbyx4ISfv5MH+uNQtPAs+Aij6cp6l3PkQ4KvdtimFM
sWmY0mq1sTPXEO7a6+4c363GDU5Q9bW9utZWrkfDLVgdkwV01TOXoQICk35bo0wv
v4/YiaVNhWBenHZtP+GOeFBbjkzfryb0k9Mlge+eopz/rxmaKmAH3xSqPZOAxScM
f5GKuawyD9VMaYnVz0CGcSEkKvi//5aYn8NI0h9LCKlbE4O8jwgalFgQ4Qe0RtoF
aqaTkex97492KlCxGCW5SCDxjs7SpdmRl9NoEmihHcZU16TfQt5GYWM9TClXywoX
ic/1IJsnj7TN+vZPy49lWSXNLzVehR0a9CGYjZei06bkorAo+WVHiE9wMUy7yaG+
YHQkL5quIZvMcDg9HTq+2YOFkN2eqwrzbdDXMyVkYKqZEi7aJGUbjCKzyPJCdNkv
rNUq/4GDLD+rQfmGBFXXbQ26EHYMdXXdLGZSwmqMFo2FiOPFGbzAtxKNWaqq4U9T
ONSVZfrOnxPTVUh8g6xx3Y4dRJUkdh3YwYaW+YmbxSEvJ9y07z3NlE/XfOaXvE44
PQZzTGZBmIguQ+d1BLKZiYKGSo5z908RkAIhbnwhOPcQJAkK3g1HHxjUbbQJSaTY
nZL/b1Pfl6FAYee9+7QnMVp3X0UZ5XGBY5I0RhTmAkq6Ffk8AT1KKE4RiGs50Z/B
3KymWHY7kEZ1R7tr+OYmqobVbwW6B3FpkLLOkIkbrOIGW+k9QPBnZkuCS49dd+LI
+DSw718In4IsQ6yPfnnhYRuiVwepEK5mEQxM6OIugRGaA8Z3ZhwC4qnUIvEthvPM
HrwWma/ixvUZV61Ddtcdf0Dn+KkAsKnH/ABnnw/9B4e9CwC+vnw+tBmQFj6qJPQ1
ZGwKvfGjCmj54FINGGwKRpKgk1TA465DaDxMBJlnUyRusPkyimwsMGeXc2so3ZNO
nLxr3YYG7iqZ+eYt3kC/cF+uEknbYz+ihMMHbFbpyjWUQLcLawjAEd+cU0bp4ll4
8td8BVmBdaqDK/16CTVGBIeFoxeLbYo5yikP4RCMUhbuG3ulkdko14HOqIHztj82
BFxmFkJ0jbeU8rJowAtdtEa48DreOtRQR3tiRwBimjVenwwxtFtTVhKUIOsgv2MO
7g8c6hqfXGnLaIDvCLBD21kWhkTdga8vivBI8ITskr0HYoz+jq1bCc6aOXBrwpLP
gFKOTV8V5jxJYRFIP9grovOyROtdOX90j8kGhLdv4tS/I8ktVzs4E1GkVHmSdGw0
iX6WwX37Pfqj6Cyn5yWGEV9FSn+ER3sDUaU86Lc0qUOXkXbAZp7fawexx8C0f8Pb
Sjf0S1oY47WcxrkH9UprnT+QDObvDtm4j42874gDAF/SiVpUu17Ir0zj1VorFn2j
10+uHcR8BSfztoo/lifGY2PfOgDOPBcMS/jp2R/ljFwupzp6v65ZQkfVw5A0JAyy
9JMbhwshUKUPO/Skw0rBZBo+A1oNLNQsRlxFqh1sReq6XZlwTIDbbZMPNwNIGEne
Wq3cO2fcEaEXdqf7Vkx2tLCRiKYCRQ6IEvvoUVcKCtJRQ/gBObeKnPAVkPwF2esN
4EgEy3vYHVazDgs4NieDt0tNLMMkwz6IcWD0mRONVApnlrkSQYxBWGKbFtIw1DBq
U/0/pfJIL5XwnKso/TvGbV9aDzkhFaei/KicSHuPQ9IU1s1af5rl4JSZ7zLLcl+b
Oc6kFhpnQMo1wOPHmF7h2Ppjzj2/YS7o5Ta3kcWq1VY5yjIQZkbJJ4gsV89q2Zp/
ZJs3dfmh/+FHtQtUdyiV7MyMFDT583Zcs5PepjNMntwuZySQA1YNIjtm2ES1WXBY
eQC1B+8qygO6yPGb5FAHlufH/c3BBqRBSCViqq3unoYAoMTU7i/rhxS9B+mptPvV
sQKSk3hV9i/32FmhmC7fuQTaBLacv+KRS7fyAaqBpqlWVjp+mXqGxkB41XvqDgcS
ceQFNKNrC7jdt8nbHBK4+iV3eZWjzKIOMl82oVclYTSpa3+2CqzspkxyiD0otDVr
5QKrD/Bx5HQ3Ks1KCCH7aYTJiBLHSVFmX7L5INpSItHxHbWNF3G9uUgh0IxpVAm7
ZLCEdFAi+n+wBFkSzwAPCCQQ6rr1B3mKSprGvQAPaAffaF1AfLjuIoB7LG4fhPAW
f+P7rx+mJknRw6cNIp8o9Yau6y876Zbc6rFomNSY3yUsUwKrhzOpcmaETc07AAEj
g43K9OuIXrsw91W2ShNewaEj3KPtXiJml1Mj9emwdqwswbqlcKOjam4J9Q6G0gJ7
7c51TazPyBuJ8VFdSxowESvtdpzDw5f7tmuShLJ1POu9/9wWtfw3BPXpi0p4WqdF
ZTVJuDDl+Ji4sgkn2ia+FSx2uTXVaAGT21p++QddC9drHpa+uY8ZNR5tsVzy5qJk
gk0qCEEPmAa9aqfdIMC/RF1x1YXBr8hritbz9cVQnvBFG3CYV9qqs97EktHzZnTR
7mOJAXyUkImC1kb/BeyHsEbj4JJvX4RxVESfmz/TxafPZDLtHbxXGDk3lBe0UKvo
i87FVG1bBiUKLLIdx2sb+NjAr/ti+JihdIU/bFC/u+aJJg1GNkHsCBFxfdF94IQf
T7ZfziKeikhetjw4JwvEMgPiWP16E7yBacYtcUwO7Q2X8p6sKW7McYLZ+LW80Q6z
MERkALpreTTwdpwxwUSmcypSa3KcDHu0JyQqKgGXThXFGoNP0qpDYNW21HbUsnxl
VuKSvGYkKquwrqmbTJDMqkujtoY3edZDTi6N1ebx65neNa0KTCLXTgPHmjSzP70q
spRNOD+34mFNiC6Ktv8jC2pcuu5rt39dVHJYPY2ALQ4LZjXhtRuOvSaQsv0cQ2KQ
+ALy+bT80PlUwD2bI9Z+RKdrElUJNWcJigrffVG1rvqjJhyDNCfY/5b4dh8/mm3p
du2106Zo2ygdlTDnzcfKD0FIyzKVI9gy3aBgbJsQwR9imTJzCGG31/CZF/7vplS0
bCry9ofSJoCZ9OqWz6mArlXOFuQgnUzA/Me+sKJVmA/siA65Gey0EeV6UYvatt//
2YxCU/h7pOKC0X9bW5/yvS9pwXHP3temkWxk0n68Es+t88+Jtwm3i0Y3ijoNd9AG
3r1u+Z5dO4dz8GzQT1NId905HJE2/LQf896N+FW8GwKGacmgOxFKYhoyt9D+y1rl
0mXHQUtu4VJHCpvdRPu5bp+D18DIH7yJkVQHVfPjrbODnDr4CVCmVCGLHs5K6pnq
Fb0GNnDtVcpL+RLJE9YrEHchPpfTPxRuShMLHRbrfH22SflffFL1HnPovj/FREgb
8h263ls2zMR7844d5fppws+PVMtCdd7tT7A0SZun6ZtqcpA+EU70Sh7RrzJpDIwY
/Zqy5in7p1Q8XtPMYCR5byZ2JSBUnHmyKa4RhdOgz0BheVNykgZU/sTMxppBt9hr
ViTNkMbfdEe+VGHv917O7YWPLs19yYQDy/ZepscksyW7Ep279ngsnp8/6AVcouws
LK7dwRZOmF441DiqIxrxML/SinO/8NiXiHDh8IdETTZ4juPn9nz0DDXmDwgy3Q71
HG/I72MFi62BmrjC/Z6kkPcq6G3glxlwxvz+PMyCrYlyzDYpXyOH2i9vvJqcvVjx
1eyHJuvfrXjkV8Dw/X1C6e+/StVqt0BPJgUu0PHXnec6GEReya17MkU00q9pb3h7
8ouPrDLGMZ0fTV7BMtZCTt1YI20DKtWu3oqHr1ZoC+2WhapFHOzVn27KdzB1rOEf
2N6mHFY2zmkMVYTB8yPH3Mf5UiwDjfllg0aT9NDIS1KoWxagGmD9OYm9bYCD6ccU
xK0CqrP1CE5MwWMTESCIxi92Ah2Vyx8ITCHyytFxs/HU+psnE0tdHiddj0UrsQXh
XfxE7jjilkhiqK65DbQ49e/b8/K6JFgxSpg4zP432xJ1xLD1b4bdQLLkwj2kfmHN
4zg/LYcjoUuEG0xXZUjfltvctcyoxxbJRqdFGjsEXK63pqeNo5yhfyZJhaWG+DkI
sOoQn+IoQrNLk8XIBfrx2VmXzf2yvwJk/fD60K+9XASYoK+DulIKkShz4yI6ITIc
hECpAn0gi/X1/p38xlYApwUzdGhPxMVuBnVm2q8SEac4i8jg3i9nOiDpujDaWJFS
rk2jVJTl3m+HNbpci9FlOG5QBPVxccKhQyJ4y0m/XwUHqk8L7pxHbchpvwczXes9
vFMmPC92oA4BPRfcerTD5Jgkw+s+B7DLlEWx+EWPNp/7v1OfjGu7uHSfRmwcrrtP
wQJceAVOJglhesd8B/LD+pJIY3rxyDTqGVHmZlycZuhO3AG1JJYhGcFRMbXhVvVd
NHgOL6YR7tmh6fFxSRLRCh4bvdvF4LUpmyLl4u7a9XJ10DNv1990ZvsZUMCDPlI3
H4hi3XTb3TzyLdQ1YRIJyA+Rc8i2i1CWIBuuoiNGo33hJipPW4eJvsNRL0finExx
TAliSu3Iu+McENIuClkmpfCHDaxI22SS+jpuQwqHtkGASb8KdUy/fdnZo1PKFb/l
q0kkwNFUU0u9F0p7OBkVdeNwruyGWK6PfAmKR7W8hBsyhmGxaJadPmfHPFQ53JNT
pGcXod64vFMA+HAugw+PqtybhbvZFm4sn+zKw/YUw/ZlYNBhTzX1j+fgH4CcKYTw
ELl1TqMoP3I3ajQx6HiTWnM6mf/qYhQ8wedrzi5nI7Gg0M1gQyVrEoE1CY2YIpCG
3K2UvGTAaYbMqtoZNjBm6xjcQPf/uuZEeNsea/F6TsXVQJZlqpHsNWYzoei2IMuS
vy27NFxz1yhEBlKAzypifsJkNhAqjaSOLhmubarY5rjix32rsuwVDRWMqcSteXvN
efiVH3yLijP6ymRrOfmNf78vf5T4O0iJtk1kMycnJqWE+yJRQBQJifEjSwBjnvMm
h5TzX+hLkDwuJed775dRdkper9mSxXW6uZaTCbadMbhJ5iJEscATysnRi9AXUITZ
TZoa5uxNqcwEoOaxLWsF9OXzxrNyyfzR/p95MtEg5tHTzBUxizMUUNf8CWNs3IA5
WmItcXsWysCXAyhhYw5DlJFLZ+xsGb+pt8kF4jr5WNsk4gfeFSXs83/TZe40YH7j
WsyFqMhnCtNG9RKt58myJt0JrYsUswKDbERWC0Lovf1mfM16/7EcdnUxLBMttIv6
pS2dV0SIxbOg8/5+CSds8zvtF3yNlgw7VfYtKAysXjNTtiKW10AEsWgRSmuiMZ4/
utfk0u//upZHoMPwzMiw8YWTo4xjwge/CogGiUzDOcrqUITAv99O0JonaRr69Dho
jBjgdSptWmXzn8jIoGpcwkPKY+4rtC6he/WfGiuNRp2bABF7oJkniuMNtZEg6IOL
TIPcalf1eI7Zt/xGm8HUlrosJRqhsazwnReZSzQSDiSZkVNZzkc/s66aUYoH/dH7
j4OgzeoeClA8bMva92ImU7HOOQ3hxseIrEuj3dKeANdFAvY6zyJpMDfAE/OBX3/A
XVqxwpyj/pM8gSaKKt5JholG0rmXCLuVNIRHRzEtdCNnJOlx7UnhszHL8LWtCOqq
W4z7/+ed4Ngjz7JFR4s5t8A+BuksQ+NqEjViZSyRhz0zzCCJAr+2tsYPQ8Xn7piH
xKxM2HT4MSmS507IRzZi1xySCgC8NMk+EiIWh82Kt2iCjRbeF1qR0J/exJu0v2gX
ghZYSMPINzozgfEsX/MJeaVcyjCqWrgF0juT/MNzWAS1qMuCAoyr2ASiHsU9tAP4
x+fnOTCblUdzynyFiK8ZcB/4FY/ArIA5+eXKBSyuIgQwQ9rYbU1MvTwKlzf4R/j8
zkzrDS2LbajxXJeNvodw7ZznVAN/Dg9GRdQ5OhwaB5dqSurgUWpqewkxS/lJEUKh
ketPpgONDcxqikuGk6FQ5RGl6p0NVaqMTZbep7gYsCxLLpWW6waHE2EP9gEuHZ5D
BemHZMVNsQwk71gAVdWZcZ41OHyt5yDCSImX8n6Z5nOqHdYQLYuxtqtO/mvgPIIS
MxYvVg+jM8lSPx8jjfnQv2wdyybfeMfCKQf1q19gQB0wV0istLONRTGlmPJp+3ny
mRgQprbBcmm3dJHHq9BMs4aI2ZxxZ26qwuY7YakuZoncWqiQ7Y9xz8BVXpN5Xl8C
HKZlnwDi6PsNfjIEuThM5q07kQqKzRHOr0/aekLsSzG6683ELe1CTtVIqq9hDpPZ
aPTyXdI9FgkZlDKbjX6o8N4sAp2XHkLqwA8hUlEl/tBwHzWiEGSCuCmPJQLqUH3Q
LBv+NynDsw6Qfk1hMGUORWkErELpptuYM+b2JOvHO8J1O30huyBl1gpyniRirc0j
VVEQ4z1xAO652MxsHeQN3U3iNfgtKTdK7I8hUh9gp/4y8tCqWQurWkwlee0DlVRg
Mt0dlE/O/Birm1HiDbv0bWCkFVICTB0xR0rpBaiJ/L4GDt2ZV9dkRaYB1Kop6cqx
bL2V4zRDwywcNXNJ3/Djn8rRhKue7HPJZ4yQ0tgWNxvSzZeSLtRmJrW/HiBPQMv5
L1Hbm/Y6Nr3HxZmWo80qDuAZkVEA2QtDl/y9JF1J4UwtuDd9B4I4Qf88FhAhGBlQ
zRHB3BRKZMy36TAmb9DAAWrBtYNLBkd5OjOBaPfwRdZihdKjicEH4Oc93EENn8CW
PnT/ATLJ9+5iaAdPlqg56pJ4yaFcd4562hZDc42JEjNS4CMctQfXQ4i+GDQ8f/ae
BuJNvknXtv/uqumlHANTnjKzIrvgjwl1C6W8eHO8F7t11SkQ7MDOJmszxE/leLiJ
RgVOIoWSis3r3fubojVq5U+T+iVchvf2Y/6DSuhE5UGaZ7lb3ppgHiSgPql9LEBE
yP5apUtEUKjics6al6t1UHLDbZuthGCRyY5mhigilLk+1lqzP8dLJPnE13OWifA7
339nw32mr0kYg3bq8Pmg6ydiKOwSqMoWBqreSKKPBQ7HjXiN+p5q5oPKlgJIraSj
MqKoKMpUG1WmgrLc5K/rIE7C6WDlm/R0yxJ6LYss5imno8p+EC4pFcmMzZrX3PQM
erKyPymX3DFJ/q7BVOBSWdQYkPER34sEp3kTxMeHJG8Ox5GQv+IGfWB7gd8Eslr9
fif4r9X213ZDX9J5+k4xsxE0FFZBw2zX34ZRDrvt/sV9+A6Re22mboPnnZavBgBo
LGmbQtCZwF3I6PFHveMvgO86pNLCLWFMbeH1JFufdxXJMwTrU9rT8pvyxTqJ2niG
hBQCyJ6TCUIlGzSwCzZGTgmDMN2C5FMt2asBKqJgHW3Bj+PNTZ0sxq40Ex1wxkuE
SGTwki/lHzWEwtXlXoSTD1m0L/aCY9XRYd30XwoOo6+Yo1dkw7DNmCClJ855jq5L
yeRA1tqt3GyMyM54tMeo0br4BifIwcJRUuZ380lrgZBaGc/pRjzN/QDNwXDDrWVG
wBRY48UJq3aSXSOIr5FkMsfuV2mkMHrbEcLvXI5yTKgN3jqA9jt1DtR/uGmBfFJV
f/O6I4ajshmV9lRX4xcGiBGkKb0+ebjYp/XRrMy1YozWFb92/Wkg1RH6Fnj8EQ2Y
ojP9YP0i7+zWxNJlgLiULTHG/Tp2euMdGR4f+ipG2VWXDNiavcytgXZG4tO9GCO6
dl9AE5plxosKt7DBsw91y1kys2eYXsLh/cuCTgfLwYQw7l4e0bdU525ZUpZw02B2
pblqQhNB32LN/nTmEzalnfEXDWvuK3Xo+qGw4uXKjGdHAnBflUuPg3n8vRuH0vcI
0Ud5TI2mfImpJ+get2not+5JpSp1gX6r5HjBNQGGwKUy4tjlrY62f2ZG/qt+34uH
1UD8C8ivDRE0AOfSQfFdUer4k+3KDrUFuvvPfaiGgdMcn5wQbT5DaHzTlXoM2Afp
n3+BTBlB0aDXKcp7JLQHu8BAf8NSajFDle9HXQMQlNzCv9EaC8hkHgaASxP/DFTl
1oLl41nhGC47EI2w7GNee7d+xh2kGEZ9cYCwjiV20vVQ6jzDPaIMk+96tklLtQkn
R6NqILYQM/6AXhis4gbuvz1N1VlLuAf3owvT84ZrXslXvESEl57JhvTwQ/KA/HeO
JkMXiGeHqmEGYIYkCvOFOU5a22a7JLeYmicDE2DrBG1kIaru4+C6pBGaM3wwjAgm
5Gh+w8HXChGdS6f/dj7JuzPomqePyBMdG9TpFYQ6SuhCLDOORgTWzETKBPkNaf/P
QmpOC/U+0cppDxiBEAyK/7qfe0OtCYmrRHnFS+d0YoB1mBsZVgvxw60MfNUiAZ8l
cs+bdvXk6HgAYgYS2PyoYmzZBNZ2HcS9Vf1frH5Pw45omUeHG4zu6+Fcm+d3WhPs
Oas799pMJo7YCQP6i8nIYetNN6HfNvPkOTlG1TABZMOPC7jIUaJrxoKbQ7x+wi3Y
xhbFGidoiq8o/NFihpxdhWdxxslSx09dfeJUTDEZN4xwu0FV8HpvbQkzr5QBEK9O
yOwGZ6o6yIgLID0jxng7mXAdlEf+9jqMKuI0mC9WY61+2npMZPomt2k+nN41LmOk
IL4snElUNeD1Fii3nA+u0Cai+MOwR93go47H4XzGzyIIhR6xEvrsKWqu0QJXgC0X
oIrvgH3MIjk5j+dzFexulWLLGvWZsac1NsFhsFkPc7YLZugX5SlfqwmaoFcAHTjH
LHuFOXv8wnClYzPQjVstW2himKPdL4SNNgXtxilwDTaPh77AhECR/WTHmQmbcL4x
ocRdO0omRaQBnB2dXR/FShNco7vNHE9fMvfMM2CHA2miq1eurI+ue6xY0NkRLKsR
4ENtFBphPfwe30ZkW/6GXEAFNmfBsLd83RGqtYEsBhx0zuPOqVzmqpSHuZdKoj8C
c8YsCBvEN9TLDDRJ/9kPOtGrTFI+tB16p68OCajWyonhXnAegHYaOWOSbWhorzey
lCXopiXsnoxShtv3WISQGKZWBS89QlgWL1vGmQs+91fsQdKaPkOq6uAD8nPl6q72
PiM+mRBdUuhz8+EBY2K4ehRiZgQSIziE7XqCVqHiM8hYRLkMtzkBo/BoqoWs8AsF
oqKWhzqTMJ8Owd4GuJ5MHDmy+8l9icdCjlEcB3FPRO+bwsrQqo6POkD8catPy+2a
ZeonCh5ES0GgegdIAEbUvFBk/rsw4LQc0xjVoEV+vJFaChQlXa7LKh1iDUOfboUZ
XjfVni0abFG30d0y22kUusc59l59Ixmiakih1joU9Yi+9grA4uOxgh3ZTHbtMOYk
fBOm2WaQo9y2jN5zfTMcGNXkzkdbxtN6hDmjdY7V1RtwHa4QYKqCL8R5LFiEV+la
GKSCBqf7LBUnDbkecM6QpOSpAoN5ia7nWkGFCeYwdPp2sKBjdQJa6UtTL5t9CPgg
0NDlbcNmCQ1dNXS29LnjUQuRcDvVaSkhhMS0zNHz+vbg5a+O+6okxjEBdi+fsoSf
PnS0R9/pzlamA50bzjtLlbta8VqZzHKJgRUkBxzurjp9lsEI/KAgKzHNAdhPRgkn
7Jf609KI38zeAnafcK8lIM6E38GloYpgA7ee/daozEDJqIOI5SKQhUao5PlKV+A5
Tv49iDlOQZb/5anuP55BzbS+3APaCMT+7NfsgD87PSFeUdGBRNiv8bQwSJPlpWby
uuw3ehb+7TEWSBeuwrLJ6aHM5AavW0z03tLGTGYBjZ8CxGC4qV+jOOomrzrs1XjL
4c+DOPJZN+Rz+xG0DHkyYCMnf9ZYU1qTV6XBj3NgMEB7uvLZzHJ/HoyekY0bQjZd
RaNcup4wVlJkKUguDEv8TYwiLgli3Nc/P3JTermDQREccv7k+TiwGCPLSUdBeFQU
wm3ibo6tso/I069BwFcW4T+me8lMsDscp8gC6c9muwC8SqPRWYT8/70dP4QPXelf
tR+2rzJH40Phk/QkylWrhVo73enno5TdZD58OyRf3Vn/YixD0zt11gUcHtW7K+o4
wkGQpobPT0IjLg+8kcQ3lwy+5t33pw8Q7tfIvtBTOvdwVBEKYnalgi3UIEdKg0aA
mXsNsrqsBhMA+yoITRAtFAtfxWX4N4nm7IwkwqS41EH0D6tIdh4vOAr5l70fkg9Z
4eb/fjfaKvDgok/gQTEbPsYzp9RLN1kO3BcrAmZOZ8bfGXZarBcE+T3PM8x+w8Kg
f46yoM/cpiAnhgN/TOlAWF+a8+UxkYwZ/xxaiXluLMs9oUD5Tx1mzwgZW4CtoM9g
dYbd0xOmJk8s/knF6fFO5OREaRI4u6H2S5plFroArbWqf8cW6Gl+ziIwW4pl6Wpc
dQrQ7PztnLcKmIMTT5mWB64+wvAU3AfTKij58Og1MDG7h1IEw1WQO3jKx1Q4gS9J
//70of3bGO5rjmfFKiUj34StWzWf3+JXEcIGx9KNUwrk5Zu7+aHUhCa4sX1NOVww
TAiPrFURuWdM8LFwlLheFwu20kkemt+IV+djnK4oj55TUmBAJaGRNuRa/W3xWDKg
iWk2zDmIE/wPBwWHsLGubpId7VfRm6zvZrifNdg6gfgYc+JNwK4+E5UOu33gxX/i
OeQSf8qNetH9uGLUzGRSh9ePcfaGSdY06SzTUNbr5uVmLLTiUtjdy6zduKbcD4+2
Y3fw21Qcnx0DbK6Dv6J//87CFRWAyeoNfBsIwU+RhC+vjpyGMyXSKNBlM+RuK4rS
QlXUdM6Ms0XRi5UP/oND+WmNgVYkrGYk6ycceQSig+ZkPLxeLPMtElUjst5yNKpU
NWKfsNfDKWCDvzkKspKnP/23281Jfdpism+NN87jnIQVMv3pBhqTpyzXAsSTFJTt
zfak+lNyvl6woRB5Bw+CqiL0dgSboGpapx+XlYwAkODfCTG8BsXxyDTJCN7taiwZ
5E8bZiPZG5SFrJb5SThZaCos1vhnaZpDtwSmYkoh3ZwvcvNuHHGX7lIsG0ks235Q
bwD/I4YCNVCQ+VQS7QMGr4vmFGdpO9sDK/M9zZaJ8d6GQ7p68Nye2m0HZS/AyxMr
eUGtAaMa3GroyId3HIbZ780Pykq2nyQFV9AUcoAl8ciVPZ+EgCi+7EyeXEn1W6T8
LKL7l3c1euFVCEV1IwgTFeTsLNbweblL0KbQQwMFfdtKoAh3L6RskT3RlB0SU8EB
rSGSChWCTabUxTntIYkccTnuUHMt2jLEF1ab+gOWFQo6ZQOT8uZYE8VBO2LTx3LX
LteNKflf8NFlTLWM2lEyM7wazPy5NW2S61oX06xtQLj0NmTIml9Ux59r/3OhXVWo
NfpJLqGGvDwOK9ir44kPEoPSnI8TKOyyhNY7Oje+QjoZe52/2STuyusmnyp6Wye5
XOdScHHUnY/NClRAkAlxPnourYD6ICgxF2xZlsMtCXYQL8Zny9goE/GeRrQ6tR15
1QIfPGDfyjS+Pha7mN830dlIDvKlOtn8Iurr9C1GovMYJN+paIJFrcujqZdMQB8z
ISXCFxzqrXtS0iajfIx8pqD7Y65MjhUKNnBXhjNRu63rwROynLKjpLBN3eKFbkVv
CTrJ6TU9jjbTp/I30BfannMAQAojVKCPkVbRaATdeRC0xwAgWgsorWxEEvUOyUa9
j6zp7nt/JqhIIJpXSzmzB85q4/y1hhWBbdOavDiR09ES1Gkp+37yMEMO6S/SPyw5
Xojn+DezLWOMlBz+2p97u+/3vYSqA16/+zfEG0fl20ExqKcjeyhGROL4Q/gOm5pK
4+RHH8K11G2Y99WM2X3Il40Y1eD9cnPzwKet7Pe6rhi49IJY9ebwswcOYK7c9lZJ
JH/YqAc5axbQYMzhlFFb+MjzPI96Mm2KgtP/ZixW8VqqKg/IrYx7jDpnHSH41VxK
jOFxG/dET2Y6336+4CsJI2HtNseUICzuL93hcrqascE8ceZ45hkQvzdE0Ar1dQVb
DhgweT3mblE5cQVclSZBGuStbvhILRNJuviALlXE6bYB8yqEc24ToCMhplinrioF
H1bpkmWZdQAMiJH3oqclDMabsht6u4AdX0fHXXD+C+c=
`protect END_PROTECTED
