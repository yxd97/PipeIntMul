`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8DiuMJ7FoT44FclCRu+YP4uVgX4/gG0nVhSif/yOn6a3qwbt2SSLfZmTFJBBURfJ
OqK8DJ23qtGdiO+y1jivzC2YCxEwNqSH86PmeWKdLv8m9SgpeNJciGEel1ADK0K1
R8TnjXBTnb+tLn/BzlagIIQvsTCBlQke0WtEsEgpeTdeFEvClFAKaIL8pGeUf3EK
QCgPPAehniuWeC0aNtGy/J0GXKsRRiR8/FK6Pu5icc+fXvdmrPeXzU/QG1tDDJMR
E2iqPD17exFlGQVQIimq+mPaR/LPZJlhv0yu5VzGOv4=
`protect END_PROTECTED
