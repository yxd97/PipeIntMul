`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9m+sVpyodZQwhW0V0ROA3wYDf16GpN16VBAVTcIZC98hTl5mgLJlRFK3LLomc0PG
57APx4Z7dQ9v2n69j1InUtzzOsDlKHObA6N0HSSli9Dy8MxkMV9xEm0FE3/zlLTs
9oba0L/ZxYaPWtlfXhrAgTy9yVSmMWRdhYU0SbEsGamSNT/REzSoVe7M8Usx4yhp
lbHnns+rFqYFpIDBMZoG3t4B2pQYZDRy1hizZryjDi2d8n+PrGYiW5eEUXy7JnQb
dCn/WSoSmtDMkp96w8vBAj+Z/YZd1rDIX+hswfzZg2j/HjXK6HLV0UfcNtAnjbhK
gzgS3Y2WxG3cRTP0SNDrr4qb2dGun2EzuJMRz3eZLhXJ3ELOuZ0N0R6SR7Qo5mlW
/goFe4+B8j3nzvjAMAplZR2U8E5KRtQjlhL8bw89HwZbbF6MqNHad/RO7tQDunFn
WegofLA+DLGdfbSA6GGWNbsDGg/UNMwws7bMv8j2OQnNlNiPzTghIMAMk/7SfhCy
2I/fWnhA57Ybo9NuMoIDOk5zr45HEDCaBiB6B87+2R0h30XLyFO4OJzOITPKynf2
KYj02rR/yDAxhMOz+REUL3G45azz0Jj/oTJIBcvT/Wbe24syCWUhi3Yk5pRo1DG1
hFGYNCAxVFPX9xJAhR4j4WZ5AkMpOBX1rpGKJxKka441KJ1dLCjwCAqgAeRnfkoQ
p/QnpppvnSbho3hPiblmeNJd4l2n9E7IuurLQ7icePiefpjvLGVz/58C0s/RQH+w
wudyYYTYaYYXYRMNmCmAUdOlc588quAgeMlPV8d0zirIDrHjBfkCiuO4mKkr4unp
PRrFozUcbhNDcCgVpDIRPyId7PLEUIClAlvrZLCecJZyCwJBHklxXmpFlnnKdd8k
`protect END_PROTECTED
