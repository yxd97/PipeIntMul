`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZAoleLgWUws33WwieVdkVX9ssOIA0paw2a9FoPSdQj3TQJxqtMhrtoufE7wEZ7/3
kvJ4qid6jNxsbvWniA1gsXTpUBynOV7jCM8dA0G0DqNqHTdRMEfasbxiEIYFBaUg
46wFq2IOvIoNGqDrs57OEX/QP12lmwWfQ9YNwiNS3SL4VBFD8f35zTh3d+kQdrHD
jSBqwoCajpagf4CNNs1OxP8wH7Uh96aLp8Or1cDcU4tnn5Y9uhfWJiH5/UQ+rr6s
icPKNG7ApMatGEtvdTcPc15ZTGComV60Z1FRohzkNGXciR1YboeLj0ThctRKEw4I
q6FOZlWZ19vyqdrkHLjnK86UYW8Z4Hghn6Pkoyb4AV/W3MIk+COBX4BzjtLG0oxn
ABuE67myre17CDv3JB92Jp7ZoyZYoroq0Ne3yZYzqR7hqkG3Y9szwiUxOaJyzw7E
2dM/ZhO9opxuQQ/rrCK5U6Vpy3QuNV+IGRD+yNFbQSFjnD7gGQ4dduj35Fh7qsm+
Bqjz+VJoeeE8niZQShnn92vbLF7D6Ung1peKEiMLQoqUkJqM+ToCH/lsNTjY9kP7
xhN6u3+xEdHNiLK1DyBZwMV7s/YZBBY3kTfx9+e6BDEyHTYj/lyzJ9jey1H2d8K0
FZGetbIQzuOm2bZIUjbLdFlQO5cBfGZT2N/U/VcM3lJczQjRYXjwYITDS+g3sVOw
LQhD/gppAV4l7t1MOsYD+Wcv30vq9GXEnhqTBXeS9kSUwQwer/aolQk64p9tGPUs
cUY0djz355HAo5QIP03S8e9DvL7oBqBOjX5u44ySZi6nkIqWskzHlGgPiUf+M9Zm
fsz+VKYeSIHAT7/26wg5rBuWcpxBgEuXmWu273mhsFWScJkpr1wQ4MX2bFnMqVDG
EagpSObGWyEpAku5QkgYKg3bpSAGXcItjFanaaRQVAbvEhx9h5SyLo53ziRAfMLA
Crr834AlaFsQTNIpdAWT5R8lZkFsgiWzDIG3gJKRBWHNM3Tibg9zXIXiqzzLPLUE
Dr6DgLVeXH4WWU9sWFPoyoyfUYUgtFJeyIBpOzHsGmzJM27TZU1L5iNicmX9CsDj
BHSb5r3+VJ0URTXOKLUdyxMdPh9fotCbHo602TwN0NzK50xtn5r6EkFYXbYe5AAJ
3ZtiAzwvola6LZEIhG86xwhGGmUExwxtvOlelBIuxyFXEEtMkcjqjcj6qn2DeQGv
PWeN17b+X/qty2zF3rhQtRpKvWBF3U0x1LylmmZ8FKQ+C1Iek98gw+mgex+ZcHoN
iYnGvKBYAsLYqBPwzbpf/vcB4/np9LeFBdB3YkSiCG2Beu5DvXwuV9YPlyef2JJn
Au3SzcwDjA1pNBi2Rs2wAufGiq2VVa/S7V+tl3X4UyYGxg7HgCnN3Nf3nw8xgaF9
fFj6jPYkpni8uaM25ZcA2+g7lyojbnuTKTe9thO3mGLQb0rjVaMkjITuzrRAwK4Z
jlkpyVUBRQvcVqqjgyad0kbCJh7QP9qTZEdUeAwrDy+Te7hTIUT9JiJvpmkeBQof
osTHhV6FUw/aUuyLxyXSX+Ctt1uaZtVzi+WkKApN0kdj2TdU3K43m8oU2paO9tMw
/1JoIqD5o1V015Ya4SX+bqqrS6CAvUnh8Ctk8c1P6lrINArgNZbOjkoVoMbg6VPS
IXrKI7bfOVpi86dZErsqdfFqmd0iyn8idmoiTcDs+PP7DBaPURpDYz0weHwWV3Gy
Vp4HqtPGXjlXAn7KGdSOTzdju0yZk3DoHfHJGVM/ysjsByIZiG7rX2dyEk8aZMDu
qk9IjTWTGOv7JbJg4mYVpd9JLF36im+LH22Tw+jm9R9oDEqSMFhIu5EvDIlHsk1w
8zIJh1nIa2281C/MqUmrpr1O9zShbNmbADpshTK5h32jOxJ1IwIJQ0pGdWpSV3NY
+FLtEqyTlbNCyeEGjP1D73/lQl7A3MPA+BUW63wv3kgYAS792/9qryvuMnVrFTbB
6Fs8TRRY/z1C3FM8QkhmiJKRefl7XG1cFruk9f8868b8bSklFvMRcMBt1eziABfb
I0sDcJLWrwIwbaEgFdPRtwvkXHZa5aVmTRUEn187bUwcKv93sVp9tDB7snNJUwS8
INFIUHaWlMn9mlWCmyvMPiBoxdW1zzID3fXBQDZ7QJ2LPCYpw1mrHp8CVIiQlcRD
MpeNpUC6V7CQTN1QtbDUr6J88DYPFK45AZlOXcna5mPSawMaAWmG76sgB2tfRRol
JJZ0wVmXfsDhojrRJPBjtavZUDwcZWtkEZYYr8glQzQcZwkOWcQlgVISwdgLYPzs
apAvnmTallwtAEUGvaOzmHvn5vBk/3Q7uHI/QT/Y9maI5Q7b85DY0nvAOc1XClgA
5wEh/ktb/t62qVIhZStrSJ5MlZDTgfuv3Li6wI4hmdQ0MMG9dxWjPRnyMGlDz1tu
wNtfh95ySUBaa8WCvU2P4phrtpDNy0OINFRapu0SI2iJFtNS2hZLpy2NkagliUXU
`protect END_PROTECTED
