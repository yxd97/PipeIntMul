`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xovevRSt1W5dmmw+kkHnhs0jrDvd2iTKCCLZh5b6MwV4ZoAX+OzLprn3x7JpA3Md
7bkXTRiQGCLjzei2hPxYPqzqJpvLK1/fYJjHxhFelqsx1nQkeuVNVbTrQTPSXHa4
ykT5f9UnlkFGaFSLxMCslJu0Qi+BxPCSKELmYtvC+lUwwQDZNrW/hgTzR0d+Wlll
jRjscONiNXXek7UFQcnHYF5dzvQgW/MdmO2JcMtEb//qnQEXqZ7fCnUbK1xE8c5q
3IocvOds0A87ZkM5mviyHBl8z4kaIPCjyvDqNIXYPHOnvsYEt+zkzENlqjy+gnMs
yyEuZ7JTv7iExpmAAQXpCD00diYoQvhXXJ3+E1NlQnznsCkKjRwsH+RCOBNPI0Eq
HYHPikeoAOB1+6ewfhdYqSUXblb2M5pyMkLdWCjPp3pKj9toBzsQMOgUv7eXCMna
ykJKAAuPL3MhVQD3ITzlA9nSZP7Qr3k59ywPLFHmGjqSxioF2nhDtiFEEPfohfuY
HwmQWWrfIIkzMiKlMH6uctu6Ssp8l6HxVELnEfezeJHhps9VcQgLchUPSB5EEzWa
rJd3+grbh4l9X/TVogzhLvXW9TqboJvS/8VPi+Zs2cjad0qzlosfeKJWHTEAv+Tb
bgv5mUKAkmLAR6PviVCKwb330GtEtqNjDZxxjZi1cYRUGASDMaxi/bmdqZOQ4zZz
XUOIipKYANWFa+nOPgUvNHQkFWNuUyewcznaJcEv5WFXLdv/bjfpO/+ob4xq5dXR
8LvefVoq5BLcd5YQZeR8S+5HjMElXmLxMALep+kZdemihRl55Hrx0iioKrMxw1S9
uogI0hCuugFOgIMNPIvg7I4jsZILfTwOzo1iwikX+oTeuqWVGyIIikvzY5Jz8Qgr
wl72VT4BEFxj5nsYGYJENvqFOGFoOH+0HRcnzwmFmEJovMmjftArAWl9Y/JhFYei
B0hvNsPzNtGaQTUqD3WAURZG2tZNeb/NEuwzuJfD+laCkuCjkEnuOW1e6rX0YybJ
fibbEWhAXlyMSTQYGM4Sj8Dxe4LA62m8iUG5Pcf3yFkbDAy3bL6tv+/m3vBGfn6e
fLJxaIXJopdaPEsfwRIqHEq9PXcUk4GQOPFXOGGvnMTXQ9RuWx0txw9pDWPk5DBF
p2DRIc6Q7WRhMK0C6y2WUPkHnd/kioEjxo03Oj2wHmr2CRIg5wKOusuDlYagic8U
+sPCMKD23uwvH4qTECejxuvmdcLzSWcxk+hqSjrQXsxZvx0x8fKEdsbvmlQa8omi
c752mmVE8fSBqMwtNHecoTh0bF+xsq3IUOji8RAateB7E/0JidY+TX756lynywoc
4rV0r6tW4bM+6tSxTnkigg==
`protect END_PROTECTED
