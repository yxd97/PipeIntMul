`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VrnLK8bKLzoetw7Ots/1dBV5n7xqG7/lIQdJoy0ef30r47zE9NdriM5rc4eehO9N
JSM4J3WQPAky7qqfkDTOhN3+MbCo3+/0b/26WXi0bVUNUIJnblhClRjuqoVk8Tkr
+TBME20eByLJHpciHGvcRZg/IYYvA1M2h2mipmDbntK4rPBSqhtY1y1szunrWD+O
kV9L+ir+j3TvTnLlQiR6TUXkRrA38AN99sIciOUnrMaXBkS1AG1kosB2Qcnq30KL
qMi4dAj1d4CGqGtUaubq1Lbh5Glo/LAMKuZJhJLnYffnc/06X8YHPOB2tAc9Ket6
md+1daFM3CAKmxsUBMOVDpj9/GOOZoA7Nf07zn29MImDMsFE3B0z6/xwhCQFtm/i
+w8j342vIbVUKfOuzWcqkw==
`protect END_PROTECTED
