`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C0GvsF9JRvGyuNqpxktbj/nxPkHnteJXewAqiKyXcI55acvaN3fiwSzXXfTR7abY
eLOWlbpY89KBrr7s0ecJNpN1mR8Dno1CGhkTEbCDi7Ccrl/FVoMIZhnz6yMIzM7Q
e48qdCXtdh/NkEqcB9mV5hVkKC0sa++fk+A0j4ppQiVEIvWTX1TRLdRxp3rijTsQ
ekMkagNjyCmUk4KxO2XxSldnQ7WwPH20B4T6kC+pmegmj4MkBN4V46ntFi7Rkp0U
W3/1CzMaDJ70pjlDFBxpkftllPFHqrTki3zTem3NviqMwsIbY4ayImfLI4LdPkGD
9YvOr4m/ZG95Z2FMoTBmAPw32GmBYRlBlbn0JJUEGqEhatwzig8r0hkOufgfHrBY
5CqOru6Y5O24nLk8AwQvVk9EtKXb8Fcya72dwd6aVg4R8aYLZMSlmZXnhCkb72Y7
LVmlbVME/wFE6UePOt8AENfc2UUm+v9heTvekeBGUolCuVRNru+rpecLLH5HLkUo
`protect END_PROTECTED
