`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jp2eGxBq/5IBY02c2fNeNNgqdkJJJHdIRtj71RROkNGQ8OnDhBGXyt+YgE2Stfhb
XKg431nR2essTK8bvcVnVXZ+vL+KbgqI5quEQwDPHIq4+sFzZ07X9II5SpOzxFaq
RfSaAhEEaqFW98OWKJjJvcc28xY1w74EYKVEYmh4zVW+MjSbbkdrmDu5icDQ/W30
JFasXuAm/LV287RbejO0uCuQXssYljMN133phpH9Jgn6e1guBtgQtzLRo2kpjsF+
j3PJMFa4ViZ/46CROU6xqRhJTgkgsyu6R+Vf1HgHdrcDgBS2RqGAEa+IuCKozZh8
CEIg/vRfOvQsD10QWylaUtgByRuYGmK/uDDzGZvCDN5LydV1+pr0BkFRxkao1Bie
DGskz32xM8aPazPLmExj1n9+HNZ8DpgWsmkgMBX0Fo3dqe8LXkqUldtuSj0KirCe
hSZLKPnJ0sE8h+UeCbErpsv6NsdcqUZbWkObZdLaKP1LskB6Nse3vlWeQvR1fSmL
LbAMgZTa7qP7+LmtUy+BTCtg/OzfQ33ZNVssaFZ6Xk6aW7Z7jfU4tpy5BNFkwf4C
uyoxQuXOTGe38dIp8Nq2j3sWlw4lZqCiUzno3ciAh/4wQqZF3AuSTwqV4We0I5Ul
Wx/DNreuw6TsqSxTZGx16+Z3xnE6npxgPlb8AEf/FhRxff/nqjWvk8pDomrQL/hG
`protect END_PROTECTED
