`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M8u0kheNnhT8klxMNr3pmOdrticzRnrWzZgt57SLjobR0OPmsORvli8jU3f6+wbT
whCTjwjz4mnyD86d3jZWbFC7WE+A2JEI0MKGDcli8i15tNttnYIrqqmZmFSgskbN
NZ66eTHQPDUc/kHuqpESwvBxAKUEDsPSTkmarTz0IXSoEW4HCFtU/hsSo3Vc3Mqe
f5PY6iHaCvU190TN88+R8+RfkbE3Xwxfz9/LrMMGW/UZxtz0AgGhRoR4ik6ScFKa
87SzShNcmJYDa8f5ePb6SNPsoFmEXNmLXqQmXQ9smFEA7lWj37kHDQNmrimUMAAa
w/ogsIVYmjLzIk29nluhM7CdIpWg0nP33HuqQtohCoEekzuTLOokllr3mEpIqK6O
K9Ig0n0mSlfC5WhYecDfKLmbBT4ClVzNeB28zTcIsPRqCXzpHl1IX0RCLTWXuTTd
nkLKTVropmlqJeEIGgzEXs55hN83hwr/3Q2m3+2B5LeoXhlu4BHUKispEbU+F4e5
W4xZWVebrrk1A/XJwg1W/wOkD8HfzQ9+q6tM7K/AccrNrdW69BRsfrdg6U5aulaP
Whxmtf+I+9oZLd83JDI8avNhicOb0zIhvvhotr103fWIic/k5M4n39fToiXNiPB8
TXWMeSNu0n4FDSpCYAa0b/kk/NbHwFgpOBa1uvRM1hg=
`protect END_PROTECTED
