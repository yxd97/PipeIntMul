`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxKk/fevbg4t7Vy7gjgxl28WVg68XunrFwtVf/ZQPueY89auilrocvlnpw8/b/GJ
b1Sn6d1SKYz5kOSygz72QM643G+oiPX04zRr0dv80hdbW7ENUk/RXOankZbwjROx
WtiApNruCl5XkyxZpjLWc0jnYY3n5Mm6CVD1jKbxou8pqwvN12zve7Yh1qiqkJId
Wb1nQCEFZv6nU3N2lBFMqBplVHH6uab87WmOqB8vGL2uTk6dO+mWQIddGHngsD6n
GdETeKzzzn63Royi/8JCTpofAles46zhcaRN+2Y6s8KFir0hF4kRfKfvaxJOvHXD
VD09rMi9TPqTasFyYQWc8qnqf6oFy78XhSWuHG8Xj7ZYoo9NX0DruAW/A0qiSVXa
9SKIjA3xc+C7dAW3SxvZIQSzlurtTzQoTbdhKdVqBe/UqptvVQ5B/yK3odad1H7i
UGiI3IKzypEGmfL//Cj+0PwGjS+FoyJ25RY56TgQap4laCFSChRXtkjBeWRAnFNy
52b36p85VKvpZg07/MQItSXIBUEN5QwMkdY5KJ1K+ZDocVWC8Vun422wj8BTu47Q
COw3fckfnfOduxd6DaVqJMdQ4XUUUODAo0YggfWqUGuW9wawY1Kmj8JAa8+8Ukge
`protect END_PROTECTED
