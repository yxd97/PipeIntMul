`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R5CVXLdvy/dfhzJTfCol6wPuluwiT9XIIWSrEn8+M8eBpw4xe+PfVri3AY9iOpPn
WT+wsx2GLN4VW14jSXWZRycWzDuQ1MUzoNqXtGkCmGMg7mCnC0MX4WMskOcgAIK7
QYa0SVDPSB2F1XlZnoyI2qs+BwyNdLy+ufSZlUkuAy0iHgRe11Wc9BMh120AYUWi
BQnnfeCSx8o0q0t473Y124Gp9KB742e+cyn8iopwdJx772Ttxz3xtBHxR2yQW5Hu
Q9wX/t33i7ggrobO82rTaEv5Srs/uDQLfNOlqaBTD9aitx4c3B3B0QHK645EJ0Tx
YlgluGAslUs+2yIV4DR2drvbb/ntoFiSQWOHreCASncYbEnrhMrKcMKFY7QQ9rW9
tzvc9OvQj63SBYSLZIxfT8Iy0JK1qq5vOZ3UYhQzoshP5P9BBeJAlQuqIXVUPLJ6
A6FFNArXOQNf9iFlDRh0qed0Dfy3ztS1JudZSkcSqiVCYlax2nwWkELfqaWZyWbK
UiBmAOYVG/gtX1W5ZowWSnk11iFRy+OHhfhXXSg/IWfWMcVB676St5+rceLX8hst
Mu+tpzMjxDEMDAETspkTZON19H8sVeHdSdw0NX6sxfmJCnOz784MK6zK4HS5FFFf
BFCWRll7RxPxintjrRTGM+gVOKyw4Da/8FS0541G7s1B18+C1gRCGPjc86zi4OPm
L/nI/we0o4d94s6vzA48M7sBEO3lx/jrTDOPkovwPJpsh/+Gt9Pk0pwtwRSmNk8T
OehV8yrq5tVKKmOxNhNFLCOyJsfzi8++DQ/+Zf9xdG0IMFfK+9b5dWLqtYfuVOzN
MRNDbiPXpCZtNrIyrTV1rQ==
`protect END_PROTECTED
