`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lNoHeQXjD+HO15M283rDiJVnyUer6IC5jTTFB46YSWbcMNhd0umYZf42c6NjASKF
6H5IX0dUv6TJMTN8BJ6MnZqanW3aZD/8cfbNk7Rr18ftujTi8ka7+9GadFnZntlo
fI/0hzTuaEYiJVWFPC/f8Vhw0i9syfGLBTMnXO/K9EwBkTT1a5+E66bmJP92Mo4H
+VSD8nMPS0xzpo6dMLKr4dJOAMdmGJATJrWbinlotM7FX2pyKt1VC1M8pLDV1qKr
UhvcxLEGEArgV4QX5Cq8Z3NMFHHhqhL3iF24vYNQMyxITSVrV8MnybKzV3c1pAQi
Q3vbwm5Hf2wjDM+ZNSl7B3DFnlMixUkS818gnZCs4nAU/lt3xYRBItWvgVUcAlZ3
6R5stVf4pqGfcW65KN8ZY4lCevbYRPkN+E12l92E/o1AdVYxhlkS1++1lR5q3dMA
6ljz9EW4ONEjNGiHaun/VnrTrZq/s2B3KLg+x1LJjlOXDa72XtqrZeneTp6tZsOi
IsEtqc75DGI8PthKDNr69wt4KeH94bPcvQjORfI5TRz0606Fs9cG8hvQgXjZ8VAR
PFM1RMH22K7X69CT1QHdYsu6AR/i9T/uV5Xl48pZuyV81QYLEfIZS09V5racG9BD
nOdSfYk3CKq04z5oMyRDKtNFMz5Z/8/q7rfeNwsf+Vf49uD72rQa8gCtt6r/KTEV
YedSjYI7i3awUoPnMAAlG7vRJx65oyuzBotoQFPkADORpK/NUVpTCMMmOMjkYPrD
3ETmohpfYu1OV6+GSt3OhzYuB9KLHHjp0zzcwlFQ5v6jUyajurxv/aYyyaT59Ktr
l7w/fTfmiLXwYCgbDjXODANjKuOT0Ie6tfunMp9rNRk=
`protect END_PROTECTED
