`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L908tvGri5j0YdxEGDL3OsN74CPFs8J6r8ehoehFwzWwqoECMmaLsMGscle4mxOe
tJpTedv3bp0QvCjtS9piksOisB+cwbxE/HrE0kVr6eahvhG7DMcZDet19fiXcj0b
2st3pOvA3JTNpLrnghW4VJMhtYrjsXmI8/ao5QjTnQQdDpDE1zrUnzonhkYC2+Pg
YClyR2lwod77rn+0y6n3eCNcQ/XddtUt2D4hvCFZuriuwf4fLuW6NYgK9UYynQ88
4L7cZiWKaiqq3JRLDFmYLHp10EZ5L0oW01R0i1hAVnA0FGnyVwl9NkngOQOUWDlK
EQKNNbjOpp0k42tgxYKAmkNNtiKdO/zZ5zmKRF2YOl1IHKnXxyMEdZGl05IKI1wU
ax83mox7c8v4eMcqd/HygTonD8FIEcwjy1YjTXc0X3DaYWH8aUrWnpL98JydHzIG
C6wshjwFVAkQvm3JfNcCFHE1DC9P/CrmyflGgSuyDKYmOilSMg4x8to0THa8nZNF
pLUjvDM3AZNiD9sZduE7nHmfBgtRs5N2GT2ZXBZ8MI94IhlwmgCQeN+/uDdW3WA9
nWkRHVRk4NwBi+JaFkTHgjeKtBT1MDNN+yqQeZXlL/av2Q5lZzMG8kdXJy/QP53P
L5ILq+msELULCP3oT35sWTW9vgI8Q/IyScqalEiN+FI=
`protect END_PROTECTED
