`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/etZRJH9JYBjVBWDo6VDxRrWjSGVh3pt8bXcpdFa7JqZ9W6yGyRRZwv0nrNkgbfP
89iOrj02nsicMZ+AXNQwSlnrUXeyMvHT42Mb9927WxhQXX70XVQCELWv7Q1gBLX9
hfYU44b4hY88+8tvbMFT7ycNt4aEgFmuRqXgb8vuILE1rOH/idV1uM6p8e0bSTQ1
IxWCbWKMb7Z/TPUdDfMVNQ67ujHoL5f6LKtbkUuowJvCF0scBhW8dr0ymJh5yFFW
eLuR8ZCVxtpLqJQ1eVSgFQ==
`protect END_PROTECTED
