`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YKHgycSZuvAnGoEP/BhI1SiLcWoSz+u8LI495AblMMPDP1wl1X6lQ+ShczkFF1Sq
Rvamc2fj+98TbgqeznB38NJpZ75zkBQDafZXo3vs2XN1845qhOYfuRo/2iBthJfs
OpMzfuGVSEUdwqI/hc/GbnW4QRlQaG2XG4V9xMGlCYJWQ+B3ktLCq6nbWYe/Tvz+
nxeuV3y6r0vQnS1rxec6KCvHYeFKNPWuwRzK1NthMppsrWzdT9XcNge0KvA4MJ0M
YqMTXlmwyHUblh0htPnQ0odhHMHjYK8I25aLnLadQgLN4GLSl4mv4AKRRTpmNbbX
aH+Ugs9hPC0SPSWTAC/Hr1dviWmvRLWnW/xqBv85VzBt72H4GJ+f6iyvslfp6ayI
94UVOuYheuuXQxdlo1UUlW3jSzXPEnVfv7xwviDwcxboBHfS6iE7WVy5Fkb93aSe
caIoedbhqVtKtH3iVTbgbfk6MyM/E/RhrBZNEgePmls+Vkm1XMKGOgbY+tM+0HUP
`protect END_PROTECTED
