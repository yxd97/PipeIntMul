`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8iaJU+H+NxYMzfZwiy/8jB+VIO/3Gh53Nl/HKMQzTM4DE7+N+Ys61AQpDmOQ4sEn
O6tjCqGQBphJ5rafH7PT8YHoAIOt7jCbxAW8l9GARVHKcQttXLFkQFT9lCuXU7po
bqh0nW/ZLKK2InmDIyD/JXHxXrnzUSaOB52oAj6KUj32JTyTIbnG460T3PDKJUY3
PMYm5HuOW+3h3lMaeoMN+bO5nm4micX/ylvF+iVdK75qZoMn30xTV688A+NroVKa
WFX+swCPjvjleWacbsiqcQydcbQgZnmB7iHZ1q740sckr+2vPf1PFciLTzmQgzqb
k6BRuDGKC67lq9AFiXDgdNfS13FHkkJ91D7VqzXasY9cVfSInTGfBRfvxg1m1lKL
eyhMKSwuJ0wIjbv1yz/+8UOrTVouYCFEZZdkszCDXnfsSEo+tihLw6Jt27Qnt0As
3qBLjs3ESjsDTSGxfygCWznl6lrUmu30g3ol02otrp031ywa+Bv1yM63O7SEOiRE
`protect END_PROTECTED
