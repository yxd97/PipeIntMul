`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+Ph4RovmljnmbE4bxJXfPJ6RnlpabK3FD8wZACtskwX9eXalMeqn/ubuO02ePc1
WIrFfBqgXpRi/N3PYUPJY4QkW1QtXROh03J4dPcT7s9ODRVi0i5uNCP+G3yo8pRt
lt7hFvOuOuoHMvgYjmKg3w3qvbAouS418loSjk57r7jBelxwlOscGdNZkkuMaHxE
8yrI5D40ABLhwRrKSW35bK1qMamE5HrOXVG+AYbrOnNOWjJJFsnim9O5j8bsFbDe
AjTkGy/jJ7kjDm5nqR0LUYaAvbvy5f/EqppKi2wikeHUQOf7WTafpjaY5fOnLvOC
syVJMd8kuuhDVYm5oOsfC/t+3YP7cXVmXOSF9VxNmTwHkprRBaFVfVJNyrqxb+6Y
QVCuQWEoMk7fPCxhg9oGzzTg90j/cV5byCFG4IbVfP/smw3oZq4FqedLIHsjG882
6XMbWQ5ra58cMMLh3ZXdrw==
`protect END_PROTECTED
