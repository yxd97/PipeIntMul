`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BTBY4285R6aie0U2m2SkhxYxAJhFRQxM3o3KNykBUEQRByQ6UOgbSAHHYEO7/P2D
REzCzD8jLCE8Ud3Xf6gsl6PgRX70fghyVUgw2Xsf86Zoli4T0yupSXgocu2ATBna
Q1/oh3F9Hhy/Z3MeyX0ehn20Z5iOLRk6547j4vmM/EMD9qHbi4rizyy8kGayCkZ8
1O63M6prjSCyW9QLAYM8y1JYHBJ8NC/k/N338Xs1rYmZqGiRnleYwuzvs8FhqxN1
tH1d1WhNpQEixuXu5ndag16aWgMUtZqYqOeTGJ/jZiahHKLgoL3ZX+S7q+bCY7aE
YNAHgSFM0CbJHjxMyOPLm0CyCrEL7jclOCwxXhXArkv0mFEsdJn2jZ0KhznwQtfY
1hsjNCejUww7ITohwSo6B3p2k/Cp+7jo4qV3G3bssH5y3/ltgeVanJJeBNVt8ILB
vwxJqvc6MD7pmRArpkCa8Q/F45C6cT7guTvJLNmol8IdmO7sCNNjLhYzRYKW4Q0K
182GjkVs0hfMipgv6/UNWLbBRzGrocAn7mkL+7JdxPGJ0ZZGKI9LsBv2bYSOAK1g
M81QYCrQmGIT3SvYVhWYEg==
`protect END_PROTECTED
