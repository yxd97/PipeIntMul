`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naewdmFSDnkNIO2b+IGbGjF5YHVy/64giaPjqOMwmOc/itcwSZ6vz33pu56rJb3v
dGKb2Nm2I5iTxLpjAOwwDrIVRoL1ee1gpWxikOw2bglgdoxA4HXLwRLys11zHPVs
ajXefYX6oE1OAxMOzm6fH+X67QCS/tAeKiN0JjR/s6JH5edPpE3Fh27awr7ReEak
oywkBlczXdvXlPS/99n1LGDB+UMzuCzVl9Vk4tut5tQ70UT5HiCA7PXMAxir4YRD
WBT4KhJiiTk+fTOeDazxnhdeQiSAUfCe6Gem9WCPZ00wUQgCmUd2X71pPIqRtE8j
BBvHpAq0ctk9pyQF5YijLA7tW8RUOk3tCon7eVj077IJVqwIDxTEw/i1q90bS+4P
oCCCNrip7gMM9zoFjMbjIUTOZdMU6Kv3nsFz3bsLjWMa3njOSJYp9XVvHLrEMG15
A6zt+TA0UIXy3nL9EDCQfI2Nd+YF30ApFcODVSA+254RtKzCwgjElNFtSaGzkblH
+0PzQKq94icEQ1O9Agg86NJnAkhv9NGcRMHtBeEdRHkdTi0rN63ruU3qfF5o8Aba
W+9VHAc6MAQWrAVnzcpUldpgDGcq88cy8A+PfZz57cveuZ0lMudpfrkZiZH2hIV6
e2ONMLw9RMA4kHe2GpT6N9WRmBTDz+jGl6oNyGxvzZHdCiK3EDdLQZfVm0vRVS5l
qrTXsc9KWljaOD2txVDIUUX2ZRMr/PYrZhF29SX0RWKI8xaIrwTrZcFWaWpidief
RVJEr0zirY2lLdX8TyoVsFd8AM30e+E9NBBJeesVznMa7nPEC8F1KGr/+mXaDIhw
kA500IHrP01PlQA04PO5xH3/XLuMh3b/YKzhj85vO6yEfg6tQ5GA60RjspAAm/q7
QdvkDp7bvPKOGxdOpOl+zIiJvjcPSte39VO9KUDdu5xihOLTLtkZUbJ4OPanPptS
brxbiWjUoTLpa1tfjl/9ejGZ1oB+XYvhn1To8flJEDNnqX+0staa/5fgHjV0UX4I
VzAjZeRX9AgNLvG4MjUiY4SNwavbi2A5MSlFZT+HMUU0OF/BwlRvFecC8VMb//Is
udzNLMKKmlLHY0G/tTJiwyumYPFJDaMajTT+6mF6ceVuEzUA9yMK7RKvy10YLTxc
Gk8N2lOTBG4QNsgICiAcSj1cU08wGXGmNe4mVhxl8CCdDIuHXlQaqsLqOQicziNs
5Akiq5SyJRp/aBTbTb3Pn5gG+aoWB0ulj2XofEmWm+Ok+dOjhTsMaz5ZKMWtkxx9
RnpKrhTiGhYGDsgd93NT3jIfr04wYPSlPePxaYv+qxUlKO+XWOvac18/EkW9YTMh
a6lCB1cmTw2mzM5d85m7u11sej1p1mKLHfuC+ehXbSvziKSdgZMm/cjcg2fzXVZs
yyKtN2S+llOJhz0eEHSQ0wVN8iJKVdjBD8BNMBJMJ+35KKBybZI+3QE90HADrWri
UvbIfYNcQZWOhlqwBYg51wuWz8gsF+5oBBBVyXU+RlZ8K4wrtujGiVAD9M8Ui7MG
eeU02VFTme0n/o96r2/uX++jF/LUiAigbBGiz9ZomndEzGi19Zy6Hgh2bjeTGMfi
Y9+WZ4ejXb4O2c5pOMMOI7MdyqZBlx1gEWsXoFDwzs6hV/qeMWDv7JzRRghdyF1K
Z9LtoaIWUXVyyVaaXCevTyMRL64tVU1FoxT0kBS/CjiXT9uEGFiG4eP9rqhfEdkY
YzdqJFYcY5DqqtGujKdzmJcBLbxnHvPABTgDL2FbGdMrO9VcJ9HRj4Xh2wVir6UB
4VPHJ0eoAfVbOXKLIDaEwtGXanYL40kWbvFzjXy9U2shh2G76R+zzazgLTWtJtpB
DiRdE1Hmigsmd4WbMgjNc20e1SYuLozLjvidoEmKOgHXmXhJjuTZeohADuWMionu
fKB8zIpZVJahacgZ6oAWjudFniqZzcB70pYbJTyAZ7PLYb7AhEaeCKd6WX9iKgoO
ETUsWSrQL7I5YXcEvYXXaz2cHdYTHStHJ8QiwXvcLJaVteoK2xff2/YQxbUMTluQ
FCMEDMXkbCrLbE/zKBp5c36Xl6dwP+ZkL0kCQTIbk0Or2qMM78YM0kAY7McZnpnp
KHM1fVbuZwwzgVmwBHQWkwALSCryFu+gDMh9Pnqnl81LaAslTODA9Ei3TqXdp/+/
H+f/xux1Z8KqKN4XtVp2BsDXgbYwo44KyK+412ZLSMZN69UMyDZDbI7IL2nUv7Ee
goMtPLVI8uv/0j1afDowZOO4R0hhBL0uwrn+ImwaOXK6sk2nnT2vU5F1GoqicL0S
ujN3Go5t4nScZZdP6SzEq3+c7zYrpXLym+9Vasg3p7zBd2SizuI85qU5LHy2DNtC
rr8mRDYIe7tEZ0HOawptRhj59e2YLXndiF/jTuHMiZ6qvrdKdKBZ9aMwe8icmHvK
EOK9WYp9ZEdd634I8NKF3gAqUJxwL7fj2up2ZjkEX8+zfy9xtRX8Np2Ow4G1vB2U
fmejfNQSmE15og7UFjBjlkM1gs1j0se6yq9sct15++NcwjHmPlJALmkPuKxZlvp1
regMqPdOazyMpiJbnTktRkagT9AlctOP0j3hCSWrrlgRCumLWiNeWi2S66fZROmq
3X+86G1GoN9oWSeq/PcDaIOpNcjc8DIHBXfBGAUs5pgwR7OE5SCzHavz5qk1JlrK
4IYzubDnxow/+PpmIFv6YQJTwQ4ksBIwUUbrHRSVMPN8IVdsz7veXbNEPfoUFY0e
kenV8PFjhOzRF//KuD8c9q/R9c+CIpFxB6FGISGXBBszh64NS9ONy5osS1fG74SV
WyUnb9EOp1aNkHQ9pcRp4DgAjhhLnhD9bxp3I0ppGsadYJcR18rXjv6Xg36xKDIV
MggKLN/Xu5uqYJfANJT/yrEYoB5aPQtlPVMLSMKqlt7p9cCaUSs/cIm2NwPeyS0T
EfHJtSn1ldkFok0FapjKc2+5i7qFTEvdWbSknqMhUEmJNz9cgYeEj0s8gXQLam/G
WeiaouUOGdd8iigMJXsrdTBgWVhkeYNowcoGN35814UA54Ei1wcSKN+jFa4K/7pF
DEpTcK4cLkigNoSfbemGBfA5k9Df1AuUc7oPZz1/GPPoJpbxbyZvicQ/DUqucL0+
Mt5Ifn2br+2vN2m/CSsJkUe0xrDTVWXcZ4awehD5oX97J3hJPdNqYWSWyBKwS4AP
NycLWa7ktecV7wh/yq4ll2cu/7iA2wLvWoWHawt7dSRmr9IKTi6uKYx2zeInyGxy
wo9dzJblSCTJzJFct66DWUToJvym3ftVh16LJRgQe5aF/PxKiZFcrucCTZmgl/PP
zczJ5sQl9uzF4uxD/wghAWI5saP9KmxrM3qTC/TY9WFC8EKUK0lTfULY8jQzjvOT
0M59+jlJ3unaXC4u6irKBmF1/7nOBIVZdHaeFHNBIhy/ucAOZYWaELAZ7N3Rt3Qt
9cAGqWM6sw1QwgpPrZbtSTshgWEykWQ4eBiL+wdEelZCi+tVXDg34LCkvE5+mFa0
TfCOXK6dYvEGA3Zy00i0abtsbWLBqTW1kDeurYbmXxDf4zW7fmaQsOkdJbsXEUJW
raCidkHq3Pb6oyWp4mbgJqyX+YqQv4qpwQ9wlOEagwnv7UTSkeV4jLU982w/H7LP
r5FSP2QIToQJT1QI42SH+0+0Gtm9ggXcBuuZotQtZ1rCi7YbnaPxB8xgOKjbuvmo
SXgQEw3aIKqEymeCksRms2p0ovfNwrcHCvT6vSFPws0iGI4p6/0iMlWzlqNCwPBd
i1WARJoDV0QmIScdWvVtc8QRFJXIHjZ/zUgvOAfUGL7dDwa7QplvCKzOcwGGslqL
q99tGCbkq1RS93fvi05/33PkLrclss3K+/DGL7mjed9A0O1JWfOzurRqa3SYws5m
Cb5/JTXSB54fZVfYFzxMdjWaOVI7EkOlQl+y4EUx/FLo5B7kHI6aP7z9F74E4kiR
Rm0HktotXgnRHofMZRPcggTCTfgbnrL/s64AVUxO9ooVqMSWTvorBA3eQZnYcs4h
3eZI1zXHu+CPq3ytf4snuEVoxIx+Qy8W0CJtXuQ7ICe9Cpaw9mSY7tOdTcj7yNZ2
MspSKr1jJMfCrzRQgGr9ZA==
`protect END_PROTECTED
