`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QERDq+xGD4leZ7fJw2WpElzr9YrXqAZ1RxrJwbgEtdrJKOg/KKQXRW5IVSF3ERlB
7V+Lkb2JgccPpUu0Z2eIURr+VifJSk1uGOx8LeDnCvWxl1ZgKdsEx/DPd5JDLbpk
gcsvbkZ8GmAyJE7IdMhvWzw7cmQtlE5egtjuoGt3OIZoa279N38Uj3z0Onn6LkIn
AzrbUbjPoPkT0Z41bydieGi2EbAoid//2exOo7R4IEh0eNdnEj6NUxlKN+zJvzRH
6sXv30keTX6k6sBuM3M73kPJHDY/KJotQoX3kSchkvLzHppsYlVZMjgBIRjfrMon
9cCW/wpHqgR8rK/NcmWqfJE/xWx69HmL7HILL7YeV14gnOrbIrcP/pfFg474SEE6
78XPZ567BOpdS8/Guf8pW2+pLdHYmOIJio4xmgdps9NQfVr1oI6CFZlLUaEsAIE+
KW9hdLruLwqrLMS9oum1cA==
`protect END_PROTECTED
