`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
An1ZsvwSm+EivCz+ZfGnPJcCQ02QDmg1EUeNWxtZI1HXccksrGmOA137GrZfrSqg
Vq8JlzE7wIe0CzTX75WJJ333B7m9IT3n/e53uBU8DtIiNpWKxOYyehJkr0/0q70n
Jxs9M/WflVNvidjX0NSFb143/TquZtIele4a5PZDW7ln2HnMkWAifu0DguVt+J/R
x0YHfwK9bb2uHqzHLf40UWx0ygMrFDLYOjx5L0r39DgIo94n/r+sJEdb0wUOhrgD
oMWLj2C4lQzFIVW6nf8o2Yxq4BAsCN/1GN7K8waP8UNUX9OH3p2zeFEb7ouwOODN
LbW6aqvxawC+s8AQjzDTssHQG2KvVxzvHqYXcwNMVFr2BymGN2/M9HA9F9YbrU9S
8ddVKsBxC1r6sHmHbi/LExpp13JwuP2GPVQmeci4y/XeLt+jSAtG5IZLuFRAqlUr
DVYlJaY5TlVg7tIzCKt73kt/DA7fUeoh9jCFsi938OmPcu2JTqbASqf435UYhXs3
RZq22c0AdStDT9BEGqy2P2aBVZ+h74EhcteJwZ8/E7pDpLZYhqK+sG0hsbcls9pS
SQOU+DG0oz5dNsYxCKyuvblYqjqqmZmawsY/Kjtgvn+nvdywF2HqdXyFTRG6VKxj
KnxbIsXZoZminS1uABAFa2carVpFmI3/d3ZlWN66Y3klkMFuGX4jFf93SkYTVEnG
Eq2KLPxp0EYn549TEc8MAnw1L+omCdmUw6tUYsTBdYRW2hb99cz8usfnblQA828B
z1qyOpqEDiHzklm7etblNwJsEmydJ6LoDGi2JmK4pyRfcHOllmpKwg7sWaxnnvRp
vWfnB2Allii4r7t2Qflk0w==
`protect END_PROTECTED
