`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FGpd3fmjrtB8D9Rm0hNhUI4UXNI+EcrreFV+IC6NvCaf0KtjTlrRVx3o7qwppLRd
Uvqtg3ulc0pJOTSZYFZ9G1/JZIyQ6iVmk4vskZJUd5WUUCstv3oOl+tckgTAqtmf
WE1G2WT5YIbmIAn0BWz0I3k3AvFAJWbB7HqOZpetrNg2mjwA/4FlXLt+8GNlAr4h
fGdnOdHgxLNX9xqkxyInmmHesfJZ84LYyoGuyu2pN/DNbzX3jgqUvF3PIZwvlt+6
OsCnMdbCbtaOjZVfV0HSpV/o8vk2OLsb3zzPBXXS7ASEmUYrWLVQBiGQqtxlyEC2
uG/vV3peQD15qWBAjqMtdXgy7fyKiuxxvy8PMO+UrXAUez/pX3vm1PKxmWClhXuN
sUIsoFvTeXFli3p6MYMv/8rJI/4d99CjzbfqgPbC6a5N4r7z/08Vuo9Kf0q3TDKR
k0bPmE5lEBbFJifheeOlrssjWkuXIS6SBl4wd2df6zWtEof0Z+2w95AK3gAWzEVS
2T5fibTpbdBbiw63WON2lNMd00H/GCI+FhHZUlJDtOl8CWbYwkkyxIwFuJlMw9vX
OKnepR4NxF1iYmh1KW+zCa5EpIbUlmIem83Qp952u/EdhW56U+pnGRclDcqLhsBR
iTnYQwjlaZqgE8GrFpWft6tji+M86onVi0UF2JfTtJGjT/hkwsMdWARhWxmv9D8r
KAcixaaRq2tjuoMMb5tl9RLTg0Gwh6gRM9yipP2h/zNIXXNuGqhKrUEc9+rYCwIh
`protect END_PROTECTED
