`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7rG/O3Val0lI8jiC9KgZLNwYNhFMOYtHyVYFV1fDJ66rQPFDcW9DOW4TgRZsLyL8
GTSinung1u6kII4YqALigKNWMfIsdmCMlJsfkxSgLPnYAVio1JodZXY2d+pa3vQH
V+lEn5Sgd1D/l/HgI7CKuLcQeo1mNNna9aPFktiKBCzuW3dYkn1twCwZA0z+Hk4i
kiWp5w/9zFLCV6UO7Qfn+TjCofPZnoLoIeiOG5CHYkmKatrRwVulr8N3+sdSIbSX
SNc3Q7EzCypmo7RCcxjRXdIxeH9g/2DoNVif+6UyN3Jag22KAeJrUaro/MRZQbTk
tuZLEgmZu/CGm4iUpmfMJUQJ/5Xu6LF+nzvxxHVJ/WSLsnvZAoZedVK8q8TtHTsI
blvA/0arsHF0lFDztTnuZ1vVailxK9vZ6pKagsnkkDdJOTI7z6OsSbgsnldS5gaA
gxyXnzJc+/kLy37ZAwhZPJh3DlApo42N+Xys4mk+w4ztv2FDHFiNLChw1eWUNbUb
Ly4lA+/DHzZ9YdsdwAuVOEL9LYyQs39FZ2KdMa07EvlqbJvFcLYL71k2GkF2oCbG
ha8TbpreDVCTCb/VTzZK53lo2rwASjksIb/5j7+E6nlS+bx+LCKvU4QKnwg5FraV
wpIqblzIz70BmG2pasy7GkQpxW6TzLDeB0muQ/ZFSnrQObG2/BwgEFDEg/AFYwH3
exTZ8R7C+oJq7Cvpp2nN5efZNOuELZ9pa1R0YfCrVajbCE8hq/Fe8/d+mcjAD47y
AbIo8lYqkOA99dJar/YvxykZM+MC1YblxJOVHDgRlaHHXceI0T4IZu9vQDktRf6L
pCy8IBOfXsyfn/S3jPYZnlRaEyM13gfEmikV8Tk3uXyRgchT1jEjVpjeketPS5cz
2YfpUfRdddYYXkXfrrWuGAPbkKwlc7E40W/7KZv0wd6uZsv5R3xwyRY1IG2zeq4s
QwuYmlXWMTRbpR9bX6eCkiX1Tmv4esRTc1JxP/23dykEUvmKD9+A4+yllSweS3OM
tr2SbC5487PL13wZxSWQMRKfdBWAopsYFIku0Ksjb+7weGamB2jZuqyZDOjM9Wbe
g/vtDlbE6H+X53yVXJ96ngwjUiEdImQdI2X7qePh87w3+foRNwWSGd1CTqeNYLBx
UM8CRMHs2MvgiJjdVkMe9QfRU+6y4A+escvVIJy0kP8rbjO58nxK4wECAUrQV07+
pmk2FmNCQ0e4gPKnyqDoCTAD0k10KmMjoW1sePlHaixxyRRgSvGaJYwv3Jkw0m+m
wqRKi2hkTbiRDsM2zywrKMCxOLM9LRxCHf93rHjsxFAsMMg2Rh3VFWuhRAZ38M0q
VPp7c47b7Ap1EiSObXaY0+IF/HSCitBUI/HD5xQJFsv1UHQRErbLqjwCrkFj+wPc
DW15BPS298AadaKGhbYAZ9FLHThtn25BBu3dFsOQXoLzAm0iw60zasCej7ghexF+
FEuxa/tru6ts2b8awbJMFVz3e/XHeRFDl4gfH6nNkqbaWFhpyax1IR3MJDl05IDY
q/rIEPo11JkVMIrQvxFhSWbXydN6Up7S6z4x5gfDtN2UM9zYAgqAxxAYEMvnp4lW
DewXCf+zoc9o/+0dtDNCWqP0DqObMEGlRGP8OlaVZWXUb1FcuvBv6lrFWBMu5WoU
fn/C5pPsaM66lin3erT5uoJ5avrIMe2Fu9HIyrc36/+1CL/2lbyfOddQZGwPlfj7
N9rsbf/tSA56Dz11/3nIvX/3iMVVbpQWmcx42mEdfqdtrTmUUPExSzFFk4HYFQ+/
Sk49rIeBvZ/gME9xtZpKRJZyqm1ylxw6Wcupd4npQMpHgC4fKcTf7iv3w7qh9LSB
z26Em0NACN8lQmXFTC1Iz2hg/ySCOHgrdJwTP4+ACTtdmdmglPfGupGFfHeahhfQ
/trQ5xJ9tp68zpPvrLJU/2YROByEd0cJVx1p+c4HHwIMrr3z2BOmyTj7eYRxe/Dz
Gd+ohiXKaGFakKtEbaEcDTKQH81avqZssuj9rVTfoiewOhmzZ64ZVUiLUcOPklWJ
HawgvFMQ3Z9gvSSSyWpYlx7Zg/iCjEtuAcJynHkNh1qka2NFEsk1vPiahVP3uWPp
Zijzjm35mexJTuqW1IzQRCUhJpSES/XVdEmVnejbu2Er9/vd+hNjgyi3NWS33nfA
p3qpTVn1RDp8j5ovBBA78xPm+mVEHX56+EtKrlJIv1CaQ/S79eDNzuD8+reKEC9m
MF8fzVUuGpKFb9knQwPsUrXCaa/2OCsXADa24qQIRsAIC5fpgHS8MY9JgEGw35+Y
p0MkUPgLYfalegjmz82PZOA/aCtYQG3IU7aZwOjQQl2cWDuERJz8w1Z1+SkdnDf6
hyZmeDQpwgxeDQOm1pmx1Wxgz7+LqoAIwb+7Z0iCZCFSYcStrnTw9uxA+qT3CegK
4/ZhMj2cfMQ2IumKC8oB41YxYrEDls/4ATlq38ewOfBvqo1J+3iQK/ntGTNHrWK9
EV44rn+yLMr+aSmeBIKq8p424IpKHjwCz+TycibSZI8fih+R/1GcCoV9lvmtzEOB
0S8dZAh7+v/43b/rzdkdfUvB9JCv0h+SVLWvnKy45g9Sk4FtKyUO9QBrtSLiDkqK
`protect END_PROTECTED
