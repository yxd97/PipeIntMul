`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LZAr6tkIqC7pSPOwCN/A3YihzjxtwSVZWpjvs7Vyzbm2mr85rl7SJWFa6+/xmIev
7TmQOTSb8fL757hfrm3VBzmKwxWNOzaWNkK4gEUYx5nO4qdKGmqnEqr9oGsOGGHa
/UEl0/ihTyw5nJFi3Yif0fSsZWRG69w+6UR0Af1sO05ohpY3w5xXC6/ywas0c/pU
ZgYXH7QlN6yhmrJHeQy7dAT7EjCYLWyYDIBU5zYPwlXEp5Sgd2p9t7X9AT6JN6pv
ofZRvXwrrzMhhmqORR29HUzLpFonZMlD5DnV0zdiNERH0MnJphTBd8juPC/sDTC9
gwIV01O4Y9H5moC+ybGVZdt1ey1PEzty+6/ebkqxttNH34xK6RaKYQf5HcB5eX65
1ITrwIfJxu/iVcEydwgXRy5aLJ1CE7NLtkOP8s1XJdj1BGOCBPuAnSqhJ7QBgwSJ
qhFExKvIgYuryfZbh7Y5vWLjjmoUovMywCREPlTJ2Hs=
`protect END_PROTECTED
