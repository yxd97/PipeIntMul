`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0JqN9goudgmjCsIN0P2IZ2eFPytCFcRyYPXcDM+X9tRHj+QQJQR/C8aNWdNfuBXc
BVoYjThN+TzUQW23PTnjCZngkhdHLJblOQNMNP3TkKbA/O/nYbJSwPtJVKe0eHBW
LFRiif6dhlAIiG+QRYC6vQ00+NEAnT+MchNXuUOeEzifAW8C4O08NuB/7CgHVCrC
Um0j1XZbJeJyl/WSvuF8jSqer7UPwy4XZ59pAqxRNaT4lvQwf//BrizHdNKEMGCk
oza3+JgFw4A41QzOxOpyPGqpr1t2Yuoz6on11vzaI5PvbmAziHF9vmK8nuinHC61
qYKh/4n0hr5mj28FqOHEHT0f6kty7r/kEevHkaWD1yWOOgrH6GW6RfJIuVrC59PH
ozTMDc2PESGXq+6JLPOzayMTVVhSuQRMLVC65SEcUDcqWO91SMtN8xb3gmk1BOEt
fI8jRnFyAKz4jO6/icYwbVMHwyFQ3WbB3cDOdwG/y155k3SSdQ7cPCmpkEibO1As
`protect END_PROTECTED
