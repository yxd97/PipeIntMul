`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Jbo5jQYryNGxQX3CmR4DZj7sd7Nm44PIUszxcvV0LJPdTlWnN+YN5eE7+glJE27
LGMm5j2jvDywX3qJA6mHLs8La+MIGzq4frF5AQ0/UCFpEdtSpKyJRjoj1aPG8+q+
iZXaFCZEncSmR/iYIXqtjMecDQBv+rIB9crpHENrHkMXhWLEcIR9KMNN97586CsK
aHBW+IluO9dzBU0b9Us8DU5ekLxiMqYAeC90WT1vEpPeOdhs4Ii70NjicZr8E3uz
JggIcWgyMnylPKW+3gYp6APPC14S0cG8pzCN4p8oUW8DtgHNOfQeWEfjjCveJ4t0
D2GXYYwsBuzdvkVb1NAaWNCiZYcr0DViRKjvED6edpoUNqVhUKLV/QgEBQH4PCwt
AR/Fs2jV8VpvMPAtjNiXe9o4lspxA5z9he++qbN/BPe4LzrCEEXoFKhFRX1/V0uf
0nqX8BWqwu70b0bcCww4rwSU888YYAeWDlrwUMKyNIKg605kcNO+CiCDg/cHwvVl
C2nf4zOCeY+nCq0NFMdYszO7szQkFNmMzNBnp3iX1In37394+k9LJ9A9GwDn9f+b
95mXYoDTcVtOKrZ8XvAAihLftbRiklJHZe4Z4YwI2Pw+pgvc5rY60LWnI/6fIfM+
`protect END_PROTECTED
