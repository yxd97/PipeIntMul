`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ixpUF1xeuYAwyGfeZOljurBdlvnYtOTi6LY2M2/50YyxuGao6bbtIjCmuPS+YE2
6FGncdNR2yIUU9wCO/L2D6Ty59adCiFoyMq81tfspuPO5+rIpNCKA5/1JMtP/8Pa
+MeRApcp7L6L5kyo4qDc5jjENfwSrD7W4A8z+3bHGN6qt1QeBpZkNkRPFGYzwP2b
QppRj31n7tAsucXVZ5iWhf/sEItzg9W8vQ2Cb6ypzw9jXI2m3bnI69B8uAafAAS8
V2dCjZZKwOEDshiAC97Ex0OqtkJbwdC20dS0TnBp6gPDkF9D/C2tXWVhpVTKJStK
ifWrLl6SfNU4yV84aNM3IaIDLsrZYPemCuuqs/Zs5bJ+t3ltCMcraoKMcWPREBCY
tT6g85qAyC4K4r3k9JqJXcnKpoQBvdxY5d5nXFAHtqngWyEla7+QBjqPaJTdm3ai
hPnlZszMhyjnZqxmoM/f8XtKcvzRuJcuxNKpzsncFziFGOfLcmasDt6vix3ElQU9
gehCSzCEU+wDOnkC0ofo1HMsn1fC+/GJ+lw32mRIhFiwYiDz/vIkJHuBOl9bT3Tu
ypQq4DtpwXxO7UHM8N5fQOzWCMDf4ym8lUyv7SWlAZUhPAoaIZloEk7MuHhDuXay
pb4DX3Ks9dr/haO3zdbylrz7qE14cCV20mXwT+qPDOTnyU59PhMT2RmhJchC/vLD
x9WnDjjDQO0xABJLx1L2XqC+kuWhfv/roBjpwXP4p9mYgdkKuqZpX0NuuPa6FmTU
yl+7ouwB7CFQfRY16JlMozZBiYoHOoADItEvMaUfPg1CdVBQk0lOEPLociKOeU8P
tXNB6+Ezt0tOz07JFSqnBIj8CJefxGo/Q+x4kcy6jgc=
`protect END_PROTECTED
