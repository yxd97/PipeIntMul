`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSTOj7TG4JHN03whB9C4UsQBLnsya6VaKiNnDMD35VD3YrCEO2e4wQixe0Ma93qj
PyFyGx9IGtXC53FASb7BKnbSEakCXb2W+eMTh9HdQThDywK41QMi0RmRkTdmHdwl
c4k9EzeXugtfO/DMsvFd1qhpCtGB+2LC02vpvy2Nm0v2KMsZDtN6yK3UqXmy9fCj
msUajWy2GuXj+GxconQSZ+jb6I6HWIgyLPkcUV5sjUkKSZCdrEyhXeLmJRDkJH8m
Q/7do/zTFBjDH0UPQWPY4BqQpDAlwT3NyNyS6alx0EHfTpUOPY1Inp1aeYE3irkV
pAYblnU4lTjH5s2FCP0QpaPpHrsWxmSjobb5XGr/X320x2bHwciEZCm0yD4XBBxO
Y9rXk7X0zhZcDlZz49Eck9mjMQQjndhSGrUSlHySyqXMVXnYJA7YjZ0Pg6qPySW1
CGOWELxDigj7D0E5BaBakGWbW0/cj7vyymXBTnuaIHMPVctLjGFWhOd87icE7mAX
/zfOH6AdCk5Q3Uv8DFDDRnrNKyajGYPpmiNyNhWgY0TkfcsysZpthKZGaGoH+Dy+
PIZKtTH3GBPdVAOqihfy8rTrvFC39873FQ4N3/28S2nMNt/eYW40WicemWzRgc58
FtCIb6+bW1hx13L7TZH3l4Dl/az5XuHN/bSch2ophaHarBvWOUzIxR9cs8q1im4z
xArhHPEtsjOVJX38cA+3hZJCWDQlUvv8LPqmR+XSb+WsvNhChTVqDg/hZlxpybrk
aRZK51t9nYQ6A14gorUlmQ==
`protect END_PROTECTED
