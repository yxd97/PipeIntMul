`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pf/U/jXhfdqYalAAz2iMZm4vXM8oXhr5epEuFCyFkoQGVfPjRwc2hpLIulLJfKw+
pNWiwi3rSlqZ/AX8yRQnF/OSU/GPh+fJv60U4GU5Fr2A8dTLwYcNSMxa7LG0vjDR
oe82Lq4lSP7g7cDUTU0tspq/pHJRd9D31Hx5CsCD3cwR+a3ggxE8qHyP6i28Zkay
ZkCg4kSTELRZATUXVRLdgNPVAQePob51Byt6kpr3kJxAOhnhdIuKqn/Uoae2te60
StJ5Dte+jWu+2BgVsH+QGXctsorWVGASkpk4eROwkSodmq+PTsFRXUaQJE7KONWx
kpHib6iSWqVhTMpSMvwC5ju6nWgZmcGYc9QMkRjNbF+5O3nl7FWrlbBsT3emmMjv
cJjoI9BtrbWbhs5rnq50ipotVMXg6N/zJQ78HmApS7oh9nyHaznTgpxoxzn/tyUm
rmWyMcOq628MLqXO6Wo7r/T4sSdPrwZpQ9lYImRQcy+XWCza9+U7VWDLoKu0K5eJ
`protect END_PROTECTED
