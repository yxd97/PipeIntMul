`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqedIHoxh05xCx/y7FVIpPwL32RLe/cl0R4MkMVcVljvr3XbOrToV/PDBHFImvGK
KusJCiKJd6ZRnsxl5lgsxluZuAjm4xmeAFsjbKnPdG73tkEiVn/v/MMOJNCn5Uw/
nYh/rFm2XXhMGBv27zxwUx85sZxZ+aZGQIAq1tWlGIobF61xg6SEQ1IyszAY9iZK
3A3/FjqJvH2AMru3DA9AqxWVCm0BdOzlK5xwI4og3Se+7LuYNgxw7Y2GqdWzJCOO
0n5G5LLQj9PPIoDWZ6fK7hPLv9n/I6wjVNQbBE47kxi8vMStvyGRETRFre94jxw8
xOcMgmmB+amNVccEg/zWtFL14mfa9GdsiL35U69IABM10aOxJhZK0j8pdAzovB/F
vZCzKm0YUuIX8p+Brb+B7WeCg4Amrla0j+ud+2oeONbS+bGZW0722QCFN8OoSq/T
h2Oz0hEDFCC++KLVQ+B1BmzG13e4p69RTHbCjt40VPAwgQW/fXPrMLE9GGXeX7vY
oGxuGpkeOUSyDU/+4MSA3rLFWhBzj/0Yto1LGSSLWg7gUyFll3qvVr7i+J3B2HGU
NcfV7jqOwP6l1t3t82sXiCZn3Y4bIuK0UvcgARgYklwAvFfq73XYQu2PFNE6Er5G
RSSZguuKBwnpW2xl/bMox8DxOh6UzbyClUR9AdvTC89MpF7pUeLzyfWH+cWF1MkB
U99V1Xjp7fyYs9L/O7z+MN2b8x2YVMbhn2bl/kfPloEMrbckF4Zo8xS7bO7dJdg+
`protect END_PROTECTED
