`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xhH2LFO4ebg2MRScqru0dQv/VEkOtRmCUwDYnfylHVyEDJUCb9XNusWLKlXTxTVE
B52xN/UU2wsEC3cOQDLCdZUG1hcFlOB1KcBupqGXEl+s2gxMzhx3+YVJHJc0r48Z
UT3Jn1JxsDXrf+yMeBRV7ZNww/tWfeqWKn9BqHU/01oRvnYeKpFTZa2fFLd4mrDz
W5b2NtrArapuUTuQrQgIkXaULg/H5bmWPHvzVMyBCGjnxoT5BAVy9jfEf8rj6rBX
ZgXqILrQN2RArbuwIOqe/8uBqSNd22/vc5i0pO69zyaB1MsPRf/gIXd4FqFycUdB
sK8+KdLNMVy3YH+pNLIkL9GO7EPoVrUxvHv/YEzXRc6laSsG/i6Fl7Jq/jyeD9qO
Hu5A6czK7aThmpAO2YG6l4IMzIhJWPqAvgpAJ6ckLbmQsrFJcG2WkbIfZ7d7/LCd
ylQD1mHUahjq6lZQWt+tRQ1qqs+qkdRa0G5wf6uStEdXOU/AJkonJArlBOgdtZDb
EQ22R+M3hjTG0P/1HKiTlGNKxE+untg6KqgFyEkYma8fQoSZHcv5jo1HzL0kQdtD
weKaIFQbWQ0P9Kb5MmF6xgo8fHyucT7TWZSM4SMSZIpzjdiCOXhqAZLsfbRAHsDX
RVZKjImgx5RwW3FswUY2ZW67Kir/eN8xYltsvpxhTn1tEiHlKUaFfAe1HN1rKsAZ
VbuuDlQVHX1FPaLu5E0Fy8YC6LrxVt7A06yktpvs7cSPuwedT183LCy+9A8ds3cY
q3Se1nvOQvkYbkbd4xdUAH1UZcZMW42t4pjoGXmOKDrC20bOgFpMHtt8PKRte2HF
msz/mqF2RSWM6PZoxYUNivlTzkfhm3N7SfWOCuXKc3qWvjiJTUPLwTv2v5EDSj/d
nuGPmRWrfjuunR5qi4Qncg1ZNB/3OadkY7ZNV6k9x0VBX+QqQ15ZbLARD0DDTZeC
cRMIwVNmQxrxa0/4y3vJSoHG/B9OhvZXGIrV+NUNjF6YUCDCuHv0lQIz6QRY5R0I
7kgoD8eHlCnQ08IZ4jiZPCXJfQPar0HpKkU65gWpkrmQdA6ctLAr8Y9TsaYNEQlP
lJA8LH9uOKQ2d2Wz/iF12vpWriuLCAOGVq18liA939OC2BRBj/kFpJE0B8suWGBL
nGUVAFs/hMUI5XWAOzfw/KKdaUk0MPkLNY6TPBESM4ASd8fkeJd814ueaj9WFUo0
nqVhKmxs30ltSX5YVsz0VAaggVMmICvS4sfTlQSo3FDI7JFul9LU8R2YLhr0nKU1
qfp9RT+G/8oSxm+jrk+FyZMYNWy3fHdqSrwLezBoeuImSIY6ZcQFDhjm1vAau9VN
5KUJGVb9CUNSYZ1nRpOOGA7SyiCv3XP6EZ7AAl+bluxYIHUeb56H17w2z/O9x7dC
Bzw/6Ihs46t+wv9EvwppBBgaA7NCea1YKFPSZTG8ndK1DGVGpJg1MVQE8h9ouDEf
5LC6Brc983dJR3MBDWudfnzAii9F8jKRBTRRmm5dHVhThM/RlIFX76ihLLClfbTs
VidhjarNwRfnR03ihCN7rpj80zyc9ymRf3z2uBRpHH3nyPp88mGrM7m5ZoTH5H4o
eyuAcRB/MnwGOF3ZcDqQ4bu6SmaKT5/JlSvQpzp8SQdGdIff1q0lLllK2jtqCPz3
pFi+TQrxoRLeptOzoypE5NNa/HCc/yvFj6zvr+iRNTNHZg1p6jcq88W7b5TUUtI0
BsPOgdhLntq6wNwGv8RsAQgBxC6t2J7LOUTXcW++3ff6uoEiAIpYxaBu9x3unMI/
Mo8T/Ezm+jvvN68djwf5x6uihlqMt1JD4qN+M4uqg0umUxt2RPu4UvAP/Xnp70L9
rNfa3IhklFRtCzQ4hLVS1swgYAmH2+mNYJqZiV5ucHtMhdeJWELQ4e32Q8DbhY1Y
eBKeqlStKkJTnxQc2mnLeUJ17tvRY65GVxA9mPS0HFSovgd4AtYRyC1m9XuV7NOq
`protect END_PROTECTED
