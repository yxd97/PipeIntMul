`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HfTNAtQZKOQqQNWTEHGJ6w1EOtxb7sFoVeaCEG6uRQ3QzS7rBb+EDcsKF7POqPx
YLiaz6PBJeyRHkafnUufhjXiNe50XeuSqDO6YjUVlLiDjN44+mC3e6rYTPTiXj8W
EJhs/EZLm6+Ejkz728uRKYqt8pSBBNGLi+9BKbzaknZAMtQxiWMTpwFr78uwqjS/
W1fWNm+OF3qvhAQOUTKTCUhIMISwG6coSVRJokYVraujFDkSnj5wyUpJDp8M58fI
F7kQAEfc6EWCG39MQzMOOwFFMcjgJsakTQOXwZ5FJuGgotSxPGXmoAfPQ1Dx+L+y
egYA7k3rp3wxtEFR2NWqeWF0yG5B1j/8FwIEwvfbwq15PMgoAHw5wofmwlMT5aCp
BfD7gPcWszL/XnAskElxTv3eCn6ULC0GLLyqewE0LKENq8Rd3nkZJrvSRjDJTo2t
3aFx5QV4VOlZKFCjqyszsDwmaqDUEbcwRm61A/EK5xJEDjmj+lpBbZI3Ik3rCKAm
J+4J6ROVSrMk77S6c1mJewiI7dnP/gsUQ59PM9EhSJTs4JBjKwjjNn41q0YlUdRP
`protect END_PROTECTED
