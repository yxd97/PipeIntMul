`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbSI/tc38BGKAUN172WGAsje9FYCt1Z5lj4e3AHlsNJjng626H8lgFD8IdAOljvc
zh08brB3CsLriy6+Ce7UMQOK50oonBVykH1+8+OJ/kzKHOk/HxrfVnJyUmLYDQ8r
jBIeAcI5GTu32Xypf4meYIb9ZiuPnEbmcD6ZJ0h6qSUGm4Nvi5Ic6TnYSjcGWCeK
TTo8HAqOdW9kUsSC32V6E6z2RJKgxeFGTN/upfpqCtUAoDtuEAEb0r5VCc8DcT0r
iz6Q4qj6MMEeWPK3Dx5EzNxpJccycDEYY9knrkOLr3Xc52vz4jpLQmDqUgG8kION
4q+dqlkmTUGKfbmSTiVGsTrq7Ec0C9m8d95mNsoTg5cz9BkBqS93+qWH6ZNF1fJQ
id+zWQ09x7BDAKcvZBdNYmprDVdi5tFQ0L1llnBtrqlecMlV7q/bYN5N/cx0FiJQ
5lkcsq7jieDrM9ngWE3NLfT5zGItiKYMCwzECVvDMjeZRm0U2ncvXcWnMkEOVzUs
ULmvJrj1jGwcrEQZAsXK9ukG9t3nkfi1uLNOIJn0LpaBaGEqC7SAWo0fTsPINjQK
jfYyr4f0R3WObrkV5P2FR0FQo6wEYt9M7Up989G+jhzCMoOQeWBBTUmDbCeIfaSZ
U3iZUjanVKOOBdcXSzHe2o1OJPDpE082w/mUOKHz4mlpHbBK1a/Wj2T4GiXPr+bA
jYKd+Q+CCAo9tsPNREw5K9Yx/VkWpZwi1czJ0GWFvzeM99/Ug9WsmmnEfYoNO2UH
JyggRbA8Pn1hVzTXjmeKee575wMZ70n4utY+OMC1167bDoadRRDbaYALkcNj6wvz
mu8jB44qBtKrzR8euCAVwy01wDoUMBvuluc7nlE9+zM+Z3Ymr9lsKFLMazZ0YBqX
OKSJiPA9BZENOcTCc+Qdh6oZjPQ67CLIm7jtg+r7VhdJnl3Nug4p3aWS5VNlmfPM
iX5Ff8uQ9zOp4AdUTZAVrNv+qNbHj1Jp3c+BHLRtocCKJUMcCQhqcONAQThAbedn
/q4/sTdZTTo4f1gzXNB7ZjMC427mqG9ELax12ejH1+adoWa0QAs8p8rMwWWvRhns
e+BeqkFmoMqYOjH0cDdMAI+cH/ydj5k43ZMI4NL0ZrJ0U3TOlvmOH5OKovVhr6fv
xSRsnGy88T465nYSN1yxton5Q9zQfPVkA4ifw+NoBUwnRnK7vjQeeMhAqudbKXXz
uxllZs0r+ieLkrL/7L8mcmrlOuaCMlgXUriZdlzbid37a40asXl0MIuXdexnXegg
KPsJT3BixcGcxIExQFoDAgpKqa27VkVW2VTpvq7qEjHZj65kieXf24zp+YQnLym6
O4TCnLV0eTNS/fiC3Gy312dJc3VAJ76SMOjwI3LJVi0TmRH4OJce3ieTLxwRBp4f
AV/aDiA0dLO1S2zLXfMb0u4iWUaFoOdrHflHK/5lG8JNAJm2V+j4CUPaOoh5gBid
UjVHIYp4oe3OkDQiWbZx6qNerBRWxb5fqUXuN5c5WqACW4GEGjW79gpFr3b9eGnb
KTzevKoFyfuk60Wda7/Q04afb1Qb4AGoi/mzWSC4odRsyVUuJjsp/UoxWQ5IP8HB
6U1beYsFJnACBU+5yHs3eMA7AXT10A83jsVQHDFxJ8wxQEvFDQJxm1JH+ipdRQdr
zIwh711FV46r/aIMxBjeltZ2mHTx8b1NCzTDD6eym785hxbedOVsCNcI/Vbysr/N
2ylxgcgKagpt86BBcBSJgZxVDzxae/L6kakOgAJKemj8nad9Rcat1wbu4O7O7iO4
fpXvhDsRAXAnpMlX2aHiDFC48eh4TEFGOr4yau7jt7Yr8XSOt3NLfsnKeCoxFGTO
qHzqDxru/KoslepTlzIp3qJV/nGBBAcixRjxoFdSNjO7I7c7/Q4Mbb/34tnbAGO1
ZOE8w/MXM+nXf8tjnX30mal0jDpC/KrUFX4m1U2JDX4fPXzqwKiODsZ245JEmqeC
UnbE5r8XG5x1tZuP3wTiHATt+hCid+KTa4AE6Gs43kgGSSV2zfMwSdGyZgcwue8Z
I3o+I6FmGMTUXx9dITZZ242iqX0uBKtTEOdAy+XTGjHJJYSn1A/KNX+CYeCiMB1Y
/+1rJD6tSQqx78jWNud5bgL0u/sctSLPM42AcipROJTCad7u0t7BNiKrCf09yduz
uDp71Xw9rn/NKEbNRSxaC26c/v3t+qqJLjHfshoqREa1XH5tluAenPhKhLN1YkDs
XN9KnPVtHCfmOOlT77We9KtJSCviHkXECyDbR4FYyb6K8CfzCXS6fm/lJkwFWqzj
cvVzxMjVXzwSzw0/S/oX/DljrTBkG/RmhBz+u0gjr+ywukXkeqFO1nBYfkpVBCnn
nBAn5Xzya8dNV89ErScYjZvHZBtSBfmV1H/T2X/w1j1SvZzPbcadVYUAjLfTmbnp
rJLnComVWV8Fatmf5K2ky60KlOo3RxqELM9RJUEA6atiYd6eyHAD624qqB9pOwYP
10uRs/SMY7JjdDPrWYVPbXX+A9rWZsZaxjXjah9J/fzPMYKiM36f/rwpHzfpXfAC
03fhGyO//erCJwAKM1rPKvmkb2Rzc+AJYyMGjpaL3m8D+5L7kbZjOwCFAdZKgCBD
44MikSKx6H46T/i703KSmXaJIviHWqKI73dCQHAj8AbQOKJWBuJYkUs5nVjMMJjU
RU5bI80pJW17rdo+i/Qgk/rs690vv73e6A3kBUoE3PNQGhXrazyB1cmOFSSYK1tD
TbiMtn1zsg53eIhCVWGhc4wAnIGL/bcq98smT4af9Io45mhAUIsi2A+BKdFOexMC
mG10ywvFWizB7Bn9HOdKMN544dvDz+mVznV36hWzCIIF6He34bjaCQosPRp8nNep
fSZgFzlg0GvukjmslwSaInZexskAtm4x1NzQyUXIo08Ln8q+pTIn2VOZGuiqJUxT
n1RvsCvj54J1qu90Ha/CUkGpEU3k2+9vTyvyNlPXHkTkxXzz/j4veLFibwhzVYEK
sCtdLXMMKR8xiwznOhToIOt1crZoTuFJ3q3hdg8jJDNW41A5GfBX7LiF7CSJFCsI
NNNRvpQBFtO44AXep3cQehFzoh2AynLLGpu1Yiw1oBxrj941ztZ6frPFrJE/v1Uh
IevYiGwNFgQXlfLEp0loJsP/q9hnap6T0uIL0izZ4/tbsbtu+mfZFCo1BT3sUdKa
68NWDzLfXSpVwgQF1FO0r4eygtgTSd+3UFZJVXE3YakDLV/2Slnlz1u6msxGBT0k
QkmW9rDcISpHSUe63yXxqQYHrTXBTqKBf7s9xUkTSf37eoRXgIVL3Y2ZYkyPbb4S
ok3Y5cMd2tPXDp8CE6MKGIpoJc3hAUimru5Lw0pN5DycpUxwhV4N+/PATfXiwjge
1qJDi6OSRz31i5RJYI8nhV/hgGQyHXtdSUbHh3ucM7T1riHCjYvtvkKBJyxAVrJg
pjo4WijYrWjdfB/DhuWoM8yYxELhbwpXtPXCXofzcrx5Vf3ZAcZRQ0VT9In8pvOu
y+KnuBNNmtLmIgETyMwtLbdvm0gF9W09Ue6ORRT6jOBSeSF2BSJT8xWD5lV4PDhw
gJCOPkG0aWAD4UKGodMLWL9IZ6j8BAnRGfeOQFwWyroISYDVDzLlJaVkn8igsKaN
fZIqHbue+fbCNNwh5EwxdHG6NDF5kmT5z44/vu5mERVvPiZHSi/I/Hv01B4xbpcO
drL+ADCOJX6Lia6yFXe05p77CZGB6js79Hqm7vnR+/K1pvpyvsIkVKC3SWur5kzA
T1aG5onhCpFWM8TcCwL7B222b2lpVb58FKRNntdS3z0ztZFNf+fKuzxwQH4T+WZn
WxcxfoLm8526iXZkFHNxiMWDTv5+OrW4SlsOKD998PkDkQnx+2ommzzSrBEJczui
coGEIE9+6rw1uEqnxeOOr3EGftcoLiykg0O/TQMQx+2DI5lhunfQSTjA67OxNb+D
LSEpBu6F6/QHrnwVTWDRcx3tXa6JZTH3BE2CPqzHRklcOzOufcsBGiXeRd0+eTyh
cdj7tE6BY8d4t567cz1IWE1tjw1IaX7M4RTI/BK584AvuQ/xUgMAm5Xp3Lbh5HQU
xyKgDNOWvemsgLuhqwIBgwK4WJQijrq87wBAPopTYxhzk5KmWPX1UDUnQ3VRUp4E
SUBiNCDfKs8i4rVAS34tpNSycc2Uily1pYI/mZrNyhNflw3p2aWe354tE8m5Te2r
UyGGXY/8c2mZtnH0EQK9zhokNaOW7nru8fmFwR4ozWfoZsp0qT1RApidlYN7ElFW
ilocWTPrue3e6QP8L3EiIS3B79ZQ/Kr1LpPGirEqVqXfiEumb3EyT4RnGkD6sA2g
UCwTMZJn9RM5SxExWszXXcF7/34lVwIdiv7IfNJaCr3OsvDcJifljSD6S4uVOBrm
BHjcl87Lqeex4x3zsKLSrA1Q2bbH2Bf71K9huPv+H+AQ4bNtC8477dywiBCdKAjZ
apdCfeWHABXPBCF30Fvoq8jMhJbJfGVrDAtnASfP3kYwYaj+9tfOe2u4TOekK83z
tyvo9x9SyB2hHpn3gspBRVmFVJLAOUZUsSUwVtQ4CUNhNGLm/B6MrGaz7aM9HtYf
DPcnefMprHM5CdiA3DBmMKskZZb4Sj89cWccvj5RbvoOHym9HWG7FpCXNM2yw8QC
k8L4Tf7b6diO8u4bMF9ieyRSGnNGlvuJwAzJljhbR6euwOhOqHVo6QYlhFLYM3Gv
EWdTzMjC7jcqEfwcxeaht4rrneAez+v4dM0XGYYkFQZGCTlePTRqXFgSh1/n1s5S
GG6tHlhcjMK7kxE6VHIvV6koxYw9iu+DQOEqUjV9b2XbzaBWEPNxuRwpVoR+87uU
7VqNFWoFdRo4nR5Cjuv+D3cQ7+SMieVjIdx+30ev7/UCeX39wD9azImR8gKmgf4j
rZ2fzMKixVGp6h1DHzw4BD4PRqGEkNTWu4Tpe657sIYXeyk5SbSRQl8EJtJRWzAA
HbaY3fNsU+o19DQfCv+Mr5cm3qRCiBQVh3yg4eHDt7qs/mip3cAB9cJxKSVH9/PR
+ZEiqZEor9ehZ8mlnhcFW4O7ZWmdAUpNcoFtMXtiZqV1ouGbSbP1sOrp8LBDcMpC
1Ppak/DRiZdg61swluwnPaEaXuKuxkavGxYA0eF5fgVdlqmq4ow8YaCL4tdSczaq
yWyxE4q7umSbHrMIb8QkOQQ32FQbipfYSlkaDaJ24IdrGyyA9tpm6TsbEueX3sCh
fEqpbCRLpAT1s+3t+grCBDWOWlkd5xSL9/++eQGietQ+zO5upJIxmLQZrkB+m0uh
+G9cX3ZsBCwppyQ9b6AHL9mvGHSXJlmpfaDXT+RAa5Mpq94v4RocPLx+4BbTRcoU
NH8MgxqFZc/cjv4ntdX+vvhh7rycOf/kome8Tazk4q/03dGj7eJ/g4M7Q7eyqQKQ
gYwt71pvpHaQ/WLn7E5Pe7ox1NcPofnXRmiL1JgvawZCl9YithUnEvplUms0OuC7
RGFxco31J/DMqWqxY7TCaIgEES5l5mCak4djvpAAJMtkEs+tcI4jhzleFTPjwqTD
pUa5xiaYRjJ661oayzYAABIPSrVCnBTibXFKbLtHdjWs0skat6+8Bo21sIjt3uwb
v+e+0WmAvyWMI8aneIKRlTuMGSMGkxozeTQ01Bpo1LhkAsZyQlxjNyzMFtO8zbRP
8VSK4pPfPaekmjQRCQJ4ZjNKUmVawMqyTqkNRGcjzBOFTJhuHXii5pkoUrWNcq3v
NNpHKYBIXMTo+xa5njb2YH3erI6AEHNunnYft/sVb/ck9VULww67ubn5KsNjibdV
8RajivZA3/PW0VJN42Ni+tmVgeHONzsXrZBnIlM3YO4sa+krFQHbjW7K2RpeZ5SW
nqUs5WIPg/nswsMmoW+6YWD7hMTq5IVcI3DI9suUZdk9QdMl4q6ysynlxc+cay5t
TGoFcq4q4mXw++Jy8K7J8LGis462VBD3NmFMdMfWEaB1CPjYGYBM/b/9/fIZsNbT
trgwg/5MB6/1GEdX1Gwmafc1rh3wnCm9vQbyF58Pwm5NVVEhlmqN9cKWi3eciSC1
nVhe9Q3AM0zUyyP8zKA3HkHyDCEnlgsOOf28DBDNNaQRWHMIzE9aNB04iHTsVk5e
leilgedfzPapWiPNU5wawNVmAqZJ4mho9T9Y7xigayXSzNKdpPUAXjXBYXV8xBLB
Ff2OCTmSIklHCU28PJg8Y2+oi+KR0dzCixqlGuFW4C/poOLAvNATs9WoYkdTgKXL
fNSNl1E0nb+dpoMdjfpAfQjYGPk0Mdj5YOW2VVYFH4Q6wUEP+B4YPHU7al2T3Gvn
HArhdIwzEShlNW2/1dCvMaoGqzWme3+oIC3AvsV1FkySo5bqb4mXY9QBdVC9nZ+o
jJl9uxiHcn+N4mf66igUC1P3FRHPWL7kEA9JroN7KmXcqD4TfMlz95/LkwS2Yxl1
KBPGq+xqI7Yad4z4ZJQ3MaSFpkZogn8U2HlFkidD1GagqwOOIcBreZmAG65zRLjl
EyqQ37Il1Yn4Va7+AJVLY1veKZoIeiVXDpN7af88LfL3kfVhITpDT+dmktNON34H
oy8wClDD8+Z6QyWQ23cRUqZ+w3dlmj82qGd11kBZggw33eCTp/0cN06JDZxYTEPP
2W/NKlYCt0SnI3IIVMvoLY8hz3kJuQRF2rXnEZPiIt47NKMzCDwGF0PPm3JXIGG7
r8YCi8+Ptxgl3NdMluA0jDY43D9Rg74e3GA8yQehsPFdfc5BAI5Z/JSMFnjJwsRf
rB1VgyUWHrEhzObmK0LYFzuhtl+uyyMgenTzLdU751JNDM8OxQ8cKTMQnv+LW2Ia
26qeK8/tWGUb0V9HJmPFlG1CXq7x6otDhTnXvaXBkstjG/1TeNZGJ+9dEx32nrT1
oJNwQxaE+X8fAzZ6Y2U83+0iTEW4GFDg2dIeebK/f3GpxMOszTydERxu53zv2Oe2
VQ6xpAOTh4lzXqIr9j8e+vyDBMxiVODWpIlTrLmTcW/DANWMFWldX1AoF9NRiDmQ
tPhx+pz8RUZjTo7sWfdTCsEHLNQ1dB/r7ZPgFr9Tt0/o73MFfB0UFV2pcilcjHT3
bTlUcn6qvZT3u6n6XAnOdVDeG+Z8GKBZidCbLw2CAWQCGMa/30BhW2cX1S+6e+xY
6rBlODgKOguW4Z61zr4/UbVqwH4S0yIJFvkA/dVW6oRn77Znf377ksgynHWrGYRy
GTMmsUc380mb7OagENIxrRg8IBy/dpz+XaPStOVuNlIE+t171XRR0jl2hZZW3LUb
mJ9RVL14itKT3Xhfeg+bchv7H+nFud8d75wlPAEaJsXSZbsbJS+TjMMxNHyJgMAh
mcp/TFE769K0MQSyEABAZqE37kL7eo2ga9eaZvr2wlj5o2pWbNaFCfkSK76okB7j
nmGXlIRQ1+TzfqdyBYl9VgAL31fjzAfRPvMOlvvtBaXndy2kIJ807Vnel55Jz7ur
phtEK7Qm7dXf/lAme+wUh/6BtH9jTAvoxxF7RXf6A0cTAN8Ua0vBnYfyMc0IUNKj
s3lnUQrhVx0dgz4bxCQcDv8sEBHZA7l1VZ6walkPs7HwTryxBEman98NpIPE5b4V
9ld9j6uS9JqkiYG3BcTRlnPOn4ofUiGzlr4DhPRlOM3fygarTGfmr+t4/isp2fMM
z81wKMzrAwAVCSfKlHTu9GaX2/mJdASj1Ex4e/nL/s0GCzyxVzFthFnNBUvAONZm
G9HkuxwF+yxyow/TpF7BafQhVSFU4BCEsXqHkWeKi+lJDpwXxyWwea+NxZcNlnNF
wL/vNM5lrX+3sxPga3gbBnqVTlNJHoujAP2sVKRkIIoH3zoG2OaQ49HQp29UKSno
7he5azHXiYN07dhI+C5eCJj9oghdA135RbgCHqb0vnbOXqfvC02FBvTiRH7rnH/a
sgvCq/2C+p9Rso7hFX2igeXjAoEUDeOJxcRNZUC/FneGSFOYkFdlPIRMRl8nQCag
aYsUJzQCpL4qhaVtTiUaTrpcLcPK+Su9UEsnqtocmhCFuyUWU8+V8ilrJE5kfwFP
U84832Y4Fo15mZyVuNqHUpZ1O/3lM7nxIXnDOa9N4U6x4TDqu0Vgy7YXt/WTMomp
IjaziA8Hl/ELOVDinV1ieGl76u9dEs/AsGc8fZE07ul+l75GmzE+Uqberhn/RbGK
6E5uqNzwNLEc14LAQIHEH0E02RqeJmIjm6hd95Ta2r5UuptSpEDZ6lnYBtY+ITms
JUfdFp5xqIreuHoAd21i9PgtpcKCzCCWhjlgqTmTWUMsBd3yEc8Hr7uUDOXQE/Ss
T/sEXYHpCW89g63P/kW7/XZt+6fZhrsjXfILL2GAOYd/rZFsnGczRMXDRllE2n/z
janjySlvzFkNhY2MkHU7n+NZYjHyvsglondIfiD+pmwkaVYz7kfur9C1JFesdPX+
hQRznJp1bVn2mSA0A1sRJ0pdtU6vNnF3LbFXoflUt+2zX6Wet0dCEVjCq9Mf+vF7
THP0FW6HdunKQXcBPs+UWTYWLuSxm3GoCeA+qo9xZ73q1bRAf7nEewC2RVxQN9qv
KpQ9lEg2vWcLKF19cgpPPk68oROGkdLwKoJSoIGzfuXzN4pKUwac7lvX/V2v9EGE
haVvqc6v8xsUBYj965/I23Q0WVc1lflczCKrwltnadUGgWU3UlCPoihI3EJo/x1/
YLTrm//u70XW+rqoXmD2tXitxZHKpzmxPeEJJvDcYurLI0dNP1a0xAugSCH6MPbX
c8LXDC9H65Xk94THVtEpeZ7g5NZWn4C4oPBqRNROnoBLxuOmzGqcuIKwqNDaD8XU
UNVUkr2kel750RH2aJAlG9r+Y3uF/iRv/22HsayrFiWjksoLOOsLDpO+9mYpj/MZ
plYOE+mhQt9PAqxyoErRfncd3fWBZtPixlUj5PaIZ3QV5yVt0//qMs7TupoLf7rz
gDsXn4sr30tKU499O7b6ZHshMaBP6gmdSVxoygRxGUfjye+h+yATYCH1p7aoZAd8
+9VyMqtK6zfKBorZ9mS1KtJdOoytIEJMS3nWBzTyYroXb9QVoSNLBBIuMIyi4wTY
ZioC/tGb8HCP8KcpxEnEXp6f86Cb7VmbGWc+WkZ1qG86Ea5AJwXEWZHHbkSAq9RA
x75/AbigIz6TDFYG/DrUOm8jDUhoG8eZ5avGnW0d8V7Lsk7pUgJ6YN+0IT2vjPtM
68DZJ8rvdl4BrEgHGHY3Te4WMD6haiF8M0YGyQepknzO3r5lyPUZniW7Ky1ro0FZ
VEWOmkNi25bj8JHlmEZwYhzSb6HgLGcRemyVZ4fiC9zTkhX4wlb6s/F7RnI22NM/
0KYd3oBtyt/lMVRooVAOYHXSVzrRsf6jyPGuutdgSDcr1GVcXENplPAuViGEbD/M
Zc6+0Ln236K8Dw5CAdP9FaezQGzZZLLJ3hw2ISknDinVOkaLCTYyTa2BhAcsJMiq
pV19QouAJz1fQRMcdtMHRj8uLJWxroJPz5pUala/jpeUE8bXSNxpSAipbQ7NtHOT
KLQkpb/fJPqlU6hfp00YsYDME584C1+otfvnwYBsTxq0px/oSFvf7q1lmjY2nxHF
tafgGSNCw7ronaTw0vPfoS86nXpoNShCS+ivVHEtARpkLM8XmYpQuYlo/iq3lbhJ
BNjyiiH5Ipv35RDwvnP7ZXKZfYqeU68PU8Uyo44W0piifWHeEyrrV69JfseFBtUQ
66JN3VvrWCogQbXz3+tfut+qOp86619pok8oZHh8j3KE9s1Sz+ab4W8IxYr5BXIS
khzdBnbzu3kJuxLOPPe0E8UBgBYQZjwdTBUHjBi5mw7XhvASIztCTlanOU4WgIVy
3xs9sNM4wS1zGesm84Nnd6wshW1LbZvFhBN5Gee6yXgBXTENTV83yQ2agootEfUl
Z1F50JXqOXiI7JKeyQy+6vVwfg0GJ/kj/w3lhV/bGG/GZ5YrnJ8+MH5eXwvFz28T
AqsN2orKZ+VW4l3QP4+SYgYIphkT3Be7aljKhL/BlF3xwqYr7yVbK8z6CBTm6CQ2
F1EWCmOfRigM0NZbtNDAwqQola8g9Nf/40QHHXu6j38+pNsRcTG9KChLSePDHDFT
rtoJW9zHXfyLayab/nncYMqXO8CqzL4zZ3eql42zJ1UhhlFPxblxWVmmlQl2UhrM
sXpoqcDgTfbanEgOHVBoU+UBE5zjR7xKlM4MJZly3mvQSDFR+cZgiVQUKgcWNmMq
Q15n4e44Mn9xfI2dUlsdVDAeMqaNUoZ1fwClaj+sRkd7Kx56xdbIWYKsK5dI0cnk
Lm70vKwbIKrie4BqE+Q9f/OzTD09rmyKQf9T2myvSspMqnShzYC1Qj8rJ2ah9mZA
+QqwNKJmJXwx4SKPf7DWhno7PNnBNZxB49fm9tHrNKE5+vPQ3usWFhlvOLwRn7qK
13x4tnnHH8kmksUQ294DArHMqVauI6uJisbai+3S00l92g77Y8fODdLTNsEw5M/H
AHcKYQXEZQ+gIl13exM1RKtVePn4Q5rhN5Rv5ySrr+3iPtPueS0qrCO5DdQVMjQ7
OhE1W2ry7q4iutkHvacBUH/pRtmo1nqZuFAlp5Huo6codQY2pEnuY33xs5VyEdgw
nfff/M5NJgZtMkXErsgcWsw1SpB5UQegfpEtN0Ufh/i+k69Xrc2xPMuJ+QaeADG7
ezmhw5CVEcOlT49fThE7YZxwo/8si9SicrMXAOHpzP1Lgz4sK5qP+OcH6Uc08qhd
l1xGA7/Ds0jOdWNVNkePtfkcQynHFLPVsuIk0CCs7QL2BKhc6Vbz1dAv7sFT5Cau
ECf33GKdfXx87fG3gE6XmKTxVsZm+0CFBVDRk5ftmjlLxEbdeTrharlG0jkBTWmh
jFT5PCXTqVe3KE1demOzZMj7NvER4Zol6ATmSzZ9NsNMhfaFvwUZqmPOTr6XkQ3B
vbSfJLnSyZiD7lN60V2YzZbdt8SrXUxcXk+5ZBEspu9OfG2kDPUYAynqVM2NCU9L
GAUbNoEx9xVmCYX1Oe7lVkS7bxjjnHtx/6IBwmImtEXeIJUqiCkoP+B9UKjYIgQI
ZOebd5xjqlrVGPQZ1yZPEvFMHMNWGuWhDWE+SlRJzCoPo9YNFPYZ/SNXgg1kQ9W1
5Zs/XWm6qBpH+9CZlOsmJqgitXBUILy9i/0P428sXYf5lBGlSNKqRAk8svE2C4wt
3aVmafmqCvodpTqSxDYCeOg3OUsL0ZbcAPYWQ9OkrU3b/Y2tfb4g4BDo0VG55tQG
C1dCJEK0lSf50WXaeUpVABGTrpprdXoUqN8af5086zTcRSnm7DeJGB67DITKdPw7
HOPe1e1TSsjn+sMTAx9d77UCz4XOlCePfeAtu2FOZjNgTeEXt8nyKPjGpBC9mOpb
lUiRVVNv6PwX+vKpS/a4AWXyHqUEQ1NpGR2a/1ypiH0k4nUqXrfWnnow56tbA+Qk
lB/Tr6QLbHW6AihsFpMnjb+1Em7oDZkbRsxXUoKTNQUZZTmzpQ166TNlfpi5AlIy
1JciXdc9JTHHXWfx4tIFoxaZ4AHueWyvaykzPrnX5xu7KZxLmAlDK0VHArBfYRj9
eDl2QDsU5o1SbONLKOYyWjtoD470gqwycaXrxytqKYfSdR20ZAGQAXIPw0lLIImH
BY22oXJ3/IrrE6Ctipc60MKCuFyT4XIk3vyw9H80hA7m545pjLwD6dEPydI+tb2B
lCaLL1LqJyPB38prDb2fFJ6tpLAnK7pZFnGZwofJWSqcm3ZMVK6yB1gAwz36bWzw
EX6Fl30UKWb2NAjNcRKdd4HvZqzmm9fIxP6RMpdfVpg0J2O7TMJ6hzPiwQtO3H1a
OcNkLtpwLmWL8Tr+aqnYsrDI9wDiGPCkSBHbsWcG2AjhfpI7rADiPH6CoiSKdre9
eyS5ojiKx2FwyLPctLCpL99GCWhHJIMeC0/6DypYYc4nayilHU9qvgEdyj8gx1xE
lLUl6zyfNwbi7YQm4HL45x7LaOeXdd8pykN90JJxgt/bSa3M+iKn7OGa9U/oIZpv
8shpMZaU2/3i2a/s1SSC6bii1NT6Y//Id5ni8oBhPdGMVE16L7UAK9RfWmlI7Pvf
CsysiDWU45NPaWx9uRD+GHr4bYgBLUlWc1XR6tZhIdj5yxh1CKou6FIuGD2WP4xR
7fkt0VhIGf9X4GKbmIsoh/wTnQgDgpjzvNbRwTm2PUqjK/dseLOrgleWkm+0V/YD
QCEGHhvIZiwCSe/xUmSt5WNLetQHER4/ldQbsdlkI+6o2MMXYVPgZ6m5McZfNTjz
RQHQMNUU3Aa9W9aufuGskc9HJJHVIe34LI/+sz8aSptDurbmnlsLAvLlJfk2qfIp
iTggCeyucPb3Fi5yE2YVDVUK8s79MSg1hvBZwPWQ78/ntp07EWRmZYbLjMp6tFtc
6OyXVyLibFDz8JLU5R21PuZLATgFOcFv6ugPa4nf5IBQ4s/FM5jOhxP4gPtYxsfz
VwpSUqeV/0hjcsN4Phbaeak/k5Pl2gM6XZwdolDxuK7anXx/s6ULCaNkP+c5zQ8h
8VMt20fIiGOBwJTJBdLwMvuZ2s5G8uFb9Pt57N1PAriGd/tMGA+5SNtLkM0JTjkE
+l8ExXuyExJVLz8e8itOABIneBhZ9fYE0/f7ZWGEkELRC6bCT1FK1mrU1kr6gCiY
v9+cyknB2oNyuaQPCIld1N+H7SDy4duS3zCgnbhYO36YHDJM/udeYXoGW4MEBL95
+ZJFAdLkAxe9K02gnifHb5Vwhyt3KSn+IFB8tUgxYR2cgthzPTt/OMlrOIb85+ei
nEC8SauqqDO4BsOu0rn5UsBIMUeZCLGoUgTWDVQw2oKs32lN59nttTvHCY9YbHz9
YH7U+NJkNA3sn6ePWUQWs6SC+rw8FZTp1KfX8r9KiMgqtVp6smVB0MDqNBiTho4g
VRrAToFQ21xm3lljBgOwpH2wXHreTNZ4XsLKRhceTnsTanlhtm7pdBkZFgRUbc6U
w3Qu9Vuem7J1iNaki5LUfij4RiihggZEIEMB15KYV6HXq8t68VOTt++xKSfSu6Tn
b9O/NICvH2IdwNNXqHQs5tUgM9W3dFLzyO1G4g7tcSkE7Py21ZE1XVe8IHLej98p
o5Glx3peeh0772DqPFhyD0iAGulI1LXQQdh9q7SaJ+HNCkSOfNIswzXGF5XHPPFc
fyUK8kYp5x/iY+gZoKX0W3laUKOd4LvTiSAN3yIalGne2VMCK0713q916yKf3BxP
/y5Hh5tlDz08EChiSnnv0c5POBxOLEopegkQ/ObNxLYK3uVUyoIRjfxy3pZBuyvr
H+kqAJWhr9T9L4OREwFwfNcS9gx/Fo1f9zJngEC6wsoNhSchCzWpJaYkmZWI0PfF
sPagzvXfwKUKsXGG0X1xF7WQDD5XdlVt5VDW/eIFnglmqDtcRVhYASutfjg8Y+JI
CDgXVNHY8OCwZrxPJ3K6Tl1rBL/9BoujYvUztiutkNpFejLCApZjy/Tad6ly7M7T
sDucT8io6qX/UQWe4SVZOeMdNWkEXXpuCm10uuNjhY/7gi67LJ5AKqqnonlMG1PY
X0IJtC8IF6BiuHbDEdq4DrtIKj/q7wKn2qxwmJ25WcjnaDC4qsRZjpQqYVwtrUv9
j11o7n7ZxXtPWEbXH5Td1JCAOWoKAurAdTfZ2L0NOQW8DVY3IUJVWD5XLlyxDr/9
8eLZFif1QXHreCbTTFN84MLeAONilZBN/RctEo4s82ar3UQTlmeHsJ9Dhy0cRBdI
oK3mJv/8w8KmHDAm27cwbyZ1bkzKXJ2wbSUP7ipdab2heWxjbxJNd6emcAlzx33d
8qkwAYJhkzpzMxlR5Fxyd/zJIABnAo3/AzQwIY/u1dVUgM5JqErGaZVkeGrcbqR7
eUGjhSCntd0iRV1xqedrNGi1XHXXtYKU7PeHI5D/ZcNK0EWeTE9Qbor6ET3C81t/
+NnCQYtCe0gVMA4swoZ51uzRusQ636TUMLYF0zZUjBvmH2TrU2BWYPmzOGY7Xyop
LWOuL3FKNShjX2pFa1tJ6XFUCd5bWnoEJJ3+bbForfpKLn3/Iu6bL+ZVx2nwBpLT
IpqCtGzPe4zUiE+pO+7F3RD5yVCcnCYOtkhKDgdLNdzmRno3IhR4PzbdKOyF0+Dc
nbz69zLnrgGDAg9SVdrKdESZYpS43Ch6n7d12U3ws4PTo8MYFqSQRUugjFIQpgX9
bCPXKlmji8vwMjdk7cVoJzRPF9JgMT2FXX72bhedG0sJQY4jfhd4kxdNOXy8tVn3
Ef9GtNk3LFBcGWpPy+WQiPfaV8XZ9PX5ow8JGRP3YUT1HfZ7YkEdG/qV8asvjGC8
bghuYzRemttRK0r3LGHx6HaTBN6v+uEXQ5UnV1puaWSecIpz8agp/pzGIvmWfrlY
Qp5qA4s7KQ8s4GZ3VNrfDeDusIuryHXktzmUJPBafgHDF9K6z4LwYk9w5NC9+hDi
p/KWUKGkyNknYWM4byOJRq2BoRCNILSpz9he0Q5qDbrNC7xbhSUl9sGxRYYFw6n/
IWvij680zIIT/C/SM8qjMXreXuAkmGW5D+m/1t/ExKMK1nWGQY3iZfJNZiQl8+JR
Z+Ph11BEBMC0u8LHBR6CsRTFY79fwO5fliIxMTXUWG5JrrbUr45wEjJcu1Wfq+qN
RGCjal742o4go+yioSdtNy5trIqiT2Yk/GPPggl6VA5xJc6iZ/0K/g+0AgL8EjEi
MWL3ZNTf5GuQ2UNWnm5W8Fh2v2LHETPk96fOZv+v2Qij+iHUGjvkKuSTrxxjGWU/
27WxAaV2JSjGRUuopcfRVgc5JwPRHVR+0DVvOshNXOx+ITuj1q/dIWF0LYlgaQ4P
WkimPvj2J9g8L2YpYpRcz65O/UyapUMFRLWkJB0HJGU/Qtad+10KFfhyuuCJLP/1
+Dg8VGRkmiqe4XxfRhf7m4fltcXvYsOJ6TDL3L11NCzu4Nonx+tFJ9jQ6/bK87tI
4P8TqI8yYwh4mvKlpnPZW4wFpChgAxHxvpY2M3xUKSj3tyT/VpFxAOpdyBRI8bhJ
ZBeVTBdsjvtCXEV+i3zZzX78t9+NoUHBc1IuuClITqrG5MVrNkBTbdw8m/gM6KOL
cHm90SMguDV/T+5HuK/mO7h4Y473ACI8+LS/n6gKbjNsRdclVL0z9ne+xQt1YLMp
dwoQ8bMDG+uPQSLFuZHP0v20+JfeUdrkIRGdWxlU4Pc1u2dwCsl5OxoILktrHvs8
MCwf8WQcXHzgAor+spAyMi35GZnGmjg1YiVdDh6yB+C9NGDH9j2dlNM87bRaeDqg
OcaRRMXRcvandl55Vwp5z7q+4N39vdTeUq7IbDzlRLyzdIZgPHqeMlTPjzd1a1gB
N8Fpk+ggfTDTcyfrJ/bbFZD6vamGtlsqf3hARfHZRzBQQjotbC9nCZLuKwgeovfp
YUKu5OIcbrnT8VsyBSTsIRE9WB652YpBOupT2p1KgHoM8I71nQP0hQEHu0/k9KoF
VlbfEQBRzaa3LsODBC/UKI2epN+qkRSAgW+C1SmHuv6zpnqWTAQWDNmW+/UpbSXu
+lqWzbP5H4W1AOrOeDMI5eb7JKgYtXy6OZKqn4Fqg2SS/ZN/GuoGrvfE5pfK0nTw
bI+JgUrkbn6GNecSVaYXECkXRUniKpHrfXiEaDm0UxtFF52CXdIEah8ITkKb+Qr2
z7AxCPGmVEcoXdyIMmrbhqPUfEZp467TPC0/cNUkNEUlGTjS6mtpLFSBYhs2a1Bv
UhWxvOUAgIxCDasUUyzaHY3KGjDMdNRfZtRkFFiPrritDyl8jjXqK4c6Zdig6meN
8/eovlTNfNEOChRgl5f7R2USIGOERNnQIxmH6y/4DFTeN0ZhDTa8Z4B9gmT+lHI6
9TbHVxboDKR+2HswQgBjDCtTc68xQ/Nx6w8jeOOpEsNgUYl0BHWHljF1V8tOCur9
FwfZQARQ3SRIsHieYN/TLzevUqi40/N8Qu3jhvTnxKFhUCNDwKBd7FogQPIcOgss
kwhhXoa2J4zgjmMY9vT3hjvqL1HJf0JkhBZV13PYN7YMaZjXeUfHwIWQI3J67Oo+
sOBKW+TH9I9Z7JUE5dx/xrH4x1cJlyfTB9cMDHkNBw/N0A6JvN+oTAV9s3dQitY5
/5iNdcuO87mChtz42k5cfFBSIzloi78TSuHMrD8kdPh3GPA/IKfRk7g1ok4a/lLF
0HbU7Kv0Synwh1er8YHc2H1OmOcLwodzAjuwWfbRjm0FR0T02fCVIQx+oS6jOahj
ps8S+aAqHTC113r5u3H0NIUhZsHNFfhJOWyl5UifzkEs4Y8KXqaafDZZdMBQFAWy
g0F4QnutwklraiuPTZSrvfgMcD2dScOvh4aYXxhYDq5eIAZRT2SnLJjR6sUPiXuQ
HPAhmxTRoKvuUDc3bUFAqqBnIR2WtOwsLfPrxMbFBrS7U1AYjP7nSMCiiCZkuiWj
QFB6wifiCE+cJGE8nGvkYu5XweUz9OQWyKJiY2VdQmie7qoRgzEik0zsvD88LdnR
nlXFHMhZ6WDurd7U2Ictx5IySE/cP5TuYH6dqxQtnoRWgHyGUik07EYx/GtA9h/x
LuTyr0w9qnR7QvSlBkhs5ObTqlfZPs/mppx79WmR50CCQ2CpHl3tBWOVrZpcYWh9
cMxRomd7dwJOS3w+vWzfPZwiRZATaIiLnQPW7MbQNKx0xfF5Oyz4CKrlG5aCy82i
XaNBp+RbhSUl5i8loNhTc+qv9CuKin10TwF1CFv+RTR1Ywaa5D84xD8QbJK8fGSK
HB3YD4A88sh5nZFw77AMcSdKOEzJO5SAx2PG9CaCpRB+xp6Ky4MmJqhDEFjs/pb3
ovGA1aZeX5ayrK9tfbD7A0jW4QdJ2OLT85dbWMiJRfr2aOmBDmoOsxHqPDVvTjmh
8nrx7H7ZUuWD8DTZgw9/+mAJFtdiALY80NYWvzqLE1dz3lhS47sFhfljE3Fe3pTa
46AVtSnpjHouGbr1SkKikgsJFpryeucUxV9EIZHZs7uab80kj3aGWzPL6ofZXoym
d5caZtvWY54WWy05hJb/cGuSe4J5dbDLs/rLA8Hi8iKgCSscEBUqejiRcVyvT/eH
TqjbT6WiukkeZaPkml+fshIIu80wv4dLGLcEyYbStnsjAhGEOtLUBgSeSPLo2Hzr
28tT0KhgiY380o1loQemIg5yIeheCcLN8An0MkNwjKgm8EvanrjYs5lny6Z5BCM0
FS+wQ3z6n6hp+zLf2bttV+bzaK16H+D6/pFaG5LRhNBPIil0psrpIipKUQYhnJDW
vxYO5DVE/rQSiDygUJXVb+tMDS855XGwaurIEJxiSpo1Z8LEg5VScdxOBUE/S+g0
60236zsZY+zO4J+UeLaSP3kLKQtojFCNGj6+gQIoLYPx7uE+XL/c5HIdnEIa5D9K
dA+hbRHQau0UZeJHyYqc66AnrkYJ8xrBou6l516Y1FYvQZBLuajAp/c9V+q1hHCx
wXhh8zVYJR5mYxT5NJ8wK2PHkmRVmGjBuvvjTJdFQ6/UNYTERgiqONuIqwMR9MKN
sNoFngR4lR+KZ9CJLIg1ZCy4xI/JOnNgwCnaj7OXOpRjQjJK7cCGZjAMWQIz50Ij
P1v9uE93AUws5Tj6Air3RBbtDKH34zvA94sPtlUY6A6VeUgmEOvEGebYQ4jQ2iS+
zkA4WQBvz59Sf9bqFZEgJcPM+ieIg1I3fAgW9HJMrT/wiBEWLIu6Moy4hsSecott
W9lEG20/Q7C12QY8Hrj3i0BeDP5oBwi9M1Gi9jdQ0hfdn0iA8dwphNKZPMQf2qny
9TA0Es1U6VAubCHKYGphlqvW9JzxtFBhn4OOtSxvxOp1miKVAlKfk+ULsiC3zC0E
nWj84xG9icoPY76eyZFLjh7dk3EbLYmS/UJB04X+pAvEZT+BsL9nBWdSS96809kb
l7ZvNzCW0fGwHOJ93jglVpl8m9Yt3n2w/1hZPVGfWGLUGO+QM2SX6Y57jmn1XNoc
71/ubDQzV4EnjAYNh50uZyt1dpOwaeN4L4AssaRYiW9nt6WcH1VMD78VgPRAUScq
0dg36m9ngt3KaZqkNUQv+H0skA6uGrpVfMAHV0io6Vv4In3yVpnK7Or9w9vbFmWr
cHQo4H+D+O1Kt1KtSsb2JIc1nVWSm8p5IkKbF0UqTLVOQZVJvq1laYRHrdbXaJCO
J0AJmZzbEKT7cuU7TdaNmw+eCxN3Z3QguosDIjtnntaEfVNr/9FOetPcASqOATK5
0lSn4U3ZxTVWCfenTulS+kSgwDoJBDfv4LHRQHiVOEe58wFpBeHten3dAz+NiSMh
72FjasUDdTgYBdvpB262BcGgaATPMyQjD+wdKcdPaXONawh52QjTZbti3DNqA8lm
TdQMSwM4i60454yAOcnLSuxAIFWZ6/xHriD/SUtkW+0dQ5ma0D9iS1Hr8h7ojsJ0
/JojvIABx3JAZNmlCrRj5KJ27PJ6oF9bUS/cYPqjvA/jEggWScS9MX6Iw385Alxa
juNMc20bnO7QIss+AhFYcTMJff1Bdq3sWNLTxeL5f8FaEdFobDoMC4SAMzKbJEP7
Z3Djtp3BEY5haoKQ00runcuVVTAJCBu0uZz4f9a+jo+KTPMBzxqZflxvXM+zTmLV
J+U024hjdXse0YR+lNpwAemWkE+aFHMjGDlaAshdi+ya/yuAqIu1X8xAIiQoI6tQ
kuutyQREm8X70ckoevVryKqnuqqDW3KzgJ8pp3f2GrtTiG2UNOGAh8UQCKqdhylr
Ic7vLZ/EamXoFiFDozhYg21IaHSsv8b0C78Cq6Sh0gSQwUhklguGB7W2PWTDxltD
yYdWyAqyN0MUmIUrfGwAzSQ7IKR61371/Miu2rQLMdzZIhejhucINqGagH02f/BO
5SSvkNMRzaaN7MKTZWlltVwYe5D/MSRkkuMz8T3iFGF8wZM8XPcN2lW0TP4TwV8K
Yym19dRHOfHLoJZsW9xyGFly8+Qvus84uoE6QIhIpQEeySMBwAshOSsySWkxZE7C
v8Sm6CPKlbLqPmKvgN9LX/SmK/2IaxCUYuRrJ1/LnTxAZpugvuBuphbT+WGgnPWz
mqTAz3m5hdqHouDQDEEEu0t7gfsRldfajhPocDY+ZGCtHleybUQK0WMkXYB+39SQ
AWBc2zkT3QWKC+WicBFj2N6lEhZuSIx6Q6uF4aqdYeJXvmqi2COy5NSl1e4WV2+i
Qyq75c+ds7uDxzocwibplztTb8aMVzh2HpgDARKhcpyjybS1K+2JzIjvFAcDAhJG
u0K22sSq+IdKzIZajY0QMzMwe679ETM9nqBged2NtdSx0GTRjX3LYdbcsdTDET3f
w0CR1Yr12LFJ2SE7p6sQtIClt96hgBhevu2yRFDZaztH9I/DSJbRwBVwltfHyetN
Xaw3xivsE7SkgweLq2jLNa+kpLertoLIo3XQg2FyApTNFqD7OsM9sraqD4Eh+mvb
VgF8SNQ6TnK0Y99uGCa9oO8WlNRGlGhk1Yp8a2MDCmTMwPt52EuE7cTpNb6twuQP
LVJNB+I7729LVz0D7PEGGA6vmVnCCKYwxkPNUnW0caHKpmIfT0H6u09csFpv7wqR
KoiFrVNoo+Ybn4xrE3UYltUZrEDT5IFI2svCC0D1RikNy1cPUBSCxTGqlvypwDqo
KkTN7nDhhamB3dk5wiAngdj16SlgGKGD5fPJA2iypniU/NifkOey/e2Jvv6lq5nR
nP01+69BEyITWrjh9K0ktb3jxrZ1WVI5nfiJlHIPaAgYYDw0tfxQcZ6uBG7c0J/+
co3rfvRawRtgDZefV8Ijj7Bgym5/Bu4JeY+8H9O7FlRWfQOjKt/G46GL4w8JpmJW
FS2wBkatfQaYlxX6+lEJRzuShpN4rPmXZFSLhA3FH6GWDiJi9b2FQNFfEjAgKJvI
okdVGJtF3DWNWV/C6bheaU4UhFkhe0GMoRiAolf2+V5rNLKpb/omnsatMgTwiLj7
dydm1sYyPzbHLS8zMR2d0ls6TXZl2cldVsVbQuMdB2YRdkJsRp6yg4EGt50VDcJJ
3pQGuQP4KHU0H4B520/fMe8i8w3rWMOjv4pTARYegMF3n1b3wgsRsVGIJhW+gv97
k2co6DyKjLoY1aVsvuKZouEl8wNBku6mC9AfMuq6TI4/0wK8tnf91urYWYIJ62g9
ymRNT9gChoj22u30hFAmr7zy93d32iukAQ1FPDWwbySUmpWNvSnN1uPASPL08EZO
R1+7LSaYx3a8DpLUfu6/V8NEBg5ReHdXNjV2hqGHHMFi128PNJuWgJOJRtEC3xOg
bQqY87+fjSzgN/2N1W2sRvXi+jcgffHwstu9b9i8zN9gfL9dnzpNI5fhuT4Qz0/v
oluOXzuHFDP2VYXACaypx69vmLyTYGXHZioxklcRhvO5NuzKJNL3Pics+wEHdD0F
3PkLHLB7k4T3eEQfu0vFq1aE4qzNiyRD02rcqrqDnmANE2YdwmhIaaxA6SUU1aSc
gE2A7abTQ1Z6a+dhb8aEmhZfiPWrilKFIgH7Um7mMnyeG1RWnNAzgktjfYZsCE6+
Sx3+urGql9ErxUrcAtlyZlSDbdpr4nAc0ieLp5oNrJmcOzJL92tan9k0rghz4a3L
wCGCwXcN02VXGLoKTVgNv8mILa/5dUX1Qj4mga3MuwoduEIEBnQ6dq2hlc9HzNz7
Rv8M3Qm9ICGgumukYhjzc4K/gi+8llvekd6EF/GgTUMHcK2lhDxSQ0cloTgwKShH
ql5+XZA+4bIvDDQ3EmHqrDjqHi4HIvw42/NAUEgNKd/pQeNErMUDCPoKXHwqmzSy
L64RWzgDsnh4UTg3tliiI+2HQtzkpE1FpOxdfp9d2iY3lP0JNitI/sr+UYFne8B5
z6Oewv/R90zBlRVKjMpsUuTxPFw+9hWXL23dJiIop7OlYzL4nXNWP44KOVX0Tf43
fDfLAX8vb4dvHSx1XGVszNUOQqcHqzGdRhTPk0ukP0Nwnh2yCykqbpQJDDiLxoMi
kGXesNgiHMeCSoGAR7S3zJIHXEhfQnn7VPZTBnXHnT+Yd7BE59u4OxzL9GhW4d2v
KpPBJlQnTPAqbGzxiYUYD9P5jPfa5BvFKLxgsA7yM2ueEQH/c4FDNUORn4V52INO
x79msQSW0vclrgo7jj7BqeUjpvhJLWzYnb/wy4HWFbdehuXDjEEtcTK9P+36C/rc
/eiaIjSPTQKK62zy/9QJYOzZ6PDmaFjyJgunyGh/4CBa/pR8Dnf/0jdNprG3Lud6
39LrUkV+0pHBb2n/89Lm4D2UulJWicFprEQm2poP58uNgOmJJO1+puUA9ssy8ylS
D0K+auBAn/y/hhzYu3aVr42TidMO7FgvSZcrwRKI9ii5l2PHinA5NeWbg/VUHxke
HP3K+qCVj/Suc3M01ViOb7BbsYjMdoOivhzkDd0Jh4AXIBJre0aeFH5jfEysS0+u
M1eTJSdmcwV0Dd5Tqu+EXY/mcqz2jCcDw5EXJ9dqZUka/kd2To1paQ1B/7bCdna3
v0PxPIG8baWhb8GLciLpeJBqr3X/q5gomurTPwvqmyf5bd/HiVIxuzJUzv9RoD5j
3yaRO3PkTjrc1epDqa3HNyZjAyuwGjSkDSKqUeMbMLAtxG6XAS57vPvzXQEcgV5I
Hm+/CIYSisyVRwzuT8ThaSx9IcHGoMEOLIBquBsiBmbHVbpc26Yl7Pg7S1OWzoQz
qEmunElCApZYgWgWfYsp5PdjrXenVhb4r4+H22ydoNeg9PXos0mnVhcQirMTi8Nt
b0fjTu5R+XIzb2XFMt4aqmtBVoAUDolwqs17BmGM2sKrJ2kNb7vB0wR1tbtdZtnu
lp6DYMZHV4UOSkUlANOkLMPWzPIH5WwlodVbVTZ5hHJ6fLl63z2Odl3972V7TcRI
4BzsM3kdaUIlQH69SKYhNN2C2cFozWs4obowmu7u+zBL87etLGKLGsFCY/28H/5B
mRLkLVWytEoiFoqPRrqS/QdB+jFe//fp6Aefcmh6iLedvqzF3bBXj6KShmluBj/f
9YnXMlu3ndyPTJo13oX6bkbTNSLV6jZoBJcBQibfUZE+wp2uIvfhId7o8HESuPC0
vlJZVuNifOTsPB32OLNR81R79Qf4+uOutD37hwV+OzL0/aIDWnJu/Oiegf46QcLj
ri/tcdUos8amUZwLsT35pk/BHBVGGq/f7lBHtGlPEoA9uAdkjX04r7xo9McZRTdO
7uQKpjzNy3lKEFov+ToirjpBoYS7g2CGfhhWtkOhKwqBMBVyvg/4X8vNwIPNFdkw
8hZYdiZ9tWf1X3DiyQBwO2x0NBA9miCVcIHb5u1d3J3BAcYc/kWbp4I4rRERe8KV
k6nfqFQeVi7HF75SqSVKZeVdbYBEVDkdb+Mz+W5Rqjpc2E5OPNNLGXXAQ9rPXYcz
E+j/mQ7Qp1tm/cVr2YuLowmioT56ppE1ufSvoqee3C6+xjMhwIsUXL/3RGjhKnCZ
y0sh6TS/gCnImAu9H0viK39/hOwis4FjIFkB236KfvdOVyWzACBgSYRPBhXG6fUZ
5ffD2ZqbkUY9yimrE6etu5kIBSmPPyhhwYTB1VezNPnpY31vKSQOKB/pI2y8eYS+
4VzmJ6EXVExUfY5uF19RLd3UlBu/YmYIP60xOgaT/5Uj2tETvJtIhjXjb10jlt5c
vHHB5+MEYNWCB1C8vpzGDZoOQzbg9h2OsbL0voDb+hnxauxG1G99XPO4q6bFjJOn
QE3djhbnkSYH5bqOBwTxbA1QaSxDbNWlh4eS6apSrsDhm2yewVh5yb69I+Kmwedh
WWimsJ/rAomV5hGP30kOZqWcMmX1NcRzTGYiIjBGD6ObiGCGcFEWzmm1Lo63dOXE
tfJ6w8uK45X7x+R6S7VQ14GHs2lOUZS7qWlH/bMlszJhtEB+KAdRbe56Mzz8QWIE
7Vh1JC1ctZsu8WEg3xdPLbc1SF4T0eK0z0W0lcnzPshu+sPz3hu3qZw4ppLGtHBu
hwaadm3i4SzKsA5yTYjoz4qSFRrQYrOMb1m4GUHs3VwEZ3x6w4KC+lvsWf4EEdYH
kkO+qtT/xXz7GL5RspvQgzF+mlMdnk8n2FS5cCxHjIb7GvZU0hQM9gKIgOYwCLAY
7DxxzrJYXcS25cVWydAvZmVjj7Z92iKbMfqexfcb9FtInL9XN2idoxj84lYtdrBo
`protect END_PROTECTED
