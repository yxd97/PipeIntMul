`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B/4GGnHwVcq5qvQ7D0tJQPL8sm9QetsD6rhlaR8pPELmaaob6NRsWZ807T7acCLt
NAMJaJYn+Cy8NMKciUc+Sa1GSnNNlCvaFl2qTatzjpybWS1F+NPzQlRlSKOfJ0xX
lnAvujXgJpewLCfBASiapZNzJjPlmw0H67d1vYq7Bq1fB1OfQMztfKCCe8s7FFRV
GL4eSI+rkq7jDGfjkdTkx3a3DA9OIClYfcleD8MmQCmL3LbwJ9VpBU+QbTasd61F
Q8ExwIkd3OUXJz4EBHnuWVi6YYgTa0omW+P46UbZDtMP6HB0P4l60HfTnI6prtGD
5Vh6yTqnU7TVKD2FtzmLLxXVVsbZBcMcRfdMqEJqFePZaO7oSDZ/P8FcwOdFctnU
6g07ZX4zzcdtazukNOmaOW1xU6if0QLnDEoYl4rbl3s=
`protect END_PROTECTED
