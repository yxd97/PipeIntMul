`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FlJrnttN2P6FEkEES2oznr9OzG4i4I8dBkdcKNKUo3/TL1o/hXuIzIhT21mIi/cu
y3ivq8rU2qtpHT+yhRaUVgS1acsW3BO/LbzdveZi8pZ7JT3rjXhATTvIgNVqhjuf
Qququfh64z2fmDC9gBvyRewxArVV6qAk6Z3H8pvuYAvpycTah7ZNHRMvI2l1KR9o
Cp8OKP/prKnwQspOgLqEoHaX4rRc9RWlnPO5f7anEL6k0E6qz0xyPPJ3epsY10Z8
ySnv/9fAgVvhORtl2la0dshS8YmY3R0kAbvRUcFDpBQ=
`protect END_PROTECTED
