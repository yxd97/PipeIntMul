`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ap9dDd2X8pk7fU5wrupkKcpt9141uyL45dsJ70eubpHx5vbR4MGqQAqlEXWwYsMR
AoARfgoX16eQu+xHWB6gq+5T5IF2RNgRvYMrCFNPJY8ExVtnM+j/ceKSbS5rlsP/
iarV6ltB2yQ3BM/ApSjo+DTWFrN2GP4p7VTXnjfPL/NrDNjYb+IUnw9qunL9UAkI
HGjKRn88dYcqn7d2wDtjJDGhB1dbsY+6MXD3KDvSEWF8c2srQQ9D+FZCH+bN04SM
9vb+t9Jss4iQFGLsOJIEppt6+mkwYsSgSKUT+2LiuiPvtGSdxeDXhPrW+A8Qd8io
U23fyEkvVUWxUwRrCVT3/7tQaYJnGOk7tqzp2WcJp4WGi+o8k0AvEb3B68SZhVM6
yR/RHoZk4/tNtxEuxKaFZA==
`protect END_PROTECTED
