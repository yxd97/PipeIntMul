`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6r/Sqgi8gHaJesudqvHFLXGHWux0xH0v58zXG/qTlH2X97ErN1Z6h3mQtZD+4yr
qyJHfdLDYKYfZEqgO9TsefenwHqaobEwfNk6U/nXan/8WPUgVSalmoSZjmED2P0S
aijtV8D7mx1cstmVzNRZ8B+4OQrKOHSj4ZjszQT2BqeDNLVqQukFkpII1QgmAQiN
E9ats/MOgpZST2m89mCOci8rx6AV+xBSfyeK4N2UGqc7r/tGSGoxWzEg4fn0Wsgw
LIvpQAn/paKrcb4t8SdPfp3EiDnCoBSpuAiGU2GUfTybHcsQk6kW1vPgydx7q+m5
QlD4xn9LGnA/27FphsHJu9vt3ErNTR5gZIBRF5dUbAzx4ivFpY4VsxRLEchjirZm
VfSz/f0b6mhKQKjMQ/e6ISDsbj1NzdToeK8KfO3HZqb3mbouQAWOd9sR3m+jF93V
lP2hO7zU1mFyrHc23UEo42DNFKoPl9qhfcQaJK6uKlBBnXARbDxJM6NpgZXhSA8L
9k8a03sq4wXYm9j5VRBV+J5s4/CDfAdrFCIqJZpUJ0HnTISGIuo8m9vRI7Jb5yWK
bT8uYc5sfgpjkhCimi35M2yyrSds3H74oz2Zoqk8Z9u2sIgwHJRWTbT2LUZJsOff
xB1Dgouonh2dYY3/RsyvlA==
`protect END_PROTECTED
