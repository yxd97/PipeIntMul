`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9R2EbHwOvevvCOL4KTEP4ZAsl7r7/kacDQHVVElLcdi8o/bMNdP2L9ubK9ktX4+
gMQm3LQY33pj+nBU7wRhz5F2UdBM2iP4QOZtQ5J5TD30+ZcBtbPUceici+y/ZSf6
rhGSNX/jRILy/vHtgQ7jn25T16kkDXd9eV06znBotGmZC9Hh7kGN/RGul+uLsuPl
aPE4NdpYoU2b/YzcWyfRTEAqM6i3rZw5/qDvw0FrKNNCWomORUTB/OzAPVG8C3Uq
bROVwYCV4m4BZeYdfpobwfJ28It8NevWIavVedHv5uM16ViDGPfWzLSkoCv7/LdH
m6PaljOiFA8Lp+Z7uAhQ8fKdCd4GReBehKv5V1PgykUwaQPTLQiQsLtuH2qavqsA
Tr2fYRju5XmqrOr1sRHHtnne3s3RGA3q/qm8psssxE6rbF/blvKNF66byx06YS/N
`protect END_PROTECTED
