`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jVMDwsYZCLwg12aYMq6duN9oin9Lz8ZtW9+YQHhvQu/BUXmgHiBpJm2W1YwuCiRv
EkrtqCoCY91G+Y6C4koEHJkCJ9PI+MQqSw5TSRrt+388Mw3G99zqwqJgpDw7UAyH
Vg8/hFmxLozrCFyfJOvHNWsUaBdRMFpKJfrUKhl9vbO8Cl4xtc1WscPl/wcOP4Tb
di2k4maqPXc+OPutnXk0QnYAfMuMYWXQeMd2yJBH8BOMKrJi+Ml2LyjjDMIeiv66
LwUeE+dZkhKikkKO+oy571zUgM/JXsi//eCnWbs/bDQ=
`protect END_PROTECTED
