`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
atsemnasA4BFIsDWmlQ8fm7+4iTeahpu27jklckwKhj3xXbWXCL9Z+ONEEM9JTuO
1wbYBMqFWssKMCLITAZscja4+xnTmIXXPIST1on++JaiMWlo26LLdKJlZAPjOuFO
Jy37/jNzE6r92j8TgkkRJO8wwtNu1kGdqZrWfaUqxOlBwMie2tEKncMt6SjE8Bkp
8ppRUjvDe4SbeKGFrJVXeRDwiJHp+R8mbAuejBD/QumYDxg6h+IKR1IQx37sFxyG
w4g7cJq88uzdFn13cwpwy/xxoHjOkUHLWp1pRQzuPrKFRHCREXoZu5gqsVl4Csqy
T+PilhpMSCZUMIFGwD20eQ==
`protect END_PROTECTED
