`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DpNl/kdpkezTqj7ptVBajmF/ewOWY8a6Y7cGf6oSMTV2YBTgV7bjrA5Ef0ba9Hme
1XTQKms9995LRVZMDDdytY9w/Gsoyc4ek+zQepWDJubAP7Q70DJLc81sLGIo3Vv1
WhlBiPYzi0qx5GpKbfueOKbXan7VFLeRP/s+iRD0YxpYYUc9tnyvZnNb+BjOA2Lq
RQCCuFVtGOgUpRW7f7IFJeszgCXMFLikDgAVZ9Ssb85qCzDN9WmoVbRCuppUzd2/
2n+UnXa5zBTV7JhnBeIRgJGURMXckDEXqtXIlbU2atlGCzy8opj2B5hWQIfaghOy
BkxK3GNNQEtI7/HkVWimNCPkTn9AmJLfo4pCMpslyp9r8o1uv7glPXWw4CNqDzsJ
G/OEbjFwdLftb/s5uwFzI6uRnp7FNaEI53/lEZd9YYL4B2IlL551YLok81lneLF/
0iMswwVtlDRDcSEDGrx/oHtrfvQtAH5o6dksB5i8ZN1wubZWLbnfLi3R2ZzX3XvO
TX1USZ/tH94GRGdYZ3M2ZruJKeuZuAWU7MUDIe/am5qUPQwQTnvLuKiHXDRAIUBT
7klzb7GU3gSRcQkm6jFyiLYVf+dAw/vi0Yytf9NburM6XJZKIH8mrhKt7L47SVqn
ISC16bha+1eIJ0VOMTJ2z8S6aREhlF8hnd5Yk5TN4WLxBVvrGo4wa/dffzF6Yvu2
yr/GLJNBuSv/o4RkFrsKX5ghsgoEGP265hSfBhDMm3N1uAri/BQglQaTBaZZ6GV+
8e8tqQVbnziUejSDe97sJV9lbN9IDSKdo+p3RfipzGrk57fyE4WBWkEak++Ndk07
hcgToPhdt4dHEHiqo3LB4l6PzIWRKJUhLC5UjGnIN5JORXJ3o5I4flyjNY8QlC4v
fs/zkbERIIzk1Wy2Y58v0fGkTqTkCP93NDM549+UPOfFqlPC5Bdvvu4pwkWCxXgG
nBd7Oo8WThY2g1qLJWu3TtwFzX6Bh+t/D7XUvM33KI6IOF96jRfm08AEoJpcCWcy
0rdz4EqVtmg9wGeIJzOElEZj+rr8AWpWcK0LSGuzTbZzjI1buyIbFTOGdASjPQnY
gaMbVJyBEVllyuGPPQMQWo8ZqBrefM5WMAWYH9gcl4SWfXOx9Jv/SGkticvEsTvu
tW0WbGBydrFa8fr+9qHnG7n1SfFUvEqKQE26rY7qtzh0WgzCQeSVOAPh2wnisYEs
eXIAQWkwUa/m40KcGvt7YMztVKFWiMHx5QxfCLR1feOB2sQ5Mzip8QuKhH73i5EI
dvDjdmr2VyUbF0HMTRKEtnoGq0bQD6hjoTReRreiX4gIm/i63zmlrdZpcmibBEYZ
/k3e/VTDDyVJlO0a1PppHFaz/JXFqnS7477g7gdxwQxz9R1YPQZsFUMt7YLrKyHp
yG2cA8P8pRyCgumcIJB8jtVY8ohuMlY7nViZM+iy66rG8Ijq6tWPWpP0GRZr3yEP
sH1RvzjKPl7Moo/cgEcoEUg6iYAB7UyhZDK0BOmAEf/ewosVbtk/TQoQO+Lrc2NL
9RTGiDztrpLOoDNSR0TjBAR5CJtVcPN0QPanKpYOjADevVmmOLvW9zMV5EFkucyp
t/umHqwOSg7zlDbfsY3jW9SO583YdHsCQzP+hKxWVtIRCUBVCyz+l09Ddpe1cNQP
DT1Amo+EfNy7LITKwOmdZKdXqNtpr1LU9muqybABYis=
`protect END_PROTECTED
