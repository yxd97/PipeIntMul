`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7u9zp/Mf+8ngtCXgMo3P8XsFs50QPm/qpl/sfyB+Ls4uLkJdU54iL4oH7xNPMlcN
r9WE6ECg9UsH0pvhMG3aTJ8x5eLGmuIUNam3WTSpIGKSZfjvkrVCQTKbza/yEEiW
LYtWeA6331DLC5WBzWy3T87/SrwP07BhjVej+s9Quhu8imHa4304yXl7/RC9acsk
m6+W0HuhCCi1uNqN3bzK8u+1JaIOr2jwraycfNdompzBUVxKwpWzCeM1HSC+innZ
zo/2eaEQ01XxWVSR+powoWl70bwdgT+i1bvlgpo6zbNqUTO2A7akE0Xy4qXjFpx3
pBt4KSLsriiFa6tVlv3ZEERVGcBqk8/gj9FyI2nnVcltStXGv2Rhq4EUvulLDXxE
xsblvpCzN22xP6V6L4POahls0aACAt+apAZUmvm20ObP6uc3YIjflnwNR3dKur+n
y2U4JFygfvhLk7D1d2TpD0waxybTqw2u0Jqy6bbhP7+VD+Go87UH7DK4uH/rWRtL
IHmjOGWHuijhMv3Txh0MJsBiNksrFvrZQJHfVyaVYpzPgMlVq1TKPnmW+1zLYBTe
qEtEnMchlgjpMB0/JeCB97rNxUFnGQ0uUPKJyQM23aiv21mjFRLx8m8XaINDORRD
LVK2jzA+BCVVsQSOnqLCLQ==
`protect END_PROTECTED
