library verilog;
use verilog.vl_types.all;
entity OBUF_LVDCI_DV2_25 is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end OBUF_LVDCI_DV2_25;
