`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nb+cfAayG6fpeRrAWiIBCO//mvi7oemIIjWyLtxvEX64Z1D72gutY99QcwGOKzSN
j6KS2qHSpuw/pNQnsIL/d+hsLTIdMgm/s5xMHo+ipxhEN1e23JvSY4slUCynsZgS
d4A1j+3Gz51hQqlSSoRG8hJ0BnBwbY/D+kb+7fiI/xANWGux1OVD+LtLIMMSwWgs
5/jKmbjipwE1+J9oV9BVhMeK4Ntuswr0G5Vu2r7t7KhEiC+HSTISH7qzldbvwrsV
IGXR4ZyHejMre/nob/6eraJtFHHxDaDp4axIxOBAcmXgANeq2eH3xa9zedhcy6Kv
uwLCylW+CgTL2Ay7OsKz2FNimalyvzoRh5HMFY+HO7+s9i4UY1owVer10rdNe3vr
b5bcIrcWIdwnbe+uOE4TdAj+Q42/ECUuRJ/WrqpRnUalJsbJfrbVooZ3rd9BYJmE
CITdL5O7XbWNHAhSxhKnBHDS7D+1BZ9gIPWukuCZcjaXU8fpYj5MMnS2+wgAQa0i
djepOjiCeWao/VSY/703WWcIoroj7GT+6JdF5G1vPd4/rw89CvbSvvooeXXLJEVR
dcM23rK00jkAE4rpK+ltsjDPaFYTHv1wmMvTz8ZUJe4=
`protect END_PROTECTED
