`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdvcGLPhkF3Xc4qt0Jqtx4b2lWrMEpGXj2TKpJ0waogrZA+7zEmG0uwaHRsctLXO
nqlNYimYlwTmInJ7WDQ5QogzAkOl6bJw8zpEAJyo43zorM5hrIMCwJ7c46INofNn
sV1jaxE/cmi/ZQQWXqKUWfcxA6QaYGIbEZUhjDZKfQZH5bqbZDVV22o+9dXkNvO3
6rg6JAC953aSsWo6veh7dxvVh8YOIvMvRJ5L5QbagopPzbwIV7SRlD4rMfGKtwm2
bojds57/XMYpD1XLCUh++8uO2FOM6tn0mSRwb7gBspoLXXf9Ta59sa7R3a1MF55h
5uUdPoN0UnkKP4Fi/8G6O8oifkDz8I+q+R6URjwQWKLiPCN6PR+BRxEKM9Ekv4FE
VLaVeEZQo7gxZmXn+lehK4tWw9lELM5kAO7NVBquxdGilEN1f7AZbZRZoRfWmLHz
sI7OtXROjYCm+OdwyulVSwwmrq2LQxOiL1Xfz2BPhRweZhekyQslb/NciL/8XA8f
22s+Jm6LrpFjxsVe1kAEVQ2I//YM2J3sU6euMTDOSc+Qs52fitRviVb6qO1esBAg
c/PSSt0ur1FkZCOXXftQzYwwgZ1CCWosIMSMRBcKgNJzpuKWLy7HNSKbT/rh1tuM
w0a7ZdoPjmc0N5CyMHuVuw==
`protect END_PROTECTED
