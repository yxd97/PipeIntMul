`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ClsDcssCIW2BJBEbqXU6wUG9+UrUs2rKs26q0DLARHLu3DhXkrEJfDhcUwB4LIB
5azZoGxsjbEocNWNrS9NyPnmeQYeAIRc5kEGpquuGQMD1hjSynQYUdl2c2JGK21I
thGDpa5mLRqDaGFHi7Dq+gqQVa5GAKaaX3gur/ji3njxOCZ7loYC2Tdtrw4CxQmf
SmcCN981fE/27gF9/mB4fK7tuLQbEP5lnBsAtzk5eCC0DMc1UMeycXd+0uGcENol
al6eV6nfmsJ22b1xhqqlxjqPlZk066cHIiNXn3dNoYnIEfQhj+BAxBbMx4KoaqdG
GH5kvy4Lr6WWDg9IpK4Qnh0s/IlMY3BHowlV9SQnz5lo2R0juGQK5rY3bemZxv+S
OXGYFOIthYWnIGKtYmfuDghG6631h6NRqrhYk7sAXXoJalqjOAN50prvbDFE6UcQ
Qjnv5PBJE525XRWnYWr3igPLSXEPdfJlPj9kmcerBT8mZWbea79xWOOUoiRtpy5Z
CBi3OdRZvuuPXjjD0TROYBs+0RpDcaYRIigwRUp2/6I6pZRynzL8bgnntqYpsEFf
D8sVHe3XtshB1jzNCa7+G4qyeRiyn3hGkU4mAc7BM/5hcxPboKD3XZPhuOZv8dX+
yUSTsIoeATLW2r2w8hhcWVm9cwIECQoNQRch930xfvQNeY+kUFO977d1Iq8QQ8Ly
LLZ1QFjR9AXxqfWUYwcxky72+Vjm3/afnCMhof2X/d4=
`protect END_PROTECTED
