`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KmGWtEiasMdN1SYp3cPJZqu+9W9AJUFC7Gjwf7v4mi4245jezrDLmMh5tPtXDpU3
zmSODMjEra881122kyzYi7acDPowvhDvndxSOIOmE2wWHsNF1Onm/PbcqyIwi30M
RtyNx3RuHjdXgQ7ubcwGTSwUiJgG9I1gLhC6/aSpkzkVf9zm+BTd/5t+TSA/5rlZ
rBo7hEs5yGkmjNX8sq0MrBOG8hlCdGAe8mG7dnp4Ee80GcnP9L4FcbPcH/9hxzbq
dRNE+r78nBpl1xnAy9Hs4XnzBxfthXyT2xAaYhdUUEcn7OmC2LrR6fPfz8RR/Tk4
FJznt/H2fzGY1vUVRpmf2s0jpnit1Q7GgqxQq75VvsqLFzPW5FBNNYS9Yw/H1eS+
kQQRRFUvTxffLlXGkB2rffvSqCFAf2rvWNtsrQ0po6g=
`protect END_PROTECTED
