`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AGEQ6wxy4q1agMpUqdgZ1PUJTizpn5I3AUmfYQGdG04dHW1Y99Y9IF1YMcP1zmGp
wR8+FOY6nPzGjDWZsMVK/QmZtqujhgK7JPfq/sBkGKGK3ozN7F079MWZtkO5Gzir
CJJiVFkB4ehjWfmhXHxS7+EYogAbq1RDVaC2LMb16IWrvI5bJkll+HCmAT3XYMux
jCdxQs1TdSfEOOTmQmhqWXcFCKn/bYmq6NsvBsaIAudH/QNOEIO7wTi19PXOxqSG
aJK6J+TAe5BuP4C0KabxM/Bwtpb6bExJUZsO6LPKCuJdnxqmH4jT5f2Cpi7rHb+r
`protect END_PROTECTED
