`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLbVTznWYFWitVKJaLivF2TjYGs9MZwNEMfCnmsBvF/lwDSpjlBzDnnKQCAlb2Hp
Gq538wFzFGdBz5klLqCBmpTKPnvt3swjSh89aLFDu9GaCJr/taT5zY3DzS38Tl5O
9L9f91eXlDIS6tUOPqIyPvp7G6nd8He2kF11WaFqEcLwhl0RSpM2mVZ9MbpKDGnw
xeYbHjjCx+U1G5QB68rKQh3+2gVIE43BWeUzQOGRfUbLYr7/xLMxCwumPJY4ulgp
yFy8KeZy1Gz0jm4TYucZjNuwV1W+8kdeLqSDSJhnY3HDJTexHYJm88DkkzOwiT/f
e0wkMq9z6u+CVKvfWF200UhD2un5w0AQ/jR5toReqP7IooxWX8paANTzq/kOZTDd
00aVJsH2XZKNrxtE0Gs3db7ORKnRmXX9gMf6dr43gZbRjnzoMfXgqRFl6i1WITDO
DwaPGSZ2GNc/bq6MNs7ItnhCQOHYdpXIBI0VjUX5XNR5EEc5NvTtSOI48EJRdzev
ZrR6XhNK0wR/GQ1OyPy7PeSGB86hgtlAQ/HF/XoQt/j8k6I3ppSsNY9uClRbXfyu
2ZIczUiF2lxqQGzPHQkgGhQPS/4dqUsTO2jPehoKYC0XEXtVg/VznYTJg1HdWGis
5wY2FG83tW+NJGbwtA7OkG/aannpkcDwxslSH/Sbnts=
`protect END_PROTECTED
