`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e5xv7WekB2RQfaTq3Hn4Fn9PvZv9hyOiWfJZlOOTHnFg3/vkFfZVG9finTkfiNvT
iwXX7kLT2c4OlvoVGx3dyYzkaQgs757dsZqvR5jN6tPCxolw4+i0NvG6AN8/MF7C
L9qCBWtpLbJOQxWUOZfac+Dcnsf+EqEF0tPqPhVUywhXzGRLc1iQmZsuxCy3qI/H
is5Rf58wCZI1qSx6wHh/sUhtU93BASRAc32oqw20JY4xS7GUE4HUfTo/6GTwudFE
cL11TC4iuK/nAGoGG53lWlgZy5xRN75hvF1vrtFryTrUonYH5hq2X2eb2Swg3HZH
LnbXMaBlfdcqV6+W5hWLMagrO88j2pn4OlT5T3hRkiFAf9MTau/x+uNyt1YzQdfE
odRIBE0x/ORrJhpR5Y3e5RS20t2V2ljjaQb6WoVSPf4RLZ+wRntW5gzjx7rbX6qw
+FWJcyaJpPxfigBJEt9/+yF1fvHkCWPcAfwBG2YGpqV0kVuuWls8QuSZ5yogg6By
`protect END_PROTECTED
