`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqZ7k8CLiNswragdm9TUvTVg0eEZUSZH1+8qomdlERA/B6Jg4AOj9XkLEif0Pe50
OXoXEoWxQ6PW4YtExfJVI1Net0wDAvHEdwYW4vxeIRwAU7AMZw4bARy18WYC0tfg
yj2b536Hy81YfqEcRahrda1bLbq28ZKixTJnQkbGiQQ9aGIG1TsEny9D4krIxfWJ
ROEXgWnMEnwyUV0e9l1XqziFIw6rj7/ZSmwyMi1i15vpiLs1jfDq1M2x3dFvCfX/
nE3DCIF5BjsjBwphjCdLooqFAqi66bVXT58KqqzWaN2VWTLUiErx1NW7q0D91Drs
ZT+oYgIBIAo4VtrvaP96EGZy0JOHrcTC2d6xbqzhUzKxU5wvvImBO5NZ+Bw+OPS6
KdfP/cRI1NOmPGHZVXj1y5A7SF6vhbYfvhvCTcicwMsumETxNwKCUkgqMWaKvgGJ
`protect END_PROTECTED
