`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpxGm8IOs2ofauMUmSvnc7YiBsFkwUlh0UTR71auZizpYGC76v5UMOy/LqDu7RcM
bMCyYDRthfHblp2IZUbh+MRPmboqwXqc+VRL1nLdUJVmQ5JZA0MnKQ3Bozq0Y7Vn
LjzcFpqH9+wNUKEW+2y/AgyB8JmMRIpK2YD9ZlJWpy8nkyIXINxnsanwrmfoFoYi
afkPXvbZqVzz9qcVYfV88VyhBlPTwcn3mdoC+dbL6fqILq3+w3RPvdfo/iIJYK5+
8ljf+kM0pEGKh95XsrO+PvvRyqdxoHKdYD10Mfp/f0EpKynCi2QEpMCMtV8X4tX0
HqgKg1gDgjEFw8iNvHILQ8CJtATAb1IUdhA8ezK0i1vLMz9ph6BzHryXBOjbh/aQ
1MgIwhedDUhAvLSqrtiKr9PLd2MS6q/+H6bkhw+QPdFx9wLNZhmoENBWpuBHyI3B
q7ssadkWhg87PWKWP+BQ/qE89IW+QolTcBzLXkZy+sK0Lvyr3TvD6KuBlXtsdpKj
gUMML/6MrDCgUMLHu8EG2BwUF9F5XX+3RQ+on1l9kusePJ+IwJPoU9wMcC/IHAM7
5qjNgOJXw9NkGjqlWo+HLcIadRF5Z8lZRYIKeXQdv9IzCxFhXAJE+yZzY5D9Voqq
A5SHU3hXDcfVol4WlsnNefHlEU++9r1KtEeggyirMZjs1cUyaoS5z6CUXV/G0oDu
FOay0p7l0HXjH1J6gTtV++8tjpsYOSqAjRkGBa2kRpjmIF3/pcc5ZyRGvkcdLHTa
T6aY3FkUzmbbtGLKd6SixeNBs+Q7XrHx3Zetu0xIMQW8SWaMwmFQZ/2vxHoqI/vk
C40FKQmCTdbx8QicvQ2H9VyYreTkqwsonkyQ6C7kSeZrjkiQ23KMz5NkYefwLpHa
9hMeik/fZFY7icHbiuILos7ces6qJJG5mfG55PS0BXDzEmuDGUfHNKFSBgRhQW+v
jZf78oP2qo+7xfH/+IBPPScLIyIO2MCGPs6V6BIhYQw=
`protect END_PROTECTED
