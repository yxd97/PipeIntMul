`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLtuJh7WTaKDEMbQMLWqtBKMJHm3IFBtx9TUysUkY50O8sKHuCY7OhlJ+GWFQArP
U4z/qyWQViFzfy5sqCAiTCOyjvRczg0307X6OQ5idxLcPaXGXUwB9MAuZhu0DatA
mWGMt46MnEUXkOuNBVo6zjgl3HYsudMFYJShvcGzE/UcxUZr2YSY/G8s0VahVDGu
GKfcLTPU8PdEJSq2BLZEXjynRTGPuwOTpuKq+/22TXUH0d1VKJp+9DJ4xYZdWAGr
jEcozbyKBbaI2mpVl031UQJWG7o1GinuXJ9M5FLBVf+06UW8oE7XRfE1DCByAm5E
sQ3NSyFUqG/OnaHBU/rMazCud9lMAq0NIblwC6gfY6eWe1iSwJi7y/aQn+2aBUax
1me0dTDalvvsqKufx6gneeetL1HA+e/lGZjVMsD2cLu8txhtHDdLrW5oTPzDiYv/
sYzn8QbgaKRGaXJ9FNb1ovTUzAFkMduUS3stU2NRpuFK35GZJLAR3QbbEKKy5Brg
QphgdP7BCCH7ZKYnWCRbv16rGXb0Ik5rjIFCY0/R4gr+OHr6sSwbra70j3a29+On
aq4CH5EoBRZqMovj/kZ2u0oww3wNEIlQj/YDLAeHiFqv29D9IY6YGK+lvRbnTmJa
2kOMB9d+v6nDIXJPwfhQm15Gh00sqa/v6kmrVrVz+jC3EzHaGcKR9kuZpGQcP/bp
x6qSnhS7QS5BL19zc5uhE666hn7153qpQT5MYLS6rkLPKlSdfbOd77Th8JjSvAtt
`protect END_PROTECTED
