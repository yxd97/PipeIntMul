`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRG8YlesBR5IpTaAMOxzRHma+ycle70U4OKng4/vIKw8hZHhj3TeuQAYKwZYMVUc
kUJSfvcmkmszkGRn+z91/o5VAZw6JKvf+qzGGya19S5Cvh1VOvFxft6BUBHVFB7H
zIo57Z15N1tlcj9o3SRcuUWyW72BR28yTNaYRlkLtjJay/M6O3y+S68YeaSN9rpx
yN9+2f8XNX1h+fD9Hq8EaZYc13prKAt6sH4KDCkJfPRA/ChXg19GPa67j8JpyStS
8Ni+gi+xxh+fz3rsRjLOy8J+y/9ytuaIBFN4JyI8h4PKaX2+CY4re2PLcY2VIbSt
LLVHqMGOfmXnFjYTt4+twpiJqWjgVQiIRrVz6w3XMC/Zp+E9qmg9s3EOc5Hrqdu3
lQKf45cp/Iris3VenaxW2WWTMGkmgmIg3Zgxvis+RA3JYwz2cgpcnSK7cWBWFoUt
6rbffdI1nWHXEXRxA33MY8zqv2dkEk8lo9bGOYV/QsK2fERQZ6LpBV5I/GamFmVk
zPEnKwYe8n4gjMMjn6NeSJJ/E93OVxfWNwhNg69Le9ZgF7y/VbE5xUhRSmi1T3bR
IwxHN1Ko/AxaFGtTIm3YxieZKv58IM2aKy4/utPTeM81gKKReQhMlF+UYPRz7UY9
fycUty2W39zlQ8BN7BASMj9rst4HNAHMK0CMF/DwMOeZlUdm6Rg3YzdpJrkvjHGb
XZVmAsLKM9ABGaJsDBZkf4IOAFPeZBN6boWcpDQSZLEVsPpuUQJdZJ9HLjHKrIa4
Iw2c8bYGbZlP+0ZDY9HqtxBqx1rr8YWxhlhBSeOanYXIQNZe2uvsN+18yGDbrY20
aImHwXf5B/wKpTS4ZNmuquZkD8akH3IUCMXBe3+R4S3OTfVYow0Q3lbVpCdSpVo8
U4Z4EBg/Uh401DbASuUS6FR5aid1jkzpasmE2QIpFJGqy/uysBOIDnoGiSHAIzyD
4ejs2XxsUFqCcsw54DS9aBUhzrE6crM85tdgvbuQAKdjM/Ssb0LovcH28eBh5SAd
uefnQPlNIdIN9c5o21HmGdrmtFOAD/uO31KXucXRCq8HuOxHLO5A1Iuv3gMNUEY8
rYr2OoXQoVVUVj+wzCIIEnMIporVXIZkEZqbuCUn/M2ilceSs+HyOs+f81QojRv/
8kFO72D3N6a8lkVD0VfhczjSSkl3KSZ/eqpDk0Cr0WFTMkCyvSJeD0lOeJoYzPYV
125TlA8C67dufGy/WA9NFH8aBn1Eno+CNN58KMk2iEDz1pA7pM1Ndsvlnr8AYPfj
pGoP4yeXDmrWvYVTI+aWg38HsODMvb+GZhmotOnn/JaqVQfWyExlPgFUu6GkZdaJ
r55f2ysiUGbup5zeGBhAKJGQG4C+dLgsUMBqkvoFQfJWsqm34RmlvspRMJtjPCYP
mOTkdrvV+vq7PtyKhA0+IqgMnBu67x9IPY6xLQgFaDg2JY6eYVzthGENskA0Bst6
Ii1FW4mwIxwT7IhTrMg+gi0xj+InA7A/VIs1L4USxkGHb2guF9Q8vtaYJ6WqwFbj
wsUnU0NqjUlOslpET0QQSXz5c2AilVQzd1JszX9vBJ7F6ofgPDlYgcprZb9ITJhy
N6VQeAGI48jNcyXgwPi7fowHFAzzOa6WtsBDelYIeog1vOnDk4IlGA2r1H4RMtXi
gWyofY4J2S9f4w4uhYnC51bKE3ZNm2BU77V4u5QRQXFG4WplGt0lFfz+UG2XMgbO
SdpGe4OCCt7i2q6acX1ocsWgxzrM/uHlgTSqX7SR+QYo3tFse/TJYp5F3fRV9lcB
tdCbYJE43vzn6yFBTH3AokjPrUlpIKyax1KB8VbDiV3QrpNmJAW+lGcX6VLkGrxs
i6gd7GTCwAP3lHx20hEXxtNQqGCHQHM382LC9yABqQeL/C/pMVXE0o1e23tWystH
pEpc/hvJh2CbNbWjRk3dXwE5LmetYOkr5ON9QZIhhol927LZFciMwvTGqfl2skcP
DSO8mB4Jn1z+M+WvUYZBpffId+l4y4hDmxrIgDpzuI0Dih8Zs6o0tk4RiJyIGNMX
yXb6kaXUMqZVbKyTTYtqUpoJoffkzGqH3R9GcqUVq9SMd7uK6HxHt29rNnDOQJBI
m1nUey3Y24Q/q+14SSjVYCJ0J91MwcxvCuvCkmDHKj2oHdDlP0d9yF0Y3q9yj7Jc
pybS6d6VQ0Q+b7aWziaN+sVBZrGnmINozkuvfBeJU3Pwg3qIpMUIFyW2JQxaSf40
KWf2ixz7BUymnsu7rRZaNKt/1rglcw6QzaDv1hS538pCwggf9BJw0o/J40pNY3fD
Sau1/QWTfr1OvSSlPi0UbN28e5L2xe5traXXiGJE09mBv8BeYmDVuaRlx8+fL2Je
NMuKeA2dCY7FK37gL5+QOhSrCNQCHs1uaq7SDQMWlGy5ySoXiE6e+eiO3T/DpD1h
0xtzm8TKp9768PMd2XawAAXlNhp8yZGoXPcjt6COjhYz6eak6laGyxSXsDdjisdL
PU+S1mUMG3U0gmuFP6zbXrAO7+6xKODasW5FA5TIXjgaH0T/c8QQQ50bX2jaGF4P
NMbxfGSQ9Ed9a7Mzz48lMHA4Pa6vmtSfJeKungyC4ij25x0czDGWI+HwI/100frD
hmXk8qHlvTgHwGx5fNOkbBqT72l330XYM7SRvlgBOP6uc65QfTUWgrfkh2Ogn7b/
0wbfCliQ6YpL2yId71vET8ns85H6RVrkZkxh2bk74m+QHjdukdf0as7H3lWm/AGI
xgDIYlV5McC55l8aPbn9aIYKTy/co46b0KiBjZSXmzRtGseOCLyb0cHSk1QqRxMb
ZhYIkHSgHHjovYpNhro4zQmZRUErcHLYjdicBRWSM9H5amxzfUkyMocVqInypmCB
PdBBBA6yLT2zW3+i+hPPli8IlE98e38wZTl6uYUQXmakOex8ilgOOlKCLOz+Ug//
8xASoUF5QDHvv18HVMtQuA9qfQxYQ6Ima1dmw2otVD6lyb5vUYAU+hTgdkPlYSxU
ZpbX1ky4bocyIQtS8XCfgn6XI0RKbJiNwSTC01U9635UiPw0U0watggN+8Lngd4L
zAohCaB2c3lIQ2Y0X4w/6Web1nY1bMwBqhukZntA2qdq9Ub3jQCqHXyPLDqhZBsM
W0bKX7mqC7DiyB/Ziy1QJIgclSEtYeYScrFMxcdCqzO0O1V48wNDhA+VlSi2c4CG
O7CanmeOEm7ZERRmgmHbwcrcdnmAG17k2OYnpG5coKKTlrNgTgtNAu6jv0tFJGFl
g7VO2csd2gO3vOa7MBcJXxFEZz4RHY0htXxKVbbydMopFkP6IzESxT3OEaJVjF0n
6nGeO8AvILS622Bibeuk+kECWQvHSc4jnB4d50aZuGm5E5OHebxNoLoFl/k9tRny
9sdHxpFDkW00YJib4MhQF3rpZZ/U3IdxgGgTBBptzYwUx6BGJGYu0j2M2d+TBF4s
s2JHNSPT2eQvnj2Kuq2X2aRrbudSnFafE5ZZZB+ukcRNsOL0pNoT5PbaAIXzC5FD
PbTwX8Zyydy4wTnb3V5qIFlVgu46tJunjh2jr/RjVejxbc6VKiD0pC/dLdWE6OkM
+9grf6xT/RnTOe8P2XWHoHVCzYFiKPFtcFYA/1fOsIuc5wjxRAQ6bk7Ub3tszXgl
5nbJn8TMLIWlOq02XnFt4vIj0RTzBx5Ghj7z+Ui9ZPwXhPpW8dIFBM/Qj3GXg/mw
iPKoZ07ON5IrelNXoLqs0/p8j4wnraV9k25EEJgzaz+A0WeauhMQYPtPd0s/Oet3
NuiENBWuXXEcpdtpMrtrFopmVTX53IONOz7PlG1kRQg18PCPBvbpAjWvLvNYYf67
6Jz/XdPuQKYMiOXcUGCTnB4kfw9q7XVhmumgSttTXiuc1N+TgpPhzHuNaEHRDKe6
jt08VORaigT7QbCSYY4h5oPQD7gSl3rA0jmn1FT3BE6cFXmetAwn9qJZI4s3kcM7
pheHRKJcC/0vUErt01HI4o9LKyKnSLtioCC0pRaz8ySUx36INRRIzcRL7NnIwoCR
KXpIl62+4CX2VD8hjuPAnyFHNh0ZRxb8d4Y31fkAf1k/bzTRo4An5JXHQhmzKUt9
qXHYgUJbk6/QBKrnulAXmWo2N1/jNpv4fRYo+k8TJDzP6wc5gW+MGZM89wcxT9zR
W82isVatF0AY5I2qryWbeauwzI8aNEqDRS4DLvit7Oq3Pll24aeReoyP2r0Wgx8D
gpbC7XTgx5WuulYMSPit/VnTmZLEFMxvmWey9PFXC0MGhuYgHWeDvjCCOVZl1gIr
5TN3h1FuA5Z+g5aDMAIOLfbL8Cp+j79GPlm9SLwY1f0mx4Ped+yS3YcdrLWaN+hK
pG2EL7f6E3ETl46cKbyagFWpewd8TfjRp5pKQStt/P/StEestnBKou8iRCDHPaRv
Jsfzmg2LyuuG/xILbsXLnqI+qeFyJUiA8jrCysKJBPw/6H0ENnRQs46UgDafU/GQ
TcYneUWzPIY/LaY4v0p32s2DNhzyhEJ/eI+Kv03Lg5ctUe+OmGUBFfJSbCjr/CbX
edQzpMo5VqAC/0vaxhV9zCLx4lYAW2EDnvrMoOTaZ89FO6CEUzE0U+tvQbhFo/0e
+7ed7A80ofQ88cWpPlp5j+nd4OxdOaxiuUvpAnCrMOilZSO0Y+W2RTxc49dfE1z5
KymXghR/7lBqRtV1mRMOwQM8GzJJM4CU7x5r+C3T0FKEA0GfghaNa9rH7OpM8TgC
wIgN3jkC4ttUKnQGZ78c8OniXjH+ECMEelNA/B07y56EfL69r40DzLPGk4IBIj0Z
D/GQzuu26FMuuTyPHUFz13LgmL0mdKlseLSHYzo8q5LIvUmPrFZ69hZNPsZK57u9
U8Yg28DkPr8wIU9lZEAnh+qyv4VRG/jMnmsIZioiy9UT2qOf4wV6trznuS7eeCMH
a4YwDCdHcjLV7okBdwtqI5Uw/2KM0954y1LJDpwfB/WbErbOi4+6eBOyZZfH6PXN
qhnqUbKogx96uzXADtKkZVuF5QSCf3o17dEU3og8DfhdXXJvhk9ZSPdAmFCeVZt1
ZPAjS7+mllrsonhrKZ1yK/h+eT7YnCnrlSgP3pITau67G2pCudGZXdsRzdqX1A72
sf2Tjl+/OP6YEO3vOk6g+UYUBhjLLRG9oRkEV9weoTJVaHuo4CusmLdk41pRG8+6
Hp71nXWYSp55id91IIanQoVCygbRAPLGMe+Ex1uxPc/heCAe+PXP8reeHZ07bOJY
MTll7ThSQfSUJr0JUtEyf7ixD7Xc7PdgNxoD+w/2vKIdzUg881OclkclobB0aj5/
53B5DWatdGTtShee4QAXPzu1OvX2JOdNjW7NzWMBivme9FjS/949jxFC0ZArALeT
0LiBVQM3iA9zqko0w5mz8O1d5EyOc2lbtGSNMefB9dyQ31YqDG9BnB4y7YcS9YwA
EFhUjCuxHl6v+GrcqWt6fbtpKcZKQO3kA9+Dq5eeo/iKFBgcfeuhPfEBSkKxl5tj
OFhmnI4jK0pA6m4OuSSsQyPZBix1mUJr/UCl46o/iDj+M9KaYm6CI/Z/bOSULyDH
+SQyN6ShCk19nFF8NdCMFbhZcb+Nm+EwZxHOfl17j6h8VyuZitEzeyUbzird9Z36
0VRAATZraItPRpEl23/aVnBKxJkXxzVDyMqR134TbcqN6SHbJl/65P1nnPcyvx33
gLGO+lS4Ycv2CCXKrfvVMP+VPJJo/+qJE80G/TFtjaBlGifKqLXthDlNNdiK5s2m
+q36EgnZbpGC97gHXjuzTIsr695pUZnJxBlhpAlF6+4eGR1a0A2RxNY92LlAHhrB
xpkwCffBWSRQzCiwR+BQbHzrVyRcKUahcuninyzXuPCkf9F8ZmFFA0eXewxJpcsi
eHmQglfybGz7l96GXNjr77yAxSrTRAg+46GTNJZ8JyK9drsL8gpMQqaw9G85FXi/
1EIHL/jE4LdAC+YmYLaEGZwd8PG+c9wAM7pssJHuBFcNep5e/bPDzOR3dVL7CZKI
aNGF3K2M5Iz8mAU/1avkcv0hUCtllKT+ydv5ptjEGVzVaKbhYHZVa1lswi63yxH3
LjiiIBg2wwei+xzjkLPFY9syJjl+qHsJ+kO3KjUmy9bStDpfWlnWjnRJ9HIjOPIg
E/tBz4ZV04C1US1CLMSXH6Dx/556TbJE9LGpE3gXuaavOTu6cHSmKOVVOa5uff+T
fUMtULxEWH21Lg3VUO45/WAGQFR3lcipgX+v0Hr6lL7Tzt0N+qfHry0WzL29ovR6
4f4HO9Yl/tRYyRJTED8a/mwxUOE/gfeTYC6h8VmatoTXdFFVXcTtkT38NW7XInYW
Ac6gTRrsdoJ4luDktt3chpOTNOsuDWtgvlXoWfyIg/9y1wEYS1GuRHjSs7lN6BV5
ewpnkAyHY9SriFNF31FeMwEgO9/0Sl5PG+tlcAgEYMMtIbXWZ9AfpeBJnS0h/7Hq
tEWXUJX/QAfBJqSjUKeAU6gu/Czts2LCMJ4jUCTtif3CbR845+d/Jit048HNDTAE
FMXJ3liJE0mQaVor3QFIVRiMeR9mcqKY34GLb+BqVo731fIPWQER+0YonbnIHQcz
i7oujpzuzVpzPia8psU1YnQ5Lynqwm6YxJyUnW0YZuIDk4BTf0SMu8n08LClTzBH
5ne/dJd52qO8AbQU4R6X4F5TfTuq3tISDRj8ba11Fc5nv7mr5nYJq61q7RqIxk3d
kMfHVPPzHhzVjJiGln1CXFRaBmPhq2EWrpAS9yXo2Q4p+zkFf23vVLrqZ3S1AWxn
mdWPhAokeahgGe+RuzNfb/HA3oQQc5L9eCrQFp4T5S/huDMlDutZx/0yPpp9xw54
yTk00kPiGr2d1GhnxwcQemTcALoS7zvd7P+trxpEE+vEcUqMBuKFvIxH0sv6yNRh
yHnFiARpluoe3Yj8F+5u7sLogyNngwiJfKW9n7FyM+aj5usONO3Ylj8EYKffE7zi
k/sLS9+FIVVVC5CGR6cvpfJqjnuviM93/rTLxvImu3kiW7c/GyCP2O7qpDWDwati
kwE64JL9gDgDhiiSR3nYRtsUsSH7R5R1D00DwSH8GLjlVfnL38Hi2RIStKBjebXr
+NF70vjyESqHXoNrdKiLoOGiJnPf0MLOvsw65iGpl1aJKubSWDXlHF5/aNA9dkAL
zCfwgSbbpIXXBRe79LIqD4Yga/GWTLRlsx1PdAl2R12Bs2Vlf/6UufynIpL4Ie0X
mm+gG2JeGld3faTGlUvytlfp3JmEHIKwuLROIv+day/KPvB4cHxtu56AgyV6oDff
rRm8Mv/syAbyjw9OlqYCLPgQUru5YYfiaGnAVVw9y1nniLhMQSDgMzSjXDLihW2s
J6Rj/62/KpmDsjVuWssb6d5ubYCk2Q4V7SEk27xbrat5/NnPhFoFqBiWKjZe9Acp
w6CVsZ3mw5TtVWbkPKnFmG2CC+6sWx3hdSiBBe2kYegsyBndLY2iqsNYBikw6I+n
nb+lOzbrtK9gBWfa4WWQo2k+k+zHlgttwFcnUv6dtPAhd3ZDmmLpkMRs57F3/Jww
yiDByLOJAwjn67H7vYa6UfKBmpDdaZJzxSCwYYtwYAsqpDN1bgoJWUtO/aN2rErO
X9/sSndW6P+7CQBZ6bOg/iweXyVwlgA4Oe9mAbSlX2dGwffhU9mmYOgMCvvY9Q1o
zflbFQy/s6gfDki4ficivDqyQLdlASyo5Atea9w3TodIz8rilpiQd1mEjOE6pN66
YLxfqA9PXPQNXQ83izRLB09Qlg8SYIkICSlEaFeHhrBtv1RNT7sMOxsC36yCKi71
JIBHTyfXc1T94xTPMQX+PeKeupZfY1MYh+Wx8oePNARWhZBJ+rBZymskaLT3Bmei
TV2xcS9NjbLDIqr6yVETkW/1j2v0yHda3jklCqP3p5Hu+L0kA3LkrkXSWMlKiRWS
LN4+TaWkRabg2MUmyVDURrFDe0Q+CZI9wRJqsgbZJGuVjPcwlxW/v1SxlaN5iUz4
mQphthoizTvY3TcE7WSgfq7WMcFHIQiBvauMUO8QUWzu2DoEs2dTeaLEsnrUbC2R
ojksXBnBG4or9zil20GiS5ATailo7DcyyTotB57wOSVbN5HW7Ta5YuHGGqcpfvS/
9i8RPXQl6+ygsey+t8CV+BNqHipnPjHAlx4YnF79xvFapYuTEG6rPYtZYQ+0kPNp
+jap0sWCU1WD7pVP1fWzCRYnRED7ux8O3BsqB3MPNIdQyC760sB0c0SE/m59Yn4w
z5RnVTsOPHAPynupKpZR+Bgnxnh5RbUtkY+wUe8Q0koTtKNBR3V2gv8T/MNAxDhS
L92v2BVLoVUhhRpiVE3TKAV4E6q/HWzRjjuK3qAMiiIsy6o3/0/3GCIg3j/twgl9
HU3uWvgUMb05CztHyRAZv3HJ3pvuW58XOMMDZFBn3uW0PhyXrehN4KbTJqDMlvyk
jUW0L6M8tk734BNqp3lIbZWkQJbZAbrPLWs9yye9w+AhBcKnR9XTcbSwC4MIvWTT
+LDE7ZDksKkKg6gtfy2XLvxRbZztjFuckfcsUGZ0Oc78m44OG2zlLXytzp2s2VWa
sBy80SVEsOsWmfdmOjvisCLNruBqXxRhkClVobMJ5pXu1HIb/iJFaOVxvc/HDSss
NynBbaH7LwgDYMFns58ZxlzyTT2BQWB82eiaxHeuy9I2rkqvh3+dVAQ6zB+76OFO
d5EOIfkmPxcUhyIKWD9s6fC2hzo2r3dDXMQe3qFQzHx9YnWMvVvVoqWmgfObQTs2
6S3ckWpyxRWeWZ6mI+JcAFUt7HvH5Bq0pCsIcu8s00/0z9cqfBAH4CXBcCm8n4I0
bBauD8nEzqTzg4FCGotHEKKbroCEmZGZATeCYfpBUF23J3DGI6XJsi1wo1Sq76Z5
qPctbrrPV8d7EABJ4sMzBnMxkTb7QPwvNcR4zzrGHecgZpYJJ9LGHDwI0CYJaEJD
oazGSmjNDLLevFecB2nIYpcqS+ml+XrX7+imLRLJGVvEA6uqSSmYcyRoWMxOs6SO
w1ToDYW4Fduy0BJfPr1PbBy6uid6cvHmJx5QyItE/vaUg0mGsdU8AVJVxwOyLiyk
2z5TOSZLLBVUhWw4pw4Mt3/DNdtIjOcVqrhAQAZC1tvlo+IPXm9e8cI95JB0ZBUe
k2wqaTmnCVzl61wqeBGvTQ/9F2LkhTExSKo7L/DF6x2Q/QI7wj3RDW4Z6s9bV+co
jt2Sq6usaPltRfOOA9FLszPFMCyNN+xtkCYgzouUyvkas+sKxOeT6Po3O6x3pXjV
iXWkhPus/NsPIMuXn8E/8I940gidWqWkuRxzCkeDXElHi3mB2aGG9OcaS3Td+CLy
dyXDBYqMCVMYZAQTp7Qro6ZFR6SD2yM58Yez4mKMhL5rc5cZYh+vALX7sGfa5LEA
hNDL8h8BUe9P9nQEfPimwZ0sKV8KLrVaNS4UTG5SOOAG6ZNORLqJ1a4uqWuUJJ9m
/ASSzSGEAa4dC5w2VLIkTPX5Lp8g5rcNbeHH8KtCBRsfeQQZzoSepTA2fi+99Tna
X/4TvTlqJdExFFETDIkKYu35HQHl/bRjv5e4imT44yTq6YX2uSvCtoaYGEdNviKN
aGAfIFyBM4BXbt6BRXrfSOypltiFNxV15e2hpetVLho63RjEN4XgGmnL+5j9GKVu
0XfU5jD/HxGC13jJ+VqMj/+pkJad4Iy+akZCBVfmQvetLRZNGzSfC4bxh7NAtdn3
TSfp4w7+VT3Di3sZKMOidOZ92LIJ1xSC834p8bt18mll4Uw2wlxPLPosP8ton7E1
7S+Juj+hF4fvjeFotZeVhKZ+45tn4zr2hlnRPu/P6MEXp1NwGs7sBFdzmWtLLX7I
K9xPx/zkfu0Gr0o6ozuatL1PJCFcxBh8mplJ6xifbTbR49qCMmxw/jN7zr1AWsLw
j3nOpw9KaV0Q4D1UV5h/ijOOrx/TttjPxssMHT9aGxG0LkpT7+Zn+PTnwF6ANoCp
3GvpzcKGVBFThFspOGpxbwXbGf8Ck/ZFuZ9rpJiGU1ClMiMzRSWgT0hRJFQpSdap
74EhPv29+yAcgmxSZFigpRlIqbJeZoJ8rUW9era5Lh8USPfJOVKL654sBoO7uBbn
o/hqKb+OEEMwr+SVUOpEvzbmUwv517y1ckresQTtRRtxVyY1cxubWNTakCEjIqZr
wir+1L8z3Ree1ZZzM7n4PmKxpMZ1Ubjpnl8T2IA7Mue9TWYmTWoqnoCH/mrm67WY
9g7YJFbjWH3z/hYanPAf6nB2YMiH6BtPxJdyA8CM+1858LmB87GqauxxmNi5crK6
13unk/PkfJb6X/UipDSCeJzAD2h9yUenr7mIQKk0t8kNdI4ktYXqD4TqArlUkVpY
qsqvIiEeQ6pcIvnhBObwYN/QWE5wgjYyQHLAwRHCOnPOE79OCvlBO8Bxh9auC3Pz
BnxJ/r0WUTwE+VTU5UvkdJXwFKx+55tCxaQXaB+9XeCYHfgvFXYl731FESMZx3Pe
uyvMVABve7ksuh7Eg+TxAULTWK7b2rOyz5Ljthpx2NJD5opskkcXf0z8EiSF4sSw
QHK4q7AOECEiDgXEJoP5v8HJKasFRJqmPSYpYRHfQfCWoEnucrSP+2CRPklmnw+P
5dd02m/w9/yRXmdxGUnaQgOiDa0WIo9zKJ9ArjFKKcubU5OObIeWcsZ1XxkZJJuQ
2bMBngQxUukOs2LYCtfqPWESImTdGpmEem6G1uIyAyvwipvJF2VOxnz4QNVJ84n6
vZh0ugydy9zYLq7HXyoTZOX17hQkLlr6xsuqMPYsMSbBy8PBeP+imtNZ15NhxAPG
AlX7atRIJTynHw3hkLN4iu4k4ngm/ewKz9xRADuJS9oFCdw7FbQJhse+hMhFRiea
XDHn1NJRaflzMSfcqikgA6RjZPsZlep7gugy7wWrNSbmEqzDZWhGnxVp6klzU8JW
nrRfE0QxxDnScKzeCGp7bt3Nttv75spj/OzLtowGrQ920nYBoXpfzXeokgNnRcES
Ucgd54GJENUQotW3/2R1LmQa+ANNs4xKFGdlCH6IBLvxR5Dr5yEus/TPPmyF6b5T
iShkr3H1PcDwOX+7QzXH6cz2uncAhXBz0RruuBPiiihuMGSJsvoG5Qh+FWQWapuV
0i/mJY794syZAbV7JlHA17tyPtrau9A+x6CVIillVx/dWExyBEnO5ru6JC2bJZzG
HEzeCg3Qn/m7lcbLz5Y0yhxjMw7P5M8+g+KrkoDngdIU4SJ3jZFxyWkfYNoqGNy1
ZJutMaiFKjjZdycN9+pl8TNdWx8NksdBhV6z/Lxeq9YHSNCE+bstZxLH1Hg/NJZD
F4eiVvVUN4sCN0OAXl7GHUI6xY2yW9Uwn+CDrVmDh9R1xSLlVKa1gLW/gyCLX7D8
V4X4i2bbiAF0nTXyrxi3cy3Lrzm8iN/Hwx+5oUtPELvpR+NHXzZ/z5BG+VdRaoRd
dIQZ6W/Qk5gqvr9GEb9j/a1zuTPjP7v1Bv0SDt7cSnYc6SvXK/IfudyQgMKmpqFA
MF5ZqdUYVSFSBAU4mtQk1FUlZtUqut5j7uZJODHNCoFptqUNHJsyytmxJ5cziwwQ
nBmyhRTci5dQ8viG0FdjXCZQZG/6+4yw8OrLmQ1ounLrnOToDOfzAvfu9iFbdGx2
Tyny6QRjvY5/c3jFY0ZMUaTLos7NbNo553kj2sWH0h6NjqeiqaDNLnO7kI1E3Yiu
RjpYGOQGZQtUGjrZl8/4KUEvxiiSTchqbrdH2F4bxG2naJ5gE+7VrI4lmxSL8y7z
ExyAlnlOP+lkWvWWzyJiMgW1X4zU25/UzqcaxTZxcLP6BJTpTQYx8qgcaNYHrRlr
BIBBYIKO7BGIUOdfpcNP5Gd3ePKRPr/Tp4MFp22fI5O8D0lVIzGMLMVwy51Bjh9q
PGzIyvPtAelOVVRm8UuTs3onLxXWCUp8VZX1pgp1szM9vdS4dVZBPx7hnqWYe3Bo
uuOJ7W5grtujBciDhdjJONDfKq+kgyhWeM8v37HPR3EvYxNgPX/mWJlwzxVPYXSJ
VwTznjXHNORHtdYnJJkQA5hidSuQRxgsacYDIUYhSP/r7aXifFGnavxDbTPXyW7f
FQkF4XXzUFpFhnzRD+O4bb/1UGy+HAn2qQdtvn2WHiwezkSNgchW9dcN4wYfvaIZ
HjRyMZM7nSg7m2TtlBP50KWcI8n9Q3VeGkP8TFLemquwr/62SnrG/mJ4h6yDD/hr
MUmaOrDLmqxb46bPCT0hNNMcszg8/Cwxerd0GmC5zgC7MdKun/NbiFk3eAX7zh3K
99nJuGH4N6YkbXgkEbjMJS3KCaiXcqVbdriMGaSiGzbRoVQjxpUBejILq3xLKluv
HEjOmjfSqOdbyBy5+4qzDUHMHOfcM1yZIVFuCxLdCy4U2/2uEvvwwzNdGwiat8XH
STZSfCRrsMMPnRRsKojZpQu+ypLw7WVI6zwMKabkJRjuJRrL29cZblEHoOtetyXU
aizwT25ZuU//Z0hFJrwmWGgKY7uCIrlyyy4/jvRUQBpwGzjH/DSf1RPv6ZPt9D+O
AKP9DChTNkvEDZTDevzA75NiDBh0370MSvnXXPxaW/Ok0zBCWEMFPo8/OkW++Wc0
+2Qz2mdeSOvKW4Wf46t3xTBYNuc13Bp1cbds9Z4oN8vxQuAMqpZPvmcWz1MlbMB3
QKo8BRGXX3U+0a1ZdGViuOpRHRy55GB8lZVMJrjv4bTfO1P0m/jUMMXzhwwC9JKv
sUo4wCx+tvnHiwKY3IOEF8UM7hB81rsHJN+rykoWM8mY8ByLl1auGhb9PIUYhuCT
+oqaXh1he3B4NatknBHVEuZ7xDOfILQiRiDC6o61bVeCc1nLMKcsb5Je7KoSYu9B
aamSyXo0bi3J++kV4EdMFDVV7AJO6hrbLYoFVdE5CO6YjaDCXxaCZasXaI5GWSwI
xIbWGCBLnDF/79UgnHkmVAzmpvuq9ijZSaxJNOAiNvdrHnY1ZUBBzUIFbQWt1P8n
bZft2KLKmkQibbllFF0RVzYrAdD4f+2nbQ/4SaTXwJfWicxTB4dk0ZY21IduCaLt
s2dSBPzxTucxiF0rQ0O+VqDe6z1m0DmM2tnoL1MQXnSRCuU2DFQt61zTKIJasbQm
tBk2YnGWoNGbrEFM+ioUr5XDV/zyWHnbY5q3YO1YeLurVrAk66RyGorknkaAh6bH
LAlSAMLeVAi+QpNQwMvVSxI6GcDQ/67x88sPI+GLHuQDVJPGyI43+np8fW9t+CFK
MXzD6O/UnXGTi5Vhkb8GF2Tzz10SQDtkkDkryDfCJvADkUi7FLAnVtVbTzSQUokl
ag4K69d/PSCereI1F6jZbYdyXl1vXNCS5iC88K0cxQOQ3+dAht4vcffbDxrk9vqv
Cnyta6JD3d1RWseDaehYEgUe4bTLnIzsrKaODhJwMnzYi3UYKihshHwie/d2ur2k
2j7ATb0NRRceZn+fCR5zgJYUINKqsbV1BtzHdOD5vrUVBbjepYlVEJAob+1CULJs
uFXrIpdAN/67j7XFr3Kvc2g1Ti+ue7MpbRlawfN/wlxyI1tfr70+eJ08TjI1ToEm
Lyjfa/coD7AJTHQu+FGdYQqL5LA6A9hcKxyORJj8nwYWYS0lkmd8xhrsVQl5C/zG
FP6b7JUUzEkaJLAdpHaGgXsXmVjsFskag3sZ1PIfYjbNO6m+Oh/WQiSt+HnxTbrL
3+amk1EhvYkGmr4PUSO21+0RMEC7jGgcx1Ktb7vdalbKHps29DedIX5TDLy3Zqg4
dnDACOoMHsifuTN4l5iViFSgWCma8HCYF/1FuVWgWt++LSh6qQzc58VC1FNPQkde
kMiw/tzAsRlxi8YIWL2Pz1L4v+7BUm09/hoe4j2iHkOL8t58V2d0TOp+5It+P+50
mm5UjtKb/YIe3yxQtgwLUhGMh/yEJDgqbPumY4FGI/0XDmkYPxxUiHrhUK5U9e1U
UAL2+Osdr4Gx1NPMizzb4Sc2AmVC+UDwS2gAVHROo9rHaNIX/wvlXHJVUwvSu3Vf
yte9HyPCSVJcBW3/F/BF4+RBrI2P53TtklCHrnqezug7qkbFDJGUE3CVykPZdetp
rXGUpcdVHT1wkMu89Qd5iWIT/lpdnB1fkVi7VRrRPNBc357xmChIcubGZqFyugBQ
kggJmQWfya77Lcyv0rdyrijFNGqC35rIJ9T0CSxSfF37cAhCGrCN+6hsDU5anQMa
QRk2FAAmn4Z5wzahGi/pxnI8weMN+oU3HrqBblxsY4ahndr3J5EGdK5nf1cOuH+U
ANZ9NdYEZzzmzOUhBp1oIwv/SIpJbNKGKgm9Qivw1gj8w5GyIztrnmZcFE9iHxpS
GfJVOI6MNT1f1PutQs7XdEO0DwE2kh4Fq38HtT5rnID0bpriQtBKRU8RcF9s9ceS
xPP30yR0FHplllYou/tmekR1B65YwiGSLMLqbedWJ2Zv7ey2n79QwTcGfSBY3kVZ
D2FZrRKCxasdazB0YRRlPn+KbyDZoSrHIid3RQ1C7LNOnszrTY9kHbhPeVkfqQ14
Mvsm6z/AA50POJfMPwDwh6NYvXWdsPM71zsB9bjFIxzu17TVfwEAZMNfTS15XzuM
OLqziODeEdOfs8vr/rOmsAlH8/g+spWTcVK48xT8cUix3IVn+VzcV8Y9qLcF4LIv
uLIH5IzshKA9EvmS8CSd0UnC/4rrhiRSrBrASkgQWdZ03cm2ez+13I3tUMn7l4za
Z5IdRuAiSd1aCc3NKINGpo5UZfCWshp0DjH9CzbSW5kC+iyp86K+v5rWiAHbNSmc
sRLLwyJshmtZVjvhveWrrKi8tV0WPsQlJQdO/F3yrKoB9JEhbW+3QvJZhliMf26E
4YuEsumuIywA4kCsjg2tBAsJrh8m+/vIg0qOp9HKqG5WFrBuK3A8TUocDxzvSCtX
754NBLl0aFUX2IKOZiVQcFmEqbwVjKrvwvtWCfyXtGbuF4FEts7X9OrRyX5FSjt0
zzwGvDAdzJCdHMqOakkRapfykDddqr9nUG3GFvNBjG6Rokeq/rbQ6/G4cmcm4BhC
JUGUA2AVhTyiil9YqOx8ZNSCNNolwyLjer0p+KAaQlm0yd2UXJPZU6RH4ymj9czy
vAT0RorTjEcyPkYci8waR9hfphnBmtU9PUm9lwJ4cswubZ0mGO9eGWCbDDnhzcL+
OF0VLKAdzqXy9Ey00NfEMYBad4ZfU7W0RlysH04jTy22SnnrtRAvj14jCT8dbIQV
NEL0o0J26rfOjn27s2bTx5HCABfYy51l/Nw3X8yHjgzffOOW3VFij9O9qP9d5xdY
MLD6a1I83ngW8GBpsaNF6UJCeHsGCfzkRg/NCnBj3WTRMFvaN3s14Jr4H8q+ww1c
nLWEdaazd+iKP8vADGlhrxqlgd1XJt3JCi31t8lPyIyylfyvDnJ7igmqCvBoSVDW
pNkBBjXK22lzxsRLIkPm/F33+vSMYveuCpYSOOU+BTtAfvrWwSa3TLXcOpLj8dEY
/tnYwIt06iYQW5eEzkxoMiPfuDC10lL9RpKdNw7ttA2RfxAffW2tEfqflAqlPZnh
ovs3erHHtd1+dR9h0cviBXxx02evCs5Rc7W83pJkRRw1erjfaXirU5lc5JE+hckg
fZczEXHs0UubiJzBlZMO5MCqwcVZHZEOrjua4Cj2yvuXfTaEXH7f5sEjy2PXwzyq
XYEil0lg5ap99IId5sD7mQtjyVdhAR6LsCcqNTaZCmwcxV8R40jKVLgExmbH1FkF
NbKU7jrZLGvieMMFI3uNZOzkriwU0wN3PDZIfwdDhBTwpB2NOorvCLRqX4FLigwU
S5cs20HHjz4FY+mRXoaf7o+2Vn4fCbi7KFrsrua797u7ufgwMbv2XwgkqS3IcrPL
Xm5TONetyo+cEJZbOAupYwFPKEr8z2zJNzvLW36ZTIx2Dz4UCpnMVR+dEOIdE541
xC2z7394yuWaf/Dn2QJJWLLkDrNdnwphLBLn/NCkehQ8CoVJZCZdinAGnijzP25l
wRZQVgOf4HPt5QkmR8sUkwUYB37KR5JkpgJ7S0PGvnoyTnFCSlEtOt6tpIz2Gg4f
J1zPsddF0fqS0HJ1hoOEzoE0r8qlzBIZMtnu1s5AYYxvJuo36JZoLs7TnC0fRiE/
5u1ow2Lp9xWuwkvwMbDIdh089BzSBxO+xoFrU2WAGbxac9JDUzOf1KxEdhqcVSeP
yd0cTQd8TWbso6Zp69BkQ4AkCIGUOgzJbHxugkVmXYLbx39Zkz4wCc2mdSbSIoO5
/kk3w0VHDOFnPh6Zrb/BiNoxrll6R1/sO0u0FHXK6Auct+Q0Hb+O+5mgtfDf6GqH
266h1ZP1eeViYoGIUltWodhVwridfsdVgpifQTdIjwDp6d06kmFadBFNnY1CUAIe
sbw1aTX//Ua+rNUdomAiDdssDBgQXFoBl2/6x2lYAxWg5DrRTPRp605nnSjDmr3Z
9rXJDbRnJnywJPS6H7qm0ROx63Ch1NyRCPtZlYbqwmAuW2YEj9LrCjKeGG+yGWAQ
ltQsXhGmag37lPAHGRneu4t+4n6e8m9udtPv0s6tjfD8ITWjwXRuqsO/hWSjfxMt
4SFSTjDFkbyVv6tXA0/DuzlWDQpHCKJ5r/1/wWR5cYTkXPMDJUhp+zJU6aXKjiud
81cNdMnrZYbWDhZkr4vDcaSJ56gs+g8LsHO3fFL43NXID7V8Qb/ZUrHZBTDP6oIp
4nfFXX+qykYPUQ04tZKbzdF0QB2eGcrZoXYwWuDg/YkUWVNwIHDCVm5DnuifIAeW
w98xL9IJzFQHyTjMzJbGLB/g90B7hbBKDR1auAyV3u7RzRUh9u9TrkmmWyMr/5FV
FThoXwIViksZ67HCLY6/6VwVwwO+RVa0NS25No4sNrHKhVZPCO5np4L9i1AST6B6
4Nb4f8eBrRIuvhhs/KS9CuznjZuhkG5R8cRlC9RdzpQX4pbqLfCDb7OPxoST5bX5
AzmKlhocWr3SS6FMcOzQ/KJAojQnPtupBSdOS10dfimkC/33/tXjXDSjrBTtFDlu
m9E/DNOVP6icYUMVyZ2Z0vYSCFKVNVfvF/APTYzKKlPbTHfkURDd8NwuPWeIHaQ8
9BfnXm/vMeGhsVzTk0XeCxLqYVItoveeqze5lsv/ck02sOkSBV0b5RelEElQx8fe
gFi0e/QqZW9lteuz+j8Vl9258FnIgnAIWyNd2hS9xLGF7UtcdxxQsdtitddPwQE/
SNNEWviozFv1G6YxZ4JoESHMnVND3b4LQl4cHsZeDRoRYB9QYTHskiumMjG8yTt8
Efaiu5TGExiIAO9IaipjHYzRF/qY2sP/UNcBdlJioPfyk8CHcU0AP00fEr2oDKpI
6Essg2Q/7PCfywlsblPlBeN+CdtL8/nFngk15P+zDomjZGdJNMkYksVFKGJkAB5y
qXO6vS+yGQY7ksqSpu0n6nr7HXIkJzC1DsK0DtqHX8uOGYzfx3dwj5kNiffzf8iw
Iw33cz8yzpTJmLk/Id3WTJnfZdg0agF8LISKCg1veAjQS7/2/TJxbOBaeU1xvnbA
74YUVhxMcu2gGBAeJNJK11b9VxeVPgM9P5AqbGb4w5kSSp8iwkfSt6WdTtT9L60h
e3fJs531hHI8pH5oEDA58Nxo1DzdyE97VYv4HjFCuvE3n1FL1oNI92NAn2EQIeBU
rRda8UkKvIwOTZy1ol4XSWYbq36XuLUVNrdlNLXQSvc1NJ1Le3KRmp0gIbyMGH8n
oLKkQx5SCGKt7c1hfN5z7RyTKJJG1MYx0iwUG1Jp4N+HjLR1VlXLLmVNSyQDX4tv
ixxaq5gYIowQRGIGjq3ZKIhjRie36M1zJsrGV/+wycrLoya1yBRw5ng+tuJAn1Zp
fV5KM9pjGuhtBScBpR2/GV5Oa0YwBevAv0JisDjRuSK8fcB5UBP7jy8kUCTn9eVF
OyZbzONnrblERrxtdogy4t2oqt+vG6bSCA3UyFeh7MFFV+DcY1Wxr7f2vphZZ2pm
wuNO+lnFAeN/hp0/1Qcpq6RkEqxpLE0e2CFrymbJHyQtFtKyg8Ha4KH6D+DxDCkm
fMruYymhiO5YAg/g5pUL4KJVxXN7/WzxZNQ06RQxu74y+ahWU9bQpCof1NVpbGaU
cws5KNK/QuF+XvZnkUhsVL+JsxEPSq8STNDaYEGQOaxsIIBww+DyVwjbsWT/CrZf
MsUivQESiqCDug7q2inPslGCB8aKiLdRVR5KFr/dW/dRjEPPklDClq9TDYD9tQFA
deQVkc6HZ1Do2QiQwI9sBc/KI7ey1enqhojR2NLX6nA+og98n2q98OgEbR8Bih4I
K/Ml2xIWeQqlVguG3XYIEzWsFj4A7juC+v5DxtSk4ACIh5rhfJ0/rm0ZeVDXHaFs
fymKBm+2ZEtgIBxqsAN8feYlj7hukXxS9loVJ/YWH2k8+SlURgas93DIldbmBoDc
Yv/Iu5W94Vz4Ch0hjRLrbAwNBxHXjVNxJB55wWegeb2NYYFdg+bcGqpmg/71F3XO
oGYeVq4iVByqXhm7kfSld9W4W5eGX7oIPKBgcDnaf62V9yecSNZaS32FFv5JEFJA
cIcaS3FyQ/VJ/IjSdKsMGdgLlSRe4d0H6LyEOOHczf2Z4GY/+zmdpb1cBQf8ynVB
yyXy0yuWUg9L7bzMg/GthpVNFNfTlI26Tg9Pg1aCu/3oSqMLOn1lQBfA8JholdCz
gxCbOZbISdO+oLEGWlQfLdIWhuxF9A+3vFpWBLkvxdtQBlWwSzZ8rFCBQ3YrD1pp
WgJ0BHUnYykJI4OjXvWfp5ofEvEjmjzcC0lyc0+9mhDvoaNZKuXQVlNDBaCy2idi
cfUwAyxRJX8RUTox2ECqMBP2qvNjfN6+jodbZ6/V8DB6tfm2zdqirZFYZ5lfbV84
1WnBVlP3dgycIKgHQe5vOE4ELm+4PWhEc9Nlxjtr9KkQXJvxfoI9OkZNfIBJv/er
mYm2sSmwgY62fdYHgCCegIv0/dI5LMMsQGK0Xn9o+1DfdqXqeDkfNVoQjgyFjSpy
N1My6GwEQl+n2XR8051QLJtLhu7us6lyNjBtIFof8Vsv8UKlZDCcYn2Ec4IjdZ5w
OBPznxCpsK7LOPFsWZ5QUTDTektnpeT4XE0nBM+qh3qxvUgn5mhd5thqQFFLTqcd
1fNHJP5agfpYM8Hk0pDuTnRQRUemGHj+xyaBSQ4kJLOyjhpTytNvy4+EpkEK9zoq
UGwdfTpr1WfMpILlhegTmGbILd3FkmDjfKnuC3HmopTJGjBFFXiFfc0Sh8BRCrnb
pMQsm3VS6Yoo1Czx+HgHJDakFZsJdQXsWua/1gu//9AE/IsRhaST7ugsKgIpJe1O
oiH4vUmRj1+wsonZUJjlnvSEhNsktu5Ke78+CZgX1HuTwpBZrCbNw/MrN/mYfehk
LEw84SgyOrIYBtdTmXirGDgZWyUUNeIGwcHeBMhmdTlKiE9t1F8cs/NG6bPk0GEw
vID247R5dV2J9XZEsLQkAFPmQbj8ZseXGYnpzo6nnRjPKzBN7RsrpWu7yBZOwY1C
egMK+FWefgD8fLHADbmKjCqDC3TToNZRS2BfYxnvJzZTraK+zt7YBwBbd+krOL/8
a7Uf+rYmGOizIAn1trrYQgvYxsJi1FSx9cMT1M4mXSrKsCptrbDa/611GqB1KaaW
toHf1eUSbKm/pXAk8IbI4tCL3IyO09nP446QjLh5gHiw6SslBXzTkE0o+Z+dcv5v
+im1v6ug+7wmtG+Y9GNTLQAZRz8o/meGz8eoyDP1m1uMe8XkX6BzAUsj0JtestyP
8mFqznJPL2ENu2kChqER9dP2AhK1EQ3rE4zoFtwV6KCArvxuGrEsECRUDcP1zKQg
nVJ5m0bG1jWXWSCggkMl9CO7ukk4NrnjTlI1LFRzIzDdJ2rXnFXjrJuNkIRffvik
lVn8xxpiVvb6xqL4+APWbot2q9MqzOyZ2p8hvIva24xIc901GjxJmUvsWUezvmng
gT3ZCDpjyxWHraB3+/w9xn1TEMtiT5e7lnLuL+f+x1+lrihRkRxBAtbwUYOKEmZ6
lW0+7bS+J8E5dW9X2fzZ85h1uxAvVMmtPEyUkFxEm0HG+udiNLMg2yI4aBphLhwb
uSVQLZbnvdygdCk/amr9pLsd4Zd8PU4WpqIwiL+edB9a0aAmV7qhLB3HwtlqABh1
mOSP0nTyVNMm76tHShnlM26wsRa2m2btPyAEbuUXWtCACqmLvaZA4cM8Ao+/3XI8
PJ63GEGA0u7s4kHYGrKyZwmZfF61WHtKiMrUxd4+ps7dQflAVDpvA/yESjINkkUB
AQhZ9VcgPJFnw0fkpMRwPZL0bWUKUoPXo0p4EO1bzID3msP1zMWTax1ATKhcQcm4
tUSfh+ZEG44gXuh14a/c9WoFvLYu4i1I2XOHiGWoTR5Ih3oIpJ7CwKPWe15U/f+c
y5HqSpaJv3nlukVgnMkm6KysLYPUWtldvEsN9rVT4WHOnel7L3GE5faMRpO06ZJE
+x0pth5a5xAMKOYoLNsgWDLAD7mR7uEM3Kl7ma3Izd2Y3IVo3BEJqyhD30OUtK0p
jHA1T4Lm5THqEziYDsbVOLLhdbL2ZU3DvVxt2kiUDCClQKla62s+m6i3c4gXe0+X
o2WZO64gvfvAL7lmh9715ApZFaCttKf2sx56ZLdH2mI3EhzHiW/iIBKn8Dks32F5
k4ipBEze0O4JomUvnu2NHB3l2RroTlHPopvVEYtvThaiepd4HyatwwShbebJRmXd
H91oCIFUFPKdzOYcWXitrWNzkLLZWPqxYSlOA7dtqkZrHi+MszL7Y27Domf8/zFm
FWNwdSkWtFal6ikFrRYthbrUjwPGzjl5TJC59/FvVubYWLFRMeVkn2HJqIGK4Blf
j9XyOcQ2LcusZLbtEQRlAaiLyEHzDOkHdceEpoP0YtRitrLLOs/FyCnxwtX9wiQi
tjnRf7KJA2jSYtbC/pBTujoiXpxNe/9FR59A5EhoVSCQaNHt3yDwBtUoKf8AjopZ
B5qUg/m+tqkcKsm6mDRC/croL+onrTCFBDgR10WsCaTPP2dGOBKP5ENO0ptQNb4p
7VAYZ7oLJJyhPu4E32NACKPJepjRLLN5vf3/4SjtwUMeIP8EbThPVDGcbBiN9H6g
Go4BE/Y420fypeeaASoAR7Bz2RJXvHmpC4tx58lbrTu0GLf08xLdLdt+isb/gbiz
aehyIua/STHSDFLstDdVVVy+yYZNk9U+HLyvqmw8US4X4Ehy2fiZSvSKbLX0YSTQ
J8g0e3KHS1Xrm1pPwEc+RdZIcPkPWQNPDh5vs0/Uw7QW8Yce2Di/yjrlte73J784
7gIbhTpAq8canyriQtwsmfqZSfm9wqI6InuU16XvBSzjwlPHVA90rdusMLFLUXh9
l4H6OthvTuzNS+C7bqv5CttaRPGDvoyXu0V+I9HZnB4+gNbKaUlWyo6fiAlVQpx0
/OF5K2oQzHHYL3a92jQb6/5/u/OxEBM+PxbaqrLS3/ReaFP78GIiOdSnrdpDJrCi
MXy0PPpNBR/pRqCyNTfVxVw2PUeg2N4GSAnNVDji63Z2bXlee/Vkg1jPjWhH5HvH
LICQtjAzTv+qBqzvvMNfRr1gQjXxzxNlovprTDq5ODqBR/f+Za1ksHK9ojAB/btS
tfnkzeWENJ4s2wuZpZ5m1urhBZxMQjgC8r1CdatLE2fUp9lZ63K26Ew9xSHAQVVo
zNfMsLq4Advsp3SpE0zZXg9t4ZfQzIUZPtWHrN6gJjp4E1cFrqBIns+vSKlZ6wfa
5Zpr7vCNTCeeaF2WLzpNBifufCjhNxkgsi5eT44AKDdekwfMpZFES522l4DG06zF
1EOGMejRrUdHPBKd0ivz7MMlBJlBkqinr3jxXaEbGF83qaJiDJHJAMkigL1Hi60E
OtAW/+mpOj9KUHIo8Mm+9sVZmhz/4SDk1qonV3KqSQ/Hbl2si3EC/D2CdWVVL6z8
INAoMGuj02lzvDq6ICHI8Ly6g11kfGHhbwXfnyemBtQT1FO2T1l6+/KLQudRwFNr
pi0mx1wQOhY9SMHutQXEiAo6cCBOu5nJLhJOJD1f3LDX7MNU2XR6D5tbtvfPoE2u
joljvxb9b5RXG5aksUPqRMGit+arQ1lgcuAZKyJPx6OlrVvOQ3KWS4CsfIEwDy1n
+pYne4jEAAYbnX9BKPcE/3z2RIdPV/WphVRag0Cu6cIcd0nUIp8Qw+sknLPxnXuc
/ABcATZM2/OfstkgsU5uAzbVlgLpm5Hnh++ce59r9lZPBTxEsqfrAh9EOTC4Poj2
ttbdKzhEhK7Edmu+Kkv/MbgwUcYBF8H06+jntVDTFpBSwr2SuxKzqcwookRWj2w3
434v+PDekiJte6nDi6j+ang1SJHgoWCNM/yrPzt0kN8fpvpKCfig/1s6uwR2QHp1
a9VMBwKExQe5htM4XTzk5h6PPRqTJLI7nflqyhLExR9KgeeyS8+P8nA7Ao9aa2zt
foQpGxE5tRDQisTH6uVp1yX8K5tXuIpzreR4cCSihpAA+eZKkGzcF8wjsq1nHENX
MRj1a3z8AKRAIFfTjUSaloZggcTmexp+5JrUXm0nUrgeaQYNLIW3pWnKnwGuzlyX
OJSaCfRXuBwR4RXGFSlDtcdTEiNXLirEwdmdUIAq2wNFjbI54U9bXxiuLqJG4c/A
FjTDVEodQlF/bISAaUgn9/V1cS72CuIPe2peBEuHA4KbyQJ29P1SHNfXhl+BnKXB
TvZru93qZ07YOL58rG5EyR3jdvPuTmVagshbjRGPp2dNUMLeaQlfflSQHLUq5zDh
h7STpqCFjVx+bA7tGACafgLQVoHEo774Z4Bi7PFT6iL0ykFofLka2WyXKwGo9j+z
xF988t4orz5YeCGYxflrx/E681n9ChVDmRWICBdJY9ty3/e7aSN3gB8ZHPq8hOCt
cW7v8S91LR5rsgL4yayTOrAl4DATYpXkgRRM4jlOSpthST8go1LwIrGKe3zUUq4M
ZETxFA/jJnXRk2gSk4yoWVK+GpZnGmrLf9RfRI6jGT6R6qUUGwt5syidMiNypPym
qpYQBsMFrrJjevEov+8V571AnCDeY3feZaT8R23v5W6Id2Atck+x/Wl0vKgEPxak
GkOqCoshJweJIOJTn4UAjk9OBxN7cW9cLHnRcW72a4LaXCaomcJg46c0ppoRYwqV
thJ48BSW4eGjkJ2PkHq+8wqtW+odlYX21+ePD300eBQFFJJpnykbBSp2jDwJPA1c
p/BPx/c/SnnSKKBZdU+J8QGqOR2xl4Y2KBl8IeT3vEt57619h1aOxdvF+05P67wC
xmmReYhlxv0D/wfF8IlpK3YC+dciZ3PO3NTgm48UWwxxb8n3RytgwujfoJ2MDIVy
yqz8JEFJQK1Drfi567+NnDcQZOUpY6miTgv/HhAYo4MlpsVH/mT/9Rwaa873FjiY
CkQk7lI+s1P6IHl7rUU/cgDaHTqbdL3fVDmcX4Fx1g+UswIS25ndTxqdX/Q4wVb1
uIUhEvTXjY9bypjp/eTxUxdzmbpI14JJbuORUXU4ENiIsfCI4cQwInbFcVzt+8Fi
79Zce7Yr8AUIEqocOZbtmB5Q689BGSwdAOLg/27qJHIEfpiJH4XUpbK9oz3crThb
dxzpeDji3TmoM45XaAJNQM7issvX3t8H9CwMdHHxUn8fHqd1cMx+vG5oWrSImjK2
j94l9TUV1iq+flLZesPgg8ceTPp/qjuNQ+cMrQltAsNXW4IXxMXqewA09He3a1Qu
S6SqQdvxcV2cobBYx5xo8aCL6ctFpIn3paga3mhOqMP+jdbQQx1cPU3hrRtGsYO4
Dv/8G9z2+CP46oht1UwOJE0WYKpSU5sJ4Tdctp6/cjfhxSPSejZ431kSOdaXeFed
btxVx3euwJ+ixf4hZwTDn3ihEVpvfZ0qBYjB3nrxRTf8bM+/YvakSwMrijshpIDJ
A8YPgN3Ra1lXJs4VVnW9VHkwr8BE6XTW3NAySGfiqUme1YZkz+2qBdplQHXvkGZM
0DkD1dGrcNWzoEEJn5WcxsD6/Fv8reToMKuqBlS8lEkr2AVAYsbTay+LsY0H/gM7
TB8rMz/Ipmw5RfHWs+igb35fDCtHQRiIoPCf4j7VDL88IJvs1+vej1tJTDeg2a/g
YGLck/9D043VZx4CvW6m0GXs+lWAmj8a1UcQ2Bfmfr++A8ES6DBJkQbp8EUcuZCw
0iKM4mbfLFwnDGzhvqc4wxUSeaoeKBqbZy0GUmjRPhFvjl8psaND4BYBLDR53Dep
w1rGPORQDDe3lFuWetAg0NA/W1XSQDWqHnFaDwzUQEhlfe8Is9m43LV2UBMI8nyy
NJb2H3l68ul7DLc4rgxBNFHUMsraMRbIiroL/ViC96ztJUVVFelFzq7UqOBok3Za
KojXD8ViMYePqovUJhGCAzN0hgwgOUQ/ZAT/ZcJvuzbxi45X5OBh4sara7JWH68G
EIAGgpmL7xIx8OW0eis1LeYsKTrSKwwg4CLT4XpQmHP31ao2PzcbV/l6jWlvSWUK
ux1E4gbwVzeIlRMzhz9KCh3XW6uAa+zwPS9fEqqQjxXb1ZI0XxM/J+ypq3FUGmpt
mdKk0ftapdlCMp8HDE2dX12hvN20d604Zhpcdbugia2FmbuHVOiMPuvm0u2DrKq8
k3vwpsBqh3lv9svydQu9HuTjVmFdgiW9tXr4LUeSYIWueLNxxkubwFqlrJTT5nay
c0Lm00MbnVVLaBKAT2DbKOWYZ1wsQmuM6irQH5kHdJQssb5hKbqFkP3uMIJvzf44
tegpRzoRBulbHXs/i0Aea9K7+KUsitwOjTHIOO2yqRYFhoQf9c3VC3OMFLg6bIgJ
sI4FmAzY1T2OLDO7SS8hEWOLKwunFLYLUnzwEOI5KnU7/W7BzNpY8kWyBnXU0NQg
tJb0qHUvKg8hbVMBQ39dEZ7M5Laxckx6Pucqe7/JeyyGiRgC4+FdN19jOXym7IsD
Ksf7rbv7MRfTCw5YdW/FYAn8P2P7mXT1rvvAaHV8L0ZID+ZHv9vTHY9n1YPN6t75
T35vHiIi/u4Fm7/VThCLjUt7ti8j7lJTq300K35p7pWMWBGLcKRM0FK7IKCRTLBw
CJJDoTtYI/WY2u8gcvY3eg3z9cFC5HTf97767ARdLuL6Vv1ZEWKE4/RAmBx2FcE+
s4qETlkWG0+lq3SRPqn3vcc+6Un4zOVAyS8AeovEoe7uXN0wWmv4Y4x1+CgAx6wS
STkNrtgC1MHUA33YoIqdmir1qUrWGmq1fV3PvamA3Ma6lgTqgXSr/6vFWMGkyVM/
mGZ9+n/aJoZcyw4pbDSB+7eHHBwV7W69ikC9ZJ9HGz7H0C7d9wL4nhT8dE6yNJBO
N7BFhNNrMgefCygjPj+5rrHOM5HKSovS2fgmR94GacTK+ulbTdoE1kYDxEZ8mQZ2
wH//GSW8OHToDFWY3a+u01F4RRB7MuZfsiiMs7ekyKQ60bUcnFmwFitJJYt76W2D
fVJMZ7mIXtpKj3FEAU/gfF8xQ/GdE7HFHYxWbThucAaCRzujF0DAQplO+heWhONg
3eoWHuPU7LysrX/C9zUbM4o2wgMxIq708VTPzqgs6cQhcf+5Ou3JSNvIHgUZhPBw
YW96llVqurdA1Ww7tQpVx5TbjxLYQPzJPWtTG83PAsmQSLI5yXEWXsCMbHg0DB/P
K7X59LgJbTk1XjhD11kcK4tfTdiCdGJ6YZyHxHnACuh+Hxr8zzeDrrOi/D46PGI4
aDH38ynjIXhODVJVC/q0BiaElol76MF0UIUqc8Jrr900/ammncCWBBrpr9mwuJeV
WnISg5akD3AouzIiNUaT5YzdP1ErR5JTFq0oCkmDHWhvthskwb2gcfXBG/OPw4ve
V0cyklLcT2uJRWJ4/G8hf39beL/qzxtsYvNaKap3eVUAWY/9rrIZ9bSi5QATZgWc
3hgCSEHQ+/aRIObueMMHnFO1TMaazXHX5xzfv7QnGk2lXqZYmj2mgDx7OsjCxFZX
OaioRMmNELObo8l4QHVUx1/IxL6K20So6ooWT6HQ5v3dFOc6KgMeXHfp2oZo0+Co
sJyOAFAm0JGaYSxrukE874kv3oT2lX7sLYJ4mIHE9DK2vuFWCqiDfKZWc+EXkTZf
fTZbj3pf071aIdXxWx7LGQyO+CpIj4lggBclp369Gif9zDBjfCrR0F9HifJ6wI/X
OdBypyKHCi5sPCYxcifjYeC+zjLb8Lf5ro0SSpCopwMmM7bF0utO0AgllwdP9ifW
TYur2iIvaRV6KZ14IP8qL7vMSOiacFfNxv3vD0cmj7ndNA7VMrtZD8fpdPkGszCl
SAKYEEnQGfPoDv7MfJGWL776Spg2f8E4O7pmsP9ZXVMWcVeZlLGfDi47QxdLX1EF
XzRa6OdJkto9WmBpJ2X86wb4R0GH0Ejx4fUV5kUOfU9qjvhfjJiOgwuSVjQ6HEwD
v8xQIKZMN+jyUYrMu8iMeBeNhNfdf0OHrPG8rvkd7LcObTUNx1Q48kUJiVGd8wqX
XesUQxKzZ7bDaCRxzm9oRZm1kDwqk0+bgv0VzVpWwDzGknmjQt/qnXE+YOpjkw32
Vzn286FN+OsmmTgBTq1ICMVwFHyL2MQQVQnfF7072SxZaZmwnwAQXr0PcXAKRqbk
tJSS3zJ9xa0U8ij19BVZOquoY5YsuR1McPaFhHJrKRkSoU4d3d94RUjfieePcr9p
CFwxgJ00clWuWIaIcdlwmSu/m4VJbH/NBelW7/uxDWltivZur5QBVc/0YfzKi3AK
yjC4lLUFES2yipNSWh7hKLNgnfnScCJtw2ViphkUyn9RZ6+D76BiA0BTzq/LLoB8
Uvql1CWN0fkqnLoV/nUbtGLCsS4cHWCYi2guNLOqVQWDjBHoFofopJrCjcRwhmHZ
2qGhHnGiZMtkskjbyD/qY9JuIQIMzsyr/sqVrcJaYFmxMp7SgBZwDIcmoinC58Rw
vS5QzRkI8x+9PF5ANwg/r8wUm3rUG+fHnXo8cCjiVaABRsxHs96T9RPKUFISyS0j
6iOyvJFkNy+X8ygZ/rkZMnDuSMiLEQWldHlja1eKr6o9xQcoi/NqR6XIDOMEyQ4P
uvqAG1PwCKp0kLrKk8OBSh86VefQMaI4YyI5T25OJaZwOVuvNS43JVFwHNjWrQJS
W1q9e5KWgByc/LRcb+zSBtgzwmZiOoyyA/wE7WnO5X5IaPGdHNLKtqTLMnvn6CL1
miaF+Tl46RmeCOEPsMxIh+VAilC8w5+f2yrhWoaENHKmEbVjt7upcSSuaLhriO4G
in0zgR9JiU/L9f2bm1sVGuGndo5qXLG0WXkzE9nuGmf/xlBISnemP24xscoJ+IFs
NZR7YxM34KDTcMDXWPF3/KwcQ1PlyeCcUkVRe7IyjEFBktOOk81bAKGDggBlvAPF
3NfrUHl7yPm9bu9wLstRikh8RcnSNzYzySj0AZ6+lIm2zJZtQcISedvzB2YhUSF/
9phDewPTcb2f5c54AIrUJqfccoCHBPJT6cUfXsASQ46Aq7ZKzznd89756Rs69ies
REOu9bJT8LxxuA5f2NRy+17EhBAFiSqspMZCR1MTJCTMN4wl2g4pVWXs1nm6RP+f
nGK+FIV6JsOjteAwmlP2M1WhHxYxClAcrg/0zsff2qgziwPhtd24mkOQIE/JGmAH
Ua9dAqWYM7Qn8nSMV7GdsOHg6qQvJ4oVzdrdLVthpHzHOcPm+X0YzvojpmWBrQIp
/n/TxGwI1DtgwXPThifw0mXEhDyXyNmA0LyFLbgEzkOngdKUxoGJyvmSW2ZdZt8E
eldRUxjEZa9p4RYEyw5RWLibBBVCtOMZZE2RLG3kBsHPZgUQvn+lW6NjjUYbK2jb
u+itjXKH2cJqN2Pq251Z3u0NGoYBz6UufT2HHVMkrAAdfnRROsH60x1Ocm9wVDhM
aShC3hjxdk/d6nSSFg1fOXtebAdxxnPdnK0pzK/yxXWlTVZFpO9G4LRhOkKz3/rI
HjDPN0EF83Ya+FoeH+F9fe8czARubGGI3QVF2xMXBM/ZzRSuNR3eEqWFoOa9OSF+
6qw3JWOcO1tmbK2I74TGWJAXLyBsVbj7dsVvFjUjoeANCvoPKQH9IM3iUOssY0mG
ROkgtFiW8aTfy6zcinlg80wsrwL0ny25oStNePRmYco+8SAvjZU/IAap14QLlReI
4VWd770dXNHe8pcgQDLnraXobSatML3qkwSN2n0d36cdFL+9OUqCTIZPPt1aN/yG
lxrOT0TBnavMvcV/vd27vNA1lHgIbGNyIpW6/Rezei79B1XURlUqLUdPhTS77TDq
hVtACKblKVziJ7enzt97dsZ+jNL/APdAcFwZ6xhrktrWoDMC/pQ6kmvY0ZBm6cem
RIKCcSPgzxyfw47g6ahUmiGXKS8wSPI+lI5lHAKTSsmxlFp4mD06bv+YggFdr02f
43cA08ZRmg6hIeyow5oOPbUz8vGnutzCwymv+kYNN6WpNa6mEcZN+VICg8RRVahK
YMV6++YMi4E805k4F8sXu05Kh+QPpgzIkcYiZK0QgTre8vSfCcFEwFga0/grMMQ+
SzD+irWqEFRcMqI4MHmfIjVWMaXYOV7Ota76uIOrLMNSrytRbzIaM/55tz18qn14
eyPF0M1P/HBXWE5S+UK6CB4M30yIz5L+PUwkG794O50AB2F3AoZCz6yJhhKhtaXT
RWktn5iJzooRC11iML+r9MFBCVenMW51ooI+pXiOlkQ4BZIEWY4bH1eMP2f1TZ5O
2VDTPpdbdEIe2xDXodRwX0lAfx5IIzZkASynUoDB61D+nrhOHS9kJhWYJvzfdKIB
tkSclXbX6yLvTPWS7/Kb2gRF5QWt4exD7D1dWEf/7Db3c2BTINionod590mOEHNi
K+Jvq/CbfWaMMZQ2T5sR/wtNX1v00debwvH2soHT0FMEffstQJNLKaC1xHA2EnSa
rY9Ury7i9GYH+Z5oY/ragttv/Nxn5JscPbOVpccOFcWrB41r42fVYLszJFA8s2ci
tfvYZZpWIjaxzf/ql5F2hrl7zX+q+5oFYuC3cCX8fu8scXJgvI9ktoYnlf+4Yxiy
PDZOEeOGCAvRqmSp/Nlo9f7j0MshM7+SR+9NhIkLZINcXJJknzeBztuaDin7lHBg
qml1XKoymEE1UCYNQRm2wcY1ySxWmN/3vs7BnxHrJMF9FmZbK4/f2ASU7aD7sKmU
MUhEdSJSrmT7OAHm8+TKTmWtXz8lgLK9USPeVA2tOVaN5Q+8W9s2bE4aTLIpWEwK
xaA1ES+y7NpBP9ZaMfWfRLC/PvfUhylPd8+XLMD7C2eL9z6RZSK+Uj77FQPZfURX
8r51D8UE3niUmRdLDa1oaxGrF9i+Omwzo3iafrhjXueLNea4fQxEjwEeNcMywfxp
7jvqHMxCpAz9ZnTtArVR3dZFd/kJJcxmy5Fj2MH6jVO5j9KYci2Mo6lPT3htjU9Y
ri3qtrfUO3SWQshUt4fg+qUqcGuGUJgtv0IMQT7v+agqMqKEbJLN4pdxLj06UGnW
W4IF9sq8F+YHKnb5SGnIqsq6woeuDU9ZcI4P2nTEc61lpr5auUPAuv4JaM2f6TIe
/FTPvnnWNpryj3mpFsWygACnb2mcSF9sZcwlidTip0aQXcyLKaJv1UDrYFJh0TWl
preanaanACsgPR1Cz49gk+sZuXw83KY184b9oCa8jpugui7xMIwng/knqk3ArlSE
fUEpN+G1SItz/U0JKw/AauAoA1F1LSlv1wufqvAsDH15VZBIVqWmJ1kYOCv8xI48
KRhNAUHR5wKl18Wgyak7PFOQ9AXC6UOqO+7mGLSI5obMyFpZUYgDdpo6egcsisRv
8wCoujIbv4JQMMWE+I/0lsLTcRpFNqQQV3dycBeAoJrZ1Gnu/cltIXvD2hftJoIh
tjIRLBqtn2fKCiJq1WFrJZ4RA78zMDb1M+Wg/X9kdeUTfXJ+KfJIjomm0oEBzDBQ
DnVLGU1rQVJRDVysHv8xJf/yGTGFjL19nYnR+optXCL4HCa8pY1w2/ZZK/AZ4Vlc
qxbyHQMRYjrZ8MYgiyJP32CFKDyk8EX5s8Uig2ggS0Ur6PGZu/yyWLIlM4923YAk
NjfZnc/KqKPFC7XKPl+uYxV8QStEUp9CjrojpT+owJHYRhY4b/N26FNFG1IBxzLO
bv4Zmw0WDX+Xu+lNh3VGvn2WSVLM9ifEz33vk4VGt+LEz+584SgCa/eh5oe96e7c
QcgJANM3Fl3G+YwXa92VrY8jp30uZ98GByZxMAPuFXSgo9JLveOBxmrPY2lAtimS
HkxtQqBuXLzU4xZyDhP8X5wq/CfLtuL3fJBIfo3/oCPntESZDqI6d6KuZPqs/ede
17hdoh0GUBebzlfwXqCqRcljIORhnglB0DSWqLfP/wub7CGw1UYsePr8J86yrTEw
3muCG9peivmyVG9VC6HBMWakSFB/uzTKPYzS/tbrA+3F3LkDlInzFRkwv34hcjIi
PYCzSOzh+dXr2Bowo9IxeIvjXTDnFNM9L81WIs4snU+O9wberzoCbtNv2ToFX/LT
HMa7vNrfpFnAWB0WalmH4IBYob3YTwNsqnenCQrQeGQUAgtMnUvSLGAbroz674L7
vDG+dU2hCUIAv5rHRzVLjFLYZf9TS5eFiiKLCmLTi1lHnYIn5s8YgcQiDRIhJ6b6
kBqMZ52rlcRxxeKadivHJlU0t5l4idlkcwrTiEs0+nFZUr6/IukYN36UD7ZTbtr+
rxci2aqeFluTbPPBIZ3sogCJ9IOu3js8wR3pOXEl6anZVuadVXJldT5/Y684adIV
ykdJeFP6PXOzb8NCIwQ4/HRxDhkqLsFfHfVgGL3u/PFiWUzaZLUMI3p65QRFavQZ
6wJqxMbyFywTQGYHSCZkp1CTQFXV85FcFIzpH97rcLfUYrDExWuadd37NToIqkZi
flwpLfLmzYVfreTTL0XD6RrYKVZPEAXxzC2K4FTsCcs/lOyAfNP+Qa1Pea1kT3M+
hs0aFgHAlIe7GHS7OtjtsCD4s4Y539vXyqHQ+xUic4+DS5puu2B3Lj/35Bg/ITQZ
Y2//cXa8ndDqJQM0V9TTobWLWDEaMqGL1FcEUlUsscI6cW1j7+qiLj9i5NUZKwbK
PtnEH12UREyqp+TlLISIPbaM7U1LEXT/U0gL6R0Z4oFMB8QOq7nRcoa7w0hZlKHV
gdtZsN0CQo+BKfFDqlxBMHAdhatcz3dcFyRpnnqgwUEG3nKiOZpXbQl4x4PeP7Ad
CNoXk/G2o0q2UqgHB5lDGrh48AMAJkizJBLvf2xr4+dbqHFDrUbX/HtVRfmv3Efn
HfhPyYvFVTLOuGaZUJt9Dj9G5jH3hgdefCkqy1z/npoXKPZ0/R+ARXBzePiHpqBv
shUCjKAGCKgLkyrWCgssQ1tWVTIrvlkNajwSoeGFvTgXMvI6sradLS8Ff40trTGS
VWNqu8fy4vUnM3z7K3lXETJq1cJlO16FEVX1rFUDPiqDDwUOj/eRu1e4lmeI2nxS
7HetabgI2q2WEVTknidxmckCUYJKKD5UO3B4J6i3sK/bDv1U51k1kPzE8ZKLKfMn
e3gu60FTvdhRnLZ9U5lw+DvrQZHxc9kQKOn07OFB9jXRLml/dhJ10oK+YrZ/OHjC
c1sjp+GaYNkFZvWVvK1s0bEpzrJKd1gztYmh+O+DGjHt8OgpxKJYc7n+L1R/E6LV
rwJUkTcZmkFEKfSOHDv4DkG51A/UXgX1cpDX1pNJnZ/FXdXgA3bQkXB8QWqeH5sV
CG/pXnyKpYu+BRGTJ7zgXfUFcZqOzYPe+FZOkVU+bjIrp2OAzzBwocv/ZUc1L4ws
0JD77xm+TJpgimGlVop137vESVBGy0dzsV7NcFp7e/Yw0lem+T6X9K41Qd4iwUdX
5NBxVswmL76oncm2DdYrht5l/5hf9h66p1kZ6R14YpGujvdNFtxF6B4y83ge75/d
u6IVRuYJwk92QCZ//Xh8at2R5NzUPItbdrob3WByyw4uD8tuqZx/pPEuQdm7ZgMF
kcI25qR+sexlFCmP/qdTWkn92SJfMZkyL48FDZT/CD8+WWLzvOcq/yQ/NbRefm10
oTdCGKKcgKZSu+7qQtii1eefsq7qw4Axb9cE2rbLSwxGtfhqEURBTuWmDnp2Dh3C
3W5Fz4kwC0TgJVLOqoNX00BAKwftzaFHlWsGbbjXNDXGI4+iYnlQ5WcPsemcPRlE
v9LD5ZDL3bddvf9baTVqKcHDQ/P0Ng/E4I5urIAcn6u/nVDOkfsJFN5ARV1manRM
QzXXu5+kNVWjtbaDZHye3LMKwMq1gEZlCt9fhSJ/EGrSSyGyqzHxASY81A62eF2y
jh0UWjMXHoUZRScyutJ1Dzy9gxRLkr2+cladmjytQ2GjwlqMoDCE3r0XdGDR9Jcu
GwU39swLCuvvzV4v1IIlI1megfnXD1TzAul3i5LegI7u0PTviLESnlNw19d6m6rZ
JtDdhGSnYGQMWNlU3G6g1d+gBhsavDNmpmIm6yiJAXPX3oMQYTqMizmOisTUhzw5
jHXnHU+OiqeLNh2u0fcoV62uEVXmZyS7mEoO5yzmpVwKrOI2GQpLBHTrCtzPd/Q5
zwLM0rJk1QTPm9LvdYJg7mx1Ueof105TgIwpMiHrpxbKjIImXOXq9PvsbRkeP2SE
wr1v1WAx1pcjII6Xkos921aC2fSy/lwm1gAvZyNIvEyGvuqm1Orq6DtRJW2DnBjJ
GOqd6ke9bdaFqE9B51/ioLI3LRvVcFis4Mxu5DPCSA1N63RzICCU2M3kTJE2R89i
vg6PQiif/FdsGhCrpNfXePlpjRVzpO/FXinGX1SX+oHLOy5nvRs39fQQAwek/HUQ
mXABf6hEMxeDqB5C8kU4ib/ILroo1GLjfh5GaxmsUn3cZNUcWUY+JvuW4ZHwoC/8
cT7AabLpdPBMtl7OLrF8/j7lUteRj0uVe5dG/O6Ed1lGQfy3U3czXHUjoOfh/P6p
AR9OiyphaXY8kxblYg0YJuYNoPVTuvA2HVpkGQ7c7wcnBmU8xnH2hQZzhX/J546/
j3DIrYocCaos+vx1/vLoJOEH4xCILFCbPVtsdhwWm06xutCK1iFTYnXXnmkM+qaP
8SkBa9mVWzjdkr5MuVYbhTEJ1jkgPCq102xeU6VjSJ8VDF+o/8QtuoWBDJklW0QM
zdK/uP6i/iQMY9P/VLOnwHT+ln9XiNUSsVr1g2rPXFwUnuFqKVfjDUubfrTztdi6
b4CFGcZYZwkqZcD4OMgcNJ5xJIuKeOGlhE3+v4sB9lccCMIo3xuXGiG3h7HF7K9a
hVYqoAnlTUp2YSo8/+iPC67FRwLPsTO3zNcZluD6xCeE/3r3fb0OoZ9fvIuMjPWF
aPg9MtVskr6M1g3s+YucD71ao33Ma03Ef58gNvyVG1WTMAmp5LewiJZA36+K1OzB
EP3Tm4JBf5GeHtj/kwVHQoKLo3Bdltk1AUiCgBPoLXVTnkPNVB4b8iwXe5py+ZbU
N1IyMSNNL0WNHEp4JRaMsq0UXwu5zGVID62NwwuEF3ROtZIDRZRoYArsuL+W0ckJ
OWmoZWuUaJqP4g7is4M5U5Al79WcqK1EjNNi+DgyQgzF1II85LjPwLEnuRIUjsZk
QuWH/TlU+ZTlE3J+0CsOtyCK2hq/8NBbB3SeAcJ/390uUwaivxi++ETDPZlhmoeG
aDhpgFP++dF2SS6tYdOg/S2ctZa/pthvD2HqxM4oUvo9ezcWS9V8ozjRC1PKsJLS
dFe6xSTZeeIDnmq9tXW0hNR5Sy1liMgEau17bDurBmHHV1wXTECkYes0CQF1yVmh
VeVwvPVikqHON9PWHRxeRlbySa8vxMMvGmG6V8U1gv88jlcGC4PiiohjnNaNZWen
a7to921trDregV6PVLYaxv3tE3elpVhvJDVMTmFWvM0FhBeYrdWv4bG+pWBYNmip
+PlaIcQMgEdySB5dy/PPFqC93Ep+4s9rnmBpjXYuagD6/KAhUoksxdNCWeseIa2V
yGxI3Lj96fkBdV+tc1ys0Y8NdI/PWEzo4r6yYLRsfXqhdTVzjSFILIqu9qwpTdwL
iurm+sCqevEKM3ttT3m6DVBLbiv/MfmeAbat2UBHAM/SslXJXTZTreS41DPdKVPE
iVVWdDMfIaYMHkBLxsXBj2QC7kmi1IJjEiK8CIq79NeecANi+VLWe72nEAK1A7SR
XhRGLQUmiYFM5Icu9bRiv95wPDw2lm1GZgWxasK3jA7OjWDFsowyQPm3aX6x3lDG
BSy9sijsqfEscslnG9+fS8+9LcalwfKQ5CswhemUb/JWce2drYk6nPZie5U+c7si
cxBaOAzhLB+gi1TDp8i3zCz2maSu2oQxamMLcVkDPyxJMVM8pnt0ljiHSLRbxdYS
nUjIBLfDvCuSDKjmbqzePTCAsrjLxqaRz/rE38HQD4A17JEqHYHbUsOQMOS77mcq
gISnZtxieTb/uebAfT61aMrCVFBAV5toY4P0jgAHGLvcmRERzkG7p/Nwsa+AyQ4O
I9VHQWThJ43sojG110NjNDsqt1O5bVxdm0fM8ElFTojVjyUSLrtbrfarAP3nVaIh
4qfsnjiNSKXOZs2Lwhs9fIHbq7yvlS4weE4gQgMEExJZzEf3yP5R0pvjKyLLYUdB
2IckqFgNV0BSlQefcCLEk318Rky76GFy3jOunnHncH+uM8VVRd2lucT/WSgejRaK
4yF4vFwqbGswHs8IY6HCHXcfl65j4cAx9q4hD0mWTnGtmH/rxfHmN5pgq/29WSTQ
wll8yEzysA5gT4/ivmunFLakZYxADPUI2ETEco4rVSvyuZqpWWkIFs9nCX5fp51g
hEbu6jC/58emcthh3QHG3pwcXDIjHhXpiKCHlDKsjh+evs6hdRBMkOlD3JOOODPl
4aqOasl730SDOZHSW0Auq/OrfMfrRiVI8AVWbYIkAbk0gAByRJlluAHjpk/oGG6M
1N6HXIDyafs0rhBb3yPgXjd2eRHOGmyXJJl4f0bRZye/ecOuXk1ZMi0d9CF3R/X/
9V+mwnc5LTKoWpmrXkSSawsjUD6eHXuAlbpTBpTBk9QE7UGbJLVYRlfuGe5mEmid
Be+U4CZxdcR2MBRzsIfgp4KptRN4THPjNLsSucYJcHwWXs8DVbfoEckkvl8jW2hb
jXd0fdjuaW+QQsDJaOZ4GXwrjsm4vgU92AoH3FoK7bKsWPWAwE1ogaBCSKWSGmxy
/IjDaEIkdtNkYdrtLfOPREjFT/rlmRP9R2XmXLy4olGO6Sn+bO16Xt+gjb0re9si
L1de2lBMLACRFkVm7GahDi36YdntFpyPAfqR9B8k5UwJF8Jz3/jrnAPAVBs+Btfk
0hRwGNkiDS97elj+pFFsxn1tysFKaK5Qdstt3hOPh/ZjdDyxMvF2LDvcpnLnRLfI
flNEXX4rIrGy72RRW2yPgem5vX36enbMfTB9PQH7oAlMoHK21pmrGG3IYkycOAt5
+ffCCjIgDdNYk+2x/pB5uNE/6CV7F4KlMX07Tao90KOnhKCx07QhPL2E+skjuQ8D
agtxLJkMxj7HzrNzasLzzhVPfBVTCAYNh4XPGLOnlyCvRsiXymD75W1LhaJpE0wU
usKn5rcrZtPQaHDU7udFPANTyjDIj/FCnSwHj/rk9T3IViBnae+W5Ji2ZzEnFPgt
0H3Dq+u77mEHAiLH8+yHfeiJ/7Xh/RKvFK8RLRHv0PDE5Wc1/tNQwpvhWptj/pwV
UyUsMsI76/61vRo+aalyrqTjQldhrKMvvNICznIrx4ymrpgQTITTVhMhQrAoRPHk
Ok8RjEHrSz5CuqYrLuzpRJf00ZHrU9pcL6bsN/yizetpYIMoBmKqjKlIlrL7hLsX
d9tT1fWD7jkbmkzyvNsdlVH2fLv503kzn4DB9f0wvajO5EeiVjwud8fvgr6yN7xM
c2wrB3f58b1Ud6kclNtlCpDdZHjOpMsaQC0FvCCSl2NA13QviqcYEpTWqNuxe8+h
FZuXKeUgJcWptTeI+Hx+zqv/5HXAUKIARHdEsL9hJIDOE+901nEaM6RbY4cj9W3n
3cHQHJcFz8lqfxsVdkh2omTWt18DGS5Wo4WT9HEORz5SCff1BPfBZSZH6HLZZBDI
KNgnh5PFEza+YRtcq2vsHBeGKKp5VVqvRE48OhGYHMcRUsrlo7gEAE5fkWURd8mz
r0GFJTekhhy2U7+6C5TlnnKCNsxbPwQ41kdQfsgioJ1/VL1xOHrLfNjs/AwtfsLU
yw6V37F0Dx8QAJHZ3G1dvt+Q+E6EaGEvAubasKlGvQJBB5Rxs2GZtaNeeVL3+17d
85CLZFs2XqFg32kHfP5IhVZr3JrPWAHQWDiMwaA5hVHIqCirfCY57AeukEKI5seF
V2txF7+FegXEVW4oxnNmQPppA0c2CgtUS5125GfueMbtdQ3zVbL1+8BsIyS0R8kd
gcGtwWhqFgRN16+yxdjzGjG+Y+H7cg2GNbgoePEcQoD+7LljNULK2Ji1MdI+UMOh
9nALwA9oz8f22AKQ6aWLlyV1UhjMFf5vNr4z6o6Gu24fysyQ7yrmx3MmFmxQMNwK
+NtYd6r0FmCMBSlRcBEsfOWW2eC4a5AHTdvG/T8Rh9V/UUhdlp2s4A73ANMGJOF2
niiPhgAV9oADoKuo3tf7+p1Kho3bK6JJQSMhsNZSlM5FRn+FiTsZ790vIamyZeKq
lDXzGxS7wTk2LTmSpKKUCmjBc/QMWyn1wC1juYRzdVHy7R0/KqeTKXcJYe4HWRt6
QY46IyXoec8u17vGMflYVk8HnRmdwt0TYxmZ11u9sX7VonDx7TeMp9G7ZLKQw2c6
Vx6xqUKlDHv8q7NFHvZXRw4Wb/b2c6F1KVitdITPfdWJ3hNsny8QPYS5VtN2y3MB
lxQf12/42Y514PuvnPDPedpItg4bUaYbUFom0KXc50J30OFog5NY4YCKUhJq5FoG
CuaTrFoSLWMzBEzhHadEjMpGJtmg8cu3WMdwp+2BFogX7T+ip7jimPbha+NolLA4
NrtvwsQzeGLB7XpvVVoSVAQ5QPCgGRa1iXqoAxFV9/v7PA6pIyB65P5UOEDzH+Q4
1IOZ/Mt+h8KTxbAjnunZtk3uqJgdK+I48WbK+gTRB8EWjqRZgiwbg0zZOLm8YuKV
9zhk7Y3hCToGBZbxk/G/TD6XPLSgKSLlsSuiyWuwNkD3a43HHecK234HhtSvPuVh
D+MJBSQqcvbZ+Tiyf4oBm26sUlzjJghDQEnKwhImXVkS39GU0oyjs48Y8uhAJ6/X
nyAE61ecIh+0OG12KD9knW1zFTvTiVQZX99jth0zOuQO5q48GkH5Xv3fTcl54izF
8MZKinsyflGCuVZZkW/3aVmvKULlj0gxO1Dd4pDpnmoQHoW3V5webr0hHRHS1oCV
19JGErWrBk4M+4cItHz/o33biF/MbwsXXPnrKBj385MVCzoswpjY9oi/msNJBOuU
7QhJcrRieyxGLJkVEEXi2++K9btd0aZZVsCB4LWntYDTZrM+yGDHlmCf7sBwQyLG
6o/uRNCwcwUDkbBTK1zDAlGA0kjBAg87oHUkuJfWDY9JnH5rzcKC2FbycHlrl8Go
yW5Kix8djZMyZZpHzdsyEhh2NQRIn9JEALiKxvrUGmEnqRFxaS3PaHrIKlJnzYo2
Ck32ozNTps+aAh3mZ39EarEfwizmuXhHTnnno7NqSHjsCckGYwWGClvt3/F+dMAa
CTUbSxzO3RmgjVFuRGPktBoWEbapg1UMF6tUuoEBS+gjvcXHwVzALFWLBwVObal4
Ow9Pf1EKAI+tNhhURKOiRr/HCArQ9ghLdhK3mexV+x7G0HGEEORF4LuIZGxRMdYK
tnfMEqbwFuNBH+ndJoflvjjSSibtPwr554a6wNT8P3a75aATr10iOryf3aEir+4t
6d1SURCrvQS6sku5GgWadQdNKnOcdQ1MkwNO2g7COApS2T/ylZIJV9WSV4m8wDy5
w2E0lF2T+VQrC+2XoDHYh6tAUq8Bkowwozg0k8bJ9I95JkcnGSlbf7XteMbkFfgw
12GNt0UI4vQ9PxH6Ujdif0cPjp4T8YsCi8LbJGLYl17lrbLqnxQ1lrQAmnfYF1Bn
v9Myt0WcOc9e1SkA4ofwUauSzmhAAvV3OoyRqQAmoQNxuhDVIL/jgH0oykIdm0NP
tv6GyVRVxX4NftoWqhfcz3GSRLi6l2VvmHsEdRh7NNY+qvay5WSxTTlilgU/KeMx
KQXovgIROXy5rNcTpdkSlKUzlzA3LZIss1iRFWba7MiHuxDpcTaeK1W5NUIJGrW3
sVDD2QtkHL4SLb+fG4gBl+3B0F4RTilw21JIQoPXIRaPG9xr2EAkJ+CamApFzKM5
Mq9twGDGFq1o58osfayFyMQVvVF95LscBi/fbRVexrcwxrQ+LADuqIO24w05rfVB
7ogGQUJt4OksIIFDINIsgmy7kS6Wl6LNL2V1KcitD8BI+5arbCiSjCG5vOQpuelr
Axqm404Ca3rAxC2U6onp9/V1iAUD6AjOovnYukDjtIs+7czpEMSDH5QlUrZuuJLW
RYRuQEHqbGlVIkepk+31fFbvDabVGhTZbvnNnH8dJeVtmA6M722sXHxd/mEJIMrb
7qKan+oj66omnujDVFkjLzL5lA5H9rMC1AG53TjwOTNHcea085sotxTlXtTGnVor
d7ivNRtLqKmIirmyUe+rxZccz5Zbw1rKIcJpvyFh7L9kOAqstoWSaaQqUpkDNIBy
KjGANFl93hkJdP/61RfhngJh4S3SWyaiNeAz40Yg9pjybPc32pcU6qvxoGBvdbiP
33s/dA2dKUAu3P54pumIPER02tPTo2vlWhGYHPuVGRlVFLcGMvn58pIHFtsFh3jQ
T5/DRAyfmUdUuwRMGdqPK1YZ9yrUFDFqMToNIHlEvk1hDfhNtkjcKVWBGmtjkgcu
mQlHpbY7rx6CyFkHCDm5bFZHLDcdjHeFfPlwGdx2MA9M4giuLCQ04/LSbcG0Ih9Y
ZCOSqdhkxagHXqxHh+XoKQXruVoVze/4cUD62g+ag7yq20OQacrcB1h4Sq+fFnsL
Q0zE6J8IwuG47WbwYnCq44apRy19IryVKZ/mE1+ld8Ky+Bxu1L0ATf1h7r2sOLgf
1c8bpIj9jyaqpc+QRT+ZFym0ICzQrIVCAIC7pDDRgPcWYcGoelHkz1+b4hI3O3ah
n3CXAVJOAxKUF1cBRlzrvPUIP09JBTJuHwYpAlH8o5Gw7ponvzzwcI2QPiZuOH5i
pADVY4llHi3jIzF9lFSTVPyqKMcejrJTlaGc8vaOWa5l9KkqB1SrG63y9IcPCcX0
TAaFQFECT70HvOuzEBRTC06Bct/40O6iIJA/RC9+RTk0FXCAQUXyg779AhyES50t
ZhX4vLvcHuB/yyXU7kJupLvYjn4xNwNOLqpe82XaAvfVHbzT6kaCKHAfjSkZv/3f
H7Wn6ZPnlR/ktk5hyBkpA5UJlArG6nY+h5sXAHmtVF/ygyehVmg/yJyaLrDW4oJN
t3lEU6FGcio+FMvkZh3yhHEr/Rr707g8yp9CgGCzZzc9uPGnthwij96wB+psFG1/
K/kMHZJcdddN7k1bQ+8SpevGkMSZv9WsnyIdPQ4UzL1WuWLCRmwF6s6xWIpK4H/s
4vbhzJq6VyRFaF6z6Z+MBJnRENBileTwcPit6VA5HPXOceF2auGJdLjekRpDEv14
D7aLVdNwSAX+bdYSm6U60DTCOn6wDDD2x/ofnZmCQA0DrOGM6nqsLOdEM8OoJ0d2
i4fT9xseeyJRCerDKj8EYCPORgooN49HDwXmvNzBhPWFgRpvuOHozBGwHc53qvc4
ZeSaGJIvQBQd5wCinuKzLRh6WT22YH1CkUxOXUhsc/1GEOv7BX4zBlTjkXFBk+DW
OUaryUFITBfgY7g3UwY+GzfOv6uw4dUFgO/NLEiTjSeF74cmrSYAi8MoL6UCi7gY
ZBVT0rjybAe8av4u1pFz8Yn+/oSpsMGon6aFSIiiM59pt3+//FSx7HngXjUGj/x3
6I6hQn5/9krgocHNGoQg/mAMRJmko3xEHytq3y9lfC/S3nEPe4UtMTRI6t0qAPdJ
B1nUAwMvUHhQphye9dHBrmDtzxZ3vH5wqRxi9mI7XPDgMWQZTjdnxDkQQr6MGPHJ
eF0pHsQREoodNQJey+hog9rtKTp6IjxxboUA8HaVAV0y7yl3iHVKvt7v+EXsiBkY
IlXlrlLBkSFULg3P47bKHwr0tZDQWR99HgaO97krK5gu4bATTnR66a4xsnP/BmzX
yru4++CHEqSM8cjqs7xIO5BfX7PSY4bcaxoc1dSRR3eO+n4mgp2y99jxGZAcPtub
O9RvXgdE4Cz1rR4/a+A7zklMarzZ3S4FniXzMUT3yBuwV0jyYkd8gb283d4nId35
XRo4xuS43q9B78i5qiRwWUC+UdiAjZ5+VWMiKMikeaaiNdhJNi/vnzGwy9q5BKn5
mvGscEg+zpAE+47rwjJhQiaL4C3w8/DVB3j1/sKfewB/Z3ZVUG9mmeJ6Aqp7zkCP
7Fm8yFTcDUtUk3dHwzSg93DQZJx80Z47hc+iSi22/lTaeO3d0lgCzvgR3NKRFyJo
N/yMqGVE/CcMa80H+kmmf8WLpOxSny4XpCRgPjjZ3QtV/JSzs5Xkh+ZbQZHGLdmg
WDfhxv7uXwpoljNXFPzU40pFbMmQdTlaKo7zReT3BonRnEN3cjh45jumdHN0luwB
+OoOmRwg++ZTUCib1024Bx73Vh53R9n52/YKY0Cue3w0S+PtjTgu/sg7ceWLLPhn
DMDqqzKzPDqX8ZRy61YiiqvMvWWoWfUVI5Yl+PucR58ssfH/F0OlE3NUcRfmiqdV
Z9LQVKDZ5aUNNLHTWe1XPG1GIxonjNFYUWDfcBD7YzMY6U0fETbPU5Z6++KHC3Qz
N7QvH3RMVagZpvD90FfAeSRN1XoesK7b+wSYPCioHUwgONReNb9JTpAl7rFyGgAE
bdvOFnjjhl60IpjODJr+Fr/Xy91PhFGy+sPiuB0kyGtYaXb80BTo+fPfpeTuZlZe
x4BTa7FYDilo1fTi1DpozWh52NL5MeVJUPrgVc8j2gC8hdju95r5phvJOpej2ltT
R+6y04qm+ResbaVqob4VmLEz+997IVm2cnqiXFSeAZfi1x6DarTS/EM5eTuSlptO
/hrbiDcx0PG0gRN0DSWRv+ou1RTe/oVyFA83mp+DWgFFSlIgjdG+wgQunmWdxnuQ
cssq25OJt1ruMBQ2qeuMkm9g8W0gWSS+LfNiIUMVdZsOB2qJJqTk2TTg7vsWWMnb
b/tZnYWY4d7uy97Hk6aAg0D55LmiDUKWcIPFccdY31/zYBl2OSgXcKBwEPJu4frM
nWuLje9hUDWz7++UKdsjbofShncb2eY8qAGuKvddgasruNV0/pb8Ui7asbaPK99h
GXPiKbb1uAgcs9CyapndkDE1Nu2o9nDp3atN/KoXG+SoVTjkyoINB3wH+ICkGURZ
VCqnQuuN8/FSICqCnFuTicAETg/+bRfzco9XqzO9DrgiKZfjQ4BElOli0anKZupc
yrDQX/KM3mZARfVc+ZrrYQWhp1hvVQeDn3yKxC/9OT7zz1GCC0x9TSd2o/NVIs//
lV2VwXyve7J5XZ/rRo+6grIlxLmxAzzjC8dE8HxHJbDqiLgUUXnetDTLaPEmBakr
7U2THmWUs0YW0W/KQ7MLXrne04/SQelmXMgCdGdXH6AK7uxJs2+adCARdxEFDVWq
jErTSfvOQfcEii1pq3fDRyuuHHAXPEW+IcBifrjd3VcNXOxV9BNBvm+bbx12ksAm
S7fvO80vXNaijTvcOhVWveNbetovL7tPGJlzHXkrgiayNAyFjmom1Udqc/bKKIee
VbXIe7zcoDLQl8WRSXoS7xLtsUlp+MQAW0LTCeCdCVhBgCcjy4fKpAgBbUN8vG5C
03jF8LvSu6yEpBUyv5yOpdfxUbsfVwhPRVm7mGUEIKOMiyvoBsCtdzEYGs4Z62W4
2nQtaLpBG4TI7vi0XSkuwsKUqHSOlPB4StHKTCxM8kLW3hZoF1EX6JgpWaBB4oZk
LX5PeO+46OZRVZOzJaijntsrHXZdwhXYmHen0AydP35feJFLboqfz70ZgiOtjdTY
S3K4pwolNAQZoCAQm1bxV5qHwnKOaBB5anBmjVv5PQ+HKHOwfw8XBU9r9Rs7AmLV
GnwX12qjw1p1uzMYUrZQmqjG+7jcUquEWS7qkGQz6Kce2uVV84jYB4bgTFCO3bft
5pYkUKg6P8tqHIiKz73dqa+Krw+LaYR93OO696s92miNG+Z6Tpjj9JPDc99ecQJg
PQhCFcb7/ZKO8oTQkSLMR4wrPZZLJ6zccyZMy+XtKEsoMDY7tn5UtVXX8XDp3Aj1
1p1yniKUaS1yjJ640lCUJvwSmElTTfeV7An8nzWExG3SBAm7rVKH8zdggE4Wrfu2
aIXpiHzUJT+bq0DSaBgBb1Qf9+rsEZS2ych7KRfmys/pkBuVJ1RGFWq2wIzT3eTs
62ZNy6KvUCI41Oar/881yDrJeU68HLNaKiTOhW4dZyNt8m9ZFlPtmHAuUlj9TIMK
8ya0Zt7QKFVb4zkg4ch3XjwVtvkKT6WpN53uy1cg+yHCGMemmfltIcHxkWn0ZQ8e
wI32tur3GkxP/5RvfdtAgwazbgs3GXaWMjqbONjtPYDxLxyC9CxHXtYeqFQUcFBa
lFSUZRzcm/KmMeRTuivDBW2C8/prmwuQ/5MsETQjsxeTxz5XHDwaZo+5sMJvtr0c
PteFKzm45ZJ/GtRObGhJNsasS7NGC03GxN11rSiAOIKdf2JU1EoL9M3D/zQZmT+/
6qtd+KO0/XZHIsMiByQBDYWVZrmJzuI5guZWJN6oUl8Yxp1JD3NYHCrDXizyQcj+
CMWxJJXqzNRi4dapY/hNCmdeK8hYyyVB+9aSng6PbZ5Zk5/6XTOUOUFpe0hm9+df
JaxZJxBKL7R8IjY5JdFr8HXtF2ltCZ4++QJAGMUoPHprn2X2srLstiK8LvCXKkle
t9c1K4hsK6e3lFMWf5qgmtAB0bOD+Udm6lzijr45GNQjIAwxN66UzPJIvdTn1O4g
0X3235u6mis2cWV/z61O8zGl+Vel0aC1M48P+ggKRnP7uvSD9bBDMg7zEo3o8fp9
/tUkCAs4x5vEz7yn2ZyYOXn8EsujSt7gq5Hob9oHtKrXOuveBehGiayo6LD467+Z
Lrm0ha05KYgmPWLQAW56tNtDTgcTBLnZWEEZ+1dHDD9pifJtHaTcRfyUZqTIfote
52+dWUp+5JrFMYDjyn0CRqaUDTQNm7xy0HxahfzzaNakxhOqzIizNomD+mekqcc/
KDtzlwA0KqzHBtaxmyQQGSAxAUvRKnx3Fxmamp36GuGP+AKmwjisKmi4LFBjxS0h
JmK8vXeRW2pDmJlG+MWT71k7c2zow9EwrZCKcibWuAxMXSecUUrvCzFkyGtgjrBP
Z+KEWoh3aOaWRnPVvbM2GBrnaTv6gxTjfok++nulzQ/UBcihx0rFdXZpoq/NkFxH
SZEC57aFXf3rtrDRNNP18XSPCmbbxcHPWgsdP+uLZoMNrHRycfzLaJQLlcqw83+X
vSTyi01MqhMm3Ftu2poXEtYLsAl5bV/r19gI275ZuaIoOs6u8PZyoh1aKhMhVwuA
YMPJ2c7TE+xctIA1DEdBn3X8zpPoHMW1sQQFQbk5mX5j2U3u8B7hSGCPMkNISPRO
ZIjbIeApJDCVAOZzlnYVlaEPWhTx3SRSaQNVgDKjWA7pK3IgGPC6WiyNkJ63Ug22
H2+ArzoDC1VWIxgoqoCafW1fSVq1KwYb7xP/5xZdxyYxBt2aAS0gMT9keIpa2yrI
LGcjmONl2rE+11k699r4nmC3XAuA07K7L42wyCptBLYsV2R3wTPx4xJ/PUT3Qsnu
0Ce5UDdqzMYa178tkLiko9UFaxC+GqcVj8MIK3YWyfDslpOJ38mwZeMl7OFgLLj4
RMLqoafoJEC3g+xgPp4dkJKe2IIornXbCqYDDqJz1rDPzQUjt48BTyajEAqNjKft
8/ra/0LfCUxFoFYfeRhmIOWRHxuWgLhIeX2Qc3P3/zOY73pfqV/t4TVie7Koyylv
HUQl4aTnh36IFbw/AOW0UlVfP94EqVUDcoJaaxTe+nf6N6QxH6Ahtapg7XBxLEnh
elTb3bj98+Rd5OVPEXkQnIOb/TdI4R20WeHWOqV3+C1ZX92lN3KdDmG4G9b+RpeX
68yySIuVayYaFHXQw7paR90sampdrmX1psKykXDwXFfi3zvx92MyFJa8AIm15mD7
9crZ8bC2wDd4SzuyWV3ApNT1O1b5eD/k5ehvRJSk+xmSBkMuJaxM2UdRYGC6mQgQ
3qrhmLvvxuCim/fhfL6IR3dNkvTod+7TorOj6+ZD0CpfYshYRWZ79glaV1uU9Bn/
3MOS7TdAVZDufCzLBrXYStNjGxNPDaF294m4ONDwIgiq63YCumFuEr3eVhD3XLV1
gWBHB8McBMKHbaVZdFyI92FNaXm5H5AQncyRo0+a7d8b913b+tNIY44Z4MKf60D1
ziBEEu7VhJ0Uf/NA/cozLAJu9MDpWDiysgeccXOMmZGB05Z2jsec8jWhQDq+iYrD
qcM1/Fs+NVsLGXN6M9RwcZC0YKxVFjMXS2A5IvOsxxctTmatX8hZ6V+zOUCjxsCm
rr9u1vl0GdGm5KMS/9z/Q5gcc/yKmkehyu1TNunMPOg0sMhY5YcmdaW/7XnSMQ1z
yN1ecX9vsCuqkfsiObTNe8ImCiq9W1aqX4k96OR0Zu2mAGusdVmZWgXIMVP5/NRR
qthdniE+DctyoL0XnPKgUq/0FX+yEH5criZNlmTW2bRNlIAVFlDT78hxZukSaAW9
Ji2tCqyYSSr7cvrvijJ0eLHd3aCywocmlTcvVNbXfJDFFWwFliWpxp9B2as+nPy0
mzY5JyIXbS/KtgTui7mq7x5Mfb0C0Y0DtwScAA38nT9Qfn/dMG5wVDVIoe/QkJDn
nWqbqWjVpPO9vBMAglMnagt8O2jF+Eer3msFDGizEE41xVNUtYoC3Wxk3ymfsKyX
WlNHt+dhjae0EB54/0Zu22CnRUGHuhdtc0N9QgkhHboW6En3kNzTwlYHZTI0BWnG
7tS0ADhhxwhkHe530PaCCXs3nHGLOcl8ozoVJ0qLpPXYhTy1uvpW3KS6YLoX0JB8
83AyN8+OTUpiodE0r8K5wiVA/29/UK951Bf3Fd6BLN8kvsKgrO3R1ydZZMOXjFh1
URvB2HJle9KEmhIory3Ohrf7EMpRCDhUiFTyixonIg0lL62qK/e1vv13ipCagWMK
U+RZH09Lb5RwQAU055qsLOYFAgTSo8cxme4stHv3QyS/LhZbKilQiXIWl1XhtBd+
oRoBRtxBe7cHDQTJ6WXO0fYpKZ5k9VUMscYVpARby2OXESGIRhs4Jf1KAJGTQ1J+
XPxfvUCoRxd3ot64g2kHECmzle9fIjlL6kj8PuUCuLxQxK8XAopO6p9SwS2bav5J
hUgVA6jgM1Cr9dkRy1w2UE/BDhtdXRGtmaBgkGwDBb0z5PDmDOxIb9U4fVUARXdx
8ROHnaHRopRP/Dfn+MFkZueSF9570ZgOiyrURHuHASOiAt1lNK6e0yGkaAHXMDeq
P74kzuO+M7nh4jgQ67AMVLVc8y9GGnjaN7xksWZzE696+W+VIrre1N1UJm85bMJ+
DMMi5MlEVSZX0jg6Tw0qJeSlr1vVplgv7uhV/Rg5TwI5fB6/oZl9B4bLM8DnM98L
XjXNV1ZgRangjXKYyflDQ2T4roEurMdzwjPivJ7x0gGpKrc74ykq6+/9zsNkMQbi
4q9OBTlEyrp3/rUHwswmJWCV25TRnxPgNjlJfofGyUVkRtfDvqLJtFyBVdXaohE9
bAoh0//TnLF5vRyROgKM89pS3lIHnm9LPvFCBvZhgIxzu/ECwKbnJK+cxy3IqjYT
zohv0h6G/Iz1Hd0rbrip6ivDtaWXxgQ8lAsVf+Zmug+PQaEreoDHl1ozsb7Uww2W
9LT1A5eZNyOlMpsZdv5QrWhzlO0i+PcWgtzAh+tQgKKn2B/eSDAyTyj0uDwOH/ip
WPd9xO+Wcmu0R/E0nLNJJuwDiTU7Svx5dIU3WvW4MupO05T8RHlmnaJJtargXaTW
DDVUDMcktiKY6CA/jMsATCzc4YFfH+fyunaAYPxA+9tn/Hdrbq+6UUNG4q0wjidL
a/LD75y/xlbGuwnFuZkAXcM+6QNsE0HoWr1PooKLphR3IlaqPgxRpxHJd2xzmy80
bkh1HUfbNcOdKfip8vhJnse3+ZbXu+9NaTwYt1TmGot1UWxVOW0oXHxNZ+kgc6Hs
b0k0eqwM92NK3kNO8i57uZWH/klF61fg3BkxRmhgy8P/eKMUdPOft5HzEpT9T3CK
QMj2K9KcM/+TyM7jo5B/x/zHHc7t1KfVetc/boCEDzGbwbDGuSd7xmXGqTm45AeC
d8e3POO2cafdMZ7+7I65PQ21zBQGlKQ7ffnNXZLPsd9JXXtzyX+FYgP9SjIEfgUo
mjWWMZ3y1EUQ2rby2THsiBLD/jp7jPj1/KrHA8X6Md2yYUk456fCo7pXR1Ya18nx
GLAYLkWUNydX6MRpKXuJXDbkNCOJXKxmaKtlsAstuIEKc8g07mivkuaN8TlaNnoF
CZo1qaHqofMCpiCHDuv+CYQK9Giv1rzOCgPfbq9D6+AYIMysJN/IAfvasano7zQ2
5ptxjnp5EV7Ao/BMwl9KBMl7uvYXRJ9IsQeTkDxBePD21oT1p9PHxNqL+na7ha74
sA0Q0I0SDsGxftFsW3A1HhUbyjmBX3y2VWppZ0k4GQEMarD/L8/cdKvxifqrgTV9
rKneFO/hI1wh6dOwrsi4hq8dso8rf0M3uKuBEJ1xEJZa7drJLMoSE2CrlgpRvM0y
byy3QbvS3Or9+RyAH6t3COf5U0eeARfocngrzJFbYUuPQl6wA45JOqv4NLxlgsJM
8G/Vh8qEMZ49BnQxnGDXuaCavYOAEUEp8xNLKhtNt10AcVU3AebTcXC8QfFZvSC4
mCAeW0+xPLJobtKWPAfksQEWOK5fIBBREW+VjTtwjxOR/4VT/azWh52TdKiVcLDH
CPN55q/zLoe+Px9K6yrSX0Fkdx3WUK7OIGNGn1VyZ/SdXE7lsHbWQGmQm6nz8uPV
I14EMzaMyGc27fuG7u+aIgsVIrBAVDMq/OvNVqOJkiW/1aN+9kGJ01YtAA7ucHZD
PRamnLscijRnHbBrokyaHqhM68O2OHctR1dK0nfdcnXhQRrF33iD/tfF9lsKdpOH
mkHSBPMdjjG4cKd3hfocHta5+yOeHG9HkcSnWbPEY+A8g1faJRZOeYa+SoU19/rb
TDEIZ6TvMqvm4/V5iIRRNsFmHTBz3pgcTlZPYEB+RHWSAy47TyNQw+rXaS1jSbJ3
uSk7rCsnT7IjuihSBRirUOVqlebVMpWwo2vbQelNWf4E3G/yN9fBA1tgSuVv7/qQ
01YhSzSuo1lgnGNKGlVe+iJlKT9fekUjxkaFbjGzDdNHhpl8LiPVDTmK1UQLwAZL
skNbEaoo2c7UPizXs8wPilqAHX3kE/XpWK3DI1i7+MCYXYx9j9eVWCHX5YPbUUPJ
QVzOmJaQRH6NH0ZOA1Tb4aybMrWbVM+dGNRNSnHG4w07DikUbOaYSQ8nwFUqPXc0
Vo+HxoJ1CEKtRTNrqvso0XCPdRcdqc5hHseb5uDtbSXkyiAj9Auc9Gzgjecfx+8e
I4XdMeVyCaszJBvy5U5vFN9zZioiMJKw1AXeBnXXGgi/Fuj6kveIBibTFeCz334W
pA9/RmC1AYWPuA3NUKYOzhsK8P1PVEE2sEDRZeAeYr4ON1V0FBRckSp8z7yAMWH9
yTyfovvobWSHWOi0X0x9lfBp5U1Uu//cFSpTtTP1NQIq0z0jc8CmE/76xX22H1rM
LQyfApTgxweKzs3ln0P0rarORJtk7eueDquOK9X2jJgfsOn9s/WkfPir7hc+t+Wv
QHFRwPcfGVpre3izdZYftHJQ7xiRcL0URxaOP/snW/OgF8M4uI4r5wycouukO+QJ
b/oEG4RM3rxdW1d92kCqRpDRy6OQlFRc2n6tfZoMVP0rxic2JYhIBBUVevtDGX6I
uICyGVcb0ueoUedavOak9El5qMt7kktAxXOpe3QpGSG0jO2GHecrLI8zi8uDNFwe
D974sWdvlRFmN2OwVXteh91hv2dI5tV1GcJxd2veZYRwqR1/09JN2XAizrgmwXEO
DERvbE/uEdRo8onWWjhvkrAwdY7BNpgNaCJjAU3QG7HOC7XEURhKRiulQ30PxcHN
kE8Q6sDhlTRGlkbGJ/LTfkNsoy6FhingoI1MKCF5+NE/WMuKdIvrevRN35WmsC5s
LOrvchqqtfI6X2H6QfElceKxZqzDcFto1Kp1eQeeevvVlm+mJaj8egxmdxcnEJrH
ENqmc34gjRSxZTNpdYiF5Ckes2i7N9ctRGe2Q/j7yYnY6kLm1arIJmphHHODgqQX
9F9gLIldQGc89yVpQ7sZg3KQHdaFMU7EAeupRgREG163mbv7/s51dJfJo5lCToc0
lmOc8fPQ708V8SzBFFoWW/bhRJqMamiWJfym23VuMYgp1f8esaWtQnSPdfHtVZBa
myl0upXPv8qPE6NkrK+/P38TbCkMX4MDOeGTLvIlxug9SjEfdG9MnYzxjG3K1twW
T3jPG7LLRj+tKOK0baaZmZMoUXVfP90Yhm4WvgjYnPf8KiYLoVKwaZiudksh+92t
IM4ZsWsas90Vyv/VhdDYllw2LhDBFC7QrxLZQjWjuCJOFezHhaySO3UL64S4YnM2
RtAPQ3HVdQTG66rKQZIp/swts2JzgvuzjwOemQrF81nwH/0pc+wvRP3hUx0+P4EH
X306FqKW1o8al3noDAsHrfF8S4AFt8G+DMhnD5/7zQ+ei9GYC4WZP+vfnUOgihIy
QxslGHRsupPuxZVI+oHONw6100To03xrS864VdEla9ayeLEEPANfqAdLMzzEvL7a
LGBWL1YbFxLAB4k86Fm+tAEjIPTzgHO5VdIG/VRJVistR7FzxBhDATezdeww5O8i
PJAEj+7goIS8g1lU4mFjLQoh9rQTYVkTXkSCDKBYLe6sBz1Xunn4OlK6LWxAGS7j
Li79eL43SasgRqI2c2DF5p4VISp18mtTpKM+8HsaM6ho8R7sieq11lg90nV8zeRC
E3iIPMX+ctYuwUKvRMFuJfeWn8t5qentbNOSjGdSfDscCLYM3klhu7Q9hh9m4YPD
5z6j8QPFSKwaYaBExknpIbr8RdIlYFAlcKqwzIbFn0A3c1kVpYMpkdHuDatdK0RE
zc5wnQln0YXhwi6txIlVhm3IUFcGzjyv4ozlDEwmSihB2L7GNryppCDCV2hcxsJX
cWpmgzKLvophRzowFNGRE/hkJka4in7nSTyFgkXO0q267IWlIMt8l6knhdhyFPx1
oou9k5J/XpByitVNH6EjLzn8cT6ya82eH5pRBiAtY2phhoz8Nr3tUTxC9c+dSYQW
qMpIB+JDj/xhoepw4ZDIU7DBe1AE1c+1m1uzJtg8vqoz3h3JvcGrsgtZtQCJeQSo
EymLX8Ia+5hd7XROnI22PpldKVmWG0h/Mi19TFOm0kuCmFGiMfC60jXGz+O9tAZi
RJpThkiuKNnfkwOlt1SAT48Z38AqW7gPsrvYjdkGDYOCTL1IQF/ojT6vinm0cCOm
ndWwd0Oio6tJG2AO9VboWbEdjNzvMW5Fho4cCa75Gz2acZ0JsJ8j3/BXv40Bb71C
ZmhzDVaA51nGWsd+dCKSGB5zMJDRaBUADsJc0DhU0cVc24rsQWmlezAUZ9HwZJGc
xPa4CAorRiiJYQpXv7ovni2ETwewx20AIPJOA9ojTboMNaiEy2T9hdCZZTj17Z6p
EseAhQCKrsPxMI15xZ4KjiOwBXrjHwiZDqWRmrCtonMYrb8mbJOv2Osg9cYfRRD1
K8gQi33c0ccG0Zrr9hZ49kRRX8ujj4Q6OovygTnidpAGNnURzys9kd4uIfy7ap6J
Qv2z38rq4KbgZ7cS45zufnI0M1iIv30jPO6akRZGs9v1nFbHjzmDLh5etfWbvf/U
uWjRlHTNxYWp0vFJQCoH3JUOmEzJFpmo35FLMzReU4c11nvN/2u4+6DDC3H3st0E
XEUZae/2M3FDhPHQWv6ZDZ3L8cpCgjeCu9dV7IKUu5W9jBRHC7Tvg3MG4laxrZkc
5VGCWm2T3Ekz7AY/2ZmjJxAfJCGhPjtbNx+9mfRqroCRb9AeYmJa+D7vSiz5RPVW
KVXa/EUcl38uG953RixLqThups/ksW7OYFNd2GeRp6Cg3MsNKRc8SQkypJci/lLA
/1trhRS0PO5MQMKts0nSxJWtaCd6ZhNZO78DaCrpMKBlHEvjwsDMO7LvW5vXzfkc
PnTf9Z2HWs2zYOPHxBmZ1BAhQV0WN+3CWLgWBwEE4CX2w9BmtJQbfiRxzCaEztqI
IGhd+s1maRsPr4UjFFtDovEQx8DbVSvAnqT87GNmXtu3C3ORgAu5DMZ6GmJUsrB7
mvr/YEsO5nr4z/Ro0EbazT49k9Db2cgXVecSlIyG6L8OSCImdNwKrqLDPilYwYbO
L9gO3L8nb6zcXQnRZcHZTIwErbV+r/DM9yeJfP+infwvAu8c4Mt697hXkwUoS9Dk
7ey7Wrh3lKgezdT1p2C97M3W/sAMu/YVNLO+A+wIJ7QC03ZBsqOH/nCabl6d29Ot
Qk4iq5ebxEoknYI1RqBL2OHtQ8Q99viIBZT1oFPO3Tv3jcI95sNfDjSsvsWx0YEQ
sIdzj4r5tM6+w0rFWW/iVIxGWBv8b/NlhNfzYRrto0+ErbsbGSx3jDwyoiDZLV3P
S5Y1zrYr7Lb6pddxt/48Y020B03FoqxE1EpartMYguVFdhoKnsT/o9vWzTNnB6EF
1JOJF+D8haE9A4nD74gLbEPf1ZSE38tMnK+T/KaKHtu56YTTlLX+vCMFjksNm5e9
1XikBuz+7zETx6FLSH0XxvyG/1olzRos3nIbLgxFqKzawMsNtsrT+CgHE2Sru6DB
cwAdWIewom1AcNXjhzQqT7WsY/kC0UlIZvkGiBNnDV5C5ckEtg/VdvmsXqBplxya
VTniZiraM71Y0EHiA4yxbaTjGfp4QmJVZ3nISc3ZIZuxodmOoXbB3yYiaFL2Dm3M
IyJo2VsbQ1g1cuFhHIDWu5QSvywAeMo0SXlnBVd3zCnuaA+llS+f2jl3Pk8BF7SZ
AkSr2JpaLYI+jC3ZUkunRLTghEwLmqcWmRstYVojx1q+jQVdXqtZ/BYmBwZO3qHt
1O+WPC0nAAhE5RRCQv8XArnlYETNaA+VCWOfBYrnMmBsDGathuSGXST+SJMuvLca
k52al0fjAMGzqmqaZUiHFsoAKL6wTwOEWKO+HK9PZsIZIaENgwZ0OQH29MBo2wSy
FeE9ospB1LFRFHKwRDURIaYzcklu81VXSTMT6yOdDv0FfZXqr5pFTUMP7RSQT7Pw
Oxo8wSz6tab2nGTAVdcbmsgQ2XHiEXYdQ20fnVgpUDOXK/mybEhvNOT16xQoeYLu
w3Gy2MqnPFSLPAqMFvJC92QfmjMLdTVDK5Ez1LCD3pA2MJxf7tKvaCZxpNruiovk
GsVpd/0qNSh9QnmNxS4WByJB/4XGErRxNwu29Hp45elffepNFGXOTeJiiresNJGp
67+stptYqUVbwVvqCIuZSG7A2Najzc6gpJ1hU7CA/kE0BeI4aVL+iISA1MjJjuGs
IzhCiLmrQPcfcTgBVIZA8JlvfQxDH8ePnKAKmdZaxoqA0C6EU2vqqA5sHl5FZIpZ
bCYEvUAIwpvwZQm242rYSG7OtEjH+CAjyZtiGRrEhXhy+fwjeybD80/yM2skDNJS
thNAOiWruC2x5HyGIjeqAO3PwjL/B+0hdxeOsHKnhbGstw3RstBB1Ov7ESn57vA7
zU8Q0ir4BMWbtwYy1Ui128nEThVj/elEWQFjEYiPIP0SB2E4iq15W8XEztkJRBPe
mfMlikoqOe/PdMDKm4Di64l8g+C5NRsBj49TqTYUYvqm4UsJltwGILQEUp/MisnT
5Kfc9B2Nr4Q+zCFtQz/I9G8/mu2F+BuGF64trA4J/7cVNxICpNt05Y+JVNW8aTtY
TJYmNUkPWl0THVfdhtawf3+SrzeTaUsTEhIDiMrjNhcj2l7yaM3TO71b1WYIQJ7e
7y5qdF+sV7CyYZK9bXbcfl0dKWjATfb+mbsR3s2Z5XIGUezAcDKoZJGr4sHwYBix
bz0/vWwIf4F+Un1hNECB1yzLvBKOrizaCZBcSEKG/4+7Wy2dzEJEX+dpufB9EVRd
yFTwqcomq+pbChPiHJnaUBEFql7CtMDL2Sfgu4QT9QD7Ac6rWmqBWZngGGb1OaIy
mQvAjqWpx/qOyMedHwSTXzFyYGEhYR0L3Ykh6iNvc5SifCbh+WVkUfMxyiYRiYII
vLSUlg+G8AGYUrbkNId/NaSw7bu001V/nEwFcfS6EAgeWgyOAQ+VMgbGAHFv3oJp
Zcjx+M2mP+Q1NJpHSJinn54YOS8DOLhk5QKIIpMXCm1gHhHLGQGOg+DVbLBE0VQA
NXbnIYwu2nEgWkszvGkSVeGoGZFOGhJUecZGPRBt1JuZv0AGkTNEE38hhAhl08ZO
xj/Euv3CQx73K3eMqV6o/AJ+cVJZllfK9oooor0MbWds5G5iX0beiNOVKBzlCRgv
EIy7ak7sk/2Zp9OJRFcC72BMmAGccte7kW5+l2B/jOcn8WwIx9QqQBkfM65+E2Zt
fc/AYeyom5oRms9eHZWPJNq3GLSL6/gfN7ZDVqzzUA7R+egwGepXwV2CvowKiXGR
ZDQoyQHn4EC+XTFl+9Z5ikV4C4Dq4lKW+Wb5avYOTiDp7Tx03Lulbne+N/KNPVc4
leloU4NgpIosqwl8yiEZ36U6/Yuu9b/hrOe+5Lz58cdtSzr9DKD4V7DgAWzmoEPP
K6ZALtvgi7FjBeF4G11mfGw9PNINuK3mmB77x0J3wbWamWJsjnrWLkPohDJB8Rso
KW6f17vyAUSW7gpA9h0xMDvJcsRL926gDvbDUnHh3ZoDLO8Z54OWb0RV0nvoA829
QpQSfP84ApXIHMt4K7s/H7zNo1y+JkefFwdkJaxIzNhjomcTJgEb5vtQRcYO7sl8
4arm6WNWVJ8CgBVbtvqKwqmhjv4y1ekRD+1n78sBN+/Nbg18TYPjpbEn5DK98Kch
1iDteMC8mcvvXtLk41BnB1DZQ2iJ4xt1M+l/YxaGojJzYCw3d5wyPkuBLEI7GKHF
70HVsOEGsWU7xSU+lM1TvowNuSpOKcczTxlxQSHqwbESL52G9pOTVxo9CpYUmW9j
2Gnilk7tiO99yRmBSt1zKTfbUF/arOtk7C9scceJRrrrj+Fwmb3rAdT/1qJXf0AR
W5pTm+6PHCykZp6a+/Cj5XGkmC61EonkrPMhCe++LJwsqkLzLiFN5Sn+zjZL+mlY
zWrAOvsye/EzBwyNHmrZAZq0TE34lfGvGWvK6x94yr8SMDacLJIpuqEyc/0frjpB
0FehGiTW22BPM7hZQtP2uyJ9Osd3oMRpaYM9kk37YuOQadlKSaZoz2z1GNvU64xi
0pPmulBKPKhhMq0h6fqGWJQtVFyV5nlEkyaFjKCRQLZW84eyWFV7ZG6/DIBAWlQv
BwlzgcaQ1uVKa/TLaMYTahpTt6lF1EhJWDssLArjsOZ1DYqhf2kwPH2BGDEUgnET
E3+lhTvsdVYtzU8tTYVLXs6IeBUHMDhoJaa0tz0xNAG7SouX9hdHoDsrumGyPGeo
zgc/z99BpJRXi+yZENm7zrduGux+3XbJIIia3omHiFMyy6LSekOdhpP/bFvpK4IK
pcLBvrbJkrTeNcWS4mOG6yC0IN0hq2EKCFWCS7Xq8IizshpVHD2RbYWlu01Xuou5
15qFfptush130FSjUUskozMmPOq3gcfnALUrzNIPrOt7kK6GVtVlVnElfqbpCufG
vdJZ6HldcqMicBLsBtY1csCq3jEsOHRdEUpqM+Kl99jmpq1QxG4FZzFUj9YL7rTZ
kqweGuUhyv9c8+yWHnz6mOPu+458jU4PhpACtWYK7Yts7aaukdqOR2/HDDxsymxT
Zv8U+Lxj9GsIRoQH3toWI/gQyeLGXw7G171jcL8pqiXw+QAIQna+5mo4Q1xmtuoj
qHBSffnymYA4QtvhAA1itrOgRfvfRuV8827F+DFfkOSqreJWNr0XoJp2ij0QGsuY
xqNhx0Q1BcNURh+52WvPARXvPUZ2MtRYDOLICwI00dEcynylMckpciQ+USYq2bzd
S2T34iYJ/PT51CHdFNa+rAVrFOCpnwm45Oait81wve6Jt9TUBZ6u2R2J8WbV4Gu4
sVGVhjO7BZqzVUpDxjOCf27MCJOZIMFh1hFu2uWqbsP/zprjsF9TL2yHH8os/SEl
iolSmnfYSr/pDN/8TysLwCwTYC41wKse9hbC0LBS+HWeojykvPVK3NVOup/qSzf1
zg/CDtKU36QrcMBXb/67WeKG5nekvlWp5APbz/nN9Qxmz/omBo6Gfj4MkWAySm48
qUPMCgBWDQ1KiETPHyHmpwEJB/SsSIFgKmNgAQ6A2TKLtHlSrZEm+33tgiKcDZ4z
clUSBLT/y5XJZgYdx50TkEkEYWsr0yzmOzSg/5W6DGwHzjFlWFDElwJ+zPy9ietI
fMAIflB6iHekhbR73FFr9vblnnAOM4P95MMy5kXdusUmRC39+eVPFcPOos2/T3eH
vfYwFiNb1G6AiB6Z/5YNflAm2O+w14XtBTV1n8deDB+4huLYgACbcPwodcVxvwUK
2OaLP1iOJTsjDDS0Z9onZzF5TtDjftInD6pc72qEqPiknrO9Bemyeary3jn41WEY
7CYhkIL7Fu0wGpG82CU0yZEEsSb0QInwVW50vHoeZqucd2jLG6FD9YxoCgwQZ2wP
cGu6VlppE2YXdlYzhqPuZBZYkozZEg0JeAMRZQ4Mw3EHIPwvrQHhTq8Pg7dVOkQL
QOI0Krt0z0Axx19BjatspKoIvzHLFhUFbK5gIjV8nbqkuQgPgDWJ5Q1YJCokCBHu
qdUoskwWVHbQhaSlP4vdUkWvUzce5B+e0G6jUx4EvYYpFsCuzN7dmRub/itPiJi/
ZwB9tfyJpnlGQU/8Jc+aPGJqUUCysZucGCNdikN2qyAmO5lZarR9aBCS/7yYizcj
TZwz4OH7qFaObyA0ydAazUD0N7uw/eKxj9TuCJO4yAx0qMOGngnQOAPIEZRcKIGK
qpEDSxM06dNGDUa9SMaE0azVRcYF1DHV6hdXPYEqcTQ6L6eXbBl6Gva2OsWTdCJZ
04vhJfYXZ4ckyED38BhQ6S5JTwMUmf1BoXxAsN+SEzHR1DGwcV8pJiWv0nSMOM0K
rRElyW3IsE2RktYIsReC4E807pNiQw/WX7SXx6vOT63OUE2WsiZ+Gyv3KQQfETOq
EWtA1dv00Gextw8u6A6CbCJrVWCQ7K4xlqU2drles+X9Ns73XdQiin49QNMPhDLI
OixI/YJKj4XHFUe/8khTMFjUBKsnrGYYqYdo7VwGvnC2wJxhZdPDU8YwM9qBsjjl
4ImvcGFngmj3rCOD/shC4s4w8X8cUfKGbY9P91VKiwRdQ1mm2ZlZYBQxa2oUDTge
dWou+pp4ktkPb7GRKNkMfpSRrYuY8phI4KGMWkmxPpi4TPzrLAbwvwopGGZqiHJR
pKBWpAMcLZ9MA2YcP2hJLjnYET27T0LuLkyO4DseBXilOCpZKiRz6AQhVzaethI/
PtMOz2N4q/uvcttRyN4gEhYCtSh8sUXmg5KFYRQBm2RNUvExXOJ34zbrHNC/b9ah
mGZvg+r+LmciNzPPHMrWRXfKUdAboFxjIxMQPw5Fw6lVH14G8Q0o7w3Jd0MnSyT9
sZwfTr0HSQrzSNHKmB5tUES3mdbACdOAqqIuUYoeGSoaec8CzuaZfkb24SfmzJKc
jUIgePljIFm3LiRhZiKfWZJwW9kojn3AmBuE8Sz0VzeTLgxcWVEGB7p0KWfWlTql
i7mrxlDqf2vsvVquk+b/ItzpglKiDVj7l0SPmoXr6rOpsIjI7VrTN988mnkJ9xFL
2glGgCpYv+dQD1Mi2l/5ONdLr7MucQYlsVjkxGNpt4AApKKuUCAX5y+Hgvv6ILtM
raiAkApQjZbpHZJsECBiN21g6jkXj6X2s2ghdpNawaMd4k+PmwPctJ5fWKUkKurt
UYCBFaELCbgQzhvvOI0+nJocZ9WA2yLAu/kj0DnFYTUu81FLhQkll88xqYsnf1OF
MTcnQUqf09Juk9Hswnr9FtI9Ko1cHDYHFfCvHZL94KF7WiLvAugHmsSE78IV0nRP
xtexsloMjUqzKnQnTTdTMYHiKwbTTpG65yn6fbuV4DPH+HDx043gA1Xi6c4BHVof
v/SkeX/Jz4XLiWgrcBagTwRJSpFWySzKfCpZpotsOSQ76uYrQS2mUB3qukCJdOo+
jMWS1bHAWyw+LFg8+PbuY6GLNEyvp+XZidS+LsbXyE3H4Ptz9/kE95kFhNHqx/ms
cELrLqXRexM8gEF9o8S8PRz+eFzXbU06YxJW/575ml7uBfzWDlw4zU7NEBCDr2eH
Xw99rUIZWKrulNCcNchP4ErgBZwmQdABftZWZsZEJ0KUxWFXhJ2jbCA81OuKzrlq
muZhoo7+w5/nML8XQw9rFGok8bMyHh9wlzR3+fEUXHgV/4cxmiP1Le0eoaBwgOIV
Hrv9hQD2GQVFRY2t6ymUrh1wnRhYXI+3+olaz8+whACRkCrpewNvqDd9bxX6qVed
EMqsUyYcU061fXXJBdQxpVDbNaDwDtnZTHUk9X/3BObc6ExC8IajR7/ZBdmuCRMz
XztfR09pSMmhLTsyDdb2yrBik/PeK8GpUYNhi9vERQHCncPjMeez7BrsC5jNK+u9
+PSvT7qoawwQ7/bsTUZuhPcUPZmZ/LtBiWXuydZHIiJ3117bwLH17nCwCfVR8wim
LZ1AmfSFEpRoXiPLX+rKQmPTwpomj+NqYCm2aZDlIL6UGqEA8/cZhKkO33ss3pu3
agZiz+bwLAlF8hJ5ZZRTiRaG/1d4xpVjS8hx0fuWMRswCX3T5CWlW6uWmb2Jtu6U
h+2/Xg+70JJeG/QpNkDbAbJOA4N0a7IYRGlHu8mhm5t1uLAQzxVEuQRqSjxl0z1Y
r0p73C1xqzOhPDXRzEp5hWqrEPXpRTP795p5c5YnosgagpCq5BitW+YO0nElB61x
GhXSU8OJqYUmFbcByMrQkBF42ZlU/VmUaQxJxAfvyiVUs1cj7EoWYIkXw1YX6Cw3
NLC1HGhzDhYYm9mzi+lrl98CY8jFmeS97ASp5wT3cm/PXRbO8Bm4BraF31NWsurP
6ixLukpbd/wgubm9HMsNBDSE8KFQ2SpRffQ8AI2uwZQ4XnwR39IeS1LdD9gYVDwX
GubSswctwYtSt6ambU2RTL9AsdVPSVYokC88aKU2s0jXhghU7tKWVEoVW0tRVT2z
zf+FfzU/s2wvmNSJQGt3oXh40g6iiTUr+OUCTSEYURVFTuFdB+z+4OB2K9pPZG8L
6kuQWTVHOnEmbSvgU+Tsrw7PKsvfG0yvr7GaBGuWrz3YZdxa1YPAoa9JhFYK/Rcm
EY5w2+zt06gjcW3CpIhMCtfkW7NCMnO+zsUMP1RuTiCRpStvmvdCVQS5FxO86sjk
LHoHjgYQ9ARaZV2IQFuNJIz5lkengm4felE8NXPnby4tu/YvhyuPODntAdCf+oxP
yU9uVU3MpXwi8LaL0F4iwCjVmAgNlGmEuygsAj0/w75B/N7IMqlliMhuiANDbgXH
2+bKgnDCkiVlgRaT47qcy2cmKpGIuDAGzn0/t7WmEIDY4FiddYClPBgUXTkJB8jW
cNyVMwqNfoF7qQA/BtKN4K/5uv/SubrLBF6glZkS3CQbE16/VOWJvsMwPKM+08qs
ri/rbWcmLxOj63rB9pPO7W+jcEZT28wZy/pz1cYsdDaVg5V4PBlqY6Ajw1z7nXjD
RPCqGv8S1uCSPcI0zupiQd8r+xmVcBw0p/cIxdgyjHsS9dtA76dk7SbNu2Su7dxv
QM5ZU6jjLtgGgAY5f+G/n4Hx9qu987fHL9IQ65rUVTKKuMFuJENMLAa0PFe9iHxi
134oirICglLY/QSOizt/D/ZaD29iGT3k8mFmzHBMvDdXSaEsC4kqqjQm59IyGF2U
NSxd/pNtQHfYEJ44kqYOovD98pftckXYFz7m/eSxkRYxpM7cFwvXIhT/hlHYMZhc
zLu3IZIp1lQJ6EdK9E5DC3Z+u7Qtpa+lew8Wlf369griRh0r3UA7zcWs0lbjzf2n
Z9fl08PPkiRpkfVz06mzZyO1rEv1WH1QHZ4BzUQa/ChQF/oqfz5Rf7KkK2tqatQ8
ypSdDPAVYA2D/HvvaHi7PiKZ6usIn2MjxTmqW7iKQK5Ax+1flzAUz6WLRFR9EDB3
o5CG7CPAqaOwe2eUaccexZQ7gq6FQam1zzH+JDeM5aEOyIi6uYqj0A7EQ+HeEdeT
SeGKZVDVlE+Kuon/8Tiws/gqVROBLlems1iVdxJyKrPzgH2Cvjq1fD8q7vBSRMKq
4GKEKG7On7JnVaGotwgInjU2YccsoCr5Uit6VxoXJs2M5GIYQgeBtDe7fFfDPOTm
0K++BApqHg++XXmrGhUkpXKtJK88yUoNp3ogYSfcvdTfq+9MLzc916ro4GXP7kyV
b3EJJFS3uSnzp9/1XmSXKzqmg6hLJggtISm6WPkzxogaTLpb4UOqyK1wCEco+4zm
gcAgUwoNmvLA3z7hR8NPhwGjy5KknDgZQGyGtU57GOFkXaYIB+AedDXU6xwMNm1t
7FTjYnRvEdo1e10RjnNgmtbrR5HT5eoh+/gJF76PMENzKdu5QIgvbquNqJdOj/IM
792MJdj6NgwyLAxHVpP4nquX1h85pUYhXA24Fsw7E4ycNZLV5U8MNoVF0mMAX/Z9
rFoRc619WlpvlP6hNIsoNgGzPAugirqKsqApu8cXiQiKeq+vWtpjSkPYW/ihrLQK
2Tt2dlU5l9aifx5OdXHwLFPkDqsP+TieXLAYsdOzzvQOzEn4QuC5M+6SkWTAgpXn
1eHLOwdAUFkBgd5yYoTZAt8d22afp0dm24uPMsl26ZmmA3VzSnNs6+afuz4YY7EW
fpCBK3Vfuy1PhABjCcHVCYPOF1W6Nc/BP8/cZ0LoANI1SuX71N7rZdRxOLuDJo6z
MqKbiGAF+lkvhXenWNQ9JNL+HoVsU9BN+xolutWowSzCMd3P5B8ZMe2wnyhfnImS
9ltdMbx0rTBXm1m+mAqQABgQAAd7Og8HDnjnXugujrWfUE3pArIt9dGBtGXJXdqS
WJoLWKiz7KblS3f75DjWk07dRB1Tvxy3bCTIvk9Mmjylm+dFLmTxDImK02vRVINj
zN08kD4Es0JN+eUcvs5FI08yCz1e9447TLUZvIrajzx5ClwEUrq9Bc37Ubp7qg7g
qq/jk/hmqO9fmnfkp8vmimK7emaPfiXhYGJboCyMGx9D33DVt4+IyeebWM95pGt8
9SMP+E+B4cA1NuQjBO3spvliMd0Z+0tCIQ0EviqoOeww73sdHHABLTTdUf0qbghO
bFT0TRDI3e3BEIFvCh0m5ULcKNdOxbto5OSWrvrhWcmJTFAxkj5ieorvI4eoCSEM
XLPqBJLC9OMoSGx9APmPSB2+ZidznhynFiAymcI7ePHdOlpDPXDWKmlzm5RrC6AB
A7RYK4Posnuw4RcGen89mqocsmAngwEoWXtaU7UaKfczKYL3YZ+21jIal7DAyQTT
zR0S/4/oe/CGFwYiCpOeTxPkrfGgl730l9jbmbBoOE2+sr7xl+jIDzRZRhfN77PK
5Sy1fQRWLz3XpgDbGTatoFpKT0kk78xbuUZaOmhMyfXrvtFV/WFApZwhfMrdVCTu
EdW1s0FfE7k++cRuvR8D4IRptBMsdUTNA6ILgM7OLWT+FDz53XtVNXLAtZfU2XXh
RRSsIa22XizGa/d64ZmRiZ6ZRCAhL5SYuqrmCC8u2ZnXc292Z1ckFSbEDNeDiZxa
LtX51+RdsPzoZsaBURJllGezOArAe5paNMYJFX1YzHwXEl35bTu18/lmDnD19/O4
oYODyOjOz4fH6fAWE+KZp5M9Hs0iKNVrSnDrHhTffrE2PVASXvcTup9VcNqb1tF1
ooa5p+WgmNaIvRBBBypnsHxNM+8X3VKze6UeQ0unoibmrxSMBHBmht4N/IRBVqND
1iNkmdR84z9Rucszc46yUBgZnyKwYVcjQUZRwJYh415CTqnXy1xsvLX8V31bltGJ
LYW4gHkf+M1C9zUdhQkU3cTuXhevclkWWmmDfiIAD8ezxSnukRxq1WKPK3TXXlRm
F9jiGSBUOiLJOL1s/yKrWccYGvwIZXrn8T7kR6RVXH22kEIbg6go4MgvwlJzokXt
kQevDWLGvD3YWCTdIFnh/UvBMmD+ArCyPUu4nVWe29xWi3wV9l5NasqV2kzOg9zt
cSzJgAyWQX1AKKh0bqvy6splNzBfjpjOejoQRZAnjCKuUDiNEjAJKtpnP8lDB23P
8wOWuzJQZd5nm+9TVAV4ixRpQ5SXITILIM0DAD/+vztYdr+OyOCq8+b5xMaYhHvk
dTWeKyVZ/jbworEtTLxQcVhoRX9X2s1SlosgA7JkkHH4lOTqBMpHw1SbxoAE7LQy
ZpGbU7jffbIOmv+eKM5ye546wF+1dmmx8YGcyKTEfx2kzoIttC4XqO+kWwAjnsqN
LKvDtmkb860j+gOVdDAjdtTLfJ7I4N9VzX6Fz8p+1ZQ39uKiOZxr5ScqclL4TJKk
KK51iSHZVK1vCxhJkjKQriFlai2yTJyIrLeOv5CXdj5/UPCbzJmOvGGi/0tLFDej
C1ZfdWMSS7IOWknobhNnGTLZhTFoMm3HebN7zN/XjzXcrfk/vFDWkQCSQgB6tMu6
HK69rYl+4Ibw1pMJb2TgdpNmuz5tEWN5N5J+FPKfgi3x0m4g6OTYRuLP5Qn+24q3
nkLwXs+5bjrMmT9g3pAkTvrBOSgwkAgof3l9a4pxBCYFCCoAEULrG56GxHnbpUQI
XJQDLmyjZhZ29fP7cJsFbHEHmYeyoqaay2TEuP8gvq9N1br5808GJR57CxkauEMc
RZmET4RaBZf++FW8B3D/9NzpJZWVOdj26U0AbKC5Rxxkr9J9CvGgNGv6ORzyutjX
IvSAkjp87fVmwcY6UUV9ublXAGuYhHhCTleTuA3ShHT9jKQUgmcxxC4RdwAFIZJL
M+5Y3XdfgcER98tx5L8Ua2eTiPDL/u0Ru0mFnOBxu2FdFHo0Flg7aosXuo6NsdA0
C8wAuINPtyXWnz1laZUU2SbM5+b5lKsXHcowCS1mRFNz6YOfqracs9yN42zhACxq
eBEOUwCqQiGo3VWTjFBeIWkptql9/ViPcD+NhuBdTAJ7jBcI8lUQ78RpddWndaay
eOidWVDymq7mNF5ag1GYg7G+qh8TQjChLnaNoIFhMlH71jJoQNImRGxsgActKZYF
Bxp1ri9/I7KSafurhgbMcVPsgH8gsZ9bXOZ8MusXDEnnWHLlJBSa6dbVaoxNzuus
rGTC07aQW7MiobOxiJtnCz7ffxJBld11iYWJ68NSW96TivxHZHe/CbmNoYYIIVS9
8Vr3usu67aaDgRMr7jARzOz3q+tizwAnHz5lF2o1JnF+OU6qn9iOp+o7xJX6Znt5
51VRmy61jusDbJ9lBSL7gtJCoZpHRhsMJKTWWjZa1wwdiche8MqgGf15ldT6PRIe
VrqQHBNa8aYSk9nwfX1A28f9w88nHmepyGxFQR/FOqjINhbNBA8aAy/55Akce0RL
6eJ2cq7s/dpGoqd4IMBrXWAMg1QONQvWwd/jXrh6djCo1NnJAofOTq8GnqU0h1wP
qRf5AhcMMoTigvn08RWVMPHQb8EzVJB3QsahgEHuaeNfV249/TE9WdE1KUrcqFhY
2BSOZxzQBMiN/07xmxkbMrq4j8Qa0gGgZrcS955EPb9QmGhPSjfEkFxsj7I67d3E
UZSK9s8hImd1cpnRuhBwjjqrcJXkQPa1ZdLip+fRV8xt7qdEwNISKGB5cO5kyVoz
HcieWzb054DooXtIuEj9sN+hX5Uta/eY/CLsLlynNOAJ5T4sLOdGOwp7THy2PnBs
AaLHSRa7/pFaowgw7hgk+5Vqq+i/9i8REkZKAF8Do9XyZooTFeqjrqOaMBwnpmuY
yA3KKkmWUggUzXWtD6gbnjh5dBKbLgR5rjo4VOukt/csR1BkG3wG1JeYlcPjtDqc
qtSN4+MN06LBXS1HBXOVQUKp+vPcfqcdVznYqkiqWfIJg/blZEBYNFvs9VWVfECf
4H3aEHbrI7hgyNg9a0S+bdPuzvjiPDU+xlpV5Umoy0yoBgyHBEM6oN4MVa0womPf
yCzcB+az74tXW+9aLg+Zv3y+G1EYAw6x5CcFNvklen+syynb0cMxeq4a9VzUS9XC
NcGobK15g9HEmQm8TggHRmrg6EU2z+yTJK7Z9xD/PUDHCABFstwGQOxWMXXgKRst
dlAsBDHz0sCz0VcM1ak3DVk4qTPtPpMgN8OPckv1d0PDU2weoF+um6y3LaxOyTSw
VJoxdRaCNpLs23Laf87U1XQldbbGOIJtJBW7WPHxeI2kEyQAUmSPBm9QFwTd5GRD
oXN1S97/PuCU8nTnQcA3kGjtioM93EFEIHlqrFLldh+vz+yiNQBUtH6M8TkG5Lxw
nXziHP3oR7q3UIzVqrkdj4trBJJ8zyFoqrqGiCWxkSWWPYwwdu5hhiVwJOTZ52im
OvXkbzHRALnFbEkAi8t0vY5q6a7//hroNok/MlNhyzoXRo4wTeaKNTzGY8RUJ96z
ncg+XYw/thkk7lONbd+udX3kAsQBzK/Ra5oM0sYG4s/nTRGBuyJM1iIaNrlNnb0f
GpcWo7C2xNsTXZR+iGs+xlO+Kc2yehl+oLE4basyM5AH/nVsNp/1oUcWBq12q1Md
UViI8yIsrpNNdSkGqywHjOpJaeXaxJO8Owp4MuNuZ1kq3ev8NhuCfgHW8xp7RvgA
SJ3TiqF+Rp2cF3ylxmIEf/KQvsaSAY9gZ96dnM3SAHkrD40ZL98gfMNSsPEiCfjU
QAgIDE5Ntq4kJSV2mpFxb18aAe9nTkikAh+fnjXNryQ9hHue6lovolCeAfENdRbc
fiAt5LAcTYG2nkVKWmzmdLsMN6WHz77vL8TlVSPyzRmUgZZP1FPnxoYAXpJkQB5B
VXYkFwyeIVH72imhx+Hg3vdDHq1RrdjshPzJtaxPZfgMUven3Mt4J4UflVDg0XjJ
u4KTH6Tx3j6SB1ixjbVmSz3IJRic7gHHuszGtWpMiP8ntMOuhGj347df7WA0Puq9
ysOUbqY01ObgoVKJ+LYBpppi3POibW0Op841kYTpklCMkaDI1v8dbBPJmjq9GwBS
I6+R+xVlhcuRQosAm0XHsFFRQcgjL2UuyksYfZhqpERbxLjZ3uMTUH8r2YHSuC86
SHlISwSL0rhniUcqXe02RLjYLpbxgLMdZOPwviTq1bmx17tRkViMZAA8F3BUrf6n
GpYVx2H9fBm5PcuYt8TKQ4Kyq5plAPq1u1QDVsioy8OEf6rlpEw16zmp5Rfoyo7T
PAUmJcOoGTYyppeRgYh1tXmKt9cnT7hTd8Mtl7n29Cz2ljDBtXnbVopEUouQhH0U
dg+iXtPJd4eH2W+sNkgYvJnQB+byFfH4Dh70YoVGNEqgon5IwuhT/wRP8JGY/h5U
/dSXhmMwv4L3zzHFiaUodonxMjPxXJPxlnKq5CKNf5n6/rA0NxmGq6UKDH+7c6Xc
KCYqQWW8J3nW4Opo+v93xZW4LA/7FXLjm5YfWsMk5MbCAGqbm3z+P3E9YpZxmyLf
4MFav45vytE73WVP6Xfl9wAsVx8ceitXyH7SZy159zbTzGoRBs5mjg8g+JfH21Zv
2U6Y/YiUgOQHkCUopRo70pL7IwUTx6Fw1iOMvQlYn3tkDlcoEHAVYM/14EMeeFYY
oXbMv1PYxc+VClzYwjtwLNba1bXVJ3GxXG7zsPIEhMTF/cREOInSHDfCuFO6oySK
p7uKcqpDrdW7IOG+HD9IqXlwLktWpFkRWy4IIfj2RpOkxgif2oSQ3YSLV0ESOPJI
CnvofgdA2SvuMe5UkhAInVf50teULAervQieVkgr/Ae3lUe9E5mb+dHmBhm0ZmNV
oSCQFiLiDmGnIwC10dkm/dgjMFFgLHM5TnGYDTetnHgQ847q43dsv/PBBOozqY7R
ijeExAs6+e2MO3mytEV+72S3bv412WxXtwFD6N9ITx1sFY7qD3pagO3F9azL23RM
rJyzWs3gG83xDgWejMT3D1pz8zX7AQGuhOji6O2V+wjCXsnK6bce/bL9K2b1fHhR
d2u0VfyAjDO+tAt/crS5TmlufmCkLUnZTEoxMttzdNwYyjZXUzYhp7tKPnWmZrW/
TzysghEv2353Zmr4ZzJLt4E1CR9G28zwkM7OXZqzujyd8JuIt+EUkyBQuaUi3q8n
b8C29S960gxh0uhBAGTDMchLJYrztoxsaZjqwfcIhKz3jpBGEcdMw32wMMgub/Qt
vWEkVno/K4BjcSl9MRao+aYRXwGJPPZeam666slnFUwsblNoznE7iFmtL9+gP9Bj
VXu++KA3O2nQ683xPZJjedT+7Tph9Ru6cdkr0m9hoX9RjBBgU6lLL8FseMwB1lj+
GehYrQzdASTcA13SL6KXE7VxXJkMvp8eWDYhTymODAM1sg0WltHxzS+3vWD98OET
9fRWJDLEVPehTlKigyszN1oKpK0qO+Cd2oTIpsDtResAmtFwK3nqKQji9tXfoVvR
gSF45QCmaC+NzVBqyGsuJ4ns8jZ0MsQPNqlsx1wCTgjgiL2IPeXJORo3iWGYOLHL
ItcZ4aOLO3Swo4dtz06MEjO5HiTAPU+djKnEnTktwGw1h/w0zwRQQgffq/4ieFC1
2pRKLvOjYf9c9PxkI4c+fIx64zQnUu5pQgKLa+WPzqanR1b6TZAAh4RQO/uyoorO
h7dSyeByvCsZBnQFKe04sRN9us4jNPcQQe8GDgEKxKLiSoGSpUFflxoPsasbqou9
swrkq+R1TzVIycqnH76YfZ3o4kmTxC7FbJLGlumK/GCHzHXfwr1V912umVolYND6
R5EAB13ywnetV9yBcjZVxN6f0YnASYK2XN/zSOSoIo/sJonZdG9pM36yg4OCkpvc
24U84/gXrAJq6vmoqX/PVRB9mXmtDR4ir4LxdaPPmXdUuABb5HPPO+UZjDLUcd4U
t+lsU9RSz7WIh+VIMA83OOpU7WFsQLe9fXx/4tsd0JhzKdZ/wSWVw1vO+fcA5QMI
Bf1au6DqaFM0mD32CdiZsKCmShbsM8Y/ZULB8GC32qwBplsz1fkKz2tJecDZSlWa
6ST73CBu2FjDOviW/v8XDWSSlkwYyPBnxfqNpRWfrK+JggiCq4DKBvtN50pyskMe
ZG7GhBhix24v4ewe7vD8q4Ad6hRGvwiZJVFSoNImu/y+aVCPBuPg9gt4uwGOlVvv
lHiRy04danjRGijP5ugiwdwgW33FbYciNzlm4PObNcV4YRWycXs0dRyEjVEBzX/m
evm4PUmSmh1AI09MWkAzx512N0/kr4kd2S24IIiJU7a6ByvweYVegZyo3q5ijHSe
JwcAEELbCq3HrxvpnBQJhTGUl/GwB6FVEoWUnyUWB2G5pyQ9QlZFUlI5+FOu06j1
r8ykKPdY43FiIhMzqGRairsaPUOmdSonwu3wjpQ2q12eKOSpD506Q2v2EjBirhb9
Xd3bz0vopEorGUc6JorK3wKhD2WPCGi2U5FCuOXs8ERWNIvhVlvu56CZKqCJxnKQ
CSfFPZpQbgKqDPL/lytkpmgEf8ZciyynamoNWg49CChk6o9DjWoYD3oY0Nbe1Py4
Bx73Qe9stBdaWyk3Tk8RCmDmGn7FBHZr5gbBQaE4fpJxrsDHmgpc6TvqehO9apwb
7+azg/Y3+ee09xslTqxo+2ZNmqsppiHvcqthqyJq77bymr0uCcjxc20wqEj36Acb
SAbmad0ZaQzzmpjtIklrPL3awenOD2jV9yjXgANSglBc76yk3GwtdXyDV2J+S/EJ
lK4K9PAnOVEhTYsA4ooX5qpa3Icr0W7o/IG1yZoN2vfkE7njE3jWhQ5sKPPU+5Vj
m0eIaY0flCK1u1SgnoSY8pWRSpPHEgK38BuvFsaiUu5VznuAnE10bs65E1ZoTd4E
18FmawTVu/VEGbqDfgCbIIvuByM3sJxOs+ueC4Iw5SFJMSLExLzdt5Aqdd1bt7HM
gVTTvscqiVjl9699WpCyXJSvyaX2oP6jRh7TFI27xpJRu3uNcCwulnPzPwj04926
JpuaAQZB6s+5hpMsJ1O2GP3Vh9+HhZfj4GdqQaSLGpvzxgaW/1WzM/dFqIB1VGnX
+Z5b+xxpx7WhKO+19zDz3d4MkxBGWIZgN2CI2+jsbiaVyuwGWKFPRsK5G2BERbYt
B9s5paqqD6mLaVK1dJEsLJzY/v0eHud8+DxlBrdAKL92jwy/wj1UA23xEkUIIyi9
gw8jxQmCjxEiWRtqmcT4oKpKDSYpIKie/i1C0jyiCYsby38eOHB21k68xAJHERX9
ZQHIMCTeEopU9U3cVU7ly8bCS6yIUPSeLlM3N2IpRC6KCQXFoqbo384JvRjKw+FY
ESC1O0XIaS72HHK3C+PX++LXW+I8piwLdmIkKl/bBnfAv8NJe/zkA6u4D3pvRu1X
ZVI8+efX/pd5FpDRR1s8UKGuM8FJpw5VbSmDqNYCqTsrGC+1O0giH8DUplYK27P4
Kin0z92bgbIMeTuKgwpLFY2zKa7S+I9JKhYz4MwSq+//ZcvmlwUUNKj4whXGxTYV
2HxLQZ1KmInan1oOESXbF2vBaPW3lD/CMCd+xEl8MIyxyoM1qxTDmYH+d5oiVpm6
RxmA7q+OmPzamVB1NXFb5gGlDjXvrm0UFJTefg3rhlhtr2fnLGnG5ugziRr2aSq8
e9thkOMERQrglxe7Tgz/tI6omzTrlM5EgI0tXhkhiEloqH3S4CV53Jt/5aA5DCZ0
uJ/4ymgaa88rwIMuEURTP43+sLihjjCqOaQwqf95ZjOZsp0PxTPu6LP4o/kUvez5
b4ateo2lv504ZepFwRD46ZwjlcPbIJE/uiXQIuLXZqBUJhIYviu2xWaCcr6s5s8J
DJKsA66+PlWU/KU+YbIl+5jIcklNXts/dCXdN2WjF+Jp6ymBocnVZpor5g8Mq5M9
Q7HfuTANS/kJzYSVlw4I7rgCD2kZwHoU8mO429cZc+iijWh3UBUCvCOc/LS7JBBX
KjGobC6vI7/MfbUiH572i+yImM92eS2/CvY510q0ug94uKYv/71K+YK862sczkHj
dETVYqdhEa2vdzmBW4r9cbi0IvPl8YjEXtHC9i8Ss2wXjSVX+hJpwytDQ2647Osr
iC9cJ4Ez5YrmSGT+uNgEOo66U95SkzcWEKUmJzvqhmchyPALGcLGj6v57utvJ/is
NSIt85gb0kNPjSkU7OzrQs443p+5YFSklPE8hdYkWmyhincQY4jLeD909aCoey9j
MyzP5F4roGTq8WgI1M9tH+sJBfgiGmOMCNeOw2JGm0wfpvJ59KvrG0OB9BKcGfZI
BdqPYPs/S4kE/tg6pz0tSI1fIWjeZU/DZJv2kWYX9GLBWjpKR2aq2rRXLWgBizWg
11Pr2jFo9kYY1ksViPeUSCBl8yAkEboYbFJ5VsLCz+rxgHGaELgos8vR9LG9+yqB
qautqXiWOUz2YAZBahuBw4hKN6824AgPci4y7STI8KyUXjJx+cBJlfkDcflbMM7u
082BcWy/uEftb672DLwwWDD6HBlU8sF9IseOWBepxIpeKvNA12228TsTt1dxbfWC
TVY8n7R21R0s36xtdG1hKy+iLGP+88Qk2UUlIDtWXyQX6wLGb2odZeEl55H8Cuhg
7A84cCkiGxANNpQZmnljRQoKU4k71eb7HCb0mCJdgl9If+18qJ7e8UmiT9iVSboL
yQZFUhBJZTRFRh+gJm8M7dto2vBAT/oWpgJe3q9BiREOCK/Q9F4R65pVusGsry3H
NJOyPJPvSOsQ+z6MAZuo83XFXOCcSkKlVDsrsFp7ib9QD78pB8vBjIgRgClKEylm
LhuTyoxiq5/jZHoCviucuPBysjwsk5j1bqEKotLY8zRUzftJsBR+8dJYx5pjXkvC
IxAujqoA7Oqcwu6OYa+xY7CCVw9aHd2TeO6MQyMlfS19ac6U0pD4tL6vTqAETRhb
epItw69PL4P258iVP7IAcOa1pS2vDlvAGkIfiGECPHVy6UFjt7ZPX174Byklp/al
DQLWYnQeFewZ/2aRyq/9BpAacQgbLiqvM6BvvP3YZTg/jt4ucSHMtY4Km6EEwqzS
5Oo+B0OM3u+/V90fTbUtigapyO+EQ5kLm3UP1CW4YI1niaIJio3TG1cEfHut2Fto
QEP3gpATnEdwUpSCv0sVNXhKhBhVn7jhIlP4kbgSTDOBoFykRv2tMcJ4HwD48oIt
QKgrvvgVGWRiOjTuQvlqI2ugdHM8iElnk46o/ikrU8BW79cfUg4i9KULS1F2Zotu
9JtVxnorZeMVi+TUln4wr6Sj6Qxu/T4Bvb21zGErCVoCumwQfpCWFReMJ3wnamJs
oce+0s9PTYGx5XBNMeguaa/TZSIQ+pEc7/8+PR4qX68irSOMHn5TJCHtY9yU1TsO
p1dK7frsNq4WiuyjEkWTLFXchQ0I5dqu/YR85iw04TAwlRL4zmKOUaBzkvmZsPDi
hmY5eYeJugLsQWymv0qBfWGkDVpT3Dz30lO25b8q/7bn92gLOG0/ZiRDOV1eXGcK
Pq1RKk6L70QWjZjBgGunuhMT1/d35yDA0GDpaQARUDifKHKDKatgA5LSJMKniVzD
DAwIkbxqxEBCd3bVBA9N/m5friwp20heY7FEjLOW2/U3/ShzqHZN4FrE5r9oQZ+4
pj/aJm4Q+9N+o4xeNrkbDXg7ghyF72Hz9qiHc1Nck8AEUXq7xB7ybzerg0l2QgCR
DIR9p2qXVmZhWmB6pQNaaSBNZnzQLIZ9aWOzdmeExPJUDm+Suz/QmNhpq51UVjNv
9hEn33KPQ1qgUdaTO/ufKOumVxDWAamlL2uZ/C/xfoUCb4hLpZq6HI6lzVrfQ5ZK
L8IzGOrzVapEITuPYxo72FIWjBYYBEEJWUwB9nfFpqOHWmrbdEhO30J9DIFs4+58
qILM2gt+gmWN54VGCukb8pJhcZFIzehuIX/rcjISoQ0R+RISvNQrS2LYkYv8lNYI
u8vVeOTbIZEx5SCfstNpSsdJSRLqsmx7fZx500OMzjQB4Z1PPH4cPC6mFz/2ihFV
qV0KfX2i3sYPHFG8Au/I6SwMHB5VaICUjWxLLyhILIKFtx91KZJjZmm4/TnCRGO0
i6lQ5HPS+ZuFFaEjwPtzumb6nJCcQEV4fj6J+TJEEWrdisGnU8ZcvjR6o2LaO1qu
OiAMsFLhexlrlxk7kgyqSnY8oPchH7A/vc3aacXJF4EZo0saHQTNJsRuFb8X6BOS
BZHWlVDLSvsD26tK9ioCTK1FO8lJ3cjXP5nvsIKqRbtyESVTLSbgoOdObwSeE22R
V/XNhFXJQ4BBpeN74aCat8WklYkH07GQ7MhrRMPmFuexHsFnC7gFcmN+OoPD4uEa
dA2MOq5A6cMWWOwuK2Bf9Pp7viWkoK65lfAy89myWZEq/CPjUof2VnUhlky8Qt+I
LjW3r33BSx+0Z+m/c1URqlpGnKw2RqsOcwxu4n9ajmHcAsmMTzVWF1Mt/JcSrDeE
r5OHHwNPFgpQlCClEup7IQwUfWvbGq884jZYhC1BC5DNmmCEIOdAfZkcLMjkfLMQ
Fct3vGI8rgNZbHMhCRQPjXWKsj5eYgq9VqQlzrN3MymFjwd4oFrnJknk1bImMyUb
FptDUSu6jtr02tuy2wesEUvjIlv0ZfwDwfDE2uOZodqEkrIr6SP57BLK05otpjr0
Sn0muF9+prS9khsuCj9GnhHLtFlw37buM610XGp9qADfvdP8vf8aBPm/FiC8EuM7
V+XSDkD1f9LsZwVHkkc6Xr4RyUB5CJzJ5Nzl7Q7ii2PYeYWUQPtE0On1cCsfcstz
gKvwcLRGcwqqY4UbO4Sb2GNC32svkWxcsX0Bz1Dr4HGTJP76qwSSkpBbIcSZEHxl
XxhfdHAbK/9ushJZWp/TSnWe3XCbPZG5uIEVlTymucQHBmCUe610dQB5OC82zjHJ
U51OUExBDk+L67lR/W0q9KTgJG6K6Ze2MLYt5BdH6JK7dMFMxRl3QfOGKpPDeFdK
aXxsCVLiLVpTktLgXjyo6tFSiEOWOq7+JHIBJMPGJYYR6CT6VmSCTdaykaMu8j1Q
GLwN/XB5Mc0JalEn9cCKOLu0Iit75Kw+Tj8wua/p+Sm2mR0rC1pqpDNn6bOyEdQZ
Ot+34W+nZHqFFQq4NGhsMNZOKUsrEZRoErLYAQJi9Z4vOCCJYuRhgfv2s5CaNHkf
0hMkTR9rF1n9AlTQN7/Pn7OGrEQmCGmKdKfQKue5i1RpINO6ZAZAu8WEfiWWWcH8
SNben4aWEIynKNg9kKTQWHESHN0nMyWz3YC9qxWBU8Hqmi3XOGo1cDm5h/6W1xAD
Tx/twj0c0+VDX15lJozGKwxO3wBx/pn71ddM947gH2iAHH95Gc5308IIw7Hfgjd6
OAfZ/eMHP+no89g3YJwACVzLq0jTIlioKquIbVEUn0fI2k4nwUhw0v2ODRjFp48P
AkC+2vIJVUhcgi98i4Iy9CMn5qKWobZ8Vp+vTCr+n1VRGi5/PtKSL8n2q8iqHq/X
P7xXwNFxNIz7JQEk/uATBm+6NlIhSTiIJ5YiqdBuqa4PttV2GOm11PJ7M31j6/iI
ZWflcMluz03ksZgkpPn4EK19QmeqoYlUV62ltXUJ1o2N1VQ2xaAKmmm8swIc0JBu
s1RFUZAPQImerNNH5cghD80yR4TzPjkWPTH0M8o8Hi2eQeurrJSguNYBRwwxtNcO
0CyhAYYgRUnSxqMyEwHj0oykxWoE4CtAwdqWgZNFdSygm4KVS/KZqXl6Nd2HU2Ed
8OvI5Nqgj1Vy4wGFJERqxW5wYFrGx2VjPvsN7yvZCePjorWHYvQyOfIbX2xrDTlV
e0aH40hckikq2AxjcFVOHe6+MklU6ZMYWtI0RChsd+x563onY1t3FwYlBEE61G+A
9dYImJOv3tRSPCoyr+OAaOx/hWgQzPa1qeczo2K9Xwlne6ncPnSy1PTYoSphfMpT
b96domTEg+sMk5piFr29waTQjvS4Vd/48U22G1rtIrBbQ23bZw5atLrY1C6sXvA7
8zuCONOkvqS22pHUiLlz7TctPsArjT+nr2r6liz85h5SEX+Jz88oyNtwKWdbVkpV
MzUlN1gihEKxWJS0pHgCbYHzMfLPWkhINEkReGtPnqz41s84OlkYtz2PM45s9ekb
Q/wy9CC90RSTEFbleeaJEuNF/ZLNHlwF6Ze6Nm3WbSGAjcaWDyUE9lVptJwX+OXT
6tPBCWRdl/AahjLCw52GBZCUlhikJqxQtTeICQYI7yGtipFN66YeBXLv4i1JYK/W
DqgyXiq7ghhM1O5F7eBRMKI6XNQnLT3I1CHyhPYLZZI7G4QMDDNPFuLyWvAtUPHd
bE9FJHwwZH8hQvRVUMKheBpcM7IOQ7XCNo4D4rnArNvnpyoXTkp4GysyeF3aN+2N
HwO4ZbSNiBUYJ5fqI865ivfimZm+usvKjQ9uREvjFfQ7jAEf6pBOAr0UuQq7DvFi
4X44HIsl6cSDN2upOsRz5xFAY6v3tA/asfPHcuOlnEUFy31Hasq/Jj06s4FFuyWJ
l/3J00zz4OPgqlFXe5G7zuoh2A4DZ970tcV+ylekAJI8fJQiQRXE6GYlENdZPioh
qv2nDyeBYejz20uWMgtQkKf66BwjUOPev81i0Myh1miRE+8a7QdpHqetijBxNVU2
Mb0rItJiXCJwhCJlcr7ClLMTLsi3YbOu2V5DjCRzHsld7Q/EuNgvs+C8C2uUAFPi
bX/qCe9vXGF19kM9hBrroGQ5T9dz3xyTbjrQy1K6HTC8bkuPuwhGYoTA/SEtnX+H
75qdZsn/gbidVVowqzTBIW4AHpXThsbYSd6XfA0ohxEpCs0PGRuhtGyD8LbYI3Rp
OTyQAK1msMlGNaiw060KnrRf17SRFhJoUQzPAQTVP0qJLlY0yv18QKI8eieNVZh1
ABm/6OxzhtYV4sySW9gmkocmUqO/vX3S1iAjZadniowigxZ6RcQ4FdBvI8hF7BBU
X5Isvx5ZnLHa9hwcPkItlkfJ6zT9KygQUJtkfas1d7nhkzEu+n1oyyVygLeMO0WT
Ueh3+gF1sJF03EyCzE8BXGngFwxfE7vo3ek6nSY/TOn7aujxqrcnHcDMVDuvyN++
BksR9jNIAZpHwC5kA8XyoPQ1dcCDyM3rjPJdFwygYYYRJ+JGuBRXtZhgtv1l22fh
x0uloXSYUyLcdLt4kpdxGwdqbjbgkN8XwiF0uDiV0hS6z89P4U4iv6ja4ySk5HN9
HylsqL8sJWQVM1oT9CWMJqwRQOfnbNr8GP7XSoarDmn1NY/qCmIlxUnb47QXq2d8
A76sSpv+5aKUer/EwSMl7n2JeWEdoSAFiUzBDrGRg6RTvh2fxwMt3IpOboEOjgq3
fnkpDLA99AfJ5nWToiECC29xSVCY7PE5bV2ZYx5mu2mpRoBE7dNcYUnKbP27HDSF
sf5lGC8mxacYWJmj6mRY3Vk0rsp1gIkd3oYHIMg2BF67x+b8UPy6LlrOGCOmJ5e9
gCq1JldfJ10xu2SkhypzAlCWwpwaw2Cj8h1DnvTONfNQlP5VLCs9QkRys1eLZgHN
aolHDrSTfr7hXSZIIRryq7yp7mYbChW+rAIeEb2Ka5lIau6nfofQXv4g7IBKyD6+
pr56OKZ9TMbhek/FF7QNob5xV9u5FkQwJSdISkclNBvQcrudmPTuPAj8j97UoGEF
XBfA67uzmjOXPoE/79u7/0mYKX24QWehvJx5FYfDpnTwDnKsQ0m335c00Yg89HOh
j5/8LVNxa8M8eL1BShdHJJjYHON+rYIP4fDGCov69ArEcwY1ZCrfu6std8/nw96f
EAoobXD3e+t/rVnQikrJT1VLryp4N4LFM0/I+d9UfxTfhIvpx04P7xglf2yCHt2Y
8QZylte9F18xGMS5gTLt7EAyr3tTFL1CQP+JDvbTFlMDIOcpI2RXl8+PYxqXWALB
aqQQ57rNnb9mJY9od21BRFEFz0IGg2LP7/M/rIsV8cPE18W1p32sR1HSSIRrjluC
56zIF9FsH5tvfJ6jlr9kl+yffpMQuZwQSqOKO9wVBsSfHQnruYirYwwO/Sc2sTo7
NIkNVvbjRh7kE7kHO4rq9kV/qmfnTEWHF/uoArno4gskShMweTJS0czLtfETUYum
behVNHGSTIFNrFtXQwe7qkMoiL2/6ls6RMsEg8SkHeL34cEpTrAn9ehKWMQMimNf
ECso+WDmXI4pttEHLUWhOvPGhVr/+fCONOGgSo9hM7k+yBVFUUm/QHaONlg8mJ04
1DG1txh81v9oDVD+RQ9HacvI6ZeXcBXm0XW+mo6Qj/H8WeJilrVxtdBmVGq26hge
useX48Leyb3A/7PdKm5YYSzMw9NcC6gSKelvRindMGuqwieSo4blOdpiOEpBW3k/
izEd6vDz+8dIj2zbze4VXwPbcFMkhXwoCTHuDcjRyYamkVM+QDoUL7nuaFZA4Yvd
DLXhMjRvrGOnKZjKNYK2WLFzbck2t7gZx9SsejHdqYO9Gehf6v7gKcTigJ+hQ3wF
wC2D/tmGvVzNy2kn5BLkx0E4bfM7PkllkVfnSxY1JHkwpRc7iy7GYbKK299ZzEcg
MwgZYQVt8V+o8MiUw7Bhy75QgdyMnceryCMEs8Fd63z61Lx2Jkpi7yCS1Max4GYT
AotfOtkLsIZ3C3Q0nAZ3rhc7jSblhjXqcbmM9loICiGdeK6QA8PLsu2fDeZxFXkp
5rYUkJRpm7HniVEluRvPf+aQzP9XfnyjOj3zKk2B4casuCd5ebgqhEUCZNofUtor
yXkFua2sPF8qrx3QIPepr4KdneY5pSkkcyv3EEn+tsqI6FyVtsFFhHVOC/WP4+LZ
zjFkWZL5/WCzamFJbNiglnSxOCRUgIui2XGXMUXWIcdhuPcHdvz/R1j8gQFDfmYc
XkOc3N4kArKYoNO2jKqA5nrVk6CMizZ6/dB46chDyK8sVv4zPf5yEZkpic+3vx+I
oaBQInRDwvy2bk9zmHJb9ckkNJzGA84O4X3BEsXaqTdzdH8tK/f7D11aedPru1CQ
TTyoMj92g7A3J8udheKDJHbMwIYyFPrrWb5WYyyCk9gXGU/wvVSKMBkVdrcecuRf
e8E+Jz7w/YiHRdMOp4j9E5u4sGITGmNMIsdS+RlGC5jFGFoK0RDw1bmnUVEyif4Y
ypR9mWH6NZbecKRB+jYVRSLhfdV+pYiyb8EP1Ie114fDjxZymycOkk0egVhRw2SB
GfP118MF22I3G+ofxHxGIkuzM6Fc50s5lOUOINyx5/DAMJ4ZpupGO5maC8bYqNn0
H1QoRKhzLJfwZkqqLN88HGvR6rXRnC5cSDvfZTkoQgiMxGJOEX25xzvRzv900loX
wnRrMlwQJ+/GCFCj8V/em+DSER2oDSpc/nEIzS55Z5yxp6MCSktM/5vJOKx/PIYV
5/sqLNDb8XpwPLFjl0WxZukVMGSIGKfqRLEb17tos3kG37H9l8JtKIR9YrdIWTSi
iM9UT5JskdgLnTJmF1NopsViKqqlD9/qUi+f8bShgkr90ydefXUVc67R27+qOsMi
3xdOVHHS3yaNeIUY+jCw3YEuUC81/qOdAEpH7itaQMSfsqjGU2bP7Rm/O/YKPcZ3
yY4h0yOfscyoziQkR4gtytQf95tovNN0xjC6LwFPV/KdKA+tTAo2P8PLHXeKpDPe
zmYou2CRa+4O+4XOjCo022RTLguUZQR/yDV2XJBjWhyFGlDoNyWNPOqPe4111GtV
iVB5NgcKhP01qJnYVvmrMWrocj+M+nH1YgOVOtGucojHrtWjBpryRSPfIRxf/1Kc
+D+rApD6AGmmt7oyCjFNdjsb9UkPggHOZqOyHT+dhWnuGqLMxyc5ZmFT/QNw0wJ7
PbNPryqFQI5N2ITZ4rV1uqh6LMcu4oNx1TF/pII6SrqXd5/A1LO9qJpdn4pxIxd4
QuTTXrrxtQbz/x4tsmIt5NRIJv80cnnt5oOc0V/lG4SG3w8PFrgheCpvv6n507Ft
H23FyIpdlZ2VvkzwInh3m9n2v3fu0ZelTiyjg8VdeqDElhRpPRsFHVcT+Kd2TDUq
goQAgBn7ztDT6DfO+s115TbmT0ZZiHqdwHa2W6Rza9MDIM/CNghMq7FnpahDmvbH
eoB18uPVBmsxx4yPHEzfhknxkFDnTtKsfpmug8pxdedNK/P+yMZKiTxqrFGPY836
2CHF98LDzEGqq9W/1pfg5NpowkYWg7K6yogaZRlV7Pz1ZKKkB3WZaQ94TTkzVw1k
lkX4d6I2z9MfDbB8i3ahQkhtgrkVajnkX1yTKiLMEAM7Ff38I4xOFaz9AFlVsX9u
MsRF9snPc90qWcrGtocQKnVhhsJMgRbeLuXTMUGca1ECPHN1qQskpRraUD5doKug
unHHIg4uUCXDTBmSqr759HzSkc7L3wAhjBzAfzvv8LB4KB6BMTkn85WO/huxL9Xz
jglIZ2b4qFj7HsUJw3mnICFpuqPKJo2gGyUEJq72HbdrwdgJ9UHr4d7OdBxuarsi
d/MUIcD+dBUOJf4aV8k6v7QiDzaVrvtwnkUh4tkVp6RK9qZUc4vKyU9ZkdaqII7g
dKp1qj/oXHJi0YkBOfYm9oe6SDiJkc4cOTZkzVyiLkpzeWq8UKf0CweZhBf7HoA7
uz6lbwWHxNbON1PQ/lxpv9MzaL/hHpuskuHwLD3+egY99N5kEG+YV8Bc+VCMZOsD
KDIta7/Q57uVUaEsLjnnwGAKaHrt/7XJ0+VJulS8sH0fSOIO76yWHdqFtaP0QT/O
4kWnbtVr7nfz9rfJJpim3xJKI0uRdcRnaBRp6RxT2l1Bz5A//UJ04xqYb0vv/OF7
WAGplgBoVuHAK1264m9LQ2BJ2iLRtjaQfgR6HFZWfXPgEW8Wbeptxf/59xKE5eFj
vp5HZIsC+vi/8LMvSxebiYwLDyezADp4ODWBZt+KZ7zkyrp67AYCyWpUpPR6htyi
folvxDBtrqyOw0ftDnaZvSGHEb+L/Ulrmd/AV22rYtwr4XyedSWV0m2vqtYodFJE
504GD/XS7t3D9bz6+EyUk6s0OWJF0tRJVeWTyQuFrU9qCwVFH2Dg0XeeWwJsDuOF
5/Y972CMEe90BXfi/4yibRfSRsXvZNppEJsJnUj/0zQCFETeJ4+fvgFXuLFqbXA1
g3gpL7nSkHsfxPwFv+7V9/vJTY5lOZfmwSLcYa3AeM4RNdO+PpsIiC/qQm3FH5/a
P28ZTLPdB5Gr2ScFxv3XDZ0YJzXQ56AM2iVo3cNTBbfNkEr0CoWOwu8sOjgtmUiP
8v+lUL1phqUPQPyh64FVDby/TLBfsTmtXAIqoKBErO+loB6yR3wdjY79bPFR3Osk
nN9SUIBlOmQAGQ7bSceyXG0QR+vI0iENv8yXqUfU75dn+Fv0Q7Z3jad0zhlOGZSr
cG9weQRUCqpzJJKHQKG2ljoep1xG8niBK2szJRowcjKQ+d1sZIq9voshYioomsVl
MDc0TXDJFfQh9NV3iOrka/0+L203tv4vm31i+Wqg4bGGcMNj+WkncdVqQyKJa8KL
sDXZR1KD1+ObO0DRneXzSanz1Bfec+KGeFu7wpPKVZLzuJMyz572UVQACaFw74NZ
mfIksIGmBz3x6OrV1HGEto4+y2IPNNNoq8KAVQQqVS9YgcjbPT4yOKgcv3/0PD23
Q3+g+IYN1osy5F5QRf99PPvDk8pw92HDk73EzbIyKbEdZRs5CzsTb8B5s82scSt5
ctSHJGxmpy1hqyGgny9BmwtlDIhB9BGVlE06CzNdCj7zWREN7LZVSMnTmGW4vLoG
wrZvnJ6x3jUiFvHmbXi341p1ws+S9Ojqzs/pQc2559IpLuFaSiUi990iErTZfTt8
lLifACsLss91dewM8cJfPMiJ2hVZZ9IVYla/EclyGabqmC9TbZAPlYidc4oTFkfw
gXbd+nwspkkI7URYI02ILRTMC7z9Emyo5H84/OyskB3PqqNmFfzJTJFfwUEyiTZf
U985cpXN+5Di/CvjZoH9Q3JL8vhsPG+0/IM1iKOX333ede6TOy0yCC/UhuxJsir3
Yxv3dDX5a8y2X0+vlOkqAJiGmgobqioRR2+7GaNCS1l8pbTSq+/0UL2n5OYXtaVl
pwIdvk9eEW4ZSk6Fjg3LLEVz2XFzIIoQoI2igq8hCOTt6agdH4h/Av/59kCL2zx3
R13fjumLFyymkSJuxLYTCqC0h28HAUMeSKP0ewiRL21W7ULYajanl5vPZQjKh03d
Dbh66nw+AgJR1fjIRtqnzQPQssDAbzhHq+RPwiHeRZTLN0PG1EpDeKOw/5QlWlB2
7zyDqJLez3lt6Qtp5BRXVfaxqHlyqWkJlUS6CHiueU/rxsLb9axbNOx4PetDTMj1
QUNXrlRY0BynW0DzRDDDX8G37EuTg1BZwDXdrMACay5Yv72HRSpe8RapfjNkKLV/
ZbgMl4s5b5MCY2OEck/WcSOnVxZHLUfguCoR9zcb3S5qQ5GxYfnyqmb+S94EfAUy
MT0wwlB1co+N1Lb/7lUAJDiegdOh5K5Vj4jDpNktGpqlm4CBF9OE1R1Kk4I+pITu
qw5ZAJmOec9iXAx2mdM6sFPa14wF4+fkwwnp508gPK8EzYHDph+WvD/u5hmIjO7j
oxN/MUX6WP0M1qRoMoKzGNI78uavcPGOA57Deml0bpkTzyquhcurvfUFR6eoOV4p
6QrtnRXy4LfWsl76t49MXKJUC74Qryx091vE9jr3+hLKcXyqry4rr0oUMBVvz95o
KDFWubi1ClRFEgBhzRgOBvXLNEeRG5gt86kXwr80YYWGbdWZBRMKONGej1dqU5a9
CTYJ8IqAFNEebfL3vB1PXe4CMBksCfrvOCs4ywVHgNhKkpa62arN27OjF2LEep8T
oNggaCyCCL0YhUrAGqShmfnPiH84+EojqSTrc/+0zbssOpLR45QWUx7aDIsmjkJR
BYD5j5SaC+0y7aWzoZEtBb4uC2dWbJiLeCiJ7taWMLGsP1O/r7yKCpATYKRUEQak
FJ3IpYJvHQf07x5HOqo3g77fAxEQuoxPPwvJuzMVJiasj1hedJbM4ChnKH3BT0km
dQ+p9oOXDDz/FudKmMsxcRD2Qlr2f+AmEpmNG6dTEC4HbU1Tp0V6l6YDo678Mzqw
RJYsy8S/3B/j2aDHsDqJrlkeLGq8iyqlNG/vLy6Ta173FsqI98kA0IW1EKodttRJ
EVFxImlS4PiV7CGR0r+3NUayaS19oYA6/i++JEExM1crxlAm2BpG5tcjiokXOBPC
XiyraMJM/KHLWs+MbKGYI1t3B/gITCsxzdNyxmnTQu3LIC7GqzVxe6n6DY+DGiWJ
xoYir1UwV4S3aapPftlL/6h5C3RFUgm2FAYZHNFbfEgNuM+VNZ+mMUreSvpAJuMb
tqr7jYVAuTAT+wJd/YwTV3WWcDfvuiuA968WsOXiB9fYtJ9v09lk3vyHzlmCcxh9
HtvQHxWeRT273uaqyPTc2l49yG7kz3xbcOuYEjhY8w8QyzJOcNw4s80N5XGGSEBK
QEsB0XS4F2ArKrwBpFkdmIHjTP8skkGppmrDKmNRbeAdY5xXIPD3QBYgRCEuN74D
pqAqgWexuflp/TaV4n2lUQAwdmoKk0/11N+fw4Rov1UNJdfYqnEZ2BI9143cv2yk
d26j+tRVqVpI3U8QBcwb5UM8c+ICcCSN5kjVrIPXMw3I+HYEwDzPWJpiucbGHeDC
nADzWY2OtYxMherUp2wbiXRB5YMQIFa6ufmUURTlDbz52CQ/qDMsfZeWJhHl7YRV
gfgcy0Gbwz2Oyy76PYbLnjO4foj+6y2E0IS9VbtVoFkx54rBc7y0nOSjmxPr+wxd
gAGDm33JWXlkW5Oir/sbhbVIsgvh00iSU9g9umeJWyp6PNS8VcdRrZjSt1zDoI4p
+CLVUBeSqYHkOmcLIQxASY1oO7B+SKpOoUyut2a8kB91Q+amgHaknTtfa8zOh5gC
ATvRURfWchwDH5hgiTGGIQzuciWZrdrMVSgYDME7YtldgP7owmK2wozAYW9dhZXM
KUNiQ1IQWrdiEyD+9i76CreGKvrCpg97FpBAz8dA73LFVncw9sNofErcsr4iTB1A
fYcQ34jogt3DV20uDIoroSX139I7dC7XUYHYXG/WRe6uTcQn08loD/ockg0E4AN2
o1BoMvhVfm3v0kvHOpWfFTf37wrFl4fu69hTpC9CrUBjclSRGgihtnDxSbrkBMjm
uOHvxKddOZmnWapX+j1AhzRqbae3SNtv9bd/t5pBcQXo8NRB4w8hsV4hgTYS1+mt
V9XZYRhoj+6/nTW6mlbUAKgLLclBCFTvXWyV4JAs7oGRaFJytiQw0P/pLwUkj2Ze
XU+pmwNR9XDGlnBpcRsPQf6jnp/ADvb4cmUdCvFjn2oSli41QpxJHn+yAUuJ71qM
+hyqKyA29eOz9LPnvbxpZ+PkH+tOYomksCbqjhcyJEQ5jKiutu+0lZeuXvxm3SZ+
ag7ZqUrqM5pWmozNI/SGZt7/4hZCP3vz6LhwsbgSDyPW3x00pv4p5XiZ9LlpbTEv
8eXbZGDO9s8YFLNNVZHEASiJLrQVp207pdnefqoa2WYeZ6SHEg5+rcLHMvqB+QaP
aTSJSI5XjIcfhU8XSui0F8vLAWHLzpBG5lT20aEGIV98g8Yqe9cQrhJHfrNIpn6u
WZnkuF6aZwqlolZ2D8kPPTRo7CP6whlX6v5SkaNQjT1NovvLItarQEVbAJ6jYNCZ
bkcranK/cPa0cXcDimpV+2MzGw7/1wLYiB3g0SC/otCHjif1gAyrBDgl9x2kwMPr
pZrNxG3x2qDtrJ+XfoC/+LiXk+2d6NrPAaRz75Es+qosxrm5Q+sLO9iN7nKOYU2t
1p5jgFlLOpNeGVP/+AyOs9Gt7hS8MlcX8EhvPxwvvFf3vaJUILR44tsu3yJfESoY
G/U2T77gtglX8rY/96OhpUelRUljS3TmHOuIbxyXJKGNvJ+w2advj7TLN+MQcfJY
k4F2bFt6fuSRBELmqAlMuAOOWTkktyn+MSWfJSCJ4UycNRyBCjoF2oZc/TNv8C7g
631VoqN7sJJyGehjpv0EGFIQMxd05vravBYditI78rq5y1gia9GOmJLNam/ZRAzj
1NgWoJ1GYT6i/XLMyDMOh0vIW8czah21cqrfwIGlmrX0smFFurQVppEnV8fSUChJ
wUYsD1UBZ306+wr/YKL/+0Q/kQclo0uf8C/cv0XMe3Hu+jInuar1TXuSTr+ktK9N
Yiea+uvIDihHCBBFwyF8CafvgXFpVfhY6BdmOJBE4K09gZMjEtitm1vtKXNjdeWH
GMtr3Y2Xet1cyhRpaLoAOw3z/egyoGf37iYFYZBFcsIPcn5ThcM5VNn7IXNsmpgD
w9091+ZEPi+GILFI9ENf8hQe7LnUodH80mzaT6mhftCNoAxeZzNNUn+85ASrwR11
UBK+1YfOISITrHx7vJJrPMzNBNJdQtHMQkxVJ50oOrhqMwkCArQFZkCyfi5yknmX
N0K0ttysuSCbwVSCGuhUxrURNdsxztdjQAsUVUitA2VYPaaZw1QShOxTi94nFKyc
82MaQWt02g0e16MRarpkvVyvZuVzA5Ew8vZSGN9fF8ZX9X0CgmUMC0aMGWrYvUOY
2UXXoJ8ELt++/drRPrIL9SMYx9CBYM9jqkV6TRYyO60v0KiTGe+Y182YT323tY9b
VZvTXHVdkRVQO/wejn1pkxznR7TYXLettfvOBlUmIDzJ0hMMgcl6HkijbGTpBkBU
rt9VZDRnTDyhmF+QaV3RGAKvm64Cn75qDsiGUHBe6OQm3qKLtUHDXMaIAFh47FZn
Ow7UJz1XUv3ZCfyhQwdyE0M2+gPBJRXR9hgj5dcsr3MIC+m4U8bjt6AEBeFgtEK0
dC7G7+s+0dDeCsCwm+8OGVHoR1dpPBknM7SeChI0QTu3AQ1qtNWS0QIE8CR/yV6y
I4gPL5pluiQeQLxezP3ey4K5dfkaa2VLUz4UZJUqBG0zEqB5dHhr3Js+A55Lvk6s
rjJsao1uVRxBXXRKwDHa2+q3GqMqxe9hiBFgZkHyYp2d7sAYUHiGL+3oHqrdv1ed
efoZP+pnb+6ObwudbPi04NMVqoVqQnrkx5/5/4E8YbRqjGW5wz0a1KEf21B30t8e
qXnWwvxz1sU8FBDFIIF6MF/G7z4cQMVa37SR5PRozRdWQEiuhfamXaM7dANAJ2+A
vKBezbP7Rtg82y2S6fpb3atSbUQKZzjvOYoftfGq1vOn2dQWjtA/WeoF4PNw8JCr
C8nkYk4KiPPhrMcdXB2a1fiCqebAhIymM68/hxSch9nn5AaVna6ydp07xrhwU2aN
LEn4donmWvS/XulpCo6mcm7LqbDwheaHNdXYbL6NMl5PWBhF4MZ5pZqYNjq9tcX7
WZyu/w2tNerSCmhIkEn3H82NQeeRRQzd3cHKdqZAL6zocEoP4ez6TL6Bx3/KP9Z2
TsLS5UewG8YaKdNKfyolwP8NSlaMMz+dQTnav1rsdAeaqnd8b2xA9Xj9HZ3VRd7U
PsqzCfcZgSoyzae8LmZrV4p8dTDO7wXmjgh1Cjt/aXUVTqfqG/C3ogao4cdLElHz
dggzHLX6QAdabP7nnHjyCfoDIluc2xB+784KZau76s/n9V/UBPV106wdlmkWQ3J4
iOYggPsy6JY6rCEQ1ACz0qqePXWKnxD9m/eGOaX65sJ8piZH87/y5QyNH2UxW/uR
V0rFbtstBl2aAi+5463z2x5wUxUgTwB2mf/QDjPVuNbVLpskQ6QJSJpdGQiTOqw5
eylLMVJIRRlAoAFN87oXSn1KX+1ruqwohPT5hCA+zCMDL66A7gGrfA3Vmz0ksGMT
79SRG8UCXYE8gL0W0yINEh4b9J5tVLnN37GXAv7GMZ9iJRoMXOcJNwXdRKIQ8Tmx
lagIIKIqLhpYdfYfDQ4QeL0qkO8DIEu1vb1zNXpgjbEBZHDlD+4h+THz9yqzV3LR
D2vq46DtUqlmM6VtP3WZ1spOnsuEqffTgu+o43ammmLpe/MWEVJsV03prwtTYF8h
ORi7FY5nTpqvBQP6s6gh/TGEtDBhttYCes0B7pzWIdmyQwY1ShUFgoJLEVuYCAk6
TssL3UVNciujdIdDyVgktiV4+FgObNBI8cduP77q2C71YHaKv/6F3HtOfrS+Avw6
NuFrHVxj0cfahW2brMItCjFbJFa6q5+4g9+fob9T7TK4bpXjSPhjIf+AXbUH4pDd
1yIyoQjXtS8xXeaNqgdxH04FAWH+IqKk7MHmA8kTGEagz4z6Eez9KwF5se+AdUsF
VyEo9XQqmfXRFXp7fnn3veoJpYnKh+xtLtsB3ePcssV1wf0JkgiRorNLdZKOfmD2
aulgKFbxyVrR8qLDb0KueqQM+pkm84VBhZsizrYR72Ird2UgafUrwBe9z+fHqt9t
ZVeJwya8Jbk0YGcC7GpiSG4lX3HpZBgz6o21ZnNVtD5XiJxtk1YbrQ+m40CJ8Oxz
7RTtx6Fis1VK6YXyO4GTa+9tSIF2njCjEwPNF8MJfkkuUtXOjOu4riwj797y/ETX
ckCraYKMNbBk9o0pD2o3V/QK1G+XXkDXy7xQKXpdTbnQegOKj8jU8O8KOI7LhsJj
fNA+qhPByAJruvTZg4t/BW9U+jp/YmkwMxRFXAo+2EtpS0Tare2cxUCfvMbBugB2
Ad/kq2/G9hyTqAS0RGMTwApJAAKuRS+zXwF5RUoZ2upL7SJng0oOsGMlbrNJzVya
JwpXrLMGA4+nsL1RSB46s2R/lOcTTSIJ6QV4MVGkmqhGV+tty06Na8jEFw4dE0do
FAwXEKexjMxOwiD5Xl/7EU8eVWWxHho4blrD4gAeUZl8hjxJ1wHqp+FX5uCtdP7u
l4NpmK2wt9zbaXQG0gFaHOteJl0P1E78yHookzKKR30QGytgjgW7po0cQ2TjRzb2
qAWT8Hqp/XdUqsKdW9LJtYTcfmdx/5M1+3qj0rYSP2yurY+O2i29fObzJv06HaIW
yN7e8r+mnxmO967G9GJRI32iq9XfBtvRAVFcINXogSRXkvf1f7KOtUyBavBQaRwg
Xxnd4vLyYmYO6/7RSI8iFi+G5yYaYwDjQ9mRq0BI4/q0m1FLudZH+PJwx/J+LpiD
AkHfK4HFuqp+T8q8cVLXsjt3aoO0p1jrr/OTyO8RMyPQXF8mSS5lOecpj9F35G8q
lQkezFG/Rud7LfMcAFHn7RxL9LM3ZOOMp4KHc6qZkW+0O7MTBoujT07I7tOGCEFl
goC7784mRl8xPFBvfVNFKwjD1eIOcfEshHoL4i/twRQV9hMWF1TeqzCxIGXeLXlN
H25X/PfSi729B62FLEPU5EADrZU8gdgJARVGxy6L7vr/WibxN8pHS3zmqlMqwRXt
yR4+LP7jkJJlC6u+2BKcruQV9KQdMMvIjQd29222jwYwTBu+BLzN1czujyONE8YF
PxjJ4JvMts8B3ZdQZMTGlW8TVDzSgNfcKmEiTbi+fgxprz98/BFPtz8xd0yKeQNd
IfUH5YGhJjvYG7iRVvTT57/1lgYmAgFCWnCg2+ufFACCBMdXpmc9f9Ld7iivrEFe
+Do0346p87JEUCIitanivkLsxignw3B8rDJI0dXMrawtw6rXFBPzwRBV2ypBOnoS
fGt5Y4jecymAKuHQ/rkycmsFhGLKbY7705N53mv7QCe2exUH+pJ1lDjXzKRU8rsX
XgaEdt2lpcMVjXml7deE5KIk1xopFG6dEBou0qjYUOgw06fEk4IlVehf7DM+9GXB
26rHjvaoayESCsBm+qMYKJKqeC8uG/D2R8Ei7eYHuUN0X8NJ3rfPIXwU39ScjDVS
mXo0iOOnmtyuirRe+Gp2eLZa/HF8Mh3VIlhRMUOZfES6pEp7Q1dmDDGWxWDJbxMa
mxp7hE510ZfggJnD15LrPgqmvYY4+hSnZzUL6agJZh0GMUDUswdQJFMCkFNRgCvW
lkptiiV4wxfQ58iVxy7YmP4YNgVqzh0TftVM77dWa9WobJmtHo3lGJHJamPJlK/3
0KOV30eIzPZeDIkdnEk/v2fHvnLCMMOeOMZ3O0frYsxaZppoeUC/TZFZg9THySvi
6K7WQN31+y1bb3l6iNeZ8ulyQjvviHEGbcw2Drthcm3D6iBRItEQo13shgKFCr1/
SdOFR8vTm6f1FBAYieual9+xgBJ2N8NHa4QZtf3CQ0RYfB+yyxZLbrhfZI0t5C0+
NukrzjPhdz/Sg99SbExKUTm7t7MHWBS45UGryq77NsQPu99sK5T4Kg3HPijpsD17
7iYEQ8zecgrdyOxtOIiJ7lgONzPAhTqaIK2aoeeSffOZqaLPPMCLoq7JNsx2AkGn
FFJ/64OzbAj8H3ZQbHhYa70u+2oTzV/eE/Wz+fNW5KfGpMy4/+CbD2ihWRiBlgS3
BghMp7eLuSEfVj1Q7pgBcHBsQFoEXyGCmpBg5ribajPlDxFA/w0uLdSuvxA6T4Og
k8OEw9aU/imWnN5JcZTRrI5pjtPC6fveaiWUzfouVxjd7MY5DQsscQtEbGjPywSZ
c04RsxTlSORxx+S4E8qalKe4sazQ+oZ7pkxtucDWWVSN7YP9HUx5qHqeuN5mtDxs
r/ZIU2jyEVIzu7E399qv5mg6mD+Ji2HFXKZKO4IlJqNoQsQgzbVcIyfQHlTirJ3r
91/EkH49v9QZWWLlEJebe5NQGKe1ONIOwo949Jd+p6i1IrNsHj4klTT7TZangRxe
F90bqZjpe/m+GjnbBhSxKuWrheECdpiea4nVjO29kbKONJn/b7NOrq4XTENULpZU
VygQHxmH0VI9xDzoyl0XCxvWOUD+GtzaDktu0oZzOyWX5xYRvDIsHc24OW3Z0K0l
NfzCEMPlTMsP8gZtuq1AmRDl4a2+x+13Cww/zpbZ0al2QWtQHh4nOuG1LRvUABVA
fxWNZP4wTWyJ37znsaPEJqYhqT6BqOlF+q2pmaSVp89G+y8La7XyKuFjWB5huLdJ
qJBNUCGHOwiOtM4F9KIaHFbza3R2anBweXTch2poTqVdVtta4Cpzj82zap3/19Lg
Pe2i36a+SOyzYXxkORx8/QxLQ/Pu3Ryg85aqASvw+RWHK3Auenb7FL5laBL/DReX
r/yWTc1CTr4dw3NETTrcYuvDxcJsrJL1UzFlf3oZvtdIKjK4QRugoCMbKxa7jZra
7m6r7OK1Qw4RNAlqeWhdL2jxZlXpMqZFzw7IRmHz7Y4MzXvv7akHyS2ugwxD6YPQ
3Hlx0apLOj6MHjzlVti/dq3ddVPUBZkH1/rvJ2t7Hb2p+JnDGN3Zm7LCOBNdQtUD
Li4mObTZd9RRiaBKjgwqQw3cZ0BaJrnuaWWnuuv4TTRrX3ZU7loIkNDCMIbe9VG7
09ctVALEex5wMJsL+YM2f4oetNpFKYzMhEW2THHl4Y8K/lZyeqnHjd3ccoj8n3bA
n9gKb+K+iRsB8/tA3l123hDnby2RZE64BydFRvgvDR5+9EFFpnDyydetDh23bCim
pEeI6A2F53vX52CFwXVvvs3tDVJlsDpB8ABcpSJUJzw7diUI3L25Ive0XvygOIkm
dHL3yNoDh1Xp4T11X0mIrQL4Gz/5Dz+FihDqTRa+gHcmocFJvtnLmAQKQKT4b7sf
vNNo0DCSpvYplPZyTskhVE0Npb74Q+H+vhWXZ1txqNlMeM+spX2gSTFxgSJIp+K0
mWeSH6r2EzC1OQGX+6RRUELi2f7QEg6Kz2wXq74BxftP0dTnVC8ztJByJmuJFCmD
EDbD93m/wlKMCHH+q6EO4rxj6STJc6AjykfbXSn/4wJlSGyEEXSevlXIVpvUS36U
M0zJ2mL1Ws5vRrfx7hGAQqVePsaZV+d2Bls6Ty8KXKvNxHHMzHd9RLPMJv5K4MLO
6Z+AfMO9OFqpoyQlXZjVgPBJ0kN24ml1ZXD5Ra8K1/wTig7SIOHXiXTb1DRyiSjL
HF8jfj3keRZa4Zhkkc4bVAB1mQAe0J5/oAtzij8Je/qnENft+504pR5BCFZe836U
XLCVYj50cyq5tgV6ZS4QpSl7uQzwwNSzfy0DixS3MJAmsseJG622JXzEMBTcPmcP
N+Bj8ojaD3HNObKSoVPa5+H9qJrSv5K8/LiE4xVATIKKgm538U2E5nTzkeMTRP7f
JtbmwUEiu1+vDkB9SkkdgCQfO8un1m9V3mr9qBz+l34qKm1KyBFDZmu+Amj9tx7b
PL82jbxa5KQ51OK0rpIbuvBAcl1ksZGXePNlVHjtxfxnm6QPPQB98i4eakGNNZu9
OaZYG5PfhvfCgYIfdnfGu6uLhmf3q0x5ZEcXI0Bq9ykpSvmBgwUNK+f1l6g59ily
50eZ+8is5llPNYbK+3x0t/eENXIfYubEswQJypwhhAPh+PfD4i6eNYG6hHewsWLL
wJKEFTjuVBSyc29IsCe0q/2bwXWKTVv+TUcx2H7MUAepfq/wFVlukIYNKGJGorXk
/tl9t0lZ+QnTTu5Xbvxq0u0MwlXIgAQQTCk2ce9Kmw0RPbR/wBVat9IKyCe922ay
GNM+SjOOiwOoRVzPvtG0mDyXLiwcMdswvMcl7UmLlRkRcrheKlSzd/XJCVD3tp2R
F+Req+FxfxquzCIHL+LlQYs9FWbJ+4GACree9NHWxzZ2pFdeOYGrN+DDmtnP9E/+
VaQ6XDq6y+6+b3wvIDccaqXLW+cEy8obX4Fp6orVYZo1H1P/alt0vX6WhelXNnGZ
0MMzwHPjAcYjbByvQHG/q7DbBOgtJRhLr7O0kGuaO4jtboF2OxMVX4fpAN8+IACv
ciVMVmz1R3gC8EcsH1224buIdOFFlLNZHaUsibpNru3M1MXBTqSxtFj1PXfVlQVM
uk+9Rwat7V0aD4QeCIlKsEsUlDkpVFj3bJHL0fSsFF4wFXzMxXh5beZD0wse2cYZ
0PaTmubK/SH9YybWmq/7HdvYLHvDKuh7FXRyiLS50einsvKwA2SGW2TKix8Ksz3l
SiyMsclykmeTajelfXkfx9bvK3i3SRLuLZvNBLNeQm2abyQPE3HULPIbA36LE/aS
WIy/UUV8COT/XzeXLLOAp8NooCS0Q/xjM4M8fuYUB9Al97r5Pr532THuoqebV+BN
Alsy65rrNrnrXt+yGTldx1w670w3ORvj1HoEhXP2uTkQSGpdc6//jIxlt2GIrHLb
Pq0NxojyFfKvH3MHAcsW+/EkEAodSG/AtHFPB4Gcr+qWXT6YhnuKjlb8Uan0+qvZ
bRd6c5nM+9gtOq9FExWccEw2s81OFckQ462ktIpItg4cYHOw+yJiTUPc0vQ2CM8p
6kQvUBzeois27iLS8A9/Hn7bKEEWgOaiemdCiKvAotoS8yqJmO+swA8yKq6bkZul
DSHkEWE7MS9bztcXfA1qR+Mvz5Az2j+moSMy4A2KVikino2YZQI17V4+w96H6d5L
CYllkdHMeG1l33k0NNX4vzqW1ySULEobkdpP9A7lV7t8aug51H7VRLGcy0s8x7dF
JjQyfK5VDEzVIJg+ek+xRxQ7gMWUW8FKwga4x1lrRH422rhb3WuL7ju2KMw+ulFu
tFQEEFDVffnFfd7hzpLvo1C2nebVhIZTQtwKWzNUt89lsmfk5LiWr4O7kl22jw8q
y5Dm9/mn0iAYxP1M1dV4oGCACK7rW4pQJl0g7fhW92ZMB5ootEU5XNXvF8fH2hXS
EaNvYMy8w/ucKe/+MW9ijp0+NwYxkuXkPk3z+lVHQA5Mrm3/30xIlcBLafzY3BOu
W5Gydnhp0R0ts+KXbyOhcZnlwE0aHrGGPi0RuL9nSX0ctkLHBoO0V6CV+TuhbfYo
kLzSOljdpTOcPjwyzk9HJASZqJALDedDbeFFAbYNEneSkOWRQQ9dOUDEIEZUpTFJ
+fwFDI+KPLzaUbxz+Uvi8aeaUA7IQ3GZhy2OLn50RGBmB5iL99F1Sut9FDCGNknU
SyqewZ5yu948iynHR+VkUk9Hy+zB/7MoaToWUj9VI6fCW6RwtSCq5eYmvK2lIfr0
c/kpUz1vLNnkJk6lvJD0YEUtx4uKAHFltSaz7/QRwQYD9ubl7JgAo79xed+B6mTK
56DAbQk+Yn1kkxI34zhL+oE/5rknU27uRhqfVgPUGobCHCowrh7fXv/3JyI4KptA
NXD4cHNx8BqgvMoETCI81+4oeuD76UfPZx1Q+Alwg8LAwkOKU6xRCkFlI2X2L40G
T9WF3pbntWoiBpq52JRKBwwSZEtXlv9z8YuiSJLK9T7Tq4F0425IZDqZzBFfyA4I
vzpBBhvG1pCO/6MXvXo0/rjpcL8h3nCTrzqM/2TOzRaf/8oLcfqaqHmcCXoFC3yY
7E6FBOAHuFIRWw9BiKn/duaGAevzpNSFJldPSkImPQ3XXd86lYoBO3nZLXbgq8CX
LDaOF+SVCm8FU+oINU5n5BeNmyw9tzavrkwlqg8pMAvR/lyV8o6o2Ny9F/MV/IkV
PTP2yk4t5H5Cd5vnglll8ZHEUEGXsMCCiI5Yse17dDtl7g21j4OTxkXF4Pb3FOCh
wk0bkovUTEdx4cmwoghSgNFr7q2vSG2RPrS4o8+SIC8D4XJ7jHz2VaI6cPYc7N37
ulTdacps5C2vmFD8MuyzFrlIG+im1awv7H4wqxJZ4DMEGVzZA7iZ+4jw9ePhjfEB
43tTLjON1GOu29DZhZD5Z9fD9Tf27uZokweLBdra4LBARmJrH0wQsoNZHtK7vymx
o1zR7ciN/8wrVHy5wBn7oz2rAi4he0hl0SZFoFt+gySd2TFVBM3U5WPA467PRmMV
laWBqYtWg/1ejzg8CKWvmR/lFBAwj1dfiUEwiwecoQr/qGlR4zuEMAq4IKI/NOIQ
gEP8hdCiYGbOPYNc9itW5fzkoc1Y11n8MOny2ZGe+zEn2xtggX5KQH1PZYSze4Mq
5fV6T34I/aXUw8HHDXSXUmvEEiHU23W5JzbzNZYPt5tbELrhGo4QowmM97x7QdoW
HPcajh1B0x7anna/ArWzyYISoF4XgLijHZqnp2+clYM+OAOo4xTXAQR4A4Ov2sXS
IS/Yzt9/7OSvZ5hWuI6usXPG+VcfYhB1gbmewN0jiOv0NQDF1/KtrSU5G5rf1bF7
tg87shqW5q0LYfQvYpJlRayLyq63GGd1XqfdWSwePtnRuPrew4DyobhZykINOFCv
RXMAQvhEDMrCIOe+kXFK1xVX8opTygxtXBQCtMKCdlLDPn+sj/TKOmB7cTE17pqX
5cbl0Z8wiegwjrZI330adyeNijfTfuhHJNsqT8EsLSfN3hPzze48NwwypzR9YLZm
Vrl/mMWB+J5DZeoq19cGCAzU1SP22QmjpYSXDbHYQtvrekr5dGOngwxNUXVWK2fP
uptWGhJAkDTQvQEZ507/+I20j7iMrHZMBNzA+9r0hsFa/H+lU/nXcixFmjQQl0s7
PwD9f3u6V2khKQDJF+kdxv5af7IZyqpLcNkxgQDdSVp9m64gwLtyxuN0TovQ3h20
7N6cMPkap1MFqdBVK99aD2jUaAnmfGIx1AloM5ghu4NV69WPMp46/ClQdlNvno88
5BxTwJrFnMX7HEX7J1L2O8eb8C1JropfTln9cB//5gVjeEjy3vbzb3dVskoUHL1t
IcK2Z/PnkDMjkC5J8L0H1DqoDHUdn5R7Q1EPdkadsY6xWwXkim+M9B2olwU0Ea2S
KotnNH0vqMiHkEOpeVdM12KBBanXLYdp8Gk4qH+C1XrrVE2p6RMf9M1TYWnKjyWJ
y4iUA+1uun90iNYUao77kEEaPcFroemVtLfFb0Y9/ZKUmSFva1fa3Qvk2H+8JaO2
DtfsMCwQNGT+pEG9rUCpyUapZCzbByqjjP10jIRF5AX6R7Tx4NH6KuG3zMR/ARtY
C2RlOd1531Chh+7E+1wjv3rZEoXxjP0nAGnmNyVIF0J2okgn5a3/G/XlCR3tWQgA
OurWy1hsy/OI3Y0eJevSRlp6hGjGVZDYWYIi68AUYkCO5Qzgji/fjn2tbsGlzzHd
usOjbCHdKENATXyFmkLzUJqEbNd7MB/Y3nhi5dvJuoaSsu2HZh4mLzJtkWCEXoZv
J1FDHs7dp6BccTNAKVPxAmOCNoCje/d4IN1jz+ojEFsliX7pYwgiy6LAQfvDgyS0
W4xzuUp9KDyygmx3JNHZHYwZeLTEJmw3aR2o8oH1QPmGr+ruHjUROMWpXyMeYdJo
MeJuXvSdVSSVaPJ8yPGMi4lFYEEpW9W+J4D3KtV2kUVxNK0ym87iYh0QqnycRRvl
Bw2g72hFBHW8ZQP0m4saCkQR1+3nqmJxSkcU3vKfg1jvMxut8qjO8nUEOBGybBRU
aDgwkxPecxHX0HF4JkXAnBl8G1KDSOahznBP7xOY26vKiitghYpdTtEuyWwXOFQp
kXPreImFROI3MmskbQJhsjSMCYOmcMQDX75B9Rr3FeSDrVJAevaP6OhZhAUzVEDS
ddli//tIbkWI/EbSGJIU88fp5yMYV6PCa23WGYwrtYG3d9niJwgEHu983cR263gq
gJ08UVt7RWUoLy5+rxHHq6/lgf7PVhavhZzthlON0UyUM85bEDfeaQ3SIjPJmOlC
6IEhwRkXCovzfrfcGg8g5WhN20ojEaC7n5K8T2o483i4Q6YqaKuuQFVB99TPdfnh
vO4TTSSBNCaravSCW6wdEjKVD8np7rhWJEzW4EMggLM2vSCoyWZD+w3P/yvfUOtW
GIqnEDUrvA26wJ48R9wQ6Rfj1HiHVXDkRDiF8Dswo5VsqV3RCM6nHchc4Y+8JgoE
d4hBvL7vjIswiY7S7HfdFGa10FIaTOOc8E7Db2s82Qa3xCjtcNE3hLDStNmg0mBw
250uHeGXNA7FTfn65PMsqDjKhW6T4BymMg6JiXpL7jJN1Z05iDsUn6o4MO0sV/Bc
0hDyk9EwJSKjdZpCt9RIS0jrL8C+SPlr51OQqcMlSaqq+Kt41jU++9GiSdeYzTky
3o21V1KiFJjVPK+dFnVKstSUkJ1IQXcGhU89y7TPl1PD4Kh3J6jOX3xOSMgkIjoL
h2Z7wB19ftePM+rRMw5LEKd+OAhJEPNMjjxNLU8XNqC9m0AAh2wK24GNhV64igRZ
ltksPuz+M+GG+CNlR8d7sjUCK4kvDPqMPjCQF0QAiVBv3wOQY0NIVHp0aqbI7PZM
eOXjvVZHMqkZb/Mi7caBxjkrrUjSU5kK71tarIBmRRP41lKJomKsddxyL49Fe8Tn
NXd+4UfUA6lyI1QjiEAfVrsJnYkv2Ls4e7Wbmrd5WKQXaXiNvrBw7NUIqCk4ukdj
263Q0E4Kc25f/QCMDswDQZiSRQaZqEzyH2ccxIISnb1y8SfuKICeqzsweZQlarux
0RqRGrP3pAcRPEomHFtQiU3mywl5m8eTEY4aScABkY3rEV8000vVUQplGT4WSkgn
NtR+4pxxHFsiG2/jrPnAkp8mqtTEGJ1gwP7SRloZ6SP54Eulrn29kp0+VgbUiUFc
U5Z1fxp+WjIBWN/K3IUer+yLCeWoN6S1jqGXrF02cr+phsRn76hYyaEGRvzeWq04
EUF7Yyf+YYUMlSZRr7Vgr6aoS7w1DwlHpBA2GpZ/f6XWCd7/6uZmzu24HC4RxJLJ
I6PYfg8GUuvzL2xZCCztFBZSoIdkqjj23VTc+p2sItttrhtaVS6IYQxNhtsJi3oA
nERL6keg2ynu+9zkhTNpyIoM0ITBGD/mbrZgs7PlmmPtwiLzPg1q4GRk6yXDnyFq
6VX3Z7I8JC3dwUUS6RC4nTUbuexTdeXdfSRKsiEJcnlCtysw+WhBzjBbZENOoOfz
Z+oyCG52W/bs8M47vs/tVgl8HG1fbqYsKJs3bXVCcBinCDXUxdfTkD+L8/hnmQpI
rHJo61VQ3taB18afYM6CijTfDsTjYxzWqGOhJcKU0ZRjUtYEOAmI262IA/nmPDqi
6bgXUKalC+M5RdKD6fivMG+PM7yQlLSxLtuKV9IpLO6OI77WLwCHE9ioAGCAEH9R
WOkBTKzWsFUhk5AsySJBxlOwuFfkbC3ssOysZlWn8ESx4OOnDytANCW2BFrWylyK
uazcq9AqP3uETnmMR00yIw94IgWaQKwCPSPi7ea2z4GAJOq2zbOspWH/V/vfxkF5
jWz3zLpci8L3HyDgVnT6TcWgzbjgstdJFh6BMsDklvJOrG88epUxF2mzVTJz7YWf
+IYh3skvzaWUQNRtHeRVk6SShEgK6Q6lqRWqASarqpc4hTGDlAUyGOqyt75eDo2v
4sUpknETG9FutjOcF5GcwXPS1wygS21lGVUZ9A3Qv98oVrSkkP6myJ6dlO87+wrb
EdrgeZLDLIMeb6AqGr0YnOjChhpgy/OaQf3OulYM7AI0CG/GZIAvkaTlPtsZQ3ol
h8kdyFVLa2radkHJG/4Tvj9uvXiXQOw8ypY4Excnpl4LaEOE1b2ls3Y0+2LyQq1l
TYPjRhKY74mwZcTUuqnArIruHWC0z+EHeqN75rwdWEs0YSXKAffSRPgsZ01MuR/S
vM2xdIWi8qCzNqENZUDGjk4M7XLzZM2x/cFir5W94nKadprTZNN2KZdPKUWmc63Q
edfiT1xI01oPSP9lNaRU/3qucEGYxe65JXMIwR+wX/dVpSopRdazY5UVl9ZalIKd
u+MfBbQin1j6w34zRgUNMg7LyxuLeWgTlcxoimqUbPJ1t7+seIye8LmqIe3RTByX
zcFi0h9ql6pyeQrvLr+41eWuka5KBkNj9WZLc3zHTx5S+fz84v/WSDejS5QnlsI9
4X8TNs/JheeMrWBqHpYNtJnAzl4ZOUaf6XwWrlrCBlKMuaK9PTG/EVeb/ro7jD4y
L+5me+X3w10g8EQ5iO6mZKPpL+0dy2SAS00IzDHYcjW56QGnmN9LYMw0aKVdTo5/
nEUmBa+w0znASZ8zgTJnW8kJfzvgACeIasEVLuRWxyknASiG18P5N6BoyKSBzmhk
uyox3KaEAhxreUsrUouGQjg5W5UYTopmfZBNW8KaWhZsZrmDNWJ/Ot5kspk+zzfD
U3RsNonVqqG3FTskcjFrc0kO8JTcYCFcTi4YP0kAQRc9G4cSnao/guUk9HKhVZSG
x2u+XduyoCXSSCCMoyLLpUO89eI9K4cNPERbuYnXMwX2fl3FiSrvXjP1bymaZkMS
uU+v8KPbkpab7WJxfrWn9cz7vLbzneM2SDJaKvvIRfC/H+vukaI0b4CVroWRnUBj
13wNDVRpyKkYMXDwiIjqEydn+1hik9Liy0yx7+Gw3BTw2gjNFtRhptxe9xWB4EAu
+uNQLY+GdQOy8a6zdAt3Y9goMq5TP+2PRA7TNXWAZnIddkgDxGOt+1etlD9tEBDK
PNGERqiyimp3twGZiTX5TH6Oi5uwg+j6xzBWbyeSTAM/TA5TYu4A9H4Tq2H1OhS7
DPL4z4TeiTTff5JDVFHDIIXrxPvTSDQd0rLTT+m80NYoqgSYE+EtnvfdQw4cv4cL
HLh+ZcihOznL46xiZtLynK84UR2TkBsCgJABnThuiW0tzT7wA2xIe0/ASQ5fhjVB
ukY22zgyrrIXhBOLY4NdzuP2dziezprZwdX+VpH/6G6QLIrDrr8DIhCzxZSvDDVO
wu+jbqN5BsG7SYbI4+KTWtuEgesDF1fjXY9xGTGz3anfoNNz/kO78C492pweNchS
ulajigwZxcWZo4ig8gD4zmwKGduYZ+TUXILsPAXKWCJsCZo50nsQU3/RHugn5ZSw
WRlgSykgo6/A6bZpH+7tFgoF1zKB04/EtUe7pFkOYDFCIRReEcNMkIam7k6ihRFL
6FMoxHEKWw8vMsdfXl4JwdYEe4oQBatJChHx4oLQSZa/9BZHNoeeXWojQ259nY3p
7yhEKo72MkzN24fTUluPX+IkE7SK+rVqlkV1IeaqxbrNipoEPZhJ1RK5Hdkgx0c4
hx5TpCVkBswj7afi3iQsyzxhuHCLpr5rPPm3wvzjiulZuFvRYTfnEb2XhVQjB7fJ
7g5sjl0oG0XuB07kAMZShzSw01AIP3Fh/l4ai7BQLleblCcXX7IYQ3edyG/mDmrG
KfyiVbLq0WU2ws0KZnkQn+3Y5YGGkZPtD+zZ4ZU+x8+csCURfKJcCX5O1iSRPDLP
zDsSIo35b4tQU4Zd8WCtj7lqJdIqdDZObHGS9aPWdZjQMkjQzNmW5eL6huGDeFhI
i0+dGAXX0UNhr6TJ8gsry0JWuaYt3yxwQ2nil3X5vOF6jy6zkKEXrbIiYp34DaKT
H9bSfw35FU4bTMeHynSk3yu/IS9OAjOjddwqga99T/BdQ5ukYlqSSt/UZqIUgAqn
p789PZijD5WWdYcXeEFMzv8aB0EgSyiy/OQ81WcjU8dCFSOov449SRww41hk2fnP
dm/d9mkSaAmlJ5BC8VcmdB/KIhq3jNLtPT32S0JXIInSsCxh9AONbhsKZDqhvQlg
QV+mG8gahyj5ID5smvcMqg1o8uXDhtkMDJDgHnzZIEti0BnyAHB0ijFS0Zxy7Hrv
lNPwDmhh36PTXHC8FeHfvM2MWNQU5nupyS7M9LXQXFexA+nC0mdT6uCOYbZPEtXd
Zx65EqJg8kFSOqc2n+i9djqYNSs/7mIyFPCFMw6KquFqgBXMmxqCsdY7Pht/Pl+Q
UXM1j5LtcyHNiREQBJMUtvmAkVSs/c7ZmEHjATkFfRZ8meQ0rR1AWLbJI7LaoCn2
LAay5yGlNhzKO78jHKiEtP92oK9joTziujupvuHEuKv04b0tQvqMdtQo26RdgFYx
e/uwJpXea9+kccZgEUHE0GxIa6MnValpIIpPHA1h4NHRFgl+cIHaJ305zBJ02qNy
96pgALKIJs02PQ8Fat8qhIyvno2vh1iUbFGvWGYCIWDz93zuFZOzfcXCyNXVmUTa
wF8zuILzppTLYSUrT1O04h/o4AjopTmNGd7SeNuiQoYzmC5c4I0Xxv5AWtpJ8mMS
F1bZXdZup40QZJ32mxb/05tRPp30zWOi00WWPEfQslFvAuyIB07i5PR0+tnX3H1g
yy+aJD34orxHzPBiZAstJLpN5QIbqVJQ8/YU0hZihg1Gv0maZYwk3kF8h2IG63uB
5oXvmZszRTJAq+DI8km6I8I9AjiHjlP8XLXfP9+I/N5BiI+5ykRkmbpm/DV49cua
t7eE+XX1CWZ4B3XXKVN+/Q5Cp7AsK7zZrOhN+duxtZ2MK6J5pwHqCGFChAYhfAIj
Ocdg389koLEKuyq+vW415VJubby+BTnMX1bvXw+6MKI3GvHOufOw8PSTW/ghlGPK
2PGqOlN0wuIzC4VJBrzPwBVndjZp+5cX6NBLoFE8eBFb3ZheCyMmLiwJPFZDi1Lr
5zCfqIYUO/eVqq4FjpUWtaM2wJorOvcGFFrKewfx8wSI0CLH5to6iAlq93qWCTWB
XahWct9zvbSts0zwCFWTkqXWVzkI+yyYSnAxbZ32i8OiCBMq9nOrbk3jDpmWYtFH
cjddpu9nc1rQ4d3/t3wiDD57oAoxUkHw3O59fENcZgM/jUKheGZPbztdfYMw4gOh
J+NHPoowJU9PkrVoiqVBcuAIOA+OgjkbZTI1Vr08HD2DnkCxvjCD2opxMnzC7o4K
Zmz7g25cebwqhC6BdnZomERpcBE7sZ+XNlrMEeipmYVfUtDQ+pHL/z3k/gIRGFI3
Yvswg4N/yTalxFxdQmLI/bSi8ZSSgHeb+ZS59EefgRqDokvl/JCw3oqdlOSRxhkj
bF/gyogS2r87qLXgm5BGN4ZyNSZ3lCM78h5jh7Cgoa+oxApwMn7c1yGf1cTXh+Ka
etkQhf0BSFOfcNBDaDy5EM02YshhBHVGxHUVIYHz7quG3AZeSR9iN2CYgDubKCzn
eUOv0eRT/tDBANMk0kidHSRMCSY1bnqgFxG+0WtAPCncLS5zfzo/NN+U1+5WTPSg
n102hOxZVcHHNL4kBrJhbiP730Iy68g200X5gqy5DNCulqUw48OYAc1a5qRf/+nt
pyKJb/MBz4GeIzRBxH2+JJ8xqxWYZOJPrTUY+PGHIXQ2EAwolTDlWrUMaBUW+fgv
HV6tl9OuavKcAwWOs6KIKojR+U3roZz3AvxL4aQLEAS/3+SfOqJc1hgm0+2WcwOJ
ns8godEtr9vNNfFfjim533dtuA48C2Rq/bPIEUCsxqnV75Ww50fWdz+2B560fFBH
4L69WrWnsEVW3widJzvXwJnRh/A2evt/AT4utxemuoVfVNwWQDOOi/Jjs799jICo
gPE5SmUuLK6ozf1E5Sdy1IO4uzVvdT1p7nbNuoxCSIiAqIqxWvvBGflsOUAiJ8ba
6dnBKGjMwbKhfBs5cbWQh5ZnrcAwa4tkrPZqsn1pxjNHyvj3t8moytf5qUFSI8Pd
NubZ5Kh0EEDj8vph0vTHZOtOlk1fVDwNV8F70oocy5J9EUsJ9dakGEyUfcqOdROM
PK+nRcyKtck1u+S0VpszHI+b+w/m61qFDQqP1VpSV6cvEdF0XLx0ZcwvAYwRwWfY
GwmJiVnETSc2+10IUd22aFqWgQa9Vg7Lm2rW3OYgWWnllhr2+hgnyEZ03E6fftGZ
Yv1wZFVgConQ7fvJi6R+bmiZ6SAKqpduXy19F7TkfcBkQ1cgP/3eoYJzfZmQjPbq
wxzpDgoAscfvJRbScUoh9bUcr/mFMB/GjqxezYbG3mkLUSieF/e3MDOUXQ47mrf1
SLELvvQT9MbUtmZhp3RpELKX6kH4n08bh5UvyS/cbP6ewq86XzXSwGaXLo+vL/Qw
lwo4LVzxwx4R05U3wKI17YeJCMZaLDRPWHq+Rgj/lUzEUBJN/qTWKifJ4vHxw4Np
G3Hv7vRlg3ozbCZnjJbP97s/ecWAzDi4xvZm+SNw6/8HD+vi695dbt/2SJMLsq9e
dKiseb7qHw4U2ajxFE4nEAhR2IcbzfWZ+auP+CF5wgDJz2NKGZo8LOs5R6IvRnml
tkT8il0K3uxlV2LEd+SvdWFnRdqaQN4UOCY6Aj9LASU5cKQk8oaW4jwhgDtMxO/1
JbEyokTLmOQ+GaPlnRGZ0GPDoU040MJLrcfwQ8TiPeD5cNBBujkNOb0IUOotlaO8
6FYYW6nSD5kUx6i4xaKrBnYXM+S6PMoXSd3rHBVkdljNuitdAOZLj42wSBsFaJ7P
yF/+FhUtqADxCS7DEzjsEgtH1CGAcM5nKdPCxTgCb52ogJf4G+4PtLdmzxzhHDHr
KChl2ZxvWjyMxnTnRf2p2LXb2TilKBWWes0bGxE0LwjSTWI1OSPcl5gsRwdkZ+ck
O57Wx4IcRxLyILHlOdK8x7Ola+6ivLYiAITYPA8/QwyF1rslEQwMdbotJ4wReodL
ec+TVCyZ4E2Tf8Eo0k+wEOgaOWFQ7G0MNpctyUo0L1CrePWahekhDY+nBHhfIfCL
iOQx+t2xcvocajgG5p8MZfV1pl9bi/emKulpM9YwZlcsrtXKOh7nM8RccEhrh+10
kN0BhmKMeOXKmN70ZFd9TBYFTJaVM7GaXoh2Zu294PkxEvWIYx4B1xbTxrOvClzH
p4/74P1oE6JKItYrtQ72CsQ95iSV/vLrr30OCg3CE9G+ZiOWSlzTfflv9Ur57dbv
zwY98F2p5LlzHWtWBzmYymVur0ZoYJ3paTLR5EmYnE8hFGMzORJH3TqZifT0vKaX
cjIhj+Ffw/HkS8yJ/jhq9luyEYaaJecnfXGqvLNxg0IyMRYvJCKkJptRDFbHJsC7
+PbhuffoaqlyzPy7bU+Cv/BqRiU3lfRY0OPf02VvBn2SNzdsAjSBF1NTy3rwxOXi
tCk8XmDwf+sLqz86cdGMWBibbZ5ZEGr8oBVA1fIZJI/rf0/Be8/gXLCkytQq+IrE
alA486ItuqWJaz6xOUeDQHs1Y/yloV+VJr9U/v1/NKa1TPw9YVM8lwwYla0qlyLr
P0kM781/mKT+l5Hj1yHPYBe1JYOikIlgMOlIMtf0eRChgNKgyXqp8txFJ03TijhE
/4c5cPHqj2Pg0WKfGRnqnClw2yvPdV3ITuZT25caamiWklK48CzngZx7RbgXVL8L
cmftzeqrjsNu+15G/CNq+IyPbdKMDeAjtwsmLCZXnikOSOziazU4QIRxkG8VoHzR
Ckf4YXi3O1n7xczFjU/2TZzzOnthDvrzlmxPPj+8/KB3miLorKFURHg5pUOpVhq9
XXobSUdasUyuPEqIfhTciKooj0zG0UGzWDB6hylI0X1q1D4b8SAUZRovgq7OfHx9
6Y7DY1HdAgW4VjqlA0x6uS9wgwj/o9Thl9zDGrzJYmBQg2CcZZAAwLz/ou1aig35
kHM3EZs6zgdH2OAVhWrCnM0e9Lwz8ReMEe1APanbC/33JaoXtfTWZzBtHHPlTXgv
EAMFpDB47idC4vB2fvAoXYQoRGWefvyr8m+RRBceKh0=
`protect END_PROTECTED
