`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
96OkiTvFmp+GmvePr+td2VuBPwMXcV8u662mKqXkJ1SQTKm7XukVnl0aOsb1KA7f
1VCrW6HpaJL3WuMHZHgmQm9OaMV/2V9z4nEg5lIMd1hwF2th5q1mrM0csMbHjCH2
EHhN4H0XW6JQA7y6Xnm5xmg4H7pqYT1k8olsfJoYB0m4WM9h/IleqbklhfH0wpg5
I8QfTUYrdIlbUszPHqTUPZ/KfbFx/ChIdWqw5eJvIH7K1EDM0iPe/HlFYmFc54NP
9pi7b4gBZ0eavj7zpdgUWwjrsSg2yccbQT6cmeIhu64awWfk72wr30X7kSn9WMNk
28FsVEEW12eKpIE3i8Zvq/eXw8EeCwrBJ0RVT1I1Xg5V6psKVjMoo54RypkbYVG4
Gk1+lEC0cuN37IqTmdz6fkHkyuEOJicZuXGZ1he50h/QvS1likVxKhw4hVmStc3g
+hN92UzXzrMZTvol20TS1mipxKXwA+ebNmdcOoeuAug=
`protect END_PROTECTED
