`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sqyOAX2kVKC3rcF33YgXeNzrMDIODa2DeUFMSYYB/QQQZ557d3GmN5LyG6XST/Kk
U/R9rizz2n3usqimZfvQGxxGj+gotPXgyuOLP7TSicHBPi5bCR5Clo6F2+5OsbHI
QvziNmqA/P3xToFwxijC9gTD4alQ2MQJt6m29GV5tT887cWWmH6y9jEmKTGeBopM
+p0hJvbcH+yNxPXK2hTa+SWHqo+kGTyQ92kITgIgUyOCgio4kWHzymjTu0Hemgiu
9lBWMvE4gBbbaECsIWf3FU5xT3N3JXu5CLefYXbSz5ON1CZog94OSjIINiNCQ8kH
rMBh7n5QxkkYTjEO7oci8ysHpWi5C4QD8drT9VoZUmEA2HXVJfI0ZrHlteQq0Ob9
kgvm7OXNccgRq8/poQB5qdDNU9Ht8zMP8rWgVVdekTwaBneSRawk5Lj/ALBzFKYw
A2yuM32On0tH8Vym2RU+6J2LhJLyAvj9XksuRSJmEPb7cCw+tnF3pUO4m/zxsION
ERJeYGy8BIK8Bf/h3VNdoswrQXwWrlTTOCRm6984GwOK1jxEF33m2yQ4lQkZ3lYA
lH7avjYtuPVAoeaHrB+noGbRLUNfjHpSDeTnjVnGj1AGfoE34Dlb2hyehi9AFukH
TM9Yrnekt2A974JnVXF5kRAHCD+4Hpa4gMsqGNasj0iGcJQKqHx11qVXaG91+bQ+
KAuU9rCAKcmQA3We/odDWZmhfPr6soql3NEuNSYKvH+sL1/gq6ifhhdIsUsKRxh3
DpilGu3eFpNXXcsLWxuntp0wl0CGC4gp1ud2WBY4I97m2JZjkgP/weE/8FVR8EdQ
aZbRAUDYSyUKBXcFGUf1zRfy8aZGNVcVtAyxmZychS2D6jx6j40qrsGonmIghQAu
mtUddGcqk+hCsTKqS1kR6vIUr1XlQVisrJRUa94Aa3d+kyipUWMS0GrapEgoiCWD
7N5GuWfYHR0FRzIZntqIIsvKis+ghf8nCo3p4VPtz+3sICclfZc+f/CJ+6Gtc41H
oXVEngUTxvQw6xjE7IDVJnYE16ubegSTvoPqiOEumNjeasrmvePWYOO4uLkx6Bov
PS6pn1162/tC3hFJ6UgI7uN0fIzguuht141DhecVCtV4i9rvP6Ya/+lm+I4pEe/d
UAUpM3X5jP3oW699uzKYiq5x8rZyx1uRgKOxa/prczofwZat0ZQWh2v6Sq7kkxtK
A5Fip5XgWlKXgSCfjT8n+DIQbyNaJeQ1EoeYyJm88fqeXXdW/y+5SrjCSqJkVBfZ
fiyROcmkY2PPberckq8pc+Pnv3saxOEzfQAJ+kEoU0p35V4eJ/8KlI2CmfhzqHYX
SyAYDT2hksSa0XL1Dp4RkTQisPbxtC39kzX0ADRUUZNtHl9Lx3JxhdzHfzQtiRYj
`protect END_PROTECTED
