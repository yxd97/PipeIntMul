`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWcibC9OSpeIojfDDZKWKTbcvIXGsD/WQ/U/PBeOj7oQsYEA0CYnI2pXeG4+8/1i
zB/lsgq1wMT5qhpNc6N36uOfupwdjWcFvYzg/Pl7Ef2uGJ1myfYPOfatqn2b9r+k
u0WHUExVVGhXBzMEihRS+y49LwZQp4n5fvet/kKe4cX1IIasvrrz8ySfSeXYwVJx
k+JR7Jz37o93Q9Sy73ImUlNzxbofPqh5pdgOAxBP9juCPI1aRbDvhAHJLqIioRvU
h8Pxh+xN+dhpJETyXEFTzeYOuUmxCajpzQbw4kRR7sZJr1XfNIpgtmqEGkNJERs+
5ctK3zlZ+hsdP7f462ipYzmIA3f3M0OZkAt4HuDY/x3RGq9o62u3xHfflbyZ28PM
rUP2EoHwNcNMmtKx9/cFoT3yghkr2ce6lp/rW0Oz4x/fMLYLk9T8CbljwPZjWQtZ
NAjQ8DM/qF3DXGrS2PR0PA==
`protect END_PROTECTED
