`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euMgGdJARsZbcbL1WbkJziwCimqBh5+TZsG6dzLSAovJen/uGFGjo3F+0CQekccr
4PP7mriOy1VEwQrHrXnMej25hES/YFVUBwfk9JXO3+whlGAkn8S1Y/WxzckxkjBW
bBgBIN11bVxAUYGEI754IDPl/iD1H8feHbpPrly/AJ9Cng+4CWS+dQjpKN/xEcZV
W8GmOym7LyFGNYNFkRX87Mr3L2vdja0UC/Odxn/DoSjNV98zx8uljXHJkePb4PRq
QDi0k5Sb1x3chXYFyOxc6UVoQYb0EwMTXNISlqDGW6EoxD8mWQCl5aTNIAxGrEY6
zaDQN/HEwIQPMqKv3aaN0gHsAj6RZY4B1zpcXyCbeUx1cpPfsoI6iMjz8Dvtvlly
mIyfmDkBuT8BkLBoEWrqImAMUO6cUiFpA1HXOOdOKh5Yw2zyjgSqyrzQeCEfYKL6
pEWVXaYqf6BKxw2UHl0NvPQCeLjX1154zKKo3ME9nZiu+UA8wFtUYLKGHkvkiScH
aehvuDKNflfbQFGaRYslxKzU0mjCz4QI+5rP8j4HNXY43G2MkyfRWv+dsGO4czfm
sqR9lhvAjqMKnaB8WCZzA3oEWzZkuQP2JigBO5K2niPqhS2Q1EVbeO0fjzc/GDvL
Q9XZVvceRqLz/d3DqEMYlFLQii14MW2qV6tUXlEQbdcjbxFP/6FqBwj64cJAdns2
nV92Q4txe1Bi7XwWlRBb5TFNX7St+vYNcQQAdt2oqpxo/9NIwtS1DFeGaR67WhNX
tLAHfGYI8dG06ZZCbpNwBK51pR7YV/TaSWMbDXDrJdadeBtCcKSql3WbFOLOtJBr
UwQvrnfhLPIZanfz8nlRiSNghodyZfmmK7f6RHfCteYl7IJDeNab7C7Hlb8vC7aL
L3WYeuTmkFT1tUd7vtT+wb828SjEj7YOrq+Gz6pmRjtgEA2hYEBaSP02deP2NT+W
`protect END_PROTECTED
