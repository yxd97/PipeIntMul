`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7VA4UBzelwUwoouIUUG4sbiCTEEUuaWQO0gL+X+7e/j6Ql8gi2RcQxHph8PYYdO
6vuoabahucT/QS3SudRmN1GKtLrFhuBa0sSLiqow2JSu9kTnJBIaFq3DgBuxecb7
47rV0u6c8aJmQ9DAfsJ8Sdmml630Ol4AuEj/5OwgagnOs9bVjj+K/SgMY6g0vl/F
WXYqY9JOIPIzZWUjxvRNMe4ge34Ccv1oEBZuXrW0FIPflq3cPOOtVh/NE5Fk/tmf
KAMVHo5aO5caqX3E593fakKqHRRVi/3X0gQJyiS5CYPVuWghJ+P1+SvN5Gtuvaq5
zOe4MnnPjE/hMXya6T11VJDCkLxQqa041PXLfrqgW2GdiqsvN7Z2f9x0vAU8+OCE
YlWCR0/tG1xLsIt8jOMFjHOkFXidQ5CerOUe2Rjdin5jGTQ6NNIU/rh9Qiuf8yJn
D5cDT7esamKu5/aHFIHbBM5dxv14l/atL7+F6m2LSqJILf89Mi3eE/o48kZyfQPV
bjUzUV11id+06bUOrP7T94swdsBQU+JW3PaAtvXlcYODl0oIfmqbnTletcegd3t3
WyUzMWpFxs+NGovpe/yVelqZlSuiLaPgaGZLhXsTIufwtnfnRH9uqjTLa0p68Je6
nKXxCCfDKJHz7Hi7aAdVLjVTD20Q6Ay137LhiGNmBRYcFqwMOINAJpjLqqQ86ohE
bZN5kc+6AuyyAHXGJvXpE90ag5lOSo2SMhxlgR8c535hwmSCYhosAW+CUfhGf/0I
lzuzCV3XaOycGfuwzjkjljQyP9QpzOQqnSMdIt1HKPr8XbI5JZoOUyrQR5suj56B
pCx3bIxoEorJac0uJDBi0W/6GfvUgVuodAy1BKcn0SyNmFF8pMfQEIuvVoOduxv3
V7IXFO93xQvB9+XSpkPjvbma4S0L6W6KAM6fW2m8k2VqGXM808lx67wGeMlejNvC
Pdzio+5zKdsW7z+PPeffPhtEWOsAvZ+ypTG59+dpn96mE/sMWR9qiiCfIrPacxrA
4Ru11ARHoYgeIXfqibvjhFe066wtDV44/+Odcv9I4AW5fDmuY7nScgYcwmWgxmB6
PRL5XDIiW3rsj6wgfGFpNDGOQVbbFBXDhIZ6PxQEVXprQ3F33+DCT4ugtn5n1ZYK
BfDddpGXDn+0yIr5MtsIYxJIsEKbGMMPCdeLl+xutXiCn8JMVMaHm4slcuag2yKD
Wj7iGAsXclJUm8K0K8+mB4D6GVIcmhsjyr9Dh1rWRPPT2rUnQJyHKqxGOtQxHwSZ
PCMpr3S8uExD8fJAExc6z/3RAyyQeXjrTrj0srT5Jk9+xl2Z/QsDWAS1plB2LoLk
ZYGiVP5FSVCxifB7ikG2oS3KvvVwqql1KHrXXMYuLJyKqGF1Mf99oXga9K5+pDL8
vpFNUERcmAhJfxW7q+nrTZGVgwYK/qaarZnDXsPsTp6Wu14NuUzkj8iHAJvHS1ze
8FDnCHKtJMdC+kPXcLvdjnpcM/b7Y5pO10UlhhAUB2ijLTe31+0MN6Rnzm5UD7iy
kl9QmVGgrrggEdHUSNTuqLJu6xQlY7iNl8zMeVq9iqptRCDFj9skIBgqkgDpGVDc
5VP1khyWmrGWCviWm8gyojKZQcPFnaTTCjX6Lh7lOjK/Eih9pp/67iU5Zdmk7zHf
dp9IfpB107RUUKrfWRHWFT4Ff2oQGLTkNmJbhXZgBja8kWVOsbGuQsFhiY+yJ/Gq
BlH711UCfHR9XTkVubxYDlkk0aFsTGotYylGywiEiVsxvGYRs3iH5IjPip309PG9
scGxtRRb1DkwWbAvhs9XZp7d2t4Knj/M8P8fd1br9hh2m7FW4jrLXzP2lBSbeA2X
DxyOcvVgacHv5FSOZle9/vGOIOIMX04J2euofwxVD59Sm4m6Vkmh3wiOLtEDtXzY
1LiOxrsG9yMS9kG/ZO75FWZ/ok2RcfMoslUIuSwiaP+Qvw8AO2+aUcycxeVfKXx0
rB1FQZcLjl4KbWeRMf4IN9jbVF6ZOn+9AF0zCPDKt01KGAMkeh+oLM0kazxf/SoA
+6d/lPr/tD4T8g54w16HEWyoMCXIxu+BUyZNyFvNjkuhXOcarXcghOEDNYIqbE9v
tL22Z2kQaraIn04fqrcQ5toWkFK1gBX55idaTpdS+G1hlj0ZC9dANBuu6ASniE6g
YoFmw6vMLhxAB37YJ06guZ6otR1jbnj1IKwvnPxVCG4cYY79Ofnusv1C+h3CUJ03
Md5W/8lxKi7aka0ed01UMOBu4dW9jM6Foc2uSKfSyhu8mSFHKOJLBCEDSC+pRn6l
zNqqPPdJaJSproisI6IovU73HuQjIT9AB0mXPVdH6Zn4a/64d/8aR8xC0S3DhYZE
JqBAigcZGv1QyUMbkLoRNqLJhgHKWwocSEVMudMuwHlTh8BiWGbbuSpKmhxZZJi9
3JUIBrl10m92YBzUN/Fr9PrSnPNRd2VPnOwOG4UrOorUt2HoYxTHm1108ouFMnLV
aID+yd0LQnQLI/t0/8OOWxl2CG7J8y5UA6tgJ7AL4C/iuQWCLex6Psoz7+wsqvkx
ggFhNEmGs+Xu+TbxD074IkxgB5htrLu7fpwK5hRvmX+n5E2KSJuhc+KCJL8KhR+n
XtDTfkOf5fSKxpdjmwHKwYrmelhi3BeRZ4H8hZP80FbqgWWaJXPZULK/vWCTGaxw
HuqjX3uvitwJEQyvfDg1/zNX5ds/sQdDjP33giUpcNpY2LoBM5d1eCujn7TLvp88
MEkuUQReOWPaBvLfmsSPBjRatjDJam9DFaGLlUWBuLzaNZq/TrSJeZRI7oM1WQiO
sN4bAfd0bzA9R8Z3dlgHsCWRAUmIEq6+l8Ea3rCPtFrISFGKfad6/3ZRMmVxQuws
klA5pUrEx2j7DfTG3kCij7ucHf718pxMcg9StJhPmYcV9VUaBqwXs8hM3/G+mnLz
pD+ssq4xlDqbe2vfak0dqYEBOM+gcbD+4LKzSTGfVhmX+osywrFi7VmvgnFUQ59D
xxTaqL4epV3YexKrQp9Cmi4G9WwdnHZUMRLVxys+b0nr25i0enRIPITy+gAEHjel
fjMg7J1MOMJ2dwMREAB0dMkiaR0QwmwS4Xnf0tqK9x3LM9haF9yQG51rUqNfz6SA
4mhM61LviIAe2zsAAaZp227a+h/yJbGto2PU4ufWkWiEbVvV8FcwpwqFwYiT8RsE
JrYmS3YcPtKlqMxofx/XiFrNjEWYpGbY0HREqdTJJBz6zzsu6QfzvwvkkWxsm1oF
uiRBUiMUq1nUHRhcsM0SJFG7LYPuUp+6HXC95NnSMBhb9n+g3ZSQMr29BVJlyA+3
pyQ5D6N4tuSEnwkFZfh7hIPWntk0sAaaPhA7K01Ten3oF0XrpYMCBRfxM/bws+mi
v/uy0rUjhqdkeokMSwgOURn1ke91gG5Siw+pJOteF8lmyu3+9rUo7JESUmVOY1lL
7QnKvgfXym+pD2hI5ECO0c6yQJLR/ArJCYnr+UsBJHDg+TycccR0nvqIHBjggCa4
vHx6yqYncEj2H9Hk8DAr34lbKhPAQNsgKXc6gj0PfBbNjW/UrMwsFCgCuOf/eEC6
7tpeyQ+zOA7r/Zts4JMvievRPzFMZb9FDTgaijZfO3MtKnYehpJ34UA+bOAVxGPx
OZFf1QoS+Xc1LxPGWJ5GFXaZCjTxOyAD5Y1DldumkXiGGyPqpCdS44WgdqNPRc8I
EYwQOcCEopgp09xcCpc39+mh0uOTnEynHRlrsyArKCrkzVcL62BscmmRDqkrnOWZ
igaVGBteY+JVAZew4NvvML6pUqPSaGPymZDMl4BgNl3y8FLu6bXcONrUmNn89vI+
4ZibUvXRGzCQ+c8h9+SSYMC7kdmAHTY0N9j86Gfx0BC9OfLkKIJiUEq0TASBtiY9
3zIY3/a/hg7+p6YZzPVX/gCjGVZRypejmQHCh/lkWhiKQOv+m3/tgvjXjdg7rufI
NCfb7genLvVZJ0/RrGdV0tRjLNZPfXNK/0DFmvuA78FonsQ4RyEZwcwzETdnnje3
OCEzBj6X/Z3tUTSY53mophQporOkmwk9lURTruAAsgamQ0ElhQIQZ/hE7oRXvzjD
6zbqWSOFbvHWyFjb9dethfVT9f8/6t+LAde8/4z52ultvS9R8kAt7O1jH/AI35CS
n3bG7f5zlaqgncYcGcSMANNytdO4xbe1m22ZbwM5DgrJIVhXLfjlQFbPpgng+itR
hhuUQCbeTfEtn2aglun408Q5yei56toddXpspdnouRhqFl4mCgaeIrzkyaWN/Wb7
dkntMHourrAeE+HHNIxcjTGYj6jEc9tTz48EATCEaVVA4GnFzC5bacgkg0qVJ609
oDZ5wGkLwqNxloOyXlafWeIsmUyNX9Erwj1N1xxiG0WZSzmOlOMIozaOJKfb62JZ
Fuo/8eVZZbEOUH2ito6rJlxMZDwIMlHEFry60nByg1Z+VMxDpnz0vz7LadDyB/mA
xt02hSEdDG/fb96i84/TZ0QTMpO70mkXQvlxQNh0AYM77b/kKgx2FNAWsNhAi3ks
5I2S1CPvyrQKFLGY5uaKvtXwrhxm6bilFfAxmArTmLKmarjhyymkX5FCs9A0ElG7
ggcZxLzS60DsjDstrI9HOhLu2k6sXOU/A+NR7hpQW7sgD1VMfVFHIdYLPWgicuOq
oqoVs9gF4O1jyQq4jv1FI3lNngU3vSqdrNNZsllFN2s+b0oSfjmE63qvJYHrkCoU
wy8f3/hi+AMys31Qt0D7mFZiFiVkS8KkDunTjBPr3zQq/I4P/FkGPj3Lg41u29Ep
NnjlD60Z6VXlzCBM2JbNMcTKAASKnysCqYrkMiqsVir1deP/XOFtPpeUBFZbouO7
0zXsUDk/bEIjtUUbBDPdkZr2dBBDB20xRbiUPN842Fxj3MS6BMcTzfjXD5LfRUOh
X5+K7U8ovKx8iM3QQUdUIY3+fToIwsMuBO0YU0qdSLzBeIFktKYVvxaKXXRbZQH1
Jj0F8V/8cINLApg0Nnctc0XCKX3RoQ48GuHevUx7Qu3DUKB7LNHabhVgWXTGYAUH
Txnn4u1vFBxkpQCRnxiaML32oGBvg66A11rQxj+h2r8rVitLDFgCBHsWF3t5EW+i
G01UfGVTIuPSTrtotGzmUx413WrkBFE6RYYjpSqMty7Bkr5s1obLozQ0ZVPaTmJs
IM2mPJfwaIVrije1VI7nFvKBuhyckC6DBtCFYI+xieEPctvtuSViKL/uF+ISzpVJ
Jvo0+n/mn934dTBe4GnxBU+MPyk1NU1Z68yLC1X157S0dsUDBSNJwB5KOAmKeqgL
BgoNuVU/lvfN391uD54UX0BpRbatzTz9bz8MXTf/O+0RFcNxOPK6PhbVWOmtn6uH
jQcAWRRL1AvYv1hdI4t+jBGEATAGAWcKXksxPyg9X500Rfr7biP+9SzIXxL9LsMq
SwSh2FQ6x550pWTOz3RCLDWQgU6MF00beqbDsJMUanfovKIhD6uzKukdIQk3xV0r
dNhYBpyulMqG1jxMHhl1B6cve+TCTRkQpk5IJPZVTiQ=
`protect END_PROTECTED
