`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
flB9Vte1uJCWB0zcSOPCYps3PBVVy4oNaBexKYSB1mRglOjPFJXjUC95eVf+gcAR
iTLVpkza+Ax5DAEUwdwSAaQqyPRz455cMjk8QbDsxdKx4sVLbaPRl+ahdrMn/HNt
sE+dddNafpuauEwthxsprMhihSBivSTSifUUona++zljPjTAKh2D7Ic7fjWoJUQ0
rJYkanerU7VjecLmTXp4H2TbbBeV819rlU8Z2GwOVJ/SZFPMmn7Ur2UIJecXy0dP
BJRfj+JG3BhIboiiCjFWfZA7FdiUy2ZrSnNyZTN9I+vROB7L+cWU0MlELKTlRQYS
`protect END_PROTECTED
