`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGME+/QUVQ/4qXJp0Kp3qGIAfqr4IYqBv7Gr1ec66MaiwMldvVq/W/240Db9ku0a
hcL8cxGwBzarEGrjAezqcnSiVpd6ymr4r56XaLXZ7UQWFneNvCIPtMJxcTewTk7i
eiyBxPChGEkNN2NtuLa7ueIOgFXeq/6YRDXj6++rzwAI832v+Rm47zlNWNLzJs9Q
hvUR/KjJxGxOZAKXb7NshoTtIyF6NbfehVnqBxZNb41GuWaTmhfdUgvvYYCU2Kxk
`protect END_PROTECTED
