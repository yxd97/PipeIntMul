`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5XS+YFWCntuzl5xbrljb5J1RMEh4OFc+Uk1BDJDI+a04v/r/LllBDf6EGNWWAKki
YjypP8lguST9YxQQeyJfx7+zsiwdPRdWnVwbXQGus7yU3F5wmdQFWn+kg1ZzXDMU
c8z/lzm/CvOlnDCGf38FzQX3yxN982HbsvEuHIVcFjlotLqTqDooOqOUZHhIWJU6
g9bCUwr5F3TzJL4yO15AP3O7gwuvWgg9gAQN3uG77s9gbnVHO6wwaCCAJNCXeTs2
HZsMPYeFY/TF7BK8Cw7NxvMDs5pnxKCZ6k+RjA1i3QHqTSrSYAeqeheoLRnjJuto
ufdnMmfANf2yl0//u4dfVGfOBDW5ip9n+QnkgfwG0vx0rcu4KocdymfNBWq3z7J3
BVtIpVbPj+UsAKoK3jJARu5L8OLGfN4Gl+Rqv7SuxVbNboaMIj6CQi3EKf04YFep
CbBcp5WTl38Xi4H8QOsDhN39/ggV5sjfYwGrVsnxhxjvjjZhC1f3GmH4DknW+rP+
D08F7B6xa6K6Coa6Vj0PGjvdpbsznihFIsvlM4M6km2XoJKQzTJzxXHZYVisOCdd
L3oEkHJM2Lm6+E/ZgbDffuIurRG5IzHTYl4FmjPcUtcqMI4Mp/SwqwkDwvhufvts
+Xa19tWtVEhB2RkiXoZCgQ==
`protect END_PROTECTED
