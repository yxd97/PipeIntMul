`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4OACrKLkc70ZZy2kKnhn0vUmmW3DDobT/aO7Fq4OJmmnhZsLLM4DsqbL4jnpBi99
TlJizgEcdhOXAL1Pgzzt3eYA5/UEPs++aItTAA7m+s3TkN8Adt6oONEH0T3sOUbn
CFRzCo3AZdLh1VWDmtGRvAPK0aBb3nIzljol2SVY/lBH4undf6c57xFplYBZ7Kg8
yMTXkcdF6cy2GT1Mz74DMLpi/JeV1DNpLtFYonxyw0jJMJqijadxAz2OPj8KLNgp
8yTA5VFh85Aga82oZB4qAqJ4q1tNmvh36Pcseee8bNwGgSJY46YaySOkr4bd01WZ
lYP5vw4I62SVcnDhfHCfixE23qDIJdghH5xMp4gPRpfaCWPd/hdw43++VC6ivOwg
O0PdNli/3yZqYTEEcmPT/Mnf+7emziXpc1SJTqwGKHfkgcUusq9ubuID3nL8IsdL
XW+ppidYass6T08grs26DKbgX4Ym70ANOQaVngKqU6jrAzIv6abaxpMlbz6rkO6K
dfGH5DXLfJ7APB484Hz6JSTysUfUiNikK0g3bjicWe2Fek0eaW5wOe4RwG7nCXiT
IWOvNxa4vCC0sfChqFziaiPKNy+/ZgYsMV4KL07ypraPLZuwwMjm1MZBK42tW+Or
Qz2wg+BnSuO8FcGuxVfOyujKybq4pBupNDzlrORM17tA4Rc0E/z8QisqrLlMLr1S
GOiBhadJw7Fax6pmsLAm8ejMFDhBbgay19DC0uyyaCpALKm9Z0qtSTB9WVnXib6J
3ZJ/hL0XM4kZyGyteWDfveFtUurGNYo8H9Ixvm4x1IbDcxripWthq60Wozt1Kc7i
hUSes2r4fApVJCO2GUKqRqf0kSaxee8xTC3KURtVLgy2GUszgKeF8TXLzgeytZKD
oPxHdcShhHpXJLtHkryGLCRoDuoNUYVWrbutb3bxP5VE4adjYx5KgQTtWT6O4gYq
yDZV+8i80LGqnqiPn2KP2isKDsOFKJD2Jqc3Luum94eXBW6IImRo5GhrV8B0nIaF
jFrAVyjeyzwU3PP+CiMYFPBEY1dOYSI446AjOxPBCGoTA93K8LAJpUq9zZD/djq8
MsbF9UfEJZXD3gpBtPycxbuwBGUKXV7wy6w+w1KXwyabf5TQAckc5lZpCRPeFm7N
WnQ93ReH+plu+EQcdQcaVohiBsuyAxyj/z1G6NXDXKaAFpxioHV2ZGzdS5nNagdk
BSM+ilDxEysigmnvPf+Ljs8psqBpxf12aCM3/GDLxjV2tBiYHSrZO44g47oqGrMB
tg2sjcxC693kYoZ9UcT3PGVLgmTJIrJa0DVmo/Ze77ifWDbhfJ7MNXFh0r5FwEoO
ivbo7jodb57aKYPzcvLu5voiwVxu0PwWOOZ5rm3WzaLin9OlY+AG6UV8w7YJzPn6
TErbigzvvSPIP7DfjpYO92O6XJtiblRj/WcF3JroxgGVMj2CHCdDl/cT/Qd4x4Xj
YvJdQtqirgw4N8B927OBjPtQDf1cw0vbbxfBMHgwslDFm/7CzV9F8rp8uWfkoNby
yCHRobmWWHQjQiTxtaqSY22Hp0689D+kCHZ8rAYs6S2Jed1f0tK14pb3jH7C57Vd
OGZqYUnfawS9ZrawwyYf0YyLyky6Du/JxbJBHixUASUw9uAcaIfKAUbfx7AFNubl
knDdso4+iUONCqjd2AUSPeUSnXJI8vPxqcusmzXIVuKO8tbuNM0vUBD8PNuJRVAY
I7PG1jK2Rz6UXmnJyJun88anIoAKYFrHS7JBNgemBR68VUqxv5pgBO3Vkl/bsDO9
FTY1wOVsoijivO2N7kt8rYH/nkJR7Qk7Q7MnjN1DQIfoH1KfSzMFUh4X3R3BVCqq
Y9Zi7z9ceWmYsOdr5qIBrFecnIuDrr1HSAQN+ZPppSwjmQBlUE3sroM0jTZVrdUt
HzR8zAOmcXmSZD9sAAllx3beZjDA9g/ePyihwa2VjBcJh8sr6AFoUk6NayWFN1Hw
Na8C9/g+XSOLKr00cWx6q6G0gtp1iqpAbGNzlapylOF8r5BJ1Z1R/BQZzAgBi3qz
/0tGFAu4ZUTEOJZP7TolNegsKcttr7Krco8hKcUBWJ158S7qxqHnItKbCiB9TvLK
JUfWwM603O2ks+D/lz6T70Xdz7PntENFkY70ZtHh12evDH1+vyd2/zsIOk5D5Jsc
8Xn5GRj+2pXLlGBD1sm1FlL+9ZPqSQ89Kf/fPRfzEnPJlcCvvXYOkjLIWFNjfheK
M+jpWuiza0C4yyswR2NP35JpBFaWQlI2AavtS/B5Dqe0MGmUaG7ezHrP8fL8lFmT
pQMUu+SA4DkcIb2LQslgJfa42UvLxOtJEglWrZzGSGfdI/8LR7ad370SYZsUXolt
T9/dhD/G8Vvji0lsQvB2howyrTDIjRCkDtyZNColxEexTSsMi30b9sCf58UMWsoN
fh2WKGQgIPR5qgOgNHp6igD7+5ftwoPo8AYRhKmbMwR3baADdrFj3nbQSsGmgMF2
aNtWxQgyp/huOFJEZLeShWp5deS8QgoGaj+k9xtjQgtufY+ve9X3kUwDe4OQzU/7
p9TahkP4YVG6J7B+wmfj+liYykdn6oiqI0djog3o3r/SA9QrkzouJCygpZ3gdobZ
LoMfwCJtAH3+8VxBj0Sd37xazGL/qyLRxodADLXlNPzUSKStMIriccX6W5R+TPxw
FBPzOC5cAKR5aPxKSYh6gZmHcBQaKcIiGo9JZyuSqCOc5wuyXZqLFOlrdlfY54fh
St9+GGuCkSr2c9hHJif7QeKUs4Hk/jr06ZXolp0Lmso4OcLatZ74oR881fzRAGDY
z2MEOq0875BlclUHWjENl8+odm5cBlQIJQOv4k632NqZxopVtWN7a2pQZ0eAObGO
TgnuJhgN0SIeuV1/khtnGHb9w7O3NAC0Sn43u9TUHeOefSVCEd9GrsH6pRV3WgYF
GgPEr9mKjSaqKwoDHO0gKvlGHDVaGOAzBX7tS4Dh1ia6578+83J8VZl7twG+U4mQ
tFPvXDIHO9VFcnMYIJs2fcFPLbpCsq21o/e2xJVi/AGtczoX+jzxosjLlmoN0ckl
huE2FhQZ8SY7uZftLeNHJpZAkLhptCo4Q53MAztCkrEcgGy/CTsuMZlwfnQnYmG3
DLxcrI568BpWmbBIhNL3W92fQIZB/rnBKcRCvoTERC2CDRtMyLLKSGYVisJlatg6
lyCUVevoxSGtnmvgczNiMPxIAxEX7KLzGxN09i+Ojs2sEgkziTHJBVaHnS0FlWz4
2l8hNs4H15ABuTuYvmARE8pNKyi11dCqKxMRkNKwPtKW2kVeuO1BFd1AfimqCyby
srvByy8KGTZY689eZu7lDAWesUE9qC51lrX6kA0zDb0wRBRER3aSp6zdx2KzDM5U
7cNiGSLRVOJwPIMtdcKkZJ+pepoCD9704jBjIEVxCx8TZteJIHWURqz5UIpGX3Kg
TaiagGWfWKpI1E3LtJH/6Tecsp0P2Rd6YwykJFcQX3eztpWaeu2EW8+GQnJ8moti
iyDpXFhjEtvsfOaAV8qY2LASdZ6KNhq/EdEKGvyUCfh1QBEaey8+csSAw1R+CxcW
33fyPTk+u69ZeHNGgpYl7c0TFjZ/07eO48vRjA7zbouT6/o/DAk8QGIN7Jrweu3C
B7QxuG1+kh1jaVqlUel/cZAXBvKzknWtkpG94l7nfAhYbSP3yJb0pq1GIKiexsId
RpWR9ijB9uwO1Dw0/qSE/N1toPGy7a4/3XELrD6AppErwYgfe07ks8FN+iy289RY
QcIx8cBQvVkj2ytssHpcrXEWV7G8NpSxrfhkL+aWmuiXf9iLwkoewg3urrBaTfRC
h1Fu39nylg75CiPu1KL4YO9XnwojbFeel2lqVeq7LKac/CWGHLJno8lvkApceAvl
tF+t5GFsDfUYQORIwPFNhvN/mtB9WE7B1b49Tp7kewsi4/KCruuJ8Y5y82EO8Oc2
GtVwUo6qz5S9P7CWTYMkbn9SFodylxquA51j9HtvPFk2lNJHtseg8/HNKBc9tomr
28CfK5RdNq4mW3PgwRnT9xXTFRtq0zZ03FEJPot0YYJup1LokYf3glyLK1rXDkoN
NiMybzhomvRhHh74YlX9OpzTmiYA8l4FbeQV71J1qta358hyqa8szm5gzBPIqfZN
O4juyxLYXP0jPEp+WHNzHk/9/WNrGtpgvjn/Ff5Isclkz6jbdJMkliYwIzEQsq1O
cbNj9eEoRzP+bdD4fxV6kZdV+0bI5AlJ1eJxTqskNZC2ofMUjlogJYZ+/ipFEJdc
FJwj3kq1ZgczLV4BQsa3Jf6WjvRWO8j0dLbZp7bZUbSKNYNn1uHOrlktbkCE8QPw
RPSyCmDHnbW1ac0DC2bf4t6YqmkQybr6H8liM6X/zHJHJQuPQ9BCV3tqcjez1aKU
Vb2hF3KYiw+6/tw8ABqyjLQNXyoacKoLFbgyAoIgzem6+3/gkpFsJsmyt5klLLZC
s0VAq8yE/hVAddCqAvqNep9yw616av3JTZUyddNoZWdw6NvhvrMRCSSBn2cb+F2C
2A0IymMbKOI3RD9/WchBUTM+LHFznc5uFpzWFkJQ0CR8MeoQS8MJZs/dqRUjmXiP
jAISo7DziiyscJ+/3+/LVYTTW5LcL2oROkvB8HEby64DWBmThyx7IFMvagQZvDzQ
iL36UGRZlKxMvuL7noNyhl8QdjPjLLlpfrTWvey1rk2ACQUVt18c/0lX/nSgPTN3
hswArE8o1iCZb3a0Rk4SyzcePsSw+XMP8iU4Wn7kd780G8Ils2qWYeFcMxP62ql2
hszaOJjFXhpb54KbTD0Vrpavn85RNoVs5gGkONIvpGScmknwwYDT8z1IODlxb69O
GjioQG7h6Eu7l5aZRApAE/VyjKmX/YjBI3ddY94LuA0pEFKVdyaksem03q/4aZS4
gJDiBTOmy02mGUTttUpC+jFTsi2c738GdsVAzcVeQwVfMtq8ELjlgan3PPfrBGZS
OnKMaiaRV7ULAcT92SVmwHvhCnVo1ZRYvVeVVmT5/wQ06AFsNMUOTWqTeTJy6m8B
eHN9Yiu4U2vZUHy5QgAImn71hL/Q8xftQ2jkLyNiZVbIulkZC+Th74ktavkiW0M4
Al/sWxj3o0lhbWcq9D+2c+qdifjOKl0tVFSHxOv984Ozl33QQMo3uhYCVcFXvVTp
O6HDYbePuwiU9TYdpG8grXTBujnFWgxn2u+zKAGRE+XUyhlXNe10CcqJZAsWrfyN
UTwA+rqEzXcC4ZJdhoP2BaCBpCTfXwASJJ639qrYSf7xIKr5bcN5wXz4ce+e1X1q
1gCaB4p8WcdJT7d1RFWvFgoZu9MZj57UDYL/QWzxU8T7mHG58qY3IDX8r96ebwj2
dDZBV+zgXEqcdlzvCFmg2VJORoZGVIkZ+JT3SsiCJu2jlTVeo5Hw0KEyPgrgcOKF
Ghvt7/Dx1jF7OIloYLr+o44xzOKwQ4rsq7mKOlH6xENgymYpnvbYqOE23LS31icl
R590GvFJCsQNGxuFAf2AcLr0TeElosA2Y/zmMfBFvMpyyymOgJD+0HMJe/2id7iA
nVKLeKtw56OWNr7jG1mAooZTdMw48acKqdnL1ichO+U4lt6EtO0wShltnPPjxjtr
jpekj3jbZze+5W2XcEfmvy8+of3jwjv0FEx3pc5TxDjO0aFqjnpq4dYlaQbwidG7
+bERaQV/CSQaD3rrh+53+oi3tvxfVT2vgCsUnwHWwgf4PczVvC7XiCJnVNSDFFY9
QiuelmIDveeU7Q6eyCLR/YFjhU7tGY4E/GoH2A8xlk0JTFmoEORjHPxSap/jliKv
+exKE3VKMVSa+7+l62TcxwnHTwombW+JIYSyjbURV2qFEHQT9Kr+csC2BUTFgrE4
EZg3Agr35U9ZOEL2A8/jP56xB4yIdJL4LNQOQU9ECD9iThQMbuh1uifpT5sAkYuh
h0eayZT8uJDfMG3ZoHBQw1n/fsU2SVbcP57DodmSxr6GefJzSjX+jp8pzzSy2K2j
doOl4tbELJvzyjnzsDk6nDYmIDQR7A+6enWumByDkhS5rb/1N2vgf2RU7JmeOTwK
Hw0n6LXR7U+iC5ZLS4QWJ7IONc97TtWYM1swfNtoogtWxKTcXx5pdGGFn8fV2FWM
KyWxsyEiITLBWlCRIS7oU/8mv/eEsGv3zBfXl2pEbLpvkVCswzCyPEknl9c2NWMV
aoorxyvhg6ywVQvJPdhOfIiDM6rYXsXY/ZVzgHY26f9A8uHTNIoap2qpVeaL+MkH
66NowAS+8JGVcGajTnrQLVL6MAcGHypVz+lg9ZihsZDBSFdHfumQzTiOFMAtaX2H
oUVNi84B3gmn+BnhqJ84kot6b//F14kHyRkMAF70ACPglt+UNKlhv6TFs8yaZFQC
MhHaEoTqQb23mprXz6wHAWryv94KgaQiSnpYpXCn8alxZf6crTWaLdrcbnwxh1OB
zePvFbaWqqT57uDvMzIaAvmWmG5uAdi40LVCj1Cx/nr0AcoFCarYhkbawjUqZMqV
XzY5uLKgEOKZskB2qSqGgzBBH48xVy1bApgYkuIOggRWwKBw5ETR5hkmgADZrZeI
eOrS3xEWVhTRD+TPTT50Mlgc+bKkUME27pDT0aOmuooGwqv3qYFNqJu4W+Sl6vE/
6ITLoDCr7ES+rsGCEFjx9f9FHpBhIMvgvecwPMO1db2rLSol5LNo7zrEuO+QBoA5
81GHvaEybGwoszBbLQ6Dcd4BvQsqKLTA5+8xyx4WuzjwIvZNHqRjwwMZLpkuP8w7
cL0rYKpaCiTIK2zMIAmoEn4DC6PTlzM4NRpXsRyjW9wrH9N5h7P69Vjyg6gZFFh7
bjG4r3qIwDmYEt9PhzoLGHdxlMjMaylxq6JGuAvNCyxgUnV1KNCTrTq/EVvs7+hi
s9ZQbOiAAxz/uCe/F73YHpG2g9x6OgXuaNPXvDpL13/sf0LVxanhxTNaAWIj0mhe
p+2QFHbXl8lpj6OONvVFpO/lsuFX37MQ92y2pLIGSW0YgUj3pejTGr0LGOpJrXTH
ve00s3JayZ318ywyukGKp2mVpjg/Lcy3JmhKjZY7ZziGIoAvSl0UHzoN73JbFhqm
VXDdx1O5Q2e3+jMBqZlEApx+CEw8/K8KAztxeV1oGeYO0UVrT4Aw1ocs3gVE5ZYz
uDcJfzG4NAQunBnfOdmAvaZ+4zHi4cNoREufLBufzGBG6AnPc88Uf9CWQ6BnWrlF
dknJ8/Vbhrlqqbrty7maqoXKl6aGDlSw6ZFDbQ3/hQjSXTM2bCEzLdrUyWexZX76
Zx+KQhJVPJyGAgcM5yaGtkEQwo1r/aguG0b7e22MHabv1GjnIvMqzHmmcdU86PZa
akCa5Dw53KZLS0fCva1IRWkSzNrZ/LN5aHk7CDcN48+Ul/FtZ94mEkGYFeUWGkRy
c5ieHXt+uTK/nNgtOOQ8eTiKGtXunhcXDNvtQ4EYu8vR5Ddlsg5eEaMMJa6LINio
R7G05nEAB3C/oG0D3Oeq7577G58UbVnQf2Ey6g8eTYvo2YKnKSAw4pCV2Ahdkbdy
vGuK6zMU+Nr1h6feexs7h5ubo8kRxK98alfOtVnPm9gBAIZuj6ZFcCHaNH09Q3op
3KGVC4O5jFC9s1gYalBe5B0DdczHBjhdGEwBqd9v79HqI3VN/7L14y051t8i7htR
0pd0RRkFsbDoTV7uS8kmVOousbxJghhds2+DXufYJn9lCF9///vGYpe04aadFNVJ
+j903tpTzv+z3jh/iJN0ckOkeG6bDZ4GcT1fK8eBn2N7EI/T1xobdSDyNjYR88bT
NMj02ycXO6PZ7dnOi3k8CeXF1mdnFWfeHfSkH77jRtXAVIimZK+z+q2uCK8mnPgM
S52whePu7/uP9IkzXdVObxY1gRAPMMkgNVkV+LfTzM2EXRbgT1eU6DVzObnVQ7gH
P/yqaBVTb9Pj4sT0mBdVWKN4hHrOiFwaxWJOtvZDVVqCOf76ZXiJXp9/zZY53KBw
wD/51O79kmMw1rXntssKkl1J8cxPDH6wGI3LF0Gsxw2RpbmKYFBncsLrB5ykC3rV
aPYhEypHQzSbPaSGiILp5j12SjO1kI4Md4KbeWfyHlbgYEhcDDfWJdLaGs8H7GsT
lSmfgjcGKf+bDMRgYwCBw3yK651ScrSh2c73LuDw7aw66+kaLo4u3t3itgGy/IzS
TL0MM14P3+2BflAkoiB44VkFvB6MDpCoA4kLeJHVWEZWdFcXKOAShuWj9vflwnZQ
y506z/3wJLUml2JfaoXCkKGpLg4DZe+YdSqFVwIr/nekGR7q1Iy1cih0Pt//ycAs
lWhmp14GvRACVIT+Xw7K+mFUvc44u/qdH/MX3+tjgfjVRRpALHXvNotiuNECLUBV
e6KPv2ImozqTJv2IT8tkZcuTC7EAzTtZrSK7ROfjrsh5XwrbKzMOfnLYHOxTwtrV
ZhM7WmnvHy2TXXmLGBx/E6tSIc8g2CKJRAvI7W8un4Zw3flNViFbH4Q6ohikud30
gq+UluxbtPqcQiB3qrcK0azS+4JoKWcdcUfWUo3Oy3w9EWJ62h+/X2RsnL/ZsbQg
9Le5OshUVyQTKLBIQ2mXwQW3ZagFcaYRmPYt0Mv0+5KGI0J/KmTzHMIn6A8TNiaQ
ev2RilvwBdSaVmZ8TLUCS+8a7NYQMP1xwWVExATgUE0pDTGoX/7bTlRjfULibR37
5b03XKTYN6Rktwx4uECGLm/jNRGGonP+3w/03VXNLltq/olFP4Uw8R4boXJtyDqv
Ewl58WB7A/VyusiRmy6AmGGIaxP4SZHQtVdXE+9YRcRjFHIor2n4yrRj1ubZL0je
6Oene7dd2vJV+YrK2gX4H07okyROkSyVMvrEFoP6xFgo7utaxdZlbn8/eugNxPfc
o+4rAt7Rj4EAkEOFPu5xapmYG6UFHBf3QGILcoHAq4/sg7VBBb/Sx7gx3LHevyBy
RLMyxc9gmWtM/hD5AcET3qFyLIVViK1e7NhKG8mYLs9jdV5a2SrOpvAThR1TYiUG
1YP6rd4URI4UpZqpmXIaqxbVUaxY/yGNsGNfw9dOmyOcN8zX87zzigqOafhFjDaC
ofeowqT754QgR3qE7/KZXacXj7ssFDIZ96LEQ9qwU8mCG3s4zQFNVda1n/ntDZtO
Ltc6p753HGLMDiScoX4IspwIruFE9Invf6yJLLFAYZegr7bSy6Lxi9UTK3+0caRS
Ti8vN4S9BfQa8DrHCu2Q7ruBvllB+LfxNQEtPC+yYUK3xnjgDLYMIBKBZAQAX125
9SxTlXkxAhOF138vaRr9g5vawZ4LwP0TO7LMbM89KOBxAjkrSgtAX2UyLWDlImU7
WEfvq5hfIVsU5seB1KN0k9m50AVl3UwyEBInvBS98JxSsbGSXXZFTswCFOT9h49w
gUFmdoPf6R1beTx2oR6F2fqH+GZELPhy7LZtC96LABdsJo3djZ8YhQal+mxJaTWR
GdDEYHSZ0//SwpmEfXZiGLIXqNu9CK8NoyokTvipzEvA4MYYVHLVJcd5EncBY83o
OaUal75ysVz0V+EE3/Yx5mmWYWqwyBCi4qJknS19xJTmLiDR6bAEEs7sacnRG/pg
Er1SpzsyOyCFI7PshdD/atDdnxo7WkhGRaPs8yt7sin86FFMKnx3GISK9RRumkzP
Zmwhw5uKwi65i/KW2+q2XCB+M815iyshaRqqBz1LGXuFdD0z8XLzCY5txrFiW0yF
R4tU0dhK0OjTya3i3Y0zDKgSZKCx0UOgAIA5Ipn+GUGxfp5p9cXUBU0HaQtZNJTD
Ab0L++bBI0rowyL2AA7egj2ajrrYiN2QDYX+pq6HrdbyVQgK8QbqDZd8WQUC6K6w
hG5vtUxBWAAoGtH7+1amINjrYKj7mggB0yWM4+bayv5m0Zxcv+vQYYRHdReqr1ad
gS39+qUFDDyMNZBMTtFufsEDa+MgbxMuwpKGX4az5+/OJUDBfTLBYnkkSaCniora
vPouMsdcTGchcS/DQq3Ogp6x72/JB7s7LI6Snlh/Hg1+X43V2ozhVxbC5BPuvVoo
ua36BLLnS0n3r0cQ29zK7dQw63Mzlo0d1un3/CFUcOWbTiHVJfy4XInculSl8zBS
9oDADKxRYTYxPoBaACWkP27s1QHcQ0XeFWajj+iK/kcM7qowfVeXOFIxsA9Ue+Il
vIVQTDJsByWgiU5+DzzRTNwVkmX8zKsmzI9JVL8qvYkK2pg1rRFMA/FhI8+VPbEu
aIUwBw574ZSg49ocyPB+QAY7qfoYRdTQrcP+DhXXnrgtVjKW0wXtngaDROKfE0dj
/GDOjroyajqiGmjSyddqdgIRlKU6uvNDHzvsu/3QY7QcYv0IJx6SimKg9I3fKmCt
OtOZqSlf2iMoQR79F/mMZx0w9PmkVR9ZHHaoi3dalKoS5JQs98VDLgzX7eKo8UoG
mIjpMjErjuaD2NWINZMd/+N7mvcy3eUDyGkdYUvOKD3u7rUpZjF9w4+Fd9x9eol2
Gp8CjOpcbGKCBmYRhhOX0h8YsdhCrQanbjFERf7oXxEYJ4RdxbygvZhyzH3ciqYP
vfkPKdLr4T79mrUkKcu5NoRGsuiYShj6+eBIJIRBvXKfwAxJqXqZ9PK/r2DvAarX
+2GHB+Pa57VIV1fMIlEa8F7gQSocu/j/ltph+Sk1eJ4QH/crrCZ8yAWYS0mMskxX
TVHJjZwuOkWJS3esve4hUSJbwK3Jl7r9CPoC2Jmdx1cxVPbyQjIBGCIIVGJ9LTQB
xF9q2pcKbsAiuKfIGOfYGyiwOzrUwgv9jWsKjIsk6eE6dZxSmP5quTUEluQ2BgQI
sH3kY1vE3ALCb6XGDkJra2jXsEUHevFMSVlo6bnHuVEEjR9fRaLkYarVLF/hgKZr
V64gBmrjrYFcRHnKZYHd4hZ7yVFy4xgM0hvvxiSiPQyXwPqjlVYtUQKx1Ai2ZXUo
lxACxKNBLiVP9vC7jaUlcUmGAO96gwVkO3vWvUKGbk7ALXb7m6/41KkBeYcdP2iD
me87y3lAm911O8JbECghYXpheaxUCPp53XW9AMwqKqtKI50KFtyoj90q1ZSCtrvV
q0H5uGifKBw7NcgUzjEuZdqa0nZr70BcAMpm04//CyW2v4SGwxXFmmVJzAoJ3OeW
gziiVW14kLLICkTye2g//jv+ig1jKejNsrSAK5I+sUIsewCw92xQPThzvCxLHs5G
UV16WoIeupnbqomaq4+MWeAlbJHyjzXEqrHqycWyTkN9aSjQwpkct+awM0euuLSY
5TUbVCj41pqKUFaqWyecJZQLze0yKVGqxCDWYE+ruyZpn7buEv61jE2vO8cmdZKX
wZxf4VO0cYIUXZsIJG4K7irdlvmcHoSYov7fE0sBHRklcQNNAZapv37AoUPjVi1Q
hOy5VtKDXeXlc8YkRGxgtS7XqVqKfilkUOsPjjzo7+3cbcFdmuNUcfMT6VEzPbT0
WQKHxMJKXm4ema6p1vu7uMiEALqUEbjGe33T5hcJrg5Bm1ahscFmUrZgp7RtM67W
KTHOuLLdG5zOQreq/0PxrEtHlvQ6MrDdAlJBfwdS0i12vbdG14+TWOfCsXk1TMGI
JiY+8Qo9Fg+BXh9M+h7m+BbgR5VZ6iDQ4xdTP6u0eFB/+XLAmVZ3auZbD83JDmnI
9r11KyKESjAUgcqKrpxyaZ4OlgYSuBHd2xSRoR3qKSeqLCDdHOt3iJZFDN8nPP9v
IUk7t8Se6ycX9Qlv9ZRe2xp1YFKE09XlDaKs5KFODSRA4rjH/trJGWdoLfo0UgFs
Trv15uc+HyhX3Tkhqow8A88+nKRsyblTXZt7LZR8a0A/nRhCzVBQimOagb8xiTex
yDb/JJgVQ+P4gmnkW4napqLYrIQ3AsL/oTKoykeKxcUoJdbEPGBZeS0gIWUDNMT0
jp+ZkJkn1gNaXEnnXkzGYGEK5esBLM1nyw7G7yssLzMcRfEoQk3vYilvJvvgp6Z1
iwtlMEW9cUN5cBc/ORrQ1/ZcKGz0Utj76vKkrgh2oTcE5mnPPOJyZ5a1GtJZ8ziP
oh2s++8t5IGj6R2eVzpKYIFz27ECfXej42kawuUY8qJ/mYyvPU+wlSCze/ju1qPS
yoLWQ0JpnsoCz9ON0Ve1aC4dprEKmwV33LAeF2mRw1cmB6+3MLk/fi6iNLVVpygv
ZpAznIVfS7r6BcKwgraxR+h+lizfkWrvuRQRUd1sUr3k9zu7NUHLjj/gTwfqNIId
Xw5sUNxnCXilcPmM1JhlqfwKzGxt6W0A/OcIGNuqNAVkT+uRKH9aMQGtAvkzoXW1
GcHG9IKz9oMrwBJn26yF4W3kHwd4/1XLb17zvo4T+bwVE+N9ij1R5aCMBGNCPOFZ
zCh9085Bhj2MLi6gEeIxLieeUM9qft8NyBEinl7ta8hb6LyzSWr1JD0H58bz6SbN
sBhlbr/7Vzfwv4U6jzaLifA5/tdoli45zgk+tZm23c1wgZDRV2Ksr4xFUtm0BQdS
AZRNjpRBW8vFkw7KjSClNDJi2vCe03pm7ZiyBscJgDbzcmlugW8hwnUTh6y0Aw4R
Fg6xTqR2M2bHeS4CQwUk72BI0UBo9QYp1V6x4bB+KLBmnTlUOJtZoeBIX4HEd9hH
/wGNgCz1EJDqbLx3aee2Fun9vG1nKjJSYgqqgnC6UWC9mur22Rtnk3TI/NFePy/7
v5D5/KYNxuTNSYI7/EH4Rs/0e8y29X/GRogNCvxO5+xAIkAeEHDoRThvtvlKxx9b
sl/TSwyRo6tiXuCtWjo2rxp9XF/9Z70irmHUgTNviDD/Egh3hBfMTK/2wcPdXi6L
iYUwhRz5cz7K475ii9XISO6w6X0YN6a7ykQFUC8FFSULXH1iYzZynTWs3EvokZub
i9pviqKjN039F69l4NDHy13IDNl9Oez/aXUIiLtshQRIyMnL+l8N4qQFPsjoQT8t
QvjcFz1Yfx1jBzq7xiqr4H0LeeGGJCSjEcjVyDO6lOFWp2xqR8860+aombeT0cre
wK+mJRcLTVOqodgDNZJ5kAXunxgdErLPS23dXEBsljFc43wucOU2zjyfE+f01raf
N+vMSDBPsRG2PBn3jO27MV8ZKWO8QhtqDF2k4zsnl2apgE3un7oin5OjhUxLNIrh
a2x+xEPNYJ2SO/GEA4sRqs66IjmslnwFI9mHaZCb0Rj1ZRYy9JYF0TgKa7Ecf1X/
UcI8J1l741TJ0Xd+IX3DhjagPTMR0V7Qu+vNxDNYFglgTIogyHRIzppdPOrg3Zng
0Q1/RXIy8AwRNR9MGfrOSxsHoyB+vf3VnR/X9KCdmURFkK+5GiGpTs3gdcixUDfQ
t5a9phBo3coAwQgxMnR6gcGxTLT9/9EMgyXF2hz5/gfySu1BRVBxGOca86elK+ZY
TIFHXMNorbp9qU77opM0LD6IEvsfuUX+JRq6kTZjcOVbS45Xl7cLS2XLqG9lPgBf
EOm30lzv6KlBQDCkIEjaBSZipEPSzIf1pbPaHHGrtr1jb0k5RL3a1hewjuME6ttN
MscjqL2K3T1+DpVRTPtV5Bckadk+6/r74OlPF0V21avisvc+Pz+/EBk3tIBa8E7R
FWXOEdt7qYtudXxUgAu5qIVf6SHvtSB4kuHLziqWaq3bgqcPH54KYn92jN4AYL+W
Ul4i2IUdVv7e3AVPEaLiYj+dnX+8SqDPuE0G9Z0KoKByZ72fBtu4d6l6KI6cZW36
v37BUWStkFanadUnA/0iNPbowh1SNOMnZww4bhRxagFP5rbdiTzh57TnV/AuHZec
8kvvrzP3cXBLbT49to9LX3SM5emk0xw37VkB4E4UXC42IQ3AvQX6sbZ1QcX8afE8
zlsMsI+fVE2pUC7fVdJX6dQ3fQXAcpyvngrbA3L3gfmOXTLr0FGesVmNYBC+/KW4
sC+Y+euWfYTeWLqaIiBhPTUCWCp/Jja5z107UBKGL2NPn2ZPOKvpsbcN2uwfR4/K
E1X570CBgcg2cBPI1WyeuEv57kt47z47hxROoW1jjG7mMyF7y+nU+rDBg1dCn3g6
Z1s4jQmBQT1UyjsoZ/1Df9QmMflL3L0f4bnTHfqQyBPzwpdFI20xBhcbB6qc6uO6
BneWbsi8PtnUgag12/8CVANZVRN785wTsCrlMwYpOdnROms0NT5U09NfGPA1TE5H
KXseVb0+QutAgyxUPaI4/4wnld2tV/wUrS+PHx6mKjVlBs7LGz+qwad35SBPmc5U
Gapy02NeFMHo/VOEgqbCsflMKR7/wkrtM3rybv9M+3NLoM/fRKl+KZMyuXNe/Abu
nNowgSJaRZ4EqaZPNmfMCnfJ1Srx4cml0OsK30Y3aGobMS9Anv5RczJ/jsxR8ttw
ulZrTWLEGaI95b9qJa+QPGbYNVqhOx0jT5/J/KP2OhLp5uq8gXxmZ1cbRimNa5uN
Vf8SabMpmv6mwR0QjMGSuHpMyJctB2KenmwilMvcsYFG5MSJFHBqhiu6KtPxNelv
ssDWMwChi1cmR4ElZuZJ8/21++b6rFoq26ZIU3DOythl7ZWZFoZn7+m4VyY3XumI
TZBLUMt0UuU9Dw1WGoF7w7jP+COcKOUppIRkrpwoyXLM9rRhMLXSh3PrYb4/W8dB
FNRiOkHjjumPsI3mNyulDDHYOtSQk1Eg2Xw9IMS7USZTW3ULiMVN0DkAWdHYcJL5
Qzep0wu8UMLQJOOuilCnjK1y/xDMyY0p4pAaqpjS/M4AFZJilajo5rUS4M090vhe
BslaGu9WbRXzw94/ow/oNbZsU9i/ZQ8VaYjGWCccF6M/wzWw18FkR5qpB1k/gyk+
OYJcf85K949nj1h0+N1RZR01b13938cPywcJAE389J1EALYnC46uijCQnNPu6smX
di+ruSyzF2IhvzmcJnwWuxFm51LOL7cc5pM0DOcHy5ry7RsHIsuE8EimKYCF1wLx
nM+LlL+rva6e0n8t9HnNjuB5PKpdaK6E5LYjufSX0wnV5YmUNH/IVygWBNSazmUp
mt6dEdVTZu/FMENov0UAdxIsD5YEGU8aH38v0Z/RjUCkYGci8qcMTlEFuReIr0nn
DLmdjuoc2oNvk0eALxzRL2yTcXY+hjFVYqHVKugRDFvJVPujTJLOaA+Mf2AeOwfJ
E9oUOdzi2V5nLQ5dQsK2RjwBBPZK228WJoXFbUJiLCEydHLMWrHX6HY10bePR/EY
Bj6Xi78adufkK+SoQgRfEoMLXKl52+wV/qr4NYk6uVECYxIY7hzf/S0g2AHFsx77
ZZVz3G0UopzS4M0ryZ96wCLnBh7Rvjlfq4IfpkxlaX65qwZo1TTEjzmM/u+vfVUX
tBcviZG4lWYvFJ7O3dbrj05nrEcPvqUnxmV9piVO66N5oysfF8vrse2nyxjmPgN8
dy58hl/kXEc9NCBlfLfInMkuKcB0ccDDeE0aifWbUbTeR2Q4arufO+w6PBP833mG
XRMFKdtSiN9tP90W6tSCcfwcJoktq+NdzjJsyzv2yF5lNS0BLbLeWrS0eWDZgOgS
VzPHeYdKWob5wRnbelzdtb7CuHagSsytupEm+bItV5pJVf3at5ppXgGdbhcmzyQu
ghJ5TPgPhSslmi+563+MH3zaI09tPBmTi23Js9fb53I9hajpH0tYh7iSvbBNKkj3
AWbGk01U4eOloyic40WMQSVVZXa7QKyYrpeDtEQzxfxbE3mZ3CWo3oTxnGZs5w8z
/Z75Q0hajTJAg6vgk008N7oVEC9n8576aTxdrJOVr2h58+wYalTR9ZuedFJNWKPU
iP0vacRQhNx8AO7JdiyoloNV5WcR6sL0TvAXkjhAYBwkwhL9ymseEWqJOqUSzvUD
gtHh8fIDyFPg/5thDfmgw3rkGoTxFK1ShLl3fwXkk2HsYMPoWnF8VopCKQLYdK1n
SlGKfb0ShBQKfaIh6Dz6NJ82VaRwaNXOD1yN6kMSY++p3TQqYGp4NMXM1NEZhIYt
QIzUE16yMTwG4dgK8RUZv6QJAucEkvP22ZwZMmC6hjPEGoEKticWwbWHLuc17Z4R
zi8yzRDL1LL8ku1+ED025m8dsw725rkhV2uhccwuHqm5a+zr2lUHXGA1q59hoT4Z
sZGJzRVLb5v40AwehvMsHk1p0xK7sf08CtUnH3Ghcow7XfdakIbY9+TEcmxvfggO
Dr7o/dVH1be1hUG3CHhthKw9YnleoovlCB3g+cfcQol7gtTXmXtYDlp/okzydlKb
yk3a+ljNTjOhdrgwAjMMtU3+aosoJ18MWXwCugRk/vzfST4DUiEgQSxGOwpZyaSD
C7p0vNA/IbyIIOtNa5KFUzpoR3XaBLSmZRbYQ6d5c9KsK6p0V4r4A3vgBAoLHl5Z
i4A9yqw7K8FJ3dp1QNwwE66rQM6y4xMpk2W+PE/t3VG06DZQPaTX+zdJgol82mls
psUXOli+kwNdif0ZMkHKuXLuEIyGwXU/d1MDGMWyx0Oo9IAm+yW6RL300Jk9DEFj
/w9o/pcdT15vxYFamqtOBXIZ1EWsqV0dgJ53+wJ6bkrTbCFctiSGk59rZGyxU25Z
hwKKXE4N0rmL+NmepsjTbPw++cysXut2Po6L87hmrQwlqTRGNbft9yaZtk76HDCz
w97l5sFIlrAa++g1SikXMDhjFFEfjlYFw/8zeRMfT4mvxJRFq6XAQUu1d33QHi8D
6HfkTn6Z0Pa1Sb6ybRDqlB5oYNZsorxYJRZ/S+vlOSdMzhH8YvrLgk8TDWjjyEGl
`protect END_PROTECTED
