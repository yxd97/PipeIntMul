`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6Otuz8qn+oxVH/WbS6KAA3isSpF0ut0tLcGsf5bTXxkGzs+aJY2RbJCETNcYxXS
sRgr6DeW8wMBzGbq4nSiw8pBZWnXAjQIHx0hVUOkDBYWzO0A3cspa1benBq0Z54E
xDnM+u6x57g3gAy3PrEzBRufEuBEzuWZXWKPQZg+0eOWJ/hx0b1zZhG7JLVtIhTQ
yFdZ9FeJXYMwlc01PJGGgjKCvtgkleqkvhoDwEXRYqZQMF5vI03c37O+3BnMMk4v
SaiOMbUB/tPmx5cMKXEcDlyTcRx2pOplbxBVhCBvvi4uuGoqUn1uk+/Matm9LJcs
+/VFHrHJYXLm4qV/jnu+dUIY8SaBsnG36716AEExl+OoHYPfUb/M2WfHXdJYBC2n
+FyqKlAUj8WFWYEnVVsHrqNfHiT++95URRSi7x6UzvHxJ4+Rl55Rp+/Qb4R+8mk7
xN0b0rELXN7OUSYE+6S2aN/rnlbWq+PdTJ+vs+KUpgejn5aa9jbKGWRO7V9DY/f0
rJytWHdmvosD7tQM2BjLdmFLH0K9rDidPsSyJxCfMszLeG3yOCRf0PkcVcEOMtX8
GE80xFV+5zL1zki3zqv6ZW746FkXrehEIfuTw+/0tMtu8PS1L7saLlpVzkGX8zBg
7z5YKsglK8ypEAjI/CKp/pohFevVvfrMaUadGrenQTtKZ7VLiHyJ453wm7Oicx3F
/Jh167xdhyDXVjI/w/p3KG6R4eWpUAkqgzEMZYXVcfer1VF11mUYdTKMiC1d6gF4
xI4+cZVDVUhIDxUJibwFbQ==
`protect END_PROTECTED
