`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HXXEscurXf8ZBlwbDwXVTfII2sdRIwq7lYjEERQ6qx+AMEJ1G/ptI9v1mwloh4VM
suj1I+wrlThYa0pPJt6LLYV6PWa55/ONcIJ2cOizl/wqkHCAMbCAIzilgvmApqVj
qAtGlHBDsYuAnaNPHZ/iAIX/a6a4xPrZZe734u0+5Qh780S6vkO0VZESzCWd90No
AZ6ncxEBexnPg4EAW7BgFWcHuSIWtzGr3mA1/iYuQUso1JxwPNziC46ixT13YNCv
veIfLfk0TcVxzpJ2dOAmBeZfVXN6vcS/2R0/1ShuGiuzlNvo1mYobBbte1cie90/
y9A1wvjsmFvOJvMmBebfdA==
`protect END_PROTECTED
