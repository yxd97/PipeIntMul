`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7AUdpufe5ygcBYV2ueIHcPl1w4N8MY+TfXjS+Tv6qwX/QqQxHx40jeE3Pbj5oTJ
SvKLKN/JY6pJDIPVUIOtJHlZSsrFLIMnL/1BNnH1l4itZUbazeJJ2s+NYluR6RRD
87t0QXXBtE8TQwRk5imfNOHp3t/51Zqdo8j+CckHx3Bhy7rrcuDnIVbalGx0OTG0
1L3vHXx2A+ASwrKujZVso9o23k69xPaqrQ9BnPg6guLjxg/aslvJ6WwIQQkF365u
KAKhg82CTcNRfqYMV1v8UH0gWmY1Va0tCbhx8pRnDxW8nLDX+S6zsRSbDqwVNrLK
lVCQSBFchblmkFGx6PgGs6GRrHig0F0D3r2ZunTYqeg53LuIX4L4b59+MJYZjT3i
H1GTdcOw6XKMbG3DpLP8gw==
`protect END_PROTECTED
