`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9OkPt8VPdEXW+FHHG8QIN1Y9UTjjZS4MAtbasntet3lTiLwULH5cwZYb4iJdm/vM
7HYO1T0LfEeVF3PQQS7sWPpnKVy12smw9a5SpXLWrFA9JsBvEkrpdFSjLHluaMtm
94SbdFLVoMMpyQTmwLY5BJnhhHxdKD66TV0AQqPY3vn6BXFfwNBjmTmEeA38+G+Q
mZtPDBD+3igbW96mfoFkMtWAeqH/9Rv5bcckc0jhiCH8KkJ4Bzptldkp7I3o0jZl
F559xuJ1owzfilF0HWpRs1PvE4F8MahAkNQ9lqOxXm2xNYEsOKvw7agsXIq522sp
RmmR2+qzizFPJHG/p7xNd2HEgDcuegEQiKu1KdorZCUMVfpb3QIR3I3OugdNzC4/
9dkry+8IXTU85lxwjjyd0igjfcG88EVIIQDMl6qtiwFEjOBRFqj0cES1MbBfAYDI
2fuJxMfufpEKWWx9eV0mR4CIOmDcnYEAO2gLJoBdvKk=
`protect END_PROTECTED
