`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWaijthcRmxCkavGbDFHi0po3WmFxp0fMAEsAumq/lL8qHys/wg2bEQqrGCSKzTs
20nnzYCzqqpVW62HzIHrlVscbWA2rfN7CI54Au+2+4Q8sm0jYZO//MTVKrvF71uG
7NQxPUXnveSlLg0XsSv9tbixeVooj4N1+SzHFzmumYovV8Td6EKwXgmDx0TRveh5
+0ZjmBcwUX42FVqzr+ISVpHWiGwt/h8goJMWLw8nsWD/3q2f6yTLcmG3b1HWlTDb
CZKjTFGa2jcamlGxc2zyDZ3BkznCDig0AoGmYGNHiQ/Im2NqhGlRhQIZzhjgaBRL
M8c4hFlmtudmHtdGmzFe/+VFFb5U1CZbgF/wajpNlvERaciqWTxy4IQ9oIv+t9IS
p+0iUhQrboJaTBCj25DIJTpgREZd8dMAWxs9m6pU2K6GRv/ihJpXb0zVXiL/+cMB
PHTpBvLjBOUeG6UVHWV91t0+GIceul1uGxKqTDoLByr3iiHFvg+6CsQ5iqqRbY1v
TzVnpBb5HmyzR7E3XqNzMGyl4tyym/ma3pWfsuXIIfZdr9VPAurCtKNtsBseCuao
5IO3Wq2Fq0TnvtIXu7dzVimJow4LiJu2X9kJh+0kz9LZ7bXyRh5p0Z5DJiy01b1G
Q5wJwSm9NwQK8GShWm85hGvsTVaGdGdG3tYJ6s/VkNjRpiPMX3Vz4AvI6OED2RPM
avMtFqBiwclwUlASeIqG+913e7LX2DLZwUCmssrSMvVhJX4FanSyvYyHjOF+7crH
Vt/JX3i7OPu+0k1ubtbmXFaeH2aZnH+Q7D7u/+buYiXQkjD107QpTd+TxRwKUEOH
YGR1Agz0IVgEAXObvaiLkgsrmVPTh9Mh9tp+1eHyfrg=
`protect END_PROTECTED
