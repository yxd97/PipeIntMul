`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GmNeKqclUyi+Zua9ffvvxqCm36wv1nxmvfvpSe82JRu8VSgkVMsYfOcotojLsfHm
kEf4YQ2VEV1iTbZ2iWrxxH5KaQOMfS901rDB/KvHZpi9J1/msXhsQefcDTU4y1Sz
Z1VMcZ0RCBIYfkhOW2TaRdWn3GeOcWgb5HPulF9+wd5lz/5MDeM1qrVdns5DB6tZ
B0PLEVbHFUaqWroPhQOQqmaoZyCt+InhHeXwTOlfKsPmOO3A8D4D72V1X5vKQk/s
Hnl/WNnSFPc27Jjl7wJ91R/D2pYF8gOoNq8k/BMvglZbef7OapkLeMTGBA5zGMVS
XB/WTJ4zCvlPLWDHBWV9ugQjizxGLcGPGyZxMOSMXzD+fht4WL8BLp000BV50kcm
5TxODa0iJHn/jt+9bdRC9V8pfyxxmmQrRH3xsVWsWEyZcYg98ZCWcIw7gP6zOCm7
UCiVQhXV9NEm0BnvTbWuG7QM9KiP+UAyW1DTHdD5OZIyfdCYvuy3sv7i33wJK2Ob
xdibQ+oFGeB4pB4SxNz6mEAtWPc4aqQXNKJqRrj1uADphuVVj+99xl2h8nRYWzVN
YE6xWlICHr6tkjc+oaVCNw==
`protect END_PROTECTED
