`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C9CJHBlohz5d8IBuWwuqpcDjFTFnjkAF+s3kh4n7+R91M+jcqIbAFNu1Jxz5tbTR
zI84/wuxcLKfoQBZQ/TVGxyEJa6YsMYK+XQqf24nE1XTXBveKNN2qLB4ZwoPvck9
Qa1we6qjMgQFVZ8NSuZkOJEI8XqQV5KaIoUpf6lMatPbqD9BlaKsKKU2c/9BCjsC
bUvOc9lnGG/EyT/86ZbDmNpIMsxnjkOaTQ681mindf8wesB4ce1Fdzze4ClsZSRb
RHy3ngqFBZRqa5IhttwlsGymvQjEseL2gZGFbCvLLlNoD70MuiZmia10QZd9Njts
/EjGUKUf6jdGSt2mIAj79zf9LdGHFu81KssW3111k0vC7u+x1f3iIT+6tICmVYXk
eELjwUAy49bFRoEV8QsSDJDCHIgtwY3OYUZ2ycQYxeusqcv2v/R96y4+5UjZdb7u
874LUiW5t2FgPAz3ihQWFAjXdPfHiG9uZ2BCeCbTzNKvhfBgaqHQVv0x0Pwx1lEe
hCJKqrTXen6QZRY+idjlc76yGm3RD2ZZH3JzE3H3w1vbIoW8D4RBhQo6dSMlHa1B
hxxgDbCqdVNLUGW2xEYFzFYmBYeHlrauI+FrDONcg//V/BrdFn20Yl/SDq4oCjLf
+RpA6lyY9rBqmHA1hq26Q+htv9IYS7lTmJTkvKNpp4VPBs0QweBaVCYh8rbkWFAM
MzaQ1EnJl4+RL8R7i58eXnLwRcHPN7EEB1HqrZAxgdeOoYV4MVlphv5G5IBQOEGF
MHBArY3YuoRKQNSM+x+kxPqqwZOcPyvu1DJqBHAAC5dHvSqDXUzPtBCBiMnd3pO2
x9ICJs8AXkY7nGxhwa4TWRxE5h23w4S/pqtDaAKGsO1/Ud6emLJ1D8BIY2trMc8M
1XlV2vkexnjMz+BhlYF+FTAWTYwiWODYdbQpw5uxINa5JpYP3pgdXZQMY0m3UK12
`protect END_PROTECTED
