`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/m1SE9e6wj5Orm+8Hqyore1bdKrEOpKJfNOIHEivdq6oJXUERjS9kHIc2e+CMqd
BoeY07asUPrO1lmOoeshu3uJrXGXTu2HNOIS6ewCi58l53CcWDbJnLjk+DoE0Bev
q1Dmlo/R8cDb25KqaxYgI8MSOYZ0Drs+IpcFAs/E3HfG4ylMf39LNHdzEnFjxGW9
FS8veJViXISGyzpDtB8gm1EnGXlCgGt9BIGe6tD9fX8q0hs5H4b1ugF2tXGY8IeF
YfwZqszNmjDeR4dc4XHPPfTOMxzNW1HuC5ciFtTuCnxzXq/KvDMoCAFheHoPZs4G
7slBc18X31frIVObD/sWi3bDn3q7YP42SIuiMY3i51K5wgYeLBzVByfSrTrP+g2M
i6mpUACaUoVNXIncOQWSozqOf+2Zf0SVth7GRwfOQLSqM1MmLIsLIrU6w6KFzEUG
JfHCMrwNE2l0/GpOrXseozjJ49eivVu7VpDq3A91B43OY5d5hNW//eBgp8a6/tPq
zEURCr8JwOjWFIiL8QLQELT2PD3x0Vz9DkdxKwV4JavV+a5ZhwOgRmgsimLUJrMM
aGhycoS9CSYhHrxQcgFNLvEty8XOn0erS/Dxxa+4xjjHqZD74CogukNCtrYa2zI0
UaJoVZCl6boJM6CKJ5aihOiCbrnbBE75wV7hndXqJH+eATEc1sgbGku3HdSRMQRp
LkWJUcmJJ1Y9fYKrIoaROFV0mmYgATCuuNpATFoTeUlWoKDn/+oGWrajYhxlywaJ
OK1tRlU+z4qZlMeXSdoEXkOhhSqoVyP9Y/xgm7MWFp7Y8IEvGAgwB25kCOvdoicp
oV59+l9/+beSkCR99NinGwVbqwhGJEMZWEWUzqsgJ2BZcR/L8Q8H9z1RwhbjARhf
jR82ZcXvYU0A4UCDbsHHNwYimLbMCzfHJv3NyV7aRz+pgQ2p9AfGIhLLg+QlTwfi
L9V4s73Fe/JF5tWOzk0TfxogbGUuakoi5D75B85bAg8JYWBlUTY+WBeZyNBypDh+
ddb2oo1UDevP1awNN9QHLt46K+GdrdEIVs7n8K8zZqOnSbxD5iFZc8LHH6mWeT7g
RzJlGrTr4o5OCCqpjox8dCorqE4++6K29slJLNXNpCSAUCj2zCUHL9SgkwS2hA9f
Ys8hq3Tube4Zl2p0XcgVnq++SNpgPea8XeUH16YYbz6fD21GQ5Ni6EhfK0OShQ5e
ZmVu+f76r26HVZlHtto8s+GVJL8kgP1xHXVWewhwsQM/0xHnwYdoeb6hGqIiyXyX
QgOM8xYEUvFBb+oH/n33VlMtbd9R8cDdMvyn53xLS6VRDpRxdmzA7EDHCOrIx7PZ
WcVRFjybKDIrvoX5/qA/C6QtpfKbRNS7E/jUMsc7uaOwYnSYXcWXyNXwjvdBRTPr
HJF6z1KKIEy6BvyVRFNPsquPSpQ0ElBRBz+W1jCqtZeMMRc3kJNuzbtiwBGhFFlk
e2dYPnib2qGmjYK+1HHKlUXw6O2q4e9vpMOozxjWv9EoQcWP/seCQbFhbg7SFtPw
eS5U+4yyljHe58omVIvaQZMMhvyx4IVExqqSrIL/JQ0/DyU6XRK8pFFgyQV95glu
Ik8pIhoVZf3J74TJtbyn2uESA2QkM5r5zLA390vSuVyxdEO62JcZnvyb+5BLrCh+
MjqGGlnsxGkqGnHY04b1BcENWdUnhiMqoxwP7MhlpM5nB9PhRJDTRPvPTpG59gjl
dMYS5NucMw7WESeFTqEY7obvl3PR6oUDly/hw3biW8aGkPwlQRZUx2PZKzDqrYZ5
xYC5ualPXaZtXLZiz1wS5tcnlVK/go2dW62/eHoFIJgVszfEXnpbkuMLoA6yVwEQ
aYyZkLHEdc/42iAJW/zC/levnbEeF3x2/V1rNMob80uko6i41iyogO7gOL4xKPYr
nrJYhnt9dNIAv8Jea4nBJY7P7OfWXrxfAmA0UJjN1FRvW3L9z4HOnrqYHuuEH6h/
gv9MEKtcrTAyE9Nz6uJaa0aMiv3FqHnd4iuxvZ0qH7WZvnSRJYun6Npm1Ss9YWW2
LQQr6Hd92L57hVpZ6gc2SXt1lGz8qlvF1PDUSES88gE=
`protect END_PROTECTED
