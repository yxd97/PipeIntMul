`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iz8Zss/F5j9tKADzpCMepjiYpnIssMgr/wkzCsBdPjZ/kkd44/AzVjpDKqJ/5DXn
LMEP1zs3f3xl7ZNgenBP7BfEDTQ7qjcPVMFBL8glCubdwvkYJRSFgDqPM9tLb1Gt
C+xul0pxdeqlGX33VhpvWbTaSRHH93PUBLfEtm9zjbka6V4kMCAeAVAU5gn6Jwi6
2rVe4ccX3QEftDzj9DE9uzdKp2tHZvwHoFuClSD6yWqM0YkBDRYs6KDdg5sKKkzD
amuX9NZMljjhgzuBOqVl2bowNZKsRy3mmkfXU4vX243O9UBidj4dOgH/1fCdQ7SG
u+BE/axRUkVkHfaI5S91Nd8TRbVf5lVYuPfnupn1tY1IViMWlNSoKe2LPDstAuf3
hO3SETTptqdU0vO1upLMcnDOqITXrnVzwuJXlVzaZPxgwt1q2DRWNgzb6cj2cs7E
fopb0l/gMktT0eTJcKPMt0Vq0Fx2tplFyPSxoB8YKEM=
`protect END_PROTECTED
