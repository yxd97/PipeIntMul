`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZ8W4Agb7Yl+C+0pk8ms8hwIplegu4lqIK7CW3po4HxzTpaWHUVrKOmuiT0mmdJm
p5TSEe5GDlbb315sad2XZmiAKk/M5kIHfZIUUO6HrTNSLEmuM3C6H1N0ncXetg6+
JlAjztqx2jDupHxCAtHui4bbJ3lzJ8npc3mjkVMPcAtphQ3AldLCr9F0AUQOtD+p
p27Px43CkSfKfwVsZPpeG7CZNiwJLzr0AHFBVWTRIo+DMvuJNEKEhiwk6gKtyV3m
Bwm98iTgaLdpcJCCf9F+4ql99zLwg88XyGDBsQCVlZBb6lMKW9fSeDHFJn1T8HH9
KJoyfFb09DjA/obwzjPfxJBMOYXg4RIMHnh4BHNYU2ei3W1grH8zwl+CB3TS3cY7
rBIpJJMby71n8Pf04JaVl3cjNf0CHP0dmOJIwFjdT4rCHK7Xu0jcyMgg17GQoIxi
ltYh8v0XhhZ6Xlp4zqieqhHXDW7vfKFUoiZV+xhEpa89GKNi1qfpg6hvwN82E0Ix
OWLrqhCzw6nKvDO9o3cWb+sN21EYi85kGr/a+DFFwtaVv2+klQUwcWuJFr+Gb3gG
mARhmucagOYCK0CRCJ4wizOi2gAh+3XblWZAIaNN7hG/3ezqhkqx7Fmruj0zr6B4
Thuc6QnkBjkyHUAhu9Tw0SCl1nId0G7RSE8Ly2XpNyr2CqKKZLjoKpPTIjUoySdw
Awe7odbksQBqnjSwI2wxjRWgL8PPW8Rc3mxQjjAV2ulEESeKXu0t1JzSvV303K0M
BXDBDjRJiC9jOXC0HE4oZ9g3G+fSdqxsXfx1dpmC3Md8ZjD4rlJY2qTNHrAv8jAs
2/B4DEd2vXjBD1IneD1oVeI2BIcc/t358HPADsbepuQ=
`protect END_PROTECTED
