`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QwdoRKIEVGrAvtEfS5DFWGEWfwkOt8CPROjvgjnGhoC428BC9p9bWpdX+QrJ3rkO
BIFLnKHIPoeKcUk5MlFjmYEmYkWNDvtJxoB1x33yVhzfFnOKcYEYXhGDbQDxGXCQ
4c3qIijuEd9urWiCj9I3YEjS/vYsm1TnDxGvdisln29ptGvdOnM3flWmpnCTQ4zX
BSx2W/w0/qpXB4lLp3KDODV2hZ+K+SSB6gBWANrW95qP2CGMcuDM6BDbi5KxiLpR
s2AZyaI7lmRzmhcnh63BDyfGvbjjStaTErEiH3e+qIppAotRwxHXevs/ZOZ7d9eE
AT+OMuJegByuHWhITQiOG5BGtVNgmZmi+zIQqvqcET31laa29ocdJr9fl9IHqYhY
tL3HfO9MDYIYtR7TxRuiu1PotAdohWPivzweQ2RunYy1harJRIyLwRDfeJ8OMfnF
S6eNQw4+bHJh4UF7soVpBEg0kf4KUAKRwNG7T/9UoYwQYfd158klFol6tYKAe4zY
Xmb7Bfs71DpadAXPPPvWL1nfphqgAKSRnRlas3wkMAbmM/ahyyeD/971X4kR8nBT
nrQld1XpXuIsrHqVukK/yQ7vXxEV8Vt7ca+BiO1f2545D82jzL5+uXWYu7iAB9xE
B3fcZ3ABbebkqTSfF8oCNg==
`protect END_PROTECTED
