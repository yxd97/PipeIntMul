`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/N3exQC+9Juiy1bVDmKnGzeESPu2uFL4AWDuZw/3tcLexQqPU2jpW3Bsniv3Ie7
Ii9Mew25R/K7XkjK//0SbeQJf5rDvXySSXwOVUxusurp62R0SRKvPJQb0+60dvs6
du5ZPq7tpDwnSlgjAnlLSG97dLwpbSfr8cOCioKMrInL2GlWFTrVwBQfMrXch3g7
hD3TudkJnABlkjmuMBhR6BaJeztkiqpyq2gusC5Aol2uFD/TfIZLwDWaGvGFxgiN
jyWUq+7gdrqcwhsSmW5qAQ==
`protect END_PROTECTED
