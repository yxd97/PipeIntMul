`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyE1mWaImdz61iFdywl/DVwJBEaDxPkUcnQ6FAUEnODg9BsXBzOPSmrdLqHc8bLe
jbviR6pugWIifPUWkN0rWHw3jiUwMCmajy/p7FbMuYgjAD0M8x2zNUHVjWrsFvVw
0eLObS3OwzJ8pqCQZGpbw0c+ZKv9UrZ5My37egt/xA+6QbGFY9hYsxZ19Sn4d6cj
LIDrVx6Q8ofHGiU369OFTxqEIXyn2TSya65gIWs0o27cqZ8c4gWdzLLNYMYFvO53
yrABYrpi0VX2k0QSig3dg+lc6ebGFdFmyCOryPTRqRGkSqOsF49buwRERvH1Nk/T
57fNgALre8LbZVxTvhLNNlropDd7uoTqlypScxjVfNFsyjbtc9Z+HIiiZeNbHtiv
Vb/OzcYk0Kq7x7lsjdVyGn8qRkivDRfyRi97Ie5dL/JE8dwc9quKND17XR0iWUIy
`protect END_PROTECTED
