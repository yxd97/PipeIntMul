`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcR4lcq4DD3e/IpOQ6Kqi5WIiSwzRhojNJuajyQcvS8Q5Il1nexgaxcUBESMlp7D
e1DG2O+FMuVDC/y6sAUvHrElLjep4W2RQNcnzV2feYaCGIG6UdFlTSnjsM7iX720
uvIGADTZ0I71VbTg2SlpRE4QUvZ2z35OtJvapJNl9XCbyAcX+gXDYZek8KF89toD
8KOCeljgWz9fEXH0R5sexN+Vb5SusqKHL+uSU6WiP5vnFuwbtgA8dViVkNH7Z5W2
qnQiZh5hUIf7H1W6IE6qG6E71kT552+DAeIGIwF65Z65en346Yjd3mhYF4CYWPg/
ozqKJKWrKXmqc16HijQGcBg0yRoonW+t7CAYAlhLAAiM0HhxtB45NmNe4RewQ0hc
26GIV6wI9jFcaZoDqSNphsPfLDEhxtDhvgNQlzr8hZAfomC0w08z4bewppLiyXG/
dLmK/c9BdO++lmfX7IvW5I6ciKTHzGBy21nVJFwwHxql2JNzTE6FfM/Ch/ev42nS
`protect END_PROTECTED
