`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKUd80zY2xYp45vo6g2yNKL2jmuoAjSHcEYvG2NnU4uCW5P6pgYZ/uUaCmNnUKbm
pXl5kjgvjtsNym7D/yjXsK4E+9fXJJdr2qamcBRuOnuUnSYMH4BgK8BpweNDLX4o
j20AbyaPMnLJcklcVa6f3thjY+pOfDYL6asLlGV+Ab0eNMkF10yxQAgR9oggFXAU
y6rQ4ejFvFUMicfL9DUzw51TGntJkInXJJ1W9aV23uXNlgbRA5WIrm1nlzU8w4nM
rrYKVSScx962L34/97HJAoqwlImcjSyGy6CU8pFKm3MK+aZC9/nfFpmfXjApDWDM
Ym50/4S0anla/8fKqOFAsgjRvxEGGmlqnTGHgTC3QZo=
`protect END_PROTECTED
