`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d05mnET774S13a7PPTwC6iUhA/7lC/j/ye2kYFQLpF07t7AbQaf80SoK3zJa3wqN
2W8JKveCWRmcghsoO9oSYPmIZ7YFMxxemMzXXyrukkvi+FELDjgVQ3jofcGFaVYd
O/EC9X52MdTx+csi+f+CVHh44nxmMpOXmMa1Am7c5PTM2yeay1TbszPvNpdjOk8U
aXaC6tRkzNl6N7jKVr64B7/UvP/v8UuY1nNrMhXCb6SGtaB5NuVU9tzsATedCo44
/L0HhyrwSAMuoDl8Tt+Io8FMjuK/vWCnUlb944roNoawS5jQjt5JyzfJ0V4iOO+c
VexGeGvmhURZLvkQGxUIIlsmJFTm7uD0798noabBRf6Ki0WTwbLuSGc1iBPdis1f
0D3EmHjC5n3hD3+F+HNer2yNlTdGDmW7Bkt2dqehYnUCZnX69xuzaZRkomH8P5GQ
`protect END_PROTECTED
