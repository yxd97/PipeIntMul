`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H4v5tngiqEVYksyWPtVx+9ngq99lvxffLAS5zlE0h7pNutrIDxo5UVOllgzzIZhf
acGA6nuIE6EAJi/Onpqas3DdYOq8W+9krwg97q1Mu4G+Bx6NLSL9Qe/L2bp2NAXJ
uqNH+/lbaE0VkWigwIFefa9dCIixOv6lc7w4FL8k0zQBt7+onRTzONBEexL7wdnu
0a+zUniDwN75nLkFZbss/euCUjUn0k8V7S+Nw0JpfZO6ElSX0Y8hPuVC0ZyR0pRH
eVshlZlTch5V78o2LbRwVCkKDiVP5Y6PskkPjoAr/4tkxYob7yyL5bwStbQpHkR4
DgNNyrhRurjJ1srQ3cvGf49Oamo7lAm8PLP/6NdwOwknL9nvDvFyKEapsFpT++6S
rr2c1TCi/bh4/kBHLdU/T+hE5bpie+uu2FB/sSQ2PauxDvq29kMloGRFtdRxOzu/
v1RBc57+eVfZslOYoJ6L8Y4W63OWkkEcfzjyTdxBz6liDhVrAltMzboLSAxPssCc
/Og1ptdmhP3n/IAPEC3GT/avCr84laX91PXnZNnU7W54QFzCLfthH6biDMGO0Qj+
3wy1gLgrQKh0BVhGRqx9Shnu51NMbetL140AviKQj6NZdBLdnDnSCzIU/AKfWGYv
2hXNOxN8W+T4KKfK0k+OC3Ja0iHfMABUBzk90H+wkh8sZnakfGBztYBdlTAOhnuK
XoY3tnozQt+h6p6R53ERfoXtNSWJYxJT5yCkZiVvyzUQ3XPHPwUvOFpKpe2uZbCT
4BxIIm11NXjIEhU4P59ff8pO4c9mm15kxb2vmPTS3oj2p7ym67W4eBH3vJZ5I4EP
e5ysU+nl5ShXCivZQXSXtG5HdMwT3jFV2Tei0pRogEyHKOeFWK7GeHxDEGaYaA9m
nvHtx3lzWM9+hnRe50a9LWVyRbp7D+ZcBMijYqd0ZCq7feGo5U+UNkn62SL+ee+w
rm23bHnQfvN4JNScDdaztw==
`protect END_PROTECTED
