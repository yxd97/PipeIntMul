`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKCRTRUZv/2otxqTo9LUXkcbwadD4NoUiOKHlQSpZOa0atCvk1H1IJdaWi4mXSQ0
nh0x0tRrIuY8Z/hCQMG4D3jURcD2BWNfhED1lJNfj9YN9ExtQ2GHUHtBoqlQeqON
CevRT2EubkSV7g1e5Wm9p8NKZfw6j6cQtZ6d5j3kUh7c8/N9vmZegdJRDnggKseZ
KX++OLKlBr6n/g3FzRfXVWm1XjFxJBPVH4uJ62wlHnIhXOnQaoxMDpIfo+0sj2G+
BIYfoq2P5lcs4j1ob1BrXdjQuOCDgS0HrQvv+7h2WCyifSrmSMPR1oCWFtyJ7yed
SyIAka62BBLXSZwEPjTsbStdWD9kJOCU64SECKm5gVSrCPIT6G867NA0gYU4RNVs
P6/UH+70d4BnuW1fy2lrbgzgRRbIvXFX5Ul4eXYzREEF6JxAK5oEUhqzhQjHEHr+
AwdbD0BA91ond7oU0VVXbXmxDKkJHOvxTFtvla4rNvzOPiFLDQeiXBKrnGE/qM7d
sRSntsVvVSZntDzl/fidRf9Q7Jid2BIuxl94Q+W6zEwbRqojHIivmeZDpvSi3uYQ
oBqvVP6gbbD4AaG31sai4/736UTnvCSHK77k+kN9o50dG+cvKMC0mqYXTnRQEL+m
z4/ThE/0HyGchT7e4WGW2vtGwlXsKPWE67ugL1WLlzIdOYQgJjnM8azoE2+yZG3G
6yklckt8WZAx6QrvbpUH3HflZqk9JavbPiQU+gls/Zjca4oA6pyaFyKl2gT3BqCz
scSgr8miEExCW7hwGhZ4/C3s54x4wt2iXSwzTwRit7zKzdO0eCsUBLDT3OCLMpRv
r9jULxCmTXrubOdvXdNybJHPoJYt1vCb5voGPn6OLZN+Elmfjo3k9y9iOi1YakQE
d8qU2XV5j1TZ44paAfF76pX9qLFLBF1Howimlu4GMu1onnIlpjIQgLzAYhmw5nD/
hZMss+SNXNBlfAnYkRVHGXKzbl1NHsP1mPsVZjAQ758nW66VXaaxKWuSSjNU/RPq
nYxmWaHaD3/TXoYhhvqz4tubPLHeJeiwnN6B1XSOMA46DVPKJOzPgV9XIVDpZgi+
Ejxafo0timHrXi3+MESmDg9+OrWoTUqimoYWaPy+B0AH+WOZzAKd9se9YGKo/VKC
eM1VszPHEXiTm+liIF6DtQ==
`protect END_PROTECTED
