library verilog;
use verilog.vl_types.all;
entity PULLDOWN is
    port(
        O               : out    vl_logic
    );
end PULLDOWN;
