`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sk9hs4rF22PfOVvTXY1Y7Cyon+r1/awiCj5Qp2hyFxCCNPaPRCJiLK4zCCAZM0dL
zcrPeiDpwzH9zQQKO9tR0eRh520yTpWQgoXeaXnouu1nEOD7oLKstQeLEJWCOt2s
hxC7eraVsiqEtOXpRiOHIE2/N6I9d2XLsS19IPScBRkC0YuCYjo3/tJga4wkqcy1
P25tfjMRAL0tcrIIwIxOPUuZvSw9zNBfZBnoBYP6/UztD+jfEeYMnVbDvrE5hvug
+qKnQyHDi/14VeO3woqZGvWxzP6JfgfB94CvzMyevV/YcUYGy33Gv6LDuyrqr5at
uTCbiOZlKwpVaPyDuR/X0UaADKA9mk1kyFXAEIUZkxhkUwQYsbdm1N86TCjdmpus
kxchL2JS4M8mvLCd8CKdKjlak14RC4nsEMo3rjRmUY3qkWu7oXkvUgB+grHRowtH
q7KJHkuZ612Fy6vca4xocd7P0+dE362ATJaFgtgjLT7ZiGH835QBdpNUj81O0Rhk
I74C7ON/jnOAewdVRra6XqCMp2zxCvcI4iiw+FB1SSJz33HQj91hI5nJSZ7h5yAO
oECwBzZm8tT7PrxzDqcMAexgUy9P63evRpovdS8CueFtpORO3fYvzjV/TLRODwpG
yoAhizPj+GMSxqcIozuHTMLwQCI/EzF2cNRY236tpM1YlhhOWIuU+YP/UsnKdZO+
3EW5tRiIPYDLWOkjXoEKqWtr2DTi0RION9uLflDXz0o=
`protect END_PROTECTED
