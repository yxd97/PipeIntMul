`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlEhPv86cZAOF7PL84Q1ZSdHnoKQqOo6Ru5S1Jqq/0hIEiIgHtQeUJrqNj9w2zg2
rqhQjVNw36X6q161FoLy8NKWl3B8Tz6NfJfhs6/rdcoWT0hCQojs/W+ndQEWb1Wf
wmGmpdDIzJR0Zz7wjQWk9QfaWC/7Lg8S866nLDyOW1aDV54Wz5epWv10MpH6RoXx
1blEyxoKTnnMcvxx1/sV1jkQa78rdm15Njdne+uXF+1mKGIAf2YdwpUT2PGjk4Ep
6wybWwgGkvWjftXKsYc65gasVIq2cafYEDEzOM/as7x8aDEKTiqztJZr0xuYhY46
Z4F88GKm+QnJ5gUmnNcXZd4qaiJhUr96yw4PNP9T98se8f8i1aGflXIkLQRTdExn
XdqxMPn33QkJbmA/67WkB8XjJINunh7ocINMUxHZNstrGDHChrbEpJsNCtR00Ctz
HnM884X+C4gzxT+aaKNVwD35z4X7vkvyVAlLG6HWiSOH4IOtU7jGrqKuipkF7QD9
Gx7vpfYiRKgK9a6Ff8UegVNQHEp2CshtWLPz67ScCOFYfaANlxHizaYARppO13TC
xmTyWQXniDKFITKhRLjW7RspRnmGSkaXJM3TDWBTXTRjulsFBjN7ev/iFBUuoLb5
M7q1iqRvo+jUEFTK4qex3CAvUJQyqbLb/kzR32LqhS+64WQU1kHXPK2QFfApgOy6
BqZN6t3IBYtGq/yfc+LfARnvmYLew9v/NMAJYW5xgkxoa9hCUd2MmCLsbBJ/7rFu
qnZrYFUmTKM+AwEYLlsDY4KU1FYISM1AErkuNAjbZscDZrGHWKg/kX5QIq1fsYvs
P1BBJlBZNdEcKO60zatre1migyTYm6Tq3ldVROATnLw=
`protect END_PROTECTED
