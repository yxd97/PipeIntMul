`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkEOz1Zn7LXb6KJGAPGJv6vy1Y4TOzvCY+hUVUxpWIeTqRWt8NjC9LfbWOFAsjqK
VzUNHTzvJOq3R5vE6ioF9qOPv6Ct6rFSZJSsdetQ+MPXWtibyYqytPmFO4EuhzzF
60B7HaFHHb5GtG5fV7QFSJbZA2vL3rhT1XyrqSof1Nd76Kdgd8cQbMvohVfymyDr
AFVHYClTnfZy6eRZaCizKkD5ePFvSc9T/Z3I6Hay45aY4GIC3yMdmH+SUfQr4O/2
4dA5rJIPm/IvLV5unXA/TdwGzP6o7m7jm6lsuv6k+0YEbraVkmAYr+oSVpBV1oV4
O3HLfP8RW2FOR684ThzpRVvCZglRet7i0ChNIJ49yqCfOlSbp4ZY5VVlxeThExMu
+UdNBJVVIxB/TNa/e6U1iJbs/Nsi4ni04TAhm9vudSxeSHTqX9dW5IJMCKTEbbSl
jyI/gNz/vv2uRUCrr1Wbt5sBfrlxFgi+xpP02tJHe6ouMb1TqZ8tNOE4fWq+UsTP
jLEqEQljIZI6KBymAmdEf7uS8uxSW6sp74NMp1ZiZbppe6OkrXWFxN2CEgPpGRsq
uCn1g4Tpr2dVqwBxfhOLi23eXVdWpyYPVt4oLto/lC5fltv7YKfQInF7gMilsoZk
8OngyJy3SMYZzdZPUrf5Clttx+e83EfKYCYYSsO/N26e2Ft3TRPavkIu58oLc0e5
FexTSRifwjs52wkdXWLGUB8MpcmAmdi37Vz7Y7hzqtOyMv2hE4HL9MxEWWq15IUO
JJtlrI5dhYVXLO96fbld4Yv4DMTrrLoy9aTsfYYKBdz6fIfscveauTqFG/1Ojtbz
P0GF30FP5bzQjjcbRl9gyMzS44rwjXBua+1HcBRhc+KZQ2dUOKpzOfjQuBdphCFe
sDSm1hYVLPs/2klLVGyD4p+apHc+HG7O/gazyH7s7hKPgnhzCt3ul8SaC4GzBFLx
hWa0xZihmML17wo/BiIafsIF62hb7z+BQVYswKN7B5Zs3N5bt1pVe9w0C0aIxdNG
A7qYgN9aj/WII/yLIhJLBCne1Z0+c0CKQei0L6l+vLFQI4QAP0Pbo4eE4Zg0V8/v
SvKDO+8fAF6A3UuQqdggy9uPSA/gER+IcEm0NxTQQ1W/AKdYRsRFqkoM+QdzpEv9
TS8Hjx8B2GPe4KerHOZiePVuCiAv7Smph9J79qprxwGWblwyScomKENsUfTloYOo
Wi4I56v9cFVDHloyZyHn/vZK0HJwwPLVPG56oBcyk6D8q5xcwJunop3Lu8uSdDZR
LLNZrnybYarGgN+KqkuXjZMPAaJP/USnaDZqZ7Nk2C7Ru+jKdpvhdDxvV3ahT4Ej
P1WZ8S7oEyYAZhwp2qtT/rTvr7gT18V69IV+8wdTwDMZrdrx3t60MdkTm62FR0MB
ZGlzujGXjhdIAhC2HT3t5hl2E7bJ9P8kGmpRGHBZP7n1ZUuCnwbiVIDZ6NE9A4VH
05UQ9hWN09wDVBf/jxxSJnrRkUI2KxSbo2YIostvCSjRs+GW2UF8pADCfYXcdtPh
5Bp2emGnH8WK0WPEjlSy0//a3EyoRERA2kux0BZpYjtel+ksSNfIhhAyTwfwg0HJ
pH7z7a/drSppItzVN/kGW78Ky8CCiKAiA7C+DlMJoXEFAMTl7pSE1yV9T18dydRN
vru06/TyYMbo2flmq6DWNqVFgUYb2akTz9Tj4EyxjMnG48jFdWGp054qnQRMCCk1
hpmG1zpGIy6PvpnwlXoZi1FVlmRXcJOKcya9qBflWcsgxeqbSvVFg0dJXy1eQQIf
X4Y6cROo4mHUYEBQDtxZ7GpCefRE8aFVMkeDMosvKS1HPuZKatyRSmldnqtL3ZEK
ghXtwx+IQfQDmd0sP+FYkg68QD2lTx0MDswHaKQewOJ6CgTm3CuDRyHDNMwAYj6s
pFOZ7CVyQEaSQ5AsYYoEGSyFPSy+noCzSnClLCug0yyylgLR0bwcvL5HOUIGWHgc
JoAbvpwXCis/924rOMQk3PtvXMu0cP2DM+gW4yacSrNkDfZWT1G39dgBNfDTiVBn
R/wPZTkohjm1pOm+Wa+w/pmggIbF9i0LKTeA/Q0oh0mf2cBgwJZXQXZuLEMrLvht
5d4kOOOEHkhz5ieqGpSRfMmsuVgtCMi2KAJFIKXY1dnjO7oew1SQ12zEovZKotFp
OhSOg95wb3nTcEqAz8xudu7CPlj2GX/2N4OqgBlLsom4vhA9k7DjBeutKd+V7Ly8
biwzsb5BvwjcKYS1tCnmsGIOK/ydDBhXyFIRul+QBxobTJiM3b7FWjuva3uNAaea
EenDb4zb2m4BzpZ0JLQb2cH57M8q4lAj7qpWCd+KtdaGUPAqQ7HtqDjV4b6B9X3T
lHX8EWy+l3LSTYJdfo9p2d71TbxOpEC4wW/PT70eJOjTKECPjzXws15MeM6wk97e
WBVj2/J00Ky4D7O2c+qn85vjR3VQ1UQE4IqbJiDLQtC6HMC4UD9i04dHZEDWXOfF
RRX4O/tAecRcfAHg+ew+PGRp03yMYZEamvNeIuATk26krpJ8g+ZIobDCI2SrMfUb
oFrhqnIZayjHb8GVO0oruv+xxQ9BDxrkzeLMRbRBiVMGAWbTsK/5im0oD99Ew7eu
8FkH3d6TPq9NrCeS9Jh3SXGgW0tk4RaoIvLyyj3IJe9tjGlGlw1qMx1tus6g7moo
qn+nEx6VneXfY7djD+sZdF/eVPoBJM2VbbjphYMs0IOxev0TPRv/JiMSx5RnGnvo
GAbNhqVbdsbEXEz0u/aiqsGGQvtkqLuBGcPp55Y8LCBfGOMJpAdgEkHzVT7TcQP0
xHytK4dGA/olY4Q2X4sMPpPnyD2z6+RVHhndip78Vawpor+vvilhKHOVa5Ze4tqD
`protect END_PROTECTED
