`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FWOw4vH/agGSe7+OaWvz7/hF9y1QAxPm3svO3HxG1qTZLr0551dmXykQ/Au/IMRh
b52xRMuS9qiqMIL70U5OwlGzjYhkY8wDx0mtd9aki5lY3b7BN3O6uUMZcVR2pSBt
k+lKSUXnJueyRZ92+/96rSW+JdWu3P5hogMzqRvSB78or0vUPAo2+RsRsnu0NDMs
xzHoC/VGlDB7gX160Swb4odlvfbJn1a144ihhMKa5OYOPA28oXSkU0FpZSIqgT97
AHncDeqNix5r0TBHY1SXmyD1QpKdVmJ5gDjeDO4tl9H431Qu7k1JIxefSsh8ZfG+
PgYs4i1mpmZOIde7OI7kCrHwIEd5vg1XCJA2fyFOQ9tuTEUEwJwxsuk+XX/9fALt
+NyOs7YE7n2HFGts6v4E3Qgshytnax5s4erOSDWu+zZvBoUbYzE6NbeAnVJD6OTt
kHgf4xriNDwJ+re/eeiyGMltnj+6vT9LEIZFDMm4iDT4oKTkExhB2cZVJseq1DIT
RLvf/L7XgCCUwo7pD7dNXrtG17LF9Z03kyrIJheqx0bougLcYx971uM4iv6nKUgj
XLIMFJrnVofF2X++BqtYmyKJigh/zSW3YE43uEx/HZ64KyXRx8MvdFO2ZZ3tKXSE
kTzDyxHmXYB8SSK43R4VKA==
`protect END_PROTECTED
