`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+38eHTfVdBz9I21lwj1ZdgO1+9ulbYHYrouhMzdIBQJ/PBe+/bsZKxI+QsLigTIa
E8OlwG0xoxubKav62E8peInPVxijhDs0m2wH0X9TAdN3XN7zWONUEgaF5S4lrpa0
qpRiXY3oO3pSqNl7/n3RBE5cobGrGAjmcY0vEJ/OvmKMtInOJU09dSJq8r544Akq
UtvA9uv0W+3JsndYR10gSaVL2/N1JwheQSa/E0o9eNmDn6AOZvxQovgc+xbV7xl6
WZGDQFxNpHFDZrcF2vUWHsXTC985JNBnNAhSGeCkNMd+E5VWERYPtde36gOapGKB
c4RqnCS92vDXsI4RduDqqhgTG7kBoWD4oN2PHEeP9WersNVeaQ09Uw2f0RkkhK28
utYpRhTBZDtKNCpLG2oxqkTvjUqujnTVOt79dAyltGzVQeI7nqlcgqGm+Hi2FCQH
U/crk6C2xA6cIWA13D7a08x89icKlw476Z4Ycrs6gS8/YWVM51ybq17vD1P4JvBS
j8ENjB/S78aPEQtRZ3Sq+NY1vXg3lnuY9DXUhL+zSpoa3D7mgxuKhaCEdrEDxlJ1
/vf5CWvA80tlDWOp/BdI2VvvzQQai/HR4gsooeW6mJIpjMryk5JDqTawijbImrki
L9KKUmBJViqS/6NP7kBkAw==
`protect END_PROTECTED
