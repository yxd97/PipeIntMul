`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5GGopGsSHhfP06aGbHVACrUndf5e9HKgvo+Ou7qpZTmtmDvcJCNoUjayf+niSCM
Pgd3WMLn4PkBBwKnR9ST0+nrZe3h7yfVy8RKSBRr1s21cz5yIQzrwulrGAQSXhJK
46bwTqKK4/u35BsW09McvWpflySDlY8DGh/lBupTkZrpCPAhz2r3XStegC4jgwRN
Q9OgmbjeyvWKDAENjQKox5Re7xh3gMEko2z3x/WVZGGGLGZYHT/xA24ejXUp3isW
l6DRIYMyMMPbSXk0rDMguH4+GZQLILGonxsySe/f141doXeg4kxTjHAsRC9+RFc9
l2T/4DGmRKyK6CMoJbo3B5IhFOZacN6g2Efv7cyxMKkb4mLChAR6KMzyNd/rc0TJ
Du8qOyOeLQIXzay/ea5L+qd/JwYHSC5gGsfT/kyeQ7IDA7lqsfDfAH5Tqt0WpsYi
+9NQAurzZPG+GGeZKqco3UY+ttxG35JEmaQbW+jRjoum/ezkKTO03sdqREDxmZ2S
lNeyKn2oUJUaGZraT3SlS4Jl/5AsisAFV8r9Yy3oA4zqRMFhefPXSUDMdNVWr86P
5BSgfY+IV/zrnLSdrqWh/gGEHhgSeqFv6gyzUjoR2VlRifGiel/QfUR/68EZaLSv
QvU4RGcILEZrx5qOFmmUnzXtXhVgvg58j7ft++fYihnKL5Zo8rBPyiDrCfldh/z7
LREm0pDm53glxsV+VX/oMw==
`protect END_PROTECTED
