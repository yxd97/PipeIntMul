`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P6QlmW0rUiJWG7JEjTTjLAhgzZGU85MtFJnAM+QWKAyjkajfaMuqvaZjxKF+Qyfj
6eTlGIrdfn/pH0sRGs+22LGv3ScN7n56xopL5Ph+O/bQjLeDaOqRttbFT3NGkY5p
Y/LX3rclSKt4vttSycVTmZe5aZJdc1Om1YgHunE7vVcgK2nc7sAdA4U9C7eL0IYm
rWJGhWo2OCxLOrwowu3gToYEy/FqhkMaZtauBaq73VCByonmP0xRFmYJmvnezN9F
oZjilyCm0t0G/cIvIUoiAQXHS9clz18JoFFHRREIEMjHexl5uY6VdrNM7Yyvop2M
5iG/reVOTPvjS3QVdZ3EqueXliGHBzeAohbYkgu1iJFQg6gSP02kC3C7DkU2n8PW
vyfIiymmKAh7ODNv66Tt4rwZk5JZjoOzXXoVwg2+ObiBERuL0W8ZFxUSKi39dz5T
O6j4n1QHqJ6541koYcI6k+c1d1vX1fzlpjD1IwAq8GTqnT+I0Nr6dSZitKH9mZGp
3mi0kRbkiYjAFfJXxveunXL66ExU+71KwEWpsuAuSf3Ves7gfu4R0GkUCjfGK6JN
cjSBjXgiTFqiV13T3JmXNMNoTt9K8Zv74B6fkY3eajh3BpvMvsEoQKfYDa7mnlyR
PDWwwlhYHcW7WTN9QiQVMDEA4XfaI0oia8Uprxqd2ycRm1ZDlLePATlBXj4iVqgT
rAzfKn6c0kXcRREZgOXcyD6qJEqTAhgNGQa6dbe7AB2NrNQw8J1pCBRLxzG9Gq7x
iFWNQijCdh4pzt1HYrO8Gicc7cyUXG0nZfmeflmtd4D0uL5SF8/Dp/GljiwgAHsI
k3I1Fp9li51yHoQFYCrT+sXjFPpFyH4rxb+ziw3Kyb1pakavTiDhejVGXtRcdTcV
13jv/0LS/pVNtxshrTGkhT+QpsrZi+Q8kizKEYFKN3VCmhmpI0m4jYVW1ynPYLkp
jiT3ZYR1g8cO02cTNbimDafuhCkNY2QRZqP00SDlcKUFyhRet4s1AcYmIZfhMvTP
cewZA6H36xblFfRcj0QVOfeREmmqFS2s+VNMap21L7myse4Gj09pLLoRZxLDlQIs
FjK6vsmMitcRRTUQFKrWEoDmdPNBFMU2f+Ix/1DMSVHAnD5mMHoRo4qSNIx1qIP1
PdHvfXx0om+Dx3UZoggiNC3vZXXmIvYLEQ2NFfiXUJm/iwZX1xzV/dy2RPoQqk/U
qr8QVsKoeyQKTLpv0cxBxVDgM+28Wk8HG4hMQYaUlA5pSdBu+t47yUYzULuJB+Z1
ouXQXuGyYxL/MUZAiFP7rhVOyo7CDbXDzvDOyh/v0pv4G/3PRJ9y9r9sGwUxSlOG
H/HP9sPCJ6oW2KDHIXlgn20J3LdkbW/FuawObgkf4mmujzvcCN7m8ZFTe7vPsDyK
JyrcvT0EO/No4YXa6+6XwwULohhE7yROoGL52o5dKU2ZdCd3JalEqM2qouz8OVQb
9J/+dQS9SqiCqpVjjPKajF3dTlr7jTfdblZfTNzhwxx1raRAQ4tfzS2PvbAOyPNW
OA3Yx5ram7NheRXT/StOVUiUn9yVziPYkYEYwTre9OT6L/jIbMKf4Gr6xFmzpPVh
F+5rUZTaEmzQWXclL5p0u5We71zcoW3neyu7FxTt1J5hzR0vqGXwza7PD+qvZDzh
dbnHCZtRJOTr7f4FQkXINeCVhX0KctnJg2gQ1vZtmGu6keF9jwA0xn28OwhTQEQ4
GzLTMNTuTMtEDvUzRS1GqY/UFHOeY/wq5A09R+vXO5AHRWFdntmuaTlGl2er/+78
X3QOfj9F2IQySAECrAHt2hs0azNRGuWHTAiXvaw93IftakSDEBsQ5Q8HCtCcR/Ch
qlH2fB16+GVCT5zaRyeSIoqLDRrBbXeAmMIWspkGOGw3AQ8sWgQA52VHPkRizr/p
Nq0D7K0ktrbzBDHFFpvBvi8xX5GB7iAalnbf9w2tma/o5VnLuAlMgx3bJeFHmD2w
WN5L5/SeQAN0h+XDr1Ylo5ncBB/NWBCByzDn0BIjw3KR2qUwwxs3JG3mxTZ80k3K
pIsr2ONNcUw6Dv1qoxH90E07DL4/WJ2kRNkoHYxD9nwKMq6XaT6nMIWjvdrDHcF3
xnoapaMQXrbEB6FuHhRSNkyEY/LatVAPqZHVewL+pEF35TWmvxsoP4DwXPIypy8j
UCQJZSW6Efvlu+ccrbpVpNNHAvuXV1qkPbFbSs8fd3+7YfPtfsYtnm4b1/kJfRwa
lPiuLpQrmBN8MY4cXVFV5AXnAR74u+4lXJzjZ1kJpKWq/hjSNxA/7czbmY8sMq9l
sqNlwiyKr94ISOHwnCoA8213/3SFNajhdEWutevH0tRgNEIsgL227xK0sjoT3Mgi
O0OhLXxtW9n6fLB0x7cKhBsHvlmlLzJ5M8NCT27BLmWTEvukcTwaCApNBY7Zx0N7
7yCRFyk+uVwcKDk1esoFvER8kLeejOrmf6OsPyeI6EeYe0ytslmCY4PMHs6GiAYj
6f4NbK+kDvw3vIF2GYIY+Yun4Nav6ec7uYAASJAPW4lWUNkvxXELldILacercWU7
s7/YOVrEAD5qif5ZmuqBiHlKVs5kEVFFSovt+Bk2Tz57iw24vrFryvp3Y1njPnX7
/wsBpHnjVLAbGRBrwbRCI/Q06WHJ0cNc3xYuDW0h8zyyrFfmT22CrJ7tGFAEKzpj
/FNWm88Q4pCNsp9b3YB4MoVW7y446J5DiGoGlxEYLjpeYPCFSOKXa/rM/RSejRxT
I92mrOWVf31M2OjPcj4oKYCrdij3u32O6tdtNmDIU7JVQHWYGYFnd7sc2Oqb6zrY
kEp9agzrcXyuLivCyQPIRWD1kJBlsTzSyX7gk6L52fMyfeI6qBiAJ6MdVriEp33w
4OSR7FPTg27+5PeAttw+IHnFmqBGgP5YbDMxBDMBoGqX39HfW7P31UgkgblCMPi6
IfbIHGjhRfBa/GuW51IcAXYwkI/yngwazWX1+ZO5nLqeib51BjfbeXqAq7ImLqs9
iI10OvC0Oe6CyVm8m6NMTomixAlrqjlXws319mT1FarhEttQEDAbUAQTKMc5FZss
rJ4JSaM8hsSzHYbaEYLCe+MJ0SUsQlT+fxDgoCYfLmtDPI0pFylftnNOTENISxTb
bjfevebFq0bZ7+An3q4XNgr2BrDiG3sYazfQZ7aJSKcF5QxLSYqJ14K+HVDvmpO5
bzwth2NdZQRp5QesivbFwCdzDB86B00KhOvM8Myru9C1QU3DaOCZnZzoZ/0Gnnp7
aASaaTjLRdDIiqwPyiTKfmc3+rZQNpsNmypFxgHcQnLc5vwcP5s3LC22uVrqSxUL
Ummp16GgzIoZ9djtQJvKdgvV59vt4OJIMTQz61ZtZfHwZt5logOgm5lW8LYYSmuk
oWRm1Z985imsysADzqobDRkJ/tgcrp1el68beahRjmW7q1+earNLArCSG/WP0ZAL
J+2iJ6y+TuEsd8+xvP8p8Mn4JB1rQx2qeZMgAQsuZQK5185SaC4UFNHfdUFGmdmG
BBjqV2cDHeZreWbD5dtQAjEZRqvy5h3it9JxJoCTJmT1p04Rmz9Q9nGqZf9QRF1x
3t8/QlIVkNlcdn+7TUD90KHhsZEpiW5GtWZHF+zM4hvT7C11ZAj+x6TjZBfcESuK
7jE5mqeVRHTqP/2mOD5FMFHKOZmdsqCX9AyZ5kyYKyPfPlBdEVQsngtdMuKX2i79
WVssA24gV4KOs0o8A5gjDgvv/xPZxmTtcp4AUF9F3Cc1wjVt+LsWmn04z5NMcwWQ
GzCrlxxqwa5mMC1V0zsiY/eMa2tjFb9OhwkEfdX1IDrkmzsQIt/1OOOZcqKfKSqV
THk25LxhxynIb+5VX/IV1nfkPrxo8LZMaj7pMmrbrp+5tveCeDl4g4Ru1ISTPQB5
m7YDTgyXKr8xGitckPxMP32k3lJBVejLWC5R05fqx3vykLTTlyMRUzVx9PE6QOyI
JWkTm4YzrT6CSvwXlKzs9dPgMI5C6irRJYqeb1wIaLpZIoa3pHtSmix1ellMh/AL
JqQpDSHf/O4i3jSkPJ8XIIxULnItinS8B3AWPOPwYAjP3JQXQ+YFxf7dD/vwfCPo
NB12BhYLkLIymAdSuWuqBjl1rplaKxBYDszgAekmJTVxJL5bTWeIFT/cO61k4ts7
SmkNrtT4guIb+OyMuGBZzllkP6L8WPb6SKbOgcKEcIs9Lu6UqUcIsLfMn1ez90Vr
G/xcVB4YUn/GSkH5N1vDkgS0jLRVVlLDd1A8jfPlbSdHEIvgN2Qq+cJ/C/Ddn7zd
44TO/okgRDArEoiOJ0gjw4S/+ZomPhax9Wre5M9mtC7txLDXkCD/ENKesBftrtaq
kFel8STEye6bNyydbp11AkIvgqH0uji/rK9Us8lWfhoOzHiaTxlppVBwXY6J05RA
uPwueF9j7/IYi9wJLIO68kJXxM7LVXxaeN6pVAYeZYu2Ax6IQ1C+5PTS4/tizuS4
uTftXnQvco4sLSYF4QL2mpPheKn6m19NlPmJcCswxJDEk24AJtfbLLIKfPbM3JUj
sF02ep2A5ZVH8w8r9f9Cq/gicuO4DAEs05RYtNm3dvGnUVf3nfRpA96bKFUf2qbY
BEcZTdEkyKTVnhHPqyvLml3XYZJMqTXEw3MnV5gHj7VZJd0wKJzP7mQK2NpQHVg0
xpi3zTIgDe+OtWYcq8MOjBvsZrAEt7UMk25/IdzB5SlRD8iFemMJgMeTAVLO7qbO
eJNaTIsKsMTynbsgWIYneOIQfwIfIBI8cZ7XXZHLwqXX6C8NP7iL3/7YG9SK7pzW
RExRNIrOWertDNCXCTFVwh/Y5la+RTBaY2VYCWY0KL8KopVZfOC7svHZiLZcgG1W
ioPSrS3OWfIlYXVE0aP20FAcX2ilqDNuZHfkSvjFc3Wuc+PHMVWqlfagA3QjkkSv
i7VXT+zPifE5fNF4VVISLu7eovMgip86/2XfvhhpezG5MZaEs9u87BJTWOSLRp3y
6tE4E+V1H02mcodA8lyZ0Sm1t0k48ZRclsUMDD60CesR5Hnzk3jeG7+NgdCre7t1
muxWB3WzPF16CLpmpYCSpl8ib09E9OqJJFWGh90Pl2IvsuQ1WWLrl5J4K8aQebAq
XVjTbReYKpGO40ko/wQd14xosOsG7L37752gjn3i30u56S+xsADyvqksbUIpXzZP
CV1z1xkobLWk6zknW+fR1IhWxf6Q0BPYDxIHo/0nTH9aDdPPVFeaDFNfUDYFLHOg
fdmZEa0yVX9vuYn+mbkAm4Jo27dvjfh46W9cBUX8WdJ6mYWZfLXuIgMxqvfHfqsS
ydHv+cmjWYjsYXm2hv3Y66dR6tW2W/HrtK+XWh95YC7a2fkPfdNY5/QF4huIA5gs
f6WELIG/VW/yFJAtoFKF0WZtc8nC4ix8B1z+cyf4xwv6cUvAm42qsWItgKdW070S
Xv3PJyTbl2GEJXHl/dYT2vaNNIpORjaE25Cip3N5fSTLK5zRh2lnP5Xygp/4vWgw
gtPCZuOGlgRR1+hOVrBgKQSZ/26Ce3OctclHRH45HYupVsmvskZfsljpqz47NfGy
Wf9k/8FWI3na7j5Tl7rqLZZ5Dv2IlGSAfmpPePwQATdVicR6GgYqmihLiYSRhht2
KUUX3VGTzGMynWrWJ2A3bWxeD8QYSyENgAq4QhlNtJLJI6OyBykK+iWAlyrfRiJU
ULAlO0JdjSk/ztCQikxaKx8coIlP4ijUjPu+OIrH2+i4niHwePBqhWrB3fzqSmtV
bXP2DLj0exdP2pxFJIvjUSc5OpZeJ8aPgQ1QopWjwAVgNUG+eZROG6KgmSPSVaED
yHqvZJk8w5Mc+quwm+cXkC2TomUoYisAG3KeZZoDiJKSSVBQv2HFZMW/gIdK9PVD
0k0e2Vdqp/xhnR/ODA4Ppse1Em29GItlJc9i2K1TOI5PhMSQqucohv4TNuq6qafQ
8Sy9lCVcFP+Q0ru9mGxegBjtukYmrQMrkilEs16SindOVbHtL/weofhDfBbeI1jp
liUdNE53msWor+3u0WWytdk/GW1nZugkOvPvXWHMI2CI0xh9L28OtTSHEpfcAMoU
Q71959yNPWFTDeL7xGCgny5OicgD8rh8hoWDVOotGnno6e7LY55GyPrTGMe4Q9Zg
`protect END_PROTECTED
