`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sw44YLyB+/ygzw8zFfNulrim749CeJtX40jsSNTIc8BnoPNfqkh9/0XmO9g59nXL
9seafX9DKtOXum+j59li+HKMpeQ94JlVKOs8Uaav0LzZQ8CLHJ0C7aU/tSGeYvvw
KrBUKeBE7Qb2dPmLaqS2AeIHnAkSNLBT1xDZujlwhKFT9wjresF3JtVMuDmv1+pN
BsWjIxa2DVO289jgGQ2j8l1deY7GjS6gAyWGBYkHCZ+n7I9szOyLdaRPutycXjn6
DLJc8kEO9h6FAntZGrAIT4fie1o4seDXfkStcNNnuksaIMzsfX5A67bHY1gUYUJB
BmlkO4iHhivcYx4VZzohnbIwAIwHc+XD5N+GlicCH8IuDjeETFVYX+oJJ6853Qou
k9LnFhhKYhsQaHihPf+94PUSAK1TxUDbfWCv1t4Ihee+RVhn1CDswwy/Cz2L/AGg
dUBa7Htsmi3UcwcYWrWveAd7/kOwzVu2g4rx2qRQUgVnyijkyr5ccB1nffwTfIHt
YWnU2EuXFxhkVFoRwPR7+e17IEYe+tAKE81QwDFmNSHOrh705s0pov27u1hdTttZ
vj4G2coL+7pJ4qhF/OCE3psPA8lsb4F1COF2xOwk0yjamELEwXCUl3C+hspRigab
B1n7vzGYdxK5cexxYyuLVG90uHxyGuFO1DDw2mTHwY/vMHCahWTWATIUPcVO3o5/
lU/EVoIZBV5vYWJSt8tek3DqNO1KMBW84eMk7kR9Q56mCbvt9eALCtjjiVebAt21
zogLxxKW6wWmraV7dJApp7kmrt0biReyQnuJFDdCJioyIyGNpz6iwtzkVYqvfR7U
YfNW0zu6T5FB+D1sZZIgh6aaFsVVBPez+RHL/F6il+CtZ03FWhctVlkOg4sEnmIT
pB+pn9x8/WrLXbLhPBbt9p1xQnt5UR/3PxWgieR+kh4KgigDpsUQ9CwaF8NM+4I7
EagoJJkXs8CdIpALtIbkR4f7jxdUzGOI66NeVz5vNbR/DucxUdAYxpC6WQV/iLWE
J9nz0FofOdrqdjMeRb8wSFgjh/NTQ+jVpLjik2TWfDx3kdIPLbFzAmBG1eeFA4yn
13h0ze4LK7odH8aJSbFhmPH2y3l2bkW9fiI3HX+RpmQiMcrBmhzcEXqxNnlqMFOw
XgcD4x5MkSZeiGS9Pws9U/wJeh6/Ss9mhzeZPnUIXTqKxtTMz80MiYTPyk9yTnDm
y2Kvb+ZuZbQ9yVQLfNVMzakucYao7Lt2H/7pijrtNb+FsnpTdtXeLn803M1t0Dw6
qAizZgB6BEa3rM7ZmZpi0jUubyTC1XkheO0EiOyHw2f2o8UpyetCmV1ih76dmGyd
7htea0VPpG830oxE8UU+yW9z4nIbPipMd/VeugQj9rRa8IJ13aqBw9D/gQoOv2wY
N4t9yK6toKcrbo076W6GmLkyLJIvwM5Ag8fHFfMsAU+DJ2zqQshSTrfUzxFCtH3U
mF1QgFhw4+dZo3K0Bje1sXp1SNTy1NvJ2wX8taxrLg7kLgZBTS9torVPQtUcGcSh
3DDX9+1y+WrGMI6xRfvOAXyeabyMkx1FrDd8iG9YkUUNePmvPwIez+oKdIw49S0Y
ENpWOfJENeHBPDRAN6lbjJApumcWrmqgwBd07fkcZ1OVvN1HJlGDrnQ0fZWYIPAK
8Qbvt7lA/HJKyIDN6KZhu+KK7cKOf5wbk0vPFIfxHnY4C0BKaLnm0y9kd+LqUkf3
sWdlypyvrVXZhZqn4Z9mypmOxNBS/2pIDJ5cNuw6nHMA0HYwEq9ZcE3kD110Lmes
PUJLbXObP4H3YxtRBfDf54i78KyGYk//tUH4vyLmbCzjYhafDFShMY8h4ZG0dcL/
zL54jRTNedM2HI83dayfUEX6IBrT3iFiZi0cmg7hw0UG4wtjOXxVEqH0+tmKdT+F
k01Y3w5kh8D24kaNeAGgw3D3+Ih4vQVC50QKXifCq+R8Cp2Q8rRyp30iDOyXPAh4
EyN8LBL9Q3B/W8yvIK+cguRYwVpKCXW7NGl/A0U55Pl5zWL/8NbM/X7fOw9O6bKX
gHUyIn5/WGfkw4EAu1wDjDmQ4V9jqRDePvkrqugRMtJvxvvfpftWUvLu1zxcKrNG
eyOOFkXcRJXzrC2PVdI5UJ23pQ5EdaizKX1SAPfQiY5l4EPOrwn1vNTUY+DUwKC2
rf+fMj+IF3ApdRIC5X0wmCXGFmuw5sb3t50ZV0p/7WP17VvaEczMC+IU4QpXl4AC
5LyOgMW26NFvuyp9b/Vgo+gp1wJsyJcq0isoUPEFKDJhAoRA5ZWK0RDGJpQ7M41i
7TTcixux5loXyWNxdCl440Tk7yYBp9jMg5U5fb8CE6u7aM29yl6Wtal1mgNtgmO1
roUFYZCuVg/AfnXrH64n745UYIWGgO50Gq+wyHdRUEHzvWTcUpJO/IHujVeeBUCI
rutiYHNhsdCfdvi9PnBCyAVo8yt/RFxaCLDcfJ1ZTqsTcpQJfcLCbIx30kElNoV8
YKhsYEXs0qcA/cqDAfQCpip1KrR5sKfY2vftuhVoiy2BH5aMZdCTcurvlWQAPM7o
18iLn4scxfD1utpiqIpGaycbmQLaaoTjn8jFO0dxmz0=
`protect END_PROTECTED
