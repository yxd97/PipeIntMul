`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOOuHo9OtBG7Si7qNlu4YI+rtnObJgIsakGC3T/9gNFXl9u113g2e/S6ACRoKBKV
nao6+LXxm26yj/8sPYuMSwXmq+otIVl1SWSaFsErBkgxOy6/pcBPWgonnGvdF796
8iAu1Fd++dkqPHTv6DPaLaCxWOnP1otBkafLMZLKybzihOFFmMslZQd5tz0UP799
ygRG1614yHKEuLHvyZYQHVTkEHINfKxp5w1dB4G03DyVGvpjwz4wLkALKc5myL5w
qub8BAy5kRaPkFz+CJ5BLor0ixjRTDaXSxY6krd2+eAV8OiHDxS3yknymywhdrBZ
`protect END_PROTECTED
