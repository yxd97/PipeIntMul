`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zzl1hH83yorcg5T2rMtvG1PmtuANHnnsNyg8NoQ+F9S6scQI6vVWtVEBgLsHsN77
QLkiRaXsNDMYYMveXQJDhYGoQ9T9WDiehxD+Hxn0sg7BMnYexI5IWetbpp5OV/21
kgoTCKDYygsR3Ob2lhOo5QtogI31xvOVlV4D73Smkqmu058vZU5rEr3qShcyMCYd
S06e1lklZSw/j6EOgE0do8CNOZwzUUYNpY69HgwzHShdKwDCfoFRZ73sO8TjqaT1
Xvn2Zx2ZUoNFEU79VDzVAx0GCUfEr9UKJDa3aCts41tfjfnlibw5X0lFAvkgLQ2G
uQ5a7p+OSoxfW81qFJJnricsQk0HoVJWWQ3R2BPLaLwJz0a3UT7rIMMQze/BXWAt
EIpsSRZPZ9/T0ZKcwb3tVvobXKcQHyzio+X+6kLDYeEmPLsFTWmzqWMwF8s5UcrM
BHhbm80obnpeJ5Upac0+0VRB2P0P22CryLlKCLRWzX56SRE4FNIAqu2AviNrtDI0
iylFQ4ONUSCgtnw1mxSmbIAZdcghBjFSZxT9T0TJlvo0WDPr5URa4pvrBJ7TEDWa
`protect END_PROTECTED
