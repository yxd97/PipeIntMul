`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3g6wHLLfM1gCvP1OEnTIKOT5PGMa4O/iP1cqK7uvyItHgN6mpIoC8AP+BSiBTND
FI8fbR6WhQZhhKJfJc5xswYAVNZ9iLQgcMnFfLFkOCHSGPDjmctGlHVmBRRXwU3I
RKq5i+aAR7Xa26ER5udukRq6hPm3o4dFrSMACe97n9jbZJnhifNft9AyeTWI1x6L
ZYuvq/11X4kq7Y8ZFEI0nvLBz7Hm5/ZLtdz1AjKvuR5Ov6gn1cgBPV7W8y6yomW9
Ehn7YK8pNLBLBmg6AKy5Mx5K8/RBmFqRn3trpDeHRoa8ih6hNq4H33JokmrwJ9RU
ZLLUNTL00Z4giYTECb5nwARIB7j9mLM1uC2z+y7Nge5Ob55NqOn2tBCLjjD06VBp
yhC2qk00vR2f+2jdEdtkKE7QlZTfBKZeEM/JdPN3MMc3Yp3AGZtRheaKzEQ0nwiz
VMid3A28/Bhgokto0KvzybrH1QulY+P6Jig5IWKoerZ+tBF1L3ST0WuoSjxi2sLu
05vUniZGSzvN2qigXWv2FIhHoyQaOR26WTHJnQHdJzitTnZHbhIxiSrrFT17agne
XMJwOxBgsrGrlMCWon6K89gP4phaZKMecDgz8X33FxKPasJCDqYKJie2g4kyieMI
Fo09VCgNxpXUs21ij7Bu/8MmNQ+z6A0gtwUYLTrd0LT3cli/GeWolOpPngdLWCdc
5PWf5KD4N+8zltyFYKk+0Q==
`protect END_PROTECTED
