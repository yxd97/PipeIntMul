`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VgjqiFl6eoQNhCVaK+3UkPklyy57fjf2K4/I2ezcDczRUqiY/DPW/NvbmIaDxBjf
xY1OVoL4xuDGPIp00slb6z+NiJGnJfPsIH06R1YADV1wuJovyQbLcJtcJw4HGbsp
bPTbrweTf8TBm5Mh0huTHmNUl6a0ddSHPRzKpZQTjsMqLiKb6+duZqSRop+3vNgx
FuBaoFswWOq42KXiY6ZYQx9qSmt4ljdmipeSRyWXu8hETi++sB75WEfCpRNo7C/k
yBK+JbYhhVAq6nmqtMwcxYfYaeHzHWPPANZEhn46xllMW3TtldVkli9enRSYBehM
SjXF4+awxtBqiP4rVpVMFvW1v/oqlwBuljWVRYKN23e1T8uVytiF6r+4RjwhsXR/
O4djBmxU7cbgfTRXQYi5XQ==
`protect END_PROTECTED
