`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mAEZ16eI8Rene8fMssCWhQUilqO7eA7sz6C4VZfWzxSEODIx2u38Otjd2BjqmAj
UOZA+7N+G4OfyS5ey+BiCA0RceBjJxfQQ5GFaG6XBIgRNbDCl11vc6XKOYT8xzpA
MatsThwLzPRF3cC2/xepykSCu25h1E58pkfTpKbWYnBZ28r9xM9frb8ZK9eomZbe
qpQuQ0Y1bhT4ZAt6WW95LkXZhLjnGSSZ2coXs0JqmZML6S4DgliPjyoLMjL7yyfg
vO2UWPiGA3dWXoiDqHGIBcXVyanV05UNiNIlehKZ9vXSANIRR9Xhkd1GEeM9ue0S
P/6LOYd0oPISVGiO2dVxfpag9iuID09OOK3p4NDElP+oNXF4id5nQV7PYz32pj7A
SW2EjFpUl7jYQSQvHJ0SakV7A0yvK6PU5wDa0kZ33tbf5SNKxrqkHQG8KsSm8S9A
r8LirUXuHGycDK8EGiCQHMf9zPDEqoiTeOcV0gDqfqWNmrQ28/EAJMwlG5aN/u9A
M71PKZKLvZMVjiIuuEB4Q9XAUWxdEiQfGegkRw0kxjauCkcOLA3AgHT/7izdG06A
g5+92pIgM+bcZGCQAd4wxMg5Cr0HnmaDd8YmZbdsdaNKF1bb9HpQggS35jTZJpDn
d5IdQ88CZDYJq/1zPcZ0TA3NaKBU0ZojxKcsIZ9fN3UD6Ljlt2qnZM7+Bhx4vI4o
d4hoaXHyutd85caXrolHGVmxnFEYfIaKoqkaMu9Dn/ZJ8mCLc9xVykm1g2UWh4cs
XoSllJNNhyILz0Rn3vYQR84FFd597E9+7sA2xAkM/zjgATp6dSDsPuW6cnQiqGTN
CzfHjEfq7DSO1G+Cp0mDbRGd/OQzXn55YDEenIt01vVexwSiZymy1mIubd5GcVsl
/mK9fn835NUw/UQIdt1kARTj8a8QcTTBrxBYwHoIqahRFKJALtmGZSZpqPIjiC3R
h7ByexCWW4eNqSz7UtKYbme41qtvbdp04NjfPAyZF/tiq3C3siJMMQWHv4ITqksx
HTPH3BNOGwHaSvMElZTx1abq7l6eugF2Gry9DKJysg/WsaGfF+lmsehpuoOT4eyD
9OqOxA7TIuFfgfJ5wX6fJAWlr/LGh/aywm35wFS9EmVbHukBhbFHCamQan+fW8KK
RZn1dc2pco4E0ls/qS5IEsJAkvPHnlkgDIZjjp5vv4EJrttdOlu6FgAKfbTaDh0+
rGA2b/4LY1Z+AsRLNf2UC67O0a/Jn+KWMZCTtDW1fIxrk2mbJYYiFdBiSGgULL2R
wdkReZ+tJp3AM4uH4nSKftHZ8uAcmcqV+OiGvQJZhbWro/PBwn1noPzTcGIbvWJB
jZWU4nP3P9SEfue+M6GlgtR09NJn/lJAb/xvBZL2JTH40XahFAngu4LKMly1DnRT
2539/d4TNSsK5Wx6wkMMWAUqp1T2RPTkxSjXB2Lv6gzRJcx5z6Tsx0IuJjZxUFJZ
vHb9+IGmIfhVYw5tmgw+SSSjAZokE5PbuRAFPMmVrg/48MS6lfCSH75Mv1hhmZnR
1AJnklurdxMhr8IRVoMQx5zricHdq30BTDg1Ck/xbKgcU3PnKFHXWZkgPVUP09Og
OAxw+pdRRfdtpTlh50TZujh2g7sEK5ZH+j/nnD8AOODIiGy7KiVWFMkKKxB4gMnF
1A4m1eJJv9ATwrwah/9kS4GKTM2GSovSEt25u63+3kXcwTIu4RZjqWPhgSlVdoxC
tPiiNE1lB4QtYA4I42A0H0FCTww22P8I4fuh2BsuPZmpIbaXvkjjDWO9JXaqYu8h
ZFFKXTRzadOWT7DSAj5ILcjaH5fzBnCUQTKR1yTcKe63l3zWIjeX/2hhiEsWuX22
XXyi41hn71RaCbWa+Kp7K9Rt1n7Xhx5vh00J23brFLjQEhD8UDaQ8q05WLHMSMfK
EUt3ksUGuHHy0ZRT4H/tPVOTmBsJaatiAgeiDJuquGrq39f2S7mBGj+7sVg3nQMj
oPZhaqTd5emfRSJAid0RRbaZeECy2xAY/lZriv23/8q51VeQIgVr8d55YDbYAz1A
OwvMK5fMyNy8h247ofc+bghfex83o2SE07zJ9seI0R0vOKPAotMvwpzRI/D46QAm
jkbB6ksNt1T5WxU1LuX8WQ==
`protect END_PROTECTED
