`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Co+Kd9NNfDwenQfhj+yyCDhOuyVQPiBMP9AHkijhm4JCMdns0E8H6LsB4klNXA5W
nV5On4j/ZJAJmQ8DgAaxGfd8OjXbS7wnZQL/KjffO2XqyL6foB196GGAxQgeH712
OzORkVoq1AtsUmaFItJl6Cjaozqrb07uEUM1AVFGIHkFQYBob8Ra+PpGHl5/cP2I
aZnBr0o4i5OecwHW19hmNgdEwUNTV/2hThueM7fXeBAYaCFklVDRFj3p0U3eSYFH
FatCNuD3FIbVJ2PXmEQRWNInoVbI/ur4ibA0WyZpeuiMLlgSFMP1OD0pUWv3a2oL
6ZA7jML4dFoez2igqDBujGMnKsST/QNfQOXJYgCSJT6ATv+2z5RfrD7j5HNI+y/9
4EDUpLQM1Tg4Ol59tkVy3YJVrJ/JnDNgo0u0HumWZiMwhtjYbWDMzNhFoc4bwrvp
r9//mZCViAeOPO452XTh1qu4kQy67J5MwcVWmtfxRvxMFbt4wsbBSMJ0szvSTH6f
BiLb0XJOVgK4AObJSij+z1bzs0LOEPigVTXJ3lTmXtHX7y1ID6T/QuI5urMnflPN
4BJlzF73v4f8gPNPPlezpyFpKRnzUPcaw4YK+cVZ5LsvRhNkJ63O6k1PTyxRIgmH
`protect END_PROTECTED
