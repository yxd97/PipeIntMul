`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XLwBXvLNUmd6IvbhORPSszPvavKwQYXiRSVzY3I56qqXy4p7C2nnv4e/eOklC9Po
Fl216gsZ7HxRyfHRM1l8Mo0/nS/kloewKV+KF2KWQYsHmDkqGgiUE09veO6pjdx6
0YUTnnTGAQHpGpKOqmBQZ4+bglWqsmO/ute2pNNOJEQFuwlIFnwC3hJGs2pa98Kj
ZXjAuKsZ9HRBH2XwzdJNGaaBXVh0+x9K8+anUX8XZkMsNW29b+UVPuFryFkvOR+/
McKvyqXf61/RwUdbGeXjd1oE2S416VGnWNurFiMLk2rDsD7nq/6q6i6JTmdijNs8
AFcWytpS+iv/r0axOLxqqA==
`protect END_PROTECTED
