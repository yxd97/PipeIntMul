`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9hg9o3JPWUvukiM2fV1XLmaYqsrZdhkANmH/T1sb5jiz7Ue6W+CApcqkn2TPdP1I
nnyxcTE76Ctamg8zncT9a4X3zysKawcudRXXOXtoydvpWLA3e077FNaEEpIEdwvm
0BdN3VUmGdg2eVCigbAFYuvzungH5w6hcDcN1swbtZ0ZTdQgEa/7AitvHIC2DsSd
2VONn+C6NcyNFUJSTNd0k0lOWgAmnyfIfO6RPNTC2K5WjaOQORABxyOfjHuRf+OA
kbF4+o9h5O8kPKuvmT5AvltkAICQk5wvozthLbwTqDyHYTfUEfdQfNnrp4KO3cfv
j9flSwoxTFD/TP+Ot8Ivk2iGtm/B5Pgs5rIBTnTLBNASb6x6PXc/UDxf5KX9Tusa
7DgVwlc2vqWKQOw4Cxzq5Iw5cf5mLTS77b0WQu2Jj6CnGUjrveh0hGRwyUlcVCfa
0yflen+Ians8//se6/K9FKxIi5z11SinBHNHSE9f87FBXy/VuoyHEQ9eR1OHwL8x
r1epEyu/ulv0lMKR6wXIldKc+6zlPrARpoK2+mB8pTlgSYJLgt+J0mab0cP+ynBV
CEqFtX5fFVjSXtCTOcWiRc3yAQOC41qjcerwvTiQhF3CnDsSVyEQNml50aQTKom0
sFWILiNzzaskgbtEvJTz4B4L1wBgyhTUZlJXubIOOOiP16efFSVA2ABHFP0X7mJh
OIRRdqkDzjRoSYSBQgpedBd0p+ILWprY1Wo3bW5xatKCyobylUGz3r0ENU/Zw3wY
MQrZcghBXabRAzRFe1pfR7QSLT9LafDEaLX8J3p5nHbXF6gzUAYImt03uywyAtAM
HmPU9GMY0qfaXS9VJ24kMTSV/7EjosQ0EoJBGhZsPyyJtuuR9zxxVfsTEn6A1MTI
ZN9ZBd28iRSmir/7izdowazzQY5uDakxbL1+Fc2AJ46o1emMUKG00hEQV+DZPpqZ
5QIYPwwn9cyf2SECAdAlw8Y165qcUnYN1hU3dEhwG2sT8804inHOzx6Pr2eNWnrU
Lc6hEteojJ42R7KylUxbNkEAqU2ve7JHSkbyxx8ez6LKjUun7ZpKtDt2Pb2cENo/
5x0aFWKl/UEiPglRhUiYR0Bh968GJANpvRmENrinKiHi2lbYpsFgJprRgZA4Bqxf
6WSMaezt44lxBvbw34I8mx1KgDjYBYZtXkcGwxAyZKr+wHp/Z+ogF9mbafVg9bBb
Zl7OH+GZPypWxgJeQD35lm2M9fLnSzwPdMwvxepecNWnHjqPNIZWdb99OeksLApD
qpDfW5dUXBc/TjjC95p//9+82x8XNTlBwY6TY+VXASxegsZmYuDB1PRj0SmeLK6e
IzVgxVGwo8peWGTLh7+uJ1aDWLBHf04Z++H+Zf3+LHG/rQzkuCt8vaJP/TNTyM9G
g23UvrAG02LyqpPYPawEd+uSFmNHfmpZIhGSdBNQbsYL+hM33c7rERLAH4HVgVJy
hcZXf6US63R6VsXenKObxZRJK3iFx79wrPqFyCI4oGxJnMMpBPWNcSQjf0Ph2MJP
okjPrYEEU98Q5rCkJd4+zEFMSC8AnHVsAHQWs17kFc6JrP8gRTJ4MCm7hprDTZZn
Byk/+AYlEemHknjQ7aTVfEZARlIk58w4h09O1ans4Bw114MIExfXQY1xKJ5UhivK
YyJUlr1wYBJZFTzFwkt6tA==
`protect END_PROTECTED
