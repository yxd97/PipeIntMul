`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gag60HNRM4sBcKszIJ3ty/E4qghOAdeFmNTG48b7rh4HYubuBq5OlVNBwQGEWH/p
7xBpKgn6aYi9x5LEQAC+no7+4/it1rFAhI+GvzGhSk2HbzLXAx8y/LUaBL3aDd7x
tMMzplE1mzgTZoiQLMP3pO6Oao6DNQbpkPVxAj/OhfXxwumqW9k38s5jR23SHf9O
LGyvmCStIn9q9qlhrqM2L9UqpPD9HAJiHZNZpY6nZqcAY6Tr2DTq/FA10bmYL31T
JjHWtaUlzj9IbqJO5hyz0q174dTHwNVpdu2vi26jmn3rp1TYMo3wIUCT+w6o0Jz7
RdBzheA6pF1fMhQ76Sf+nqiM6A4m8jLp7/IwlvOJzwG6z/kPRrxL/bgZEgAsCgAV
JwlBvUXo4fDijBzAi4GlKCmek1UQQxxFJmmDkblbVwQ0hrW303HnnF6+BBqPyELA
mEbMeH1SfuDlzF0fmfu3leQ/LpBkiFF4RMMa+lTA+wIWJOgsLUJvSMAXGp7mkHSx
JA+yMgdz+FiVGnpIw0beD4QH7zW8Md5DhHL/RsGypezGZCRhW5K6N+04LbSewsN/
KOIIoD6ZLjDP7rAAqUhtiL7G7rj9E75lPWq3YV+xfi96TgYsZUZ4sHFxNCL1CQid
vLcNQUuGMC3peJ9LNmRWqxdLgKUzwOw4+5KEPELeT+Uon4Hl59z5eR+iyw3InGwt
A5ouaokAJfAC5iEIhVtDxGviFQrAnIEOFj6sM+kHMYeR6yPz1p/227BPFCQSHffk
mu2Dd4PxWu7cIDVaxwscFNXzMGtl0zN/WJ/JMsuD4RtEZG31Kmfmt+1tylIQdIfY
YtSBlSp3Pmn0XyH/OZ2iLDVcXxeKpUzdGJMTUzzQaWZk9P4DyowGMk4yaCy21WW/
5Cw0iThnpSFR1sh1ufSWyuSngf4uIZ65zDk8heW6fzlYSkoSUMZy41Kl5m37NDyU
sVpDUePMEeYwH2p7u+ytrX2gtbQIBYuM0T9PubIYktk/nUIykABIUe5CRxs3UUq7
ajMh7Et7A0S7dQ/lTFxs7he4uHQchzZFRlo9Tm0sokFKNBltv3kL1BFeHmDybuQx
GQd3B163KmHzrGjjHr+y7g==
`protect END_PROTECTED
