`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UYhAu2aGgwdV6n9ord80jKlYjf5YTvmcFsC0Q7mCvKVURJ9boMGoc+MPw8uiHAjL
6LyCShnwVWrpeTezR9lQijC72dslLgdiyXPeVoVE9sihg6NxESag9xepJwcdswFU
JySUD4l66z5PtKZehUUCsYimOwFIewYFMYXk/ihnl3vJpkS1rej1WId7DNluQocm
W9wlAFQbJsqU04JepVvzC/rKoJiradOuUe4EgbVv/qNOnEUo1urVr5hkaWwzZD4H
v4YGiv8cNemUy4j0BiosRlLvwnQoHd5Ekfj4dyeoNh+ytWnzAjfOe7sAPUcLW9vI
NG/tOY+aLktBUyhyLFK3s5SodMga5uoHcLA15O8UXE5T6SrFkUdoGjYmF/NnkOCx
csOjlV3gPzhkRXb4ihXyXBb1xPsYeDPkn3LmkwVyBLjpsxYk2hBZDFYNo5VmQMT9
GTMTQZ6MkoYx2F5qd0EIF1rzazc4KaCVYcGfMckdpBwUyQsjHPM827YudjplYY1L
iAfathNZmufFFArVCY3IstlWQMMMjC9A7k+dL5dPpf5kdKWV/MckBS/KlDk1M1CO
MEIjV31OvTKcqrwrXDIPDf228J2hlG5jQzhWlZNOE02beqFIdvaMIp5oNXoq55PZ
`protect END_PROTECTED
