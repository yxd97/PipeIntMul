`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rWHmvHxup0voKLSKdNrry7O23YrmJkRp34lo0NllZk5+NXF5Bb6U+mPJ+Ow/ZJIv
nerG6MUCDVot24qfSpzoBLT/1RlthkIKB8K1XGthN58XcbCG62nHdnEqJc3vcZbJ
hvT1Xf/yLm1hDZhnMtWEZe+1DIFKSL+jnfanN7CODubx5p6pPkOZ2kNDMhPkHyhU
DLRmnvDZnVt52lkOaRiBOwJNHBTG4RiQVaPfpGOjRGv05tWwti/LVwXm5RPiVI4L
CWkYt0j72wtn9X3bQiPTMt3onByjh89GfFNv0prX1ziIOVvu7Iwat7FLZ66QLTFF
7K7tKCRiMRXksVFH9/Rz94/rapdzRfk9g8Am2lQeA2uyAlszfl4Kab08EzVNYlZ4
uQ4gy4ltJzd0hPgNvwEd0eKqXsaqRIEGH4Sdrs2QmTHYPZjXuxgZ32HMyT8ZucPc
MmFQ6Eoxp4/O7fRMStXhNHl8jHwmpAVaGb4j86nlJ9lS2ktWMvBwOm9rQ9X7wu2d
bVpEBssK7HCN275UElud+1QSdcWBqhpYxz5JTUYJLWzHDqZ974SRnXzNbvZ6QW2a
KtF2GFmnUviYYoL7VBt+bENUqlZw2RPCyJWxu53juhY=
`protect END_PROTECTED
