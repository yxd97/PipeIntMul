`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LlBcqhwHhVmcSFr76dabuABd3D4IVdeSUKH0VhQJ10kGfjxmwU2YMYPWpotDHhlV
BppopIDHkYyPTC8sGSfRE59L/2Wqug6QzgrtPidpdw88olyior+voIN+1o6qJm5V
N+Ju+Kb7EtnBJkPvpkA/vvqgD7H+X00c8qg3Spi7CZ9yXiQ3nsHJw1SjJpEvZeh1
X4dbkGXu9+WYDq6sp2KnVSSAYyDOfpmmXPobVCGsmrahSTdE94Ba9vinXc78UwuO
awB6cIWU065hHuwcXXaDCThyKLcWbxzr0g02k2EB/3tyMwOXm+d56PhenQWCfhuw
RLcx/Y1Ua6RJP/brx0FtlWy6zMBnTxrD4/NWgx5Q4UAfBAgxFC3mBoay8WfpwlvQ
2INagNmrDvrIXpSs9LmA3AQrKuzkw/yliHZztkI/7sSDiCcfAS29p4oUSVkSlXep
1eyN7cZb3Vp0zm76Gsi56NhbArdCADfXnBXyGlyiy/6s1VTzKuAM2823DZou4ODC
eiZ+cJJ3AyvFmXjMFKWGMomgtZk/c/sCf2hjDRuQI7pmiFaiYWlg/zfMwF4DtMo9
XwXpcGN3qJf6qrUxPOIW23Fl6apYskEfiJfuMmaERNe7tKBtX8JTb1lLfIwuP71g
D6+L3frfyYBPGXr3Ap2xwlLFypgWfojOFljsRZpIR8asr4gvnRW2tZaOhX2o3rGT
s+GF1AiewP/6jpvH9Z+XISfnRqMVlllfG2agcbIeRaxwqM478/I06VekxzVnxVG3
FPQz/uRbNJGYaWa5nxH5/g55m7cC/9ejopPrr2eizuCAptXoJQo3NzTNV6LTCx1m
nkJrCwMmFfBWMDREa3qzOVoRhFjwgm9cKq3KqIMyqVCtaeFp3z9WzRGwQQRFH8uE
6z0DbSD+S1a5d0WVVcguKqrrTJNaFJXdat/bPBaPgSBTO7+n+uHyppQIjCRIRjlK
B1CqQODqtMoObGpBZFFvpph1YNIdVus/SdYyEHfx1UkvqEHs53Vm45vH9g3+DkM4
t8odC904WGlbmEd4NAIdmKL1EdeELdpjdNSgk65/8njG5a4fdLx3CN07Y6QnjMBD
irezxDlmIU4W9+Wlzqy3ObRwIWP+rVNUAKogLOyJ4ZD9+uIbxrOf/PW5Um6okgBb
c3WaTAdLOe3cc630cNIe07PtnL3ljZwAGYSZYt/5quyrbtcxd5dwbERoTUCmjTEs
mMDxXXwC2WdgEsmERdnQFvQjJOuMvEHFijLbFuy8KFbSGwxx4UbFWvQnpQ0iy5WN
NeBO5zmcmVAa1lGAYEPB+28o5c4fLfG3FDEePZFQuoLbqa8etfxGZq/aVvi5e7Hz
qdrlRc7tathDxssSdKYTu9sDeJ1Re7Cjzk58kafMngKOWzL9SowV8JkfMweJw8q0
DQApbXn2ZCOlIfjvgRqU9GDkgsSwmdm/Q7JHRTdaf15yj8Gzc5ghrsIsvQpscwJ2
RoFr9EVt9LE7FScz6Io14enTtGA7zQs/4CbFBA4GmNPcCpYJS94r1Is/NvxRW8A+
PDsW8X+mA4diKOvozjJ02qRxUeUs7N/psyXH4B7I4eekn+QKDziv8c9A4Xvg8LXY
HcKCXVvST6TUXqFK1Ct883zYlFIDAO01UmwvfoAGSnkmvpi9HHdJpAYO1buiKGEl
amJMma6YeC6a27/oggOlLFxsMYFhyq5ncaWCm7F6qZrMUpMt1095cgCNpOsjaBQH
odTKMQoji5f2pLUHcE7nIxGHtvApGNXlZxq2ioD7QoCsheREObdUkiNNmR/REQJC
uCN9S07BN86TaRK5TLtTqvYOioq9P0uQXFJZqkfvAcXCe3PNFqUHIupSlbkH/URy
AylHOkx1QLTxevQ2OYzO4Wf8NWlOZfbkR+UPB8DHDgZ3XItJZDHUPdtWaT896Oaz
K2HyOWv6ulKy8hBQKNFqP21gaQU4q4g2ADYlwQNPjmNOgiq9TrbilYfZElmPlsIT
6XhMEFSQSAlCcMhxtaGZIv+O8Qbf4DkQF657ij/dB0WLZ0kQ2OitULlg4pV0YwXH
tFQ7O0V2gcqA7scMk6wE402aherkiPBoR0JJR7Y5Vf732a9Q7lplyT2kkqi7D1Wg
rzGqUQGb4G4XF5RRhsLHqYPGOwCqj0sZfgLea6eEFYpotAzetWx/gIYDwnNhQjMS
6VQTB1JLuY8f6Dqfoy89+eGb3+n666x6wOCoEm0TFWeunsEDtzfPtaPD7rd6WhBq
eE+VthZizXNhQ2mAzZhPZijckDAT8G4nVcJEHYOgv0czEBXrHF04JKkXBL9RNxwt
Mfa9oVklnyfQBp8stQdMupKrFKgquHgzdl/VHK/4STQZ87m8jwxjM8eR4nAZA8YD
0bBj5RwrqxTutU4kjIqGoTDLa0hxws5KVexDZ/mIPwIXF9KuVTet2UMubeoPQcGe
Xp/0WpYDcUDUUjwGZR56HVKHhdIu9b+IpyWZzlX+v/SMtRHRHZacq0UoEZRc1Csx
OC7dHv1QiZZpgOiZjv8CIroNElnoB9qBysP+rfAAj5XYb7ktHYUhPGklLdQq9Ex3
p6M/+dxJUzDThku0bxb8vbASD/x5PgZndEnR6DxXUIbYoeqtnTkPTUeqDPXtdoq+
1SwmsFBnlICnNArqYDunD6uYi1Y3TJSOq99M0zmTxsD8hQL/GODxVGCfVBzz0PzH
FZP8ZU8I9w34L3HhTQFHWRp+KSqG9uDF/177Rlo83pyR62aqY7bx7cTSMbLaNiMs
hVCZ0Znch+YsESlXEDoD7WOQBQJ2prrYwhwf5bb6SMZsSfgIUhKa8Hg+EkRO+nvi
ayUtffV+xnz6nSIG7F+GD82pIf43X6h+ASLblLDJ3X8=
`protect END_PROTECTED
