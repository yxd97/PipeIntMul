`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rkCM6YAB/OCXfahNzexeKP3lFx5TNjQrwwco5v59YDR6UNuima3RERvl6cUjXjv
Ixe3LBfcU1HM5LbbaVByfgR2gvsmPaf75jNWoOVMD1T1TH1Pd5xvsVcwcy2OroDH
E0udarDXT3SMqXATthlBVf6MECcwmeLw81Oknm8X1H910niVYRPlXCSRGE4MafdP
YA9/2s0kQ601iohANjVtY43o8Z3RIuLYixA0J8wIQqZ/OTES6l5RkJrwXPi9X/qB
4x7uhLdYqvaBN/SIJY/r5Q12M55wAIzY3hjwj9fgVHJPaSw8FeHT3+I9PIjb9VGm
Jk43AiW5Hntp7FFvlFQZNB9yOZeqEYHrauCj46k+tYdDk3i0knskdOFa0vWKNY/D
1XBGyQIq63vtdoNiiRI8XhGdPuQEOVhha+vx8MXCmPzQErmPOSxR6t9I8SWme+Tq
5yi0uW7weXqFFah19NMj8qTRdd6OC3rZYZT+jp9ky6bKvSnyVo+Ol3jc6AkExgAl
`protect END_PROTECTED
