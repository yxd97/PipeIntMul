`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kvis+9UTYJEC5hrrxGwJGbRGY2iWsyA8LwWtHR24ekVqASBwduQPsoWotCwtcMQQ
NpK13rQYHr0OUzKj2q/Cvdu415qxyjt18+QlQ4vbSrwk+rCc9PG+wDDjzjMxcxU8
l0Q5yy4myjfCfDDk60PVVoNsLW6WwAk5He/7QN+AJpMOFvovwgHUzBPO3A3rBw3I
zI0LLmae2S8hjBSFkNxhBQGysd9Sbumbp7RwrYV3hMWdb6kWZdwwblaHQQ3vJhxj
TEkcZD18aSGtjRakVPivlJuYDAuRIv0baNIWEOvT25L+a0rgP/E0GXQxCPj7jXrp
VRLMKvRjsM8EjL6NgZS3+ponPaZGfvNr+qRpQJc34UWOi1ug5MHaSlVi0C/Qnp4v
Vdpq5rDjTFjRLj+utFyOBnMDWblcDTwpFUc6BNXCghpHqI9O29zi9BIVNIC1mD7Z
MWTp269SUXw7KSDYE34n/MfXEaoVg4s9jsKE12+fzb+6Q9SIja75wTfWU3C2LNOe
LywffwfOEa/k2zrdnixMa0ZVq+yxIxJYofuiDJRKi5hNcsNh4XpwaCn5tITJY6V6
hZ800SlkolE7CuPL+d8OupIebjVMsLmdhRcO2g3oI3+VtxWoZisuaPQ2PA9vm67R
ET/dKKqFIW035MOO6GWwgOZQtLSf5WwlrbsukSvozsMUCYyL91pQuonh9UtRKZ1u
mriAeqr/JRtjtB+05mgM2vyaR5UPrbC3nNX+bzWpuz6LNGUpOdseNUKIb+flsiUq
4HEjZ8QjGbqickBT1ru6WCAaWphCGJJtjTdnLkk+7kbiR+vOnX2HA+QtYt0aOOSG
QN+EmpVqWD0xrxrZWu5BJg==
`protect END_PROTECTED
