`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZYwD6u6IeHAxaaAw65k2j1aw7+bza+201Ut1NkJ9BD+bweHagzyq9LVG9e68Fadx
tmwaLxdjHQSaa/P7vLN3Cj+KZ9q3WQbDI79t9EA+7RVlz2StM2NOKiOC/Oldb28Q
rVhHeMiSqOyDTElrESER6rPl1YrZTbkqT+FWm2FBxpsxYt/dUHpiH9+98RC5uEoI
0JZ92v6V6UlvQXKZ0UerbNDfYvsptYg/v2pBNGUSIIV5N66XIjabi0mMw3bvLHRf
PU5tO01r6OrZdyJLtgfe6w==
`protect END_PROTECTED
