`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dLhhpX5YSNtKXw+VOYXMYo8nIZqzCHWNDEldOE9UK1Ebuo7oF0KVdDS5dfjKKylp
GJ5qQCfOHDZNED0x23RUNnWvIzvBw3FYp+Jm+nIKSDjVB9yeLETG7EfplZ+qdMUK
2IK+1AANcBOCLx575P/7cr6PPTPQYKqvVdjMCAHYuhvK7u1H+irs6YyRxV/za8It
zsoV0AMgITsxFI8oQuIDzevOIxz69UElnR2JVOGi9BtYagIQh9RG/qihHom4s19a
eZmmPjEsdn0bJpOssBF4P/15NIQj+jRCccqDIb6NfqXGJgJWy3cPobnC0iwQrUGF
obRMvd1Dq4V3Rva6eYX5TyH+srs2Gn9Nx4qugFj/jlY3P8/zs6/xaDWCcG69exgk
Ubgh2mBtJ+HzIdb2Ug3KGSRzv9RKhhvQ4gGj6r2I8+W8JGjUUQdvG2qtt93QWs7H
4ZzsVjIPH5BpJjlVl3ShxOMBnq8+HbsIbgY1J52lrBu71HxV/Bxz9aLJG0akPCY1
qk40yfiIy5Xycu1zLw/WiVQ/uyPwj/SqAGQAw1Ug3jxHRoGcwpuLdSt0HXvNUnEG
kYjSPoq4Pu2D9eIioiyH0lRwI0OGbTlqh5NGIaaEFlLlQ6stGnCUAK47Y0h0AToJ
mhWQ8jp/LyafWRqJTXVA9ISsZCMe0gf/fCcVKz6rMWMXX65CBB9Amap6HASbDfcb
4q1bBjhj/GL32txz5GKR2A==
`protect END_PROTECTED
