`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5w7Qd9u0dkPwrjM1PlNG+NhLDNHTbtnXApQVFuVEhLeSjaulkpkp9POTidsc4vBd
+47COIVXT6GzfsMmeCdgz6Ta3E4gMni+j434kSrVpPB9DAEVmncQBlcSovPJfsEo
8/iaFCixwRLrVuEsTcgv3l4EaCcbkJ1MZlkTWA0Ce1NLDKuv0gEpkm8A53MxPpV6
f2rpJpRGxTMrFegcZuoIVNUY1NTZiZXbNzpnxPoQhUa0qpNMv5c1Vui6Kii5iFmd
vFCwIhHdecgHrNJ5TMOlAVeFNd3KrUBqKbtJo/CVdwrrNU3lJDQgJDD2Bxhamwb6
IPMWL0M5GMufd56ptpgyJ3RU0+y8y92lAYR3HOzuS0zd893bKZXhy6ZzHaEWTNvs
4wEMXWpQK26vgkGlGBSvTr0ZKgh8kR8+yrfSx8/lYPmOCfOdTx5u7Jr0CO+vvrBK
4YiAuEM7PtoQ0p6LZyXzag==
`protect END_PROTECTED
