`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0H3WKneoee0DnTu21Xb58tSirr7ZyFoxAPJsPeILCDPABZDIO3VZd+ZfdBhgC5s
FEvUQpvoCczW1C7MhlBzr3Wen6Mols4G+UWvaMeHwOkKx4/FVuTzEBtlUtinML5K
sovXHd/oWd6fSbu1kRbjnLcfBXgdKG6kPw8fMkM2OIm8OY0bKb2U7BCBkDfssTu2
DH4kG9lyzTaKC0DmLa5uFhqJpRymZPDKUlItAN/eMde91J9+3XvnxUUxZfszvkPT
pDI48KfX2v3qvdZT7RemDXVwYvBwzjCNtNLJs/EZVx4RLBcXMalQgngrMttCh96R
QT03AiEpNkGEXasNEi4R97JpLdzOAyCCyxdTXW5MDrk3k+zxByv2QzncCojbltGf
MSnMyWuWlBJApOzPY44mCEtJTUmoSHgRwB6+0lg0tbKVmjMHaPOv1PgiVKdONoPU
`protect END_PROTECTED
