`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ewgK0d14jBFrkkkJvH5GMIxYkxA0DasilVF3p3p72GKb73BNLiOCha7+pA3ExRWg
ijseJ19PJ9SqO+kGBdphHU4mYbbiAZst9knt4Q8OyZy7PDQEAbQ+OB0E2wvawCjw
D/mR08e1nPipKakjC4HhZ0xOBUNzBmJ7JeSBGJS4pTIJ2FGVYJQ4cJ8Y1/dDTJ4f
Syg3pSPnhJZ/4qvjcB7gmxMNFBp+q2Oga1+Zmtqi4M+ZU7s1DiIlQnkepOwiW3Fi
rwVaX2Qs5Odji6VSFcZvF7RV8Ada24uiiYmgoYPPsNRxIe1bydkyfyknrFcS9+7j
pzWViPa6idRTBgf6T7ehkQfWNU+zY9XUQBjsMTxoBszzjArsuQQaZwi7DUFL8pdj
N6rSjQL1E2uoehDljKr8Vd2x8R6NPjjCxxl383J9d9I=
`protect END_PROTECTED
