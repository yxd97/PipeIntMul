`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CD9rWZiLsO3ABow+6M/5rsMveHZUUd2DxE30dFFCIK+0tKFbeP5F+8Rbm2hebia8
49y5Rd2RoCuKv/k/EG3jG0EM5h9kjfJyt6skoai4Q0zF5Hq2UTQgXEKblY20kUoV
DG1l4KRMUk/FnNDFf2y+vDDHehCXHyoCwES70c0Xg87DZBY2lBNxDtgoU0iA8nNJ
xVPGu9wcsRslAczL8CLu9vHZuf1WtfIWy6Rg1+ADfwnHA4J06++rDRwjCMbCGpTK
IyyFuEBJyt8zsdhHVkXse3qMOfMDpx0l5zEc/PvFBtMygk40JfMFGLGTTmr64wm3
8j/LWm9TOze5EYu1mT0v9Tm6Kn49ODx/8BPyFAD/mNFYvuApzzsootYJMR1xe1fG
6EkHrobTvAZGE4S1hJAAyg==
`protect END_PROTECTED
