`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHjIhKeNa8AkBUhz897YQouH8+HEkcdo4KoKMADNuvKr0jlvlm2pkbwiPkErRaHe
9a2sHSZICdkHvgUAwBYyMdMBQiFo6W9houfUoA+pC+/dSqKMyd6khc10D3eA5Ncu
v72L7l7PuYzviBOysbi190uh82ZHBIbLX9Y2KrVthLCTfGFgXx6iFZUrUZtzA7+9
JZuXJwqddTiEO48xK6yMreWIt/2/sXOQv0uWG0RVFa13b0ThLAA9Fd7mPTHl4gcr
sSI4io0uBX+pKDMFbLH2z2zX8HX/EW5ZBYkP2ekN7REIl+V12o13k1ud1dYwBP/9
gLfpaidNakvxZXZ38PKYvYL0anZet1/tlFciG5eImsYoAqPg6A2MXDm33uHU6Fic
Wnn/11r8LYXltS843uMr46DoneRFwVRobqJ5hsgsnC5Lc79rX0cVGRScvxhO8Lo6
EaTE4EcbENOCta94BdRa85Cs2Pi8dA5JTCz3EwGgUyzRocnAZUdIkOejytOJTSfC
6lGaVJ/Yx7DPNzmFM7U+vVXTdEFbtt4Tth4yjw5zgRDsVX8UXmTDaiYl5wtIqcbC
rU7WRVv5xp07ZCHh1VdQKqTFGN8lnrk6YxpJMXyGHIqQ8BlLT8aQOFmhcV7NiY+K
MFbjfTtnodZk6JKrYd/c6t9wAgd6m0jDpPFHHfsf4J1wAbevuXLhY42FfTE4HmMY
G2FMTUR2UiN09QTaag2KdGkvusxbUVI2CD/clIm5o7PCNUe/ynxvo85MrfQKI6EZ
M5U3xVqLWmGmvvNLWL+9VyGsWOJy+Izmxl7CIhgeqlwLs5FsFDJ0Oh9re3dNN3Mk
6EGN96oJidjVmWPe4pwnHfv8c+lsWo90vFHzkrhv9obXvCLITJM68pGPdV/YXS/V
cqHxSw54Jitjn7pZX1N+d0UXqC3aCnCA76DA7QSkJaKDlvCPhv97iqTNFLcwFSjx
Acd7h3X5udjj9v/IY+Bqy/SkZrk5FTRyiqoVGCzPHIojbmTXQvXxOZZ3fsCcMA5x
PSofR3XUSK8SHb1DyRk80TIIla0/eD0bSbdpsBY5NsrIbzjLYazbPskht74ShVRm
1xriPCj0BjwbvhXRZEvMV6IBr/NCHXk65+XO94lhxotfpOLcqVKFav6AwFNhFrRa
dxf5ASVjlzQQ3ZuZQB55O37S8X5ru/cdnxdx7+bwAhER5z5X7fL8BeXfMhq2I3ro
kqBtS2zgv63ndIy9pdYwWkYcPD9ij9KyC+GoPgR8C2HdFDA8xA1lJ61vXTlHAaZC
QgA2xu0KxFuZHkeHZSPlf4dDZBUw4oa2vaTxjtkQIWEgFumiPtCuFWC7XzrnHzED
/PRVU1N0TnnOZmS/jn31vzaDD6n5NAW5FkiACZ8WvGo1YtdXMVI+NDM4bL3Ra5Wd
BekILq/Bl+WP1ByMc0hk/+rouXF4ggnuweV8blZOQj7/ZnnnDxxlMz9ZWS4CtNbq
MTtIjrkVo14HFxJBv60m/9nvyKPspIBMpDxKxhng2KzsGx032sIBCIw41qhdhhpi
RWZ//Si/m3+zOiCtZnNrzV8+w0gKYQBqE9DA+j33eJuwrj/WT7kGflF7AyvFVakJ
ZJwlINhbPcjZXy0I1RFg4zzB5fje3S1gixiGHpC6q6fU15mBE+25dSfpdfkyZoFf
1aySynnxW3vRiwaGkoNAd40R0MtxJMov6wxCvl4cJP60AnDUcgYjROMKew2jMbPS
0VYr9qXCi6lD8jEeLNhrlWo4o433JiTFXIotWTaZN2gBoK1xm76DOffOrujv3FEB
LmGQPbaSSLoSlTI7t+Zb3iMPbwgrsWWbKd8hAs8fFHuG9bTTbrf6prEFwXKmrrg4
+7FH26nZe/RrTzV2JDigyGzGvIwYIhos9G8+ZX8BAtX6xgVyzNHK/YaleH0p2r/D
TBHyaUgkTbgSUd06jF07X4thsOI3Us3Wv7++9MPvvS8JStFMlJtdqKMnyz/bwVa4
DDOFhRgr5mwZQ2OT6IpTCXZClZgR2Fi+he2AUcd2YxGH4oIv7w8LQX6fckSQ/qdQ
p9xbawRW9Uhj1+2XJhC/c9NK/lw896q26g3uqivWst/899o+ogX58aOVWMrmJUSW
IkUXyO97SZOpILL+0SwiCWW5KNw+AY2zCn/ZugD65A6CBbakdm8hSRhd73krvjDc
9+iQtShqmzm+QCEmBrT/6iGCQhA5XQ7MJho+XZCtcuCOyacSAP6S4DnXovkacPKa
KxW/ivNVxHUCluojVzPTsz5g/1jLNHrKO0jCqvY7Hd937anpkOpSKOdR4mASxCCy
TltC/kRVkothKNpCnJMGODAip0l8jxUiCBKML0o/1BctaUYTYHrNmu5SFbutjuF1
14si8h/qXhwaxPKKtY96tU8745l8RFCmIVY89sgfgDcbjuTGmP2lYGYe9+pxliar
HdprnfqfFgYTNnpsPmOA1dz5foPu7ZtBAZGIcEIC+QeW86hVQ2dzIKQnuu1Bthtd
rf4sfMUMOpc8oc6N8OVCJWAZFo9kORbAmjUyraEAJ1c+yTj4JJLf85coaYwxXJLB
BuMy6UmIUyvR0hxF39dJ7jV+dUE1/GAQsfup2GW/668ftD9FQZCHLblEcBKThCDt
kDjuus3sV4LjZpFLezmwzXxZ7VE3DjH3cc/YG1gxTCR/7KzYkbUKWtM/yM28Xh9w
WHvFSgpQGcizhF7MFUfx2akdJocuwIR7ilyKe4KjsgQJftnw2YNE1yCD9PuxoHY2
8o9v5ZafPTqjzXlo4L8ADMJB7wsXnRpK4lNl7YeEFDL2fnWTTrnBciXKCuf2NlwX
4tr2c+TTOEeux96wKtvLajZpZDcZmOoWtxuWti8acDLCek2C5crjoQKDv5C4YlgK
dmwf9gUsbEGlU4gG2TmZa4+zbChtif/ztDq5uuKTfsZ4AqSebzUPuwa73MqQ6XOw
XN5yDtI+XPnqS9pVpP+aLi6rdCOG+GY6DXhcPioAGbQCtpjZUGz2Vu2NX1Bio4L+
ASwAswrx2ES10knn38hhFoArogd0B/mB4arqFTL37M6Kg1x8hiKLOUkkX6SkIqes
vikKct04pJ+/LVVB0/sSETL+vT+fyijLiEDVClJE59HtyoPUSXLF4YeFkxF3QLx+
bONXrnbE70zBGB9I9dzfa5pol+4z8Kj0PoPu4uBoB91EQtt4tyS4zZ9DVaj45StB
z40h9bT60XztTNHMc2qzE/wgnuQXcIQh6WLbHtBesCnCwpYDAzmmwXjq8JQGFtzU
HI7DO+WRUiEDZLoTrZZ3crhaZ6PTRrjpjVX+bmjhYo+iUxLQBqEbr8HJcCJdagb1
9ZbV3hu3KWq+1KwNsyfX49ht6+hKVmvPSmORORNHy8HwkCguHtZbZitWH+pn+SYm
w1/a5r1Wvr7kBZ5uIeaASG3fNAqgZ9o4gyCuZ8qOamYNcwOsz3874qBMlsfhIzL4
O8vVBE48EZ2tVoKNQm/GOhP29Tarbbe8v7vwTlkWX5kNMVX9uwZmTXH2xhFC9+XA
zmPAVuaQiy6sgHgD8LUMf5TdeslkA4RkJu16qiFWliYXjxD00xdrUKeLO3fheC0C
hHO9leGW2q9c4o8z7U4zIZHJEYWxCPjitgUPDfj3bCTD+50uPcL44Lhk8fXIOuwS
f5eZ77GO6WTBRLAucEbai70DF68w3jMD/Gv4/XtPVSX1rZDOx2GcueygvRZoRMU8
KVtrO53IXxbwAj8gI3ycZ2U7HUpd7CYWyNaTZGtHVSGhx4HpEsPPk9mzs2ZWRJHH
cx8IocKLI3Cr79e0AuhR7/enxvuskgb6vkAwhYwLgWaneeh1McyNDl6ovAFcj3Gm
wUUJpMZW7AmG09942HRmSgnFq7tX1bzNNBvP9di8ILIs3SdymicUYfvANYT9M97P
lj2NqKG5MA7Tm0NzRdS10OCS1RxGyF8lxfzczVWEsDP5fE7HLPzqp3puGNLSXDAq
3Fzy2i/ajnr20kCgzdeJwkvaGgOpkvpS2pcNoYOlkcEoKRQujPwA7562qgRDcETV
s+sODjQvG0AR0ofTVrIXBu4RRuKhxQu+KBasdcbNpebMGnUPsI0BgBBlQBWFFC1O
mqnZpycUQW1qYkXsIX+tmWylYBlVOD9mra2PwvH/aa6snH3tgxBD2Fb4VHYF1CjW
PDi0TsgI8Sy1hSJ7kHQiZTKjW5vTjfHxJuN5ey7Z4e+0UkxhIrA/0WrsFKzq8DEg
1d/TiF8foaBAf/GXIG8GTl/lKLYLxd1RDHvSDxzhTGtqUliJBLB/tmgFuP4w44Wv
UNzvGS795FNybDbiSYOp1PUUBop1yjQ5fsgk3qbGRImqSfckK9lEq4E9UDv80RTu
D5/ds7tTib1kCUhse8iOdAR2gaMGCPB0k/T7ccJHRd1LSQb4Cnr2C7ManyS5Bbqb
MlormelEO3Eiz2z5ewQwtgTrNPmbmdOAqxQAE1/C4efhYVt4BeES1tW7NNitLX58
fBcSr0eyBuLAVf3St4Q5u308yu3dLqL3x/pPOFcKIqfRza7F00vpWT/0ZWrgi7Vv
xO2kMUYJip6wwPOu4OXkohSphJZ4LccaJB6Jk4esBBY2Ku7xb2zuOkhBPJdqbOwT
vhr7LzwSal6cgruDv8Zt6Gn3qP+3s7FBytlYgMUv5xJ4N8IYBGwoEigtxEDRP8Ch
rBy4ZSSlXm5QoFWHROgmrFhJyj2ptXn3BXN7XJdh8G0q80jwbpZJ8/fCRKkpawhF
TtT6uawaLvawZ6tl/iJLiBLLpUUw5qdvkBSBLiVzdR1vwBnyIdw+53kpT851Xs96
DjsXjercarpAcPe/nOdfDj8sBcffl0rn7rTSCHtfNTDimfRGr30C7iBqsuj+NKP3
jmcZ+eQWc+cjGsOxBvkADVcJZhPPpuJWRYY1m94pdteIYCZi+bWixFH/Bi691oqj
nAr+ERT0joEJpQioCtTKFfp0ytZBXKr3b2/876aL/NKsSPj4J1kFxkPBqNqn/M19
ppCUYCp7cfVeAileBuFPv5S6/l1qBxnX/G65jSl5lChzRqYNPE8P2vCwCCBjVs7t
ZJ/WqRlz1o3B1TFCm3LevcMLFNTHiqjA8AXU5nFceSlHGW98OaZ34X4Ir/1h3AMR
YZZBip7eONN56fEXnjnZtQ5038kFYxykvfayPKxN79yv9iFhrmkuUv4l52IZKZiX
g4ofN2Xvk4S0/GuQhsZKkoWbq4pqt20X5ZVIgy4eudycYvEzQs0OQEIMEnTdieUN
9bDNjd61vZVn2qd/3hw+QK2efJ4dasw4fzDrKpoTcAOLhwV9fUSswDUaDGSicJJQ
doEXwU1hL5nl32mJRgVf8Ftiy/ijSAUdmIIeEGRjR9U8UlX/XxLwMwVw4Pxz1bfO
YP2TggI6dZyTyoPkiY63Bq4wk8apDG9MKixD5zQEXTJDwoZBYFEoAo3WDMeOY4YN
Ol9w7GVWbFV6jviwgc1gOILlysA3dszMlc846AKPqR3/k7qbCUmQ1zSeNC/Vkgff
2WpO/M5nGYGijyhD12/JIB2uQSI9vGwNbHR6BdXrXb/SzRsYBqOy2lN1DU9Zv6oq
1D9wst6FGZDaJ/A/bjnF1KmS4z0AAyjAqzRFprbXubDpuLPgDLLkQfOwZdj1fOW8
pyopmi1fbH9eXpHesq1/EkXbLEyORu5SncIkJ5UU1de/cwz8YSDUPZ6tSpol53+W
YxF1ADU9VbxhFo77ciPJ+TEBslRAVSuPxCvKiybumx8zwkgMW8Hw6CoBekHZRBJ2
B3Yzb+5egTOjBoRfVZW9PKR9b0NLZcc8PuPt+ais9x7bzUqNgBahdQJmz9kgBcyo
j0RPT7GRdOphQVjHOmV4ernjcH4i6y2XKcN/TnQctr10EEGkJg96GoFKiksh0Gjv
JGq47w5p/lwRrbCctFarSX0zNefNFCdhFBOY3AtAb6yK39tR74nM3l713jJud1jd
WKGUY5DF4aUnATRgB3Zs6oU1qidpPX5GgjPvZOrv49yZwCTBWaHAJM1C37+/LbNt
8wL7h9HiZf3QBHDv5HStPEICiYrnl1ijOEs3ExwSmKl3vdYNiS2egYCiqb231ecm
xqj9YKf3kcM1VB79ABmDXE+jXFet502jdEShCpKODEy2ObIyJKKBxGprnvyxUaHl
LUuJFqqyfVFIUpsJON8E+14iR6neA2kbbUH5XOG16cALcRO3hifW6jr3nUScvs8w
Gg4M9BjThqEIDv5RoB8GvYvnUo1mDEZYd/j6cgQHg5tJNA0JsZJrFj/JWvwsh0EW
hDd6S9ZbxWKfKRVSlEhg0l2h00vpcmbsThG+zKmQ9EubKRKAKaSJoTSUTkDRkSQd
fHoDl2GcY5MZXOI/7pIWfwAGsLDoVwTx0vGppl2MMw3LGFoIoSRJ2wSf/OA+SsJr
KJYvBmy/LMk/xR7S55T1qpJZrYz6Af774WcN3TDuiMgLmn1EiB6GuqqSgsHiAHl+
nJabxkYVj3qgQNMVNT7OKDbNGuZV1TrpjwcGzMMTsD0iY+B3TFtZ/c1bA6mEFKzd
VbGWYJHQn3NamPz1taweJuCgkk1au522Wol0f59+fkmMHtR4dgAhaDfLT1p8wguf
X/1lvI67ECsZcnA5NiIJgh6RbhQk64w8uB/LNfJXzCeRBp67R1lO6HGZUfZkaW/y
sTbYyxPVovATd2tj8bhNrQG7iXnNMdNMpIvsy6o5ggHJZb5VQWPjiW5x/0yW5jnP
OikiLKO00dW2DP87hPPngZUrsyZtFZ6ILC/acocUre2lTXtT95gv875l8jWQsSP4
EJOFX7ygMjDo/GuqpwLG6RTEhqUvQwgreNffaNk5XustBWq0v8QS3/PZjDewRDwh
6I6Q9NewZJPrjBpVCYx3llO0LamatKg0QU3EGEzL1cCnNttBA9l8MRlsyu5/tf1z
xDmoQUKI/WO/CrdXfffx7bbJeH1Z20UVrATiZjYtX2JTtvlVPhMnlWU/Nk2dcyqz
m/yId6XJ8AZyMsk9/AX0U4e9SEJIJQQ9LfYI92LZ90zv9xmbJRwp28Ny42BR7n1K
uoAJEeEPSO0kBNr9Cvy+/F7QodIPrS76I2g1yE5eE7YgO1cFjaXx7nsyw5zC0559
l3yR0tTpAmQh3RiLG9MwcihksHxwqAdAItnT4zcK7rtTz0fkgMogBbxaXCxO7Hiz
qFo+eNY3Zus0WNXoWdPG2P+pL49rifvJNyUkBpuM3daPP/g9xX/DWl3Lq+sG6Tjo
y4nTUVvnV58QFq2GBAX2RLKd9XT0zvzgcVhIvfsFvhDHd0NwOu9UcN8SyZPG+NAq
xUZezOfyzW0CUHn26Zv3AyU9lmFhT85LAJqYncm8eSoO43M9rW9tXqDKIa5aPrvX
ir2T5C26iqyLvXlDudtskuarDkBrz40uEjMTepsa77m4CTC4f7cb36LYFU9/almV
60GoHYfDeg9kG9HlrweZoqab6j0eTHv0oxajh96sNJYeQqYVE4E9/4DAmJX2XHib
0DJQkokibLVRfKmTBImaYuww4aydxZbxjzv6vHe3dJtNYwq1kI/O0b0nNamp4H0P
08u3oxCdCsVmta+m8Ol0ZXGrbtUX6PLemQnKaJ8IM3foRXYAebQSMiaykxHVYLHI
e2kUm8u1jiRgtSKumGLQqhbbrdn9QzTmZs7n728MeMi4yzXstpuGNPAA2adaeW8t
GIkrn9Wjl3S0ZQqHTbRADxFaUgQIsILberQ+/uhodSJ9CJd4w9+6gcQvuPJygOqj
Vu4JJdG2GhZoT8xoHb9vCIUJZ1mWFvpZ2gLAh0YnicyrEQ3tN0WG/ael3pRHLLOT
bDeeOKz4rbz1NCui+E3/wjsWa46kNZtehcZa2UW93FZxs3j4ebvEsQ7YMK/OCv4S
fCNwwr8Ne+FzOzELiLwAGWPC480cE0sHhCGwPT1GgtYqbfSjcrpKqmHDl4OYKmT+
om6Ybi2JSFCozaoXg5Kbhm8iDVRbtiWZ3rmTUVCCCQ4WtRuPnyuCWwPn7Vx7Z8Vf
gd/JLZB6/Tz+AiWgioGBYbQh912o/9hV1CS/d0Gu1Ycahv+4UzjjfpzFIBDzLG35
oABlx1e4VIZUTAFgWVqDcGZHJson5hM/I2Hrshk/l5q3mu+wjtwnZmJpC/cmsacG
AAbnjmxkNviM6NwB1ODdS9ixR+URM/z/cGM4/Bq5vOrUOvDWip2yJRl0Y10Fac9c
IMPdZn9ZVxiRx9BEXYetyl54xiaptt/9EeF6xav9A53DElOV27V4qCJpk5Hojz6s
fOiNDRcm2e+46OLgGFujXvdrkC/ftqpT71csQcouuzkaue9MYpy+OE7yVA87720l
K2mS2eWXJnm+OEz6ytHUITwrW3tATq2buFeSOfyuz2I74QgWO1GMhxpqStS9dFFg
RU3vxxuDZf4WAKSp8zstzOw9akpu6MwaQQt5TGRB7IrEm+KXUHAOj/MARa+2Zs/F
q44IDNiniJsRHDdAC1eS+DIPP5RMG2rREueRKgpk13J0v+hP4nWiH9ObZ/1uqz6O
JbK/Do859mmi7iYiJMSC6c3Opn2WndkXpM87bSGYvOHSw75vd9O4gElNbSKzWycg
nnsPdfLZX2jq5Ig26VWNKKnLJbu9SV3NLM+TYgoWo0BFL/yYWvuF/fX1geKNtlDH
XOjeHhQeF8uM9ZC+oUssuzuogXm28A1sx9Qvg3KWRxyL9/6oXy2SJ00+TOWK7aSc
VeSagCXX46EjwUc4/jrm3m9EeQEyJZEKzuuE+XK9rqj2Wu+MMr82YCWly14Md6Op
tmgKA+yA+DDQUDpPJOTQq8Bgu4OeQpWgl1nJqO+Mgsp7obC6AUd6noD1cB8CXqRM
SbqL1shlL47/FZZKgpDIRZ2/q1iu10KbBDSN440NhwwyzVqWPeWZ9pmUNOCq2046
gAGzI95ZEGkAkb9vYkRwXP9+/hsaI6Qtjy9IM//omO9SXvNUHrc0TGRBcTnehNAc
0n+O42gVPmv7mlm0ccCdP69SwC0NQ4590I3KEh4Zm4opX+ZrrJrmJs9IfBTcgS38
GYHPhBGJivxHfFWRGjuUhlc/wa2G273w+m2HYh1gMlf+iKuxHr8VIvhGc2Am9flF
FjSfbhaNlS6LgrcBN3qccU+ieeXMhp9tU3j/XRMfJqjS6stpk9uIkxc926I16hFw
2vd0c8GwfTcPdOUFxsfew8kSPLfrXLUSVr7LO3f6h1q917oebMAuG5gDYaMG6BaW
sXYvt4LjtyOtZ/5n9tXIT7/HU3jyqGcKET8LVoSqJwOBaES1zrNF17K3MYDDC7l5
yjA0l0FmXUaPhws7HFZ0/vGm5Oio/Pu5ikRfgsjMajOsL6YKh3tYQrz+HhTLlg4V
qa/nxMzJcmuHWFt1CPzpAN9NvY643ZKQmRxgd7djPksSN9G87MKxTSNSjlb6Uxd1
fxqW0i1WqB9ix77Ve8597OAsve6/46VgZPvRmvPwRSDBETonhPBC9AgKQTOONmHB
vl/Hk02Sd88o0kvynDZ5HuPu35Kc7SSaub6GWzpevUdcqHDjlmRMcvzjtkypHjht
GbcZzKUVdnlRiOYh0wBu7v3iFOsn95lD6qsy44VbYFVlmVqdQmmTeHzhP7qCif+2
ekx3LogUVvTX6YyKs2tEju4BkW2ue7TNEYXXROBKXSKZnBnfdRiaBG0u+J1eCooS
DYCBhUQVKiCjTYxOfFbo9GREyRPOqb3bwu+onOyOXYnTTgj3lWQfO5623BRBj7GJ
yVkf5MfiFy02K2OrxxvGYY3nt+IbuZ1MgYEsRWlYMjAvuBAw9uXTjmOxKhdCodDw
6lT6k3r1fLr61Ul9NIqmn5hka8SlpHTGL6J4vW50jrYAAqfOEA7CP6RvccI19JYF
G2unlnHKpIKRrtZdLNIvU73LlKZXHlaWZp3iczEmwTLejCExvGYLt2sVbCfmRPSE
ppuWBh4yNaBE8iIw0dc8hFEvOkUGuR4DdvFGoLBqEQ4U7Bo2jPp02ejDaKmJjLrP
0ITuyjodKPiti/JwistTezGom+ahiWrxqW0xn2WhTEZdK68GID3Uwsn143xWwqoT
YKO3efjYTSt64RR4W5gZTF3P8G3vA/t3qCosvEqFAaRd5yv6zr8kGEXfW2hghViQ
eqIPb5us/lVH3D+usBNLGQqSTWxEc66+8YXESZlzgAL09oEzk5YMZ30yLgaJYKiX
7OxL9dOn+Xw5Ou+hZmuhyLuuRx+TKFF6ljBC5tTgCFM4nXwXFfOUDOB9e6p+EYDU
/dQyyEUICP/nG3ScuhQS29Jal7+505FRJSB1JABye9p0bDswlSz4aHRUeTmjaGId
CGqtC/0JgMyoPDKyyCgkaTS3Be3y7eBR539Aes2ZigD/LuVI6G5d8St9KFdLPD0P
/DPmeRbkKfCP3fU5yXfHoT2DPl26HgyCBsBLjtz6J/PPRDtEZ6saDKEoww0Kgy/E
HEd9DpEsKH3Dt0IuSs53n6We13L4Y98tlKo9L7ZuyPZJ4o5gR1L99HZsdmqpOuaq
z7uK9lr7vHrW74oEqIZ7JRJNk6JVL2LwHASFQ2lynm5bSSPssuzO/ZUy6dffYmdU
/93AWT/id3iUBnBDDW/4Z6ieG6oE6cX4J2yWafkxYkMd5FjtvH1G21Jys3e/zk48
SNtGt1Qv5ocrTkZ2MQ0QzuvXvn4Buw+D/LnxGIi7KlQ9X++2whdHMNNQqCdEVY1G
YIZbkhxWSIBj/XKNGIJVY2nxKTXf3kPlbdBGfujvXtVlQgXZ58s2NPsALPWJhSam
ma5UxnZrTq68kgfjjZcPJAMRtR21A9zcNQVHi8EOFKR4q6EzkM145jFfCi+i7pei
qOfHQAdAwU8k5ztlDEW6YebhcfjyVR4T16+JOL1de/nCYafsW9W8ansCaY4FWDyI
4/Dr5XJd23nSChN7sxAFAwlHFqkfsjlEKrcmBOzwyqT+EklCGCe0iRfWyZD6JydL
s2ANz5XaCozQw82b+46Lk88UoI9KmxoXBTBzxFFCV4UbOYENqNfExpmgH1Qm5jhH
SqN2KlY/qC98Yp3k96vMw4rrm50J5oNVkcjbyIoZDPXvqPREwppJjbMm6gbOuy8/
2fkVZ8uJ5rZI/4mBB+KQh7s2bLYcm0sKq6WJBlmJXqfmZ6sSpZtxyeWIunmZHKK7
YUOXCp+h+XhsAM+tmGbhMuO4hANgHNgJ2dDp8RxpjZzvQy30V8npLalIWendzhOy
rM8NsKG/+XKPZD4WqSzH1RHmlgoJzYJYOB1TpXD4hyffrVHXOt+3YVQU/p1OSRy2
o54Lr9M2cNRjZmCPWTAcj5IEMqEXi05CptgXLiyxusjgEYQvxnKM5BCp3aaai5D2
o9h6Qrr+OlJ4FWF7abRlFZy+9bV0SqqxN4wux3vWLkpDawYQ0BrQgV9HSfTJEvzL
7SiLQAfriKtSyYbaTdquDEeIvp5pBlIUBUOw0+9HyVQc4RXUE6S9A2g4NiAfU9t6
Jqn70OOLMF7JzRTjOHG1bFymIAjP9Drm5uIDDUkZqO4Le3kGa9J25LqpHEK+e5lH
j6YFDTRQq+TBDPFmnkb/zKTyDTZKGl8yUn2yMQNPcme/mkOiomMEwC5bmB+zcknI
y4qGJLm8tIyH774oiDgWfH8ytfq04zdYOSwQn8HMVsZ/cFgHC+U6AbXlOSb3xJ5K
akW0IQF0XpIxX0ZjklcQAHC8ylXQaPKO+9ju3uFibnzxfaznUj6xRud+Sbk5mh1c
9fVzISHcwWaRQvqa02vdqjohx6apL08VriteznzFDJtbxOVI8NBlb1NBI/WSHdEu
EvVUBKoswCQgNwDsfxA6mGbKom+NjlQx0tkrcudZLtpBMOjcb/gmA0JIz9YhAro5
RQUMy7Vt4rncjcHVuPTJxHO5kJDIVr8ycJkX2KjPE0vOTV1tPfIC5HXYGsaHW84x
4ZSVjHzYO60ZqrSU/xR5ziyx+Qc4lcVqYhEeXSVYdWRs1lgywQdYGAlulcPSn3cw
IcZCYxVDRL4M5tO74XYCkKxV4+M+G1J7UQ17vubGPxNzBBXgFXGXbYU0b0vmZGRA
HGNz/q8LN6oOwk1JF98B6fBdpdFWWLRaL+6dT/KsrhBckFIKuyBd7Nd6GbvLkd+9
bE5s2tz56towpd33ZV9TDo0xkHXN1lq8EMBukgSnh2C3NZNuioXdjdgpTgBA1mMl
qIAjn7MV2LAyzuvp/tfx4YfwwOKB4re30dzTqvOfddBJYOvXFnFOWU/25Vb4V8bj
AOHYKgPPSQRBaJVQz50FgjqzXg6YRyxt9ou7BZYFYBVwLo9cfm8IO1LOHQJVQpz3
Cf5VThcZWCQM4RBRmuinBWoVKzHAg7jejPqW7M0N85qs8cDJgEVm9PiISfmUJ0g0
WEs8ocen0wf38CqeJDQd2a40KHpmy82qGrig+n6Ne+W0i1nQ56ICvebfxaQ7mGzn
/qQNUyGw4Th/vpbvdEcQ43k5ayr6PfTEJ4MIdKAnlqQ4nu+ANA1zr2t3tcJRkwQa
4dM1sJEilYzHNbmFLTeH6Ierq4F5awqvzlsEyVm8GpHhasNoSilA9WBfBb63khLe
t3+I2DiYVEcG1wABpWYxr08Xe+Vk+ZsQfM0T/uNlpaYkV58Rgsqoddvi+FCUYv7k
VacUNjSp484qP/RwJ30wOMVqEutgFXhjncdSGad8/2Rksi5I+43tOFhk2ZdUZvSj
7bMc5aB/YQ58DEqnsuwxQQ2ISk12TQTp3SdzaRdKb6uiJUoPHlVSH3SEL35DQUV8
NinAab6z+aATgnBBqirKMKQU7027dq4iYuLDccfeF1QEY2bP0W3U416erOqgU1RJ
FuiWoYTfm698zJ3qrKyJ/HWkQGxeblODiqONLJGgbYi/KAUBbGqZyLFsRDyvSG8y
FBKJ3BGtkDOdRhBgSlx5AI6T8DcIZdJHcXHEpb15x+sMME/ltLqkrPqeR+GdP+GO
GsI9peL+DD9ktGll+SIbq+SZxTHGDWq99cX9963DoTLscXTrOJq8wWBeWos3yYG5
6JmC7pWNpDMMXFvw7DXQdC42dZDnOeEq+Ok2ruL1VOJXZD3oPYeROe1/1gdMEJ0Z
cOPELILLg71vWPk4X+BwYMEFikrNImiU3xinGQLOH5eWj667ZxxJ4GEp5i1RgDXf
tM2egfxhkAQ7TstP7kRnSsaiMBK+D3IBmRP7vU8CMtppVumzgmm7kpEAgeeeItg3
HXlt1MhwtR2X2RKg7nbI1SkeJGiBIou9z7a7vZF4TZGA9qDsJV4yK5Md1Zz1aZFI
dSFjUm9d9K9l236mtTLvcRcTAzSymgtg8Usyb/ufRF2B4zGTZxrjcXQTX+pv4jXd
VSmZppQFVfYgwtCdNBpV3JKijxOhszqyw9z4YubOxXvGPOkCrZdEA9bFlL0VHJRR
sjNMfRwCfPVduboN9OkYI76/yxFptE30YXsZr/8T5pAfz8LwKdHvUuFWXi1tHHuG
JO/dchnqqx5LqSJMNaYncSShPRSFcddEyXG7Zhn5O2Gy+U/7nFVbRRHUvc+Bt/Wr
peh/NaW+bQgIroryXxnV7UOIx4buCtOeWe6au2uBmzChQRbwhxfso532t3UcRumH
3yXVpNBQtXsZ3sA0Jpp3BZ55pdQm9FT++9yKlMbtXp8LlwnQYKGRLAYVhc89WJHM
/31MnRsZVq1t+NA820MMtHWZQ3pV9kguRbDvRuWsbRgOoCzR05OHdCqYYKgkachi
dBsTNGYbK8EtIE5ux9j9etna2NxdY3nUy3rQ3bIOVzZ/+dlJXrL+a6EVkqe51jue
ZQJ2cmu0ZVhBQQqi9gcPPYvvBVM5FUQKa4WwGsgHlTVlVO1+FO+LYeFr+P6sKztq
BZpmo8PVM+DYPSNXbrr37jhGzWSBbjA+XuhDY6Zxv2Ta7X/+oWJQGW94w5wkKb6Y
crapcq49qraXwoS+VWCqwBBVPbmH5XV8FlnysKlQ0Ko=
`protect END_PROTECTED
