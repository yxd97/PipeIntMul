`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+uMlgwMrEPj3/j9feQZsIZAWkqYfrfx99KxLvVzRQ59GYCbzxXPa4R3lUYTx3nf
RUbB7xRFMHS5dgpMu35gu6uu+Js+aVpIFhJGDuRINclZkrSP8las7+D4ZXE3wb2B
DgUXpTKCIJwTk9NjQWPYJG7X6PZlDLkHo/RdRuqRknOB08uN8zq46FvsGhUxEa4Q
L6pypBV7hml0M9JIK5/ByjBZSaCCDVIlXLW+EzYhv1tmQyHbOFJpF6j2e10so0A3
a6Yh8l9/to06+nnhNxKMC4tyMiDKm7VANuLyDhEVFDfNSno9B02bD4EcPX7zuwl1
yPz9tgTrCzYDF6wdnc1ARXYZSgs9WHPTXdHZHMHUSOzIBEvy225b6Fe9pBwUnab9
crKwRxDxQoYyEm17Lu0/zPd7xOQZnGNlBIktWYf7DYJLrBS0HCNXUdrb80+L2laU
2KXjv2+iwgl2sdyATqW4EEgNVEYPSMkpx5V+WEPY7FoqPiUhPqyhGRH28A5gIn0W
x/TbMUlmF7HOdmItu6kBluV/pyoV2Q7Q1Jxq7ll0aOMpZL+pGyAYtGcTslM0efGL
0aMR1Qd7i8TNqnjP58GkCWqHcoqtLVSt5QyGQ1UzeskABqoP2SW7O0Rw7GeJGMJ4
D5GQP2F/Y73pQ9s4NmuWnoiTPPxEG6wUaLn6tYMT9IAWvBVX8bLBP7E3W4nu+kIN
asWWaI2fgCDCCiCAOAc/b8g2bXdCEfgVLdxYSBIBTTkfpwxM5JmbciPbhlqmiMTk
RzC2x8y1M1prQOsLjFjUfs1epvoeRTMAMYTmfa2v1xdBjwYuVmoEaXmlzSHacDwe
fyEJw7ucfjbvhwn/7iJOAr8ok4JJX/LPSOx1/SoSD7Nany3osQbtxC0tLKJ1Fiph
yaoA6njLaairioN+vW7fGfD8znPezNBA4+PkXS6pwCsKQ9Soz6eoAm11NkVQVNSa
4/2TA18aGvJ6Vwgs2oboTw==
`protect END_PROTECTED
