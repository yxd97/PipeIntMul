`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHLZJumFKyPBbRYK/Lk65PFU926VMxnNau2sFQF9X8hYnLtrhx3kuwIGTngmzGm/
jm57iDJGLr/bvZXqwsU5M7X5C5Cf5TocyRdhAwsTECOjUv/ADQa64HeNlDxHRO23
OXYsQlHfD9Op3qyqq5VKJmbyA8EsEIObUZUdcnyI57TgyU3Xx4B6OL65SF98MstY
31HDiAsP1rWgmcDG1kKaCrEktzzcnF9hS/EKWfY4s9yB48rG9Er3NIdEPc5/qGM4
gtpl+be3Z2x8AjwLMeqSWnZLuz16aFv8gRlMJnA2vvFclZ3mJxZxI/ess98uT5zW
u21Y0ktAwn1qb3nKUB5Ij00btkjuk/SHX9ddS9yMp91dcJNbdOOxdcl5FNc0PSyY
`protect END_PROTECTED
