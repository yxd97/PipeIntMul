`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0biJCetZJlhhM7uZprf/NX24EVui//7zrKph5BRdGhBq3M9JB+uEIcdI7Ol/3Nid
dOe0akkKAYQgf7Huog5ggONW29xg4Lyy5cndWQHmT+cDXCJuPE3he1ZO05Clm56R
8+X/1IvQe47jUFhfVdN6BNFfsY7TRlmjcVJz0sxO/v84prNLVDbr8AP60bJLeRYH
jmPfKtO87YAQXq9XtywnEpA1udtq9h+PhiHPRo/swndUF3cm7ZHVATDay+KP721/
PJ1/jJBW1/zqI36K4RWXsjdhMde9nyUFTHkdJuDGSVCtm2AQiUtkjNE1t3Sk9vio
41BXaV+PFKKayE3y/q1JUEVr3GWbNpg1epft+DeLDKllkUspfzQglEwjjt9OYIe5
RuwA52ig1iOxntVhvzj+lw==
`protect END_PROTECTED
