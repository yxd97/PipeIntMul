`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ss1IsnhX3iCr3F74Koyx9HP6Ao0YU8NudylGQ/dAtug7Fv8a0oTspZOo5bbqzWsH
FT+gov7GKFad4zqr28ISpwl5c9LxjCSy16V4tjQ4hg+cFUrdqmeOHoyW196I95Wq
mKQOdWGXgdZkzVBRhUharQMLoY3qdjuj4MvT4CxunhW9I+5dVCvuMzUJNFX9eYV+
h2ehZL0wDNbnDCFjn+P4euPfCZSbjvTLh0/K0TQtwzNjujCjDZw9x8OA6Hn1xXUP
e5A7SyU9ZquR4HHnbT5KxYlu4WrbrofYPc4xjvVYs85uJW1H/AZ6AkP1xrZ2jl2k
81Gph6eV/JF9mOd1ULZyamNm4phQQ3qexzzocix9QN5W6kz7+sXgMS6jHZInQ329
tT+7Fcfxy3mY9VH2jC185hKIVTK3IcAKvdjR9xvmeQOazo6sUK2n6UhYwr5IVUmM
JxRsa1/YVFYATQG8DF5B7CR36lzIIu5fifC7BEcJ5GY=
`protect END_PROTECTED
