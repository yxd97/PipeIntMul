`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFCalaHyJVa8te3Mw2RhlxgnSIJwIGHoPuIeecDBZt+h8AI6kCc6mL1QO21ym9yA
Km/H6cUCIYbZzcw16e3zxp6BVVkBKVI6hQrUMZlqqdLJCHJnj2xi81mSpKBcVxUI
pQ/0Ohxo2eZzfXAym9loVaop056h+EYi76R//DCZ4c6+N2aLPgS31rYVdmxl7+Bh
PnW37dFq2QHxK9fmoVCaSURPU4xLq0iC1UGFrVu5GyU/sqXp5ZUBljZm6JdjH3Ji
ru+HMmHjgzol2+2tCQYIq0qQXHfn+amTMonyc8G29C8dPEHuqscqtk9qIClzEEC4
uFR3OPrB86qETWrC8x9RA8zZ83O5Eu4nQbcawLZCEjeiyB+ASchKZ9rHZZcaOP+d
OjshDs6TtgolSISCr5Cv3eShle96FAO8HNnU002tJqPJFkQQW1iJo34tJkmCuzre
O9gAiZbX4Bqddo3/FsIb2XCUb2SrF2AgzP+7JRsNfZAWj8NuVrUXX5BXgQXlHTUy
uUoILrpCfMGwFOMOL2FwgaGCw9mbxYYnm4l2xeNdrYyeJEJfMo4laa8dG91rokQR
tLaXKLuRQzyYgTPlut84tmSxpAAi490v1ZqZfRdCkcW8RKEqHdg2aiowK4H7uyGz
9Cv88HrzYE7W/d09h+vcvybXJcL88zP0swqLRf5Bdr6XeSLNh0RpV/X2dLcGv7w3
IbTZJiGdKqrLL/bMxjpY5USmCj2jahbqsdn4gh0j7YuA3n0UOB+JjP1JnKevdrXh
b8mvyJG3yQriEnFHSYiXcGz/UUSJrzy4xPdKMVwSxJEY6Hb09jWS3fvCIExeS2d0
ME+HyuUZNi7B/yeX2i1qhLnK31h9BTlyl1gdyEAMw74F39TJZQghoVbgN4CdefYy
QgsGrzWVSRwoF6ECUbzQG6dFU0tCqZh8KlyDPlJQ9Z2B90YUvEqR3A/4iwnkL+/R
Jd5LBIW3ms45hnLZHMJwWTskRc8Y03ZIYKTNw81pnfuqMIn+Y1pMBI/BC5Vy2J43
`protect END_PROTECTED
