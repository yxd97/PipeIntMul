`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
brEolTSfnofz+darz2oAWf3GC1h82uGo24UgL5X9ds3aDd8rCvxWjweEOn3/0Iq1
rDuVjUHEybhXVdx8xcTq4hOEd70BGwHhip0ZsuXcfeD+pwDz7LCwcqz7syatM9CT
QPV3t+WcCB4dYbxnl0NBGHIX+ORF3D4YLQxQYO4hVjZH3JakNi1wDOTKrIEf5HzM
ohDR3fyllqQuHcA+DYxBFJG8+64pVemAn76l8caaDh7TI4Je605dGM90+fJRIBC5
E9muXyc7ptEnoixp8l8lxoyueczygXdOFWrezMBuy6BrwsgUxJEi669TV+eGN/XS
3C4L/vJrWLEb6k8+NHOBNo8QmTVWdWPgMDbvew6p95R675w2QrY/+BWCR9fYc/ej
U2ypoLcAYD2t/9LdyAn7RCYdcCsMxw3P6QjMDkd7oYQ/6TE/Hpyt5Qtxry9UhGkc
WW6wk0igW+rUoiQIBrrwbg==
`protect END_PROTECTED
