`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYFi3jcdA7xwbwp9Sv6jUdciVUygfN20JE9m6StrM4IiigtbBmcM4tEteMoRz7vW
ivbCKcXYQGxHfaLBXH9XgpfPAEPKJvxO5SX942BFWaxlyVZQJlgTuq/b7XXflG2y
4yA3WUd4apJtzSND5aAJkqg4/S1CtMuiaUXsf6yReYWE7jJQ2/gP+or2DknF+/9Q
eIr5jZaeukCEdh37hsdUNuSI/EdcE1ZB/hHKkBr0Fzqr5NnWU7IkOWapWG5aG4E2
jJT/0peZftjXCnuGpLsZphNBNPWRO+tkN40XVdUWnq43UweRy16O2Er+fchZnvtp
6p/K5+eppszt4RA7gb7IK8u0BeV06qnxbb9kPsB26R7oL5eyHkcVRhvcG6r/cT9d
fTOc2bFbohK8XuUq72VVNVGFhkeGKZxKxhwOh4gMn6LTUfKpmslVYXPOAHr1vL1D
/RfReUGaCTHqXbmiphl2HT/EB/N0QF41XXg9gq9OVeo=
`protect END_PROTECTED
