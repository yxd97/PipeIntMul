`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nYoOsmgG3Eo/dkPT+A7k90beN4vRAfCIDgzyF+wSXOJJYaJV0XDJnClyCt16pa84
ekNgqfzlTfoZLfBzawgjDziCqocxmeN3k7BS1DGIeAFaoxH3WWSXS0sYOFjl9JDj
+kryNBXMhATKCrVYzBN0lM8heI++XZMXcyjdi95SEm9ifb/srRLr7fWCjDneOU4v
oSGh5fuUj3z3DE7ZmO/YQ0ILgBHo5Hp4kzxW+opSgJLO1hmCF+kuQC/9cigd2ef8
NG0UoB6sg+sQwnYNDIWkqBP/erxDoWA/nnecL/PIAmcrQV7aQc1BSvqK5LXC4Bzn
8zcantxUPC4nmKHkIhPOOQ==
`protect END_PROTECTED
