`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
93vacoARHcg3zn3sdj7MXCaI7F8ZyVhGDYMGs/7dJL9j8vXz2cKkEEwoAHENAS2C
FJPRufK1u7Lwp7cF5OwUo5iXhhiQazCfLZ22H6XsyYaR1y5CtL2vY/Io+5meDqfN
KefXB2yiFKjT6it4edadyMPIl7Jz8YVFIx2KYPH06tAXY1jICpp5QfQh2JfgCGFQ
sghN+sZTZqbj6vsht+TMeSC7adEQdh7diwewGH9wZgy/V8GSXmyCy7Z78JvWxbh3
J3p6CIe/D0x3rrmLAI7i8ciIdSxZ3tpeRYKxaaiTc1Gebq7hlCe+kt8UkrYNPoY8
h461yABo56DHyNWq8G7bHjvN86amjlsgmVLi+7s0WcnrvSX/eYBU+n8Rh2W1Fm+M
CzRL72jwCfgu9cGIZl2y0SDq+WmWeVBLlIH10cpSie12tJ4SriDzvb1YWRWMvhzg
l2P+1kjVA/yvj2VxDD9/CKuT1yDPoEHdHC7K7U6HsuWdX9B4wlSlgETuxB6kwjFx
mPmDKfrTRpJ30X0wSkXf2OAzPZ2WgGvxv6JPaW6YREJKpLsgJ1xL7f7wrgWHz3ka
VpaZ2EtOT+w6eqPRkebCAwVn6r9wz5B2cCuyv11lEVs9IhZ+B8o7CXMXOe4NQoQq
Upi/5CTjOS2CBpoqTisIF+5KKPaNlMsmx77wWL/Pg34Sy8L18pvRiFzmIxDNIzMS
zCwYLwEedBIhIcblb64vDYuVPYs7oevWRq2U7yv+Dzvk8ZU1LQ9dEkF+vPWkf2p4
4YEEYUH0fganoCJnNym+gasymhM9eSTUp4zSS/fOs69CmoNlXNtuMToDRSXJ3vI5
1asB99livyZKLjQjRefiUUIlHXzn9Uq1p2bf2bIXULU9SZg5nNOW5CORbMFuNLDp
Nb6sa/piKTcrCjWA2Z5nSamr3vRH29/SG7mWFYfGem8Bo0mMdxBGGe1Dgtcxds+4
KFqe2x3C3qlsb7hhf1GXv5lGkLFUq/iNtrq9L2a9aZf9H5Vze+jk1478n3CyZjaj
ZN+4JeICzRI0fFt1vmhjYZ9Z+veJgWKPWsM9oBHV+PrzUbOl92UH0Lxhi5iPhMQg
ywlJBEhd4wkXe5rsulyT5UE7Ct2U8FKc/cZgTGIge4PKhYU8Vw108kICdm93B0/B
1LV6mfUup/7Sm0TcMJ44FnGujn9E9H2pNGVZMyaSKNvwz6QS2xalo78ua4z/z4vC
uhjHuaJAmntNIRgdcQ91sNyfFpJLYreODcDSQ8hQmXIo6NfpGw62gA8a5LfCsf2e
X9U/9NWOaVH8LRv6W6VBBtSoBrK5QYzxdS8FYvVUC4jwK1FRkzbS3oj2N21ZeXe8
IR12aOdQYDGu8wd589gFu/aGYru/Nyqf4RrRjcF5J4fokTz6pM1uIKcUwtV2giAg
bJz2qeltsfQ0IXujQnTnWcs12xfdcS38ozrfusZxTXGyw6p1VYjeikvdlV3cgQnM
L78v7F+P3M4rK0SXKglu9JZ0/lSjV/vSoOnPhrYpk12NgUG5LY1TdgKlw86nqpqS
VWjVsFWrnzepPsyoLiXkbmhgVrfB81BCtfAPRqZJgQ1SzMJpxbQby4u4qRnFH29C
A4C/dNLtehXcggZMc8AaOToAzF1GYCmE+hesK+mHrUUvNmz94gxbqSPt1pbZZAjM
p3h8MNXkEmg0eMl380RWH9PEdl6I7vrVsLgGFTJrwjqkYDYCbkcLLPW6tpUm2NZM
gL+1BUKGOL0/I6OL9vQqhN2yyJT5zRj1Xm1XeidccDmD3RrihgtBe6H/yN6ipC6y
6k87ZGHQUbSL9a4u+fsmpZN9fPTKyQFKmeei6sw3V0HKq4gNrAEy0i276w/82ScG
o6aT2xDyAJT//9UDHxUuXrnmMK73AsPnnBpMa8okBYK+9ZKGbBPzy4BaOWsiJfSX
YgBFwwG3dfo+mzHFxRvvR2GEktr86jjg6h7yvJdLesl8nkPDietOiFUkSirqOW1x
CSRInj1uWEqwVDwopNe/8BaMCK/na88ZPa9sqQ1uvRvMpiS4yw9IkLI/xK1a+rzT
9QpiVUnKN8q+Rm60Eb6j85ENb/OFkQTEZyKqqqLDz0Vo0k6zCGrg8xoBFUy7w9BM
B9+wMiLRNOQ9/dNG7N0Lobhg/Sy9tYT1mV6byI0A6/pXj5DdBJJsJzkHtfsAt5EE
bH7XhGid+gv/pgM9w9Th1EvLXnvHwro1NJvp6ziM5GHJ6lTNh09mPH3wkxrdgknk
YTyIXxi3XWSgWLdVyYz/n2pWVK+ewzzH1yeKsjWPmY0/NvsBGQaMokXBTtxFUhka
Sieq/WXYwtEb1nMKUypUVLcg5vcNOrG54Ix//I5Ce9m1O0iGoKudhvME1gfJHdCU
lGImu/mAbKbbUN6OsyGs5ppcN4qA9laNNIG9TjbcuHAQQz/wEobYk1fP/2xyXh0B
LAPDzP464S0fst2lz4DZi4m7/gIN4/F7wQni0LdhxERpKoyRBOqmf0xuh2JeITtP
G6oSCDbTNszMbble74CCrbC3ifYqsGGn0e/hW30TCSrDfNcUU2nEAOCWFsFb6VzE
hPxAtN1WAPz/RfxK7285jGYpi0AGr2ggBak+pOcBpVYDhusRcf4ozW/5UhT7l+jm
CJ5AZXrHS/ElA30BFJvGV/0WAEeWHOIzTOdLtxdsxwkEy2wJAg82B5qnT+aRivSs
NX5Scj786v0s9REqlwO0zs/trUqUzsORtx6OM3VLBqEjxVsnwaRRMCw3sN22n+6r
c02dRCYUePFZWuHGIuSaX4T1ZU+fzPj3lRSsAoOs7jXCO5FDY4Dj/FfM1FwwaIE2
mIhypwoewtZ8hn0GBZH/bguuUTpJCCv6AFb0VP+7I5wxvPUOV8aPM06yQh/oahYH
BptBIatdq5z5flpYEN/R9GUKAgyNPHzAh3dvBJfI6/zEUQkuxffsMEUXDij2racj
ECoXxmDIcSGKKiksYxFRs7XrD1+aX723l9tXv+2IuVJ95HiW04p2b08WPIgYKm+r
+bXGPAh88+YxWETF16cp9lPxVyLlv2JhIpxAGphGpduHaX6Wg2+lR3XBrLaAvKsM
lGvUcIB9+9AVCamp1Vei1wr6oJPL8dX2v+6Etx+z43JkLhC4UTNDFvqX2/5Vd9SY
bwOfIbP3v+snNXSy8O5+l1pYk7T/xK4sThHOscO4+WzQv/eI2CmHJWyX7FJyPLYX
NzqJYEnMCRPw8OaDHoo62MBokO0cqEU5frlIvZuuLKV0mlME0ZgqxaOrEaZEBogj
1lYtkaJMTOMaVbVhlo85iy7uqkpxxUCgWibhTzz3hvre/ULKMnaE8UY7g/fZG1up
bX2JDREeLHwtCwcZ+Nw3hdvzP8iQf5r2kq8UC92m3YjgTrj0ttspSUdQVOjhzAxO
EXVq3xzgYvfODTZqJ0uFHOMfV+1+muWHg19Xus8Yj+V3ioRcBsocj2udOtMJSyr7
ZPGqCtCOmxsBgjpbpo5Dhzcl5UAW7Tj2htkMTDC8sKq21uBeCUzEF9gPkCQAO/Tp
H5/Zv4t7foIz7FVe5X4qW8Qv9uPd+oxPLQOG2ZVfgi2OGDiI6x8KAOSNSLB4NYI+
STrzaRpRRNJ5HoahJZi5D3shaZWnzu0BemNOyDtxxQg9pYO+/nL+hqINzbkBzjkW
9+Q+1gz7Ci1Lzwe6d7S9ptz7AJlAgeAqSVwM6Hbn+wnh1QBnaWdHTrySRwiNja3s
1zWnvuYSnh4zqkSg2pvBOHzjULlcll6xv6K3wFxnTQn9xr61egPIA0DFLOzL5Cmj
RaCfQ91k84DB2+HaJfBtaA==
`protect END_PROTECTED
