`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viKR+jqkFe+Jl0vqU56mwhkIKaFqECq31tksOreIJkiX8GbZdGCswRxUDMQLN0H+
7yGrvoyS7PX3hbKttSDi+LUCbxiLMCbeyWpZ/dXEeVa1qCPqae40xI8ywliXxev9
7MBommqWfhRBhsDn2ctqjVHAPNVG7/a6ZwFwEFTaPQHiwcvPATlKpAcJ1u3GuOF+
EN686qf9/bX4IdxyVHKkv/gEtsHaCARxz3V+ehWBDeFkoAHUDYm6jIB6QUzifur+
kyiTo5RN12ucIioiqMrQiEbvBzkm2+0TTKIE5w+f9unhqbMoTCwR79wzBrBZMJHa
5GhkH1v3BK1SiEJKL+hrAw==
`protect END_PROTECTED
