`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PtnQhood+7KFbqbezY3YBXE9/gaShweuUa1OJxrJfsets2TgULo/Kx+/sFIRaGjn
wSL+VHI8JV8Wbif3YcIDvl+nguQArN0rHPl+ixLyuLwqN/kBUS5FzWJAtzRX/OEm
xh7DghL4CkaESRq5MExy1R91DXPWX8ksl9OBHcWL7Mk16nNA4W+uGOBOWEilCS/R
12unhMeP588jE3uK0jXk6Tu1ZXCkcQyZIlbLJ/NJSNXV2mUHvL2huF/llA06inJa
X4U0zN6m1FSTqVqLho5nUUb1JS1c6jZOHEacViPjCwTRuegJOrOMBbsPS1EzGbtB
gA2fDSo91oabiz2IUhmH/+2CImOiSNO07B11WEQlaxHSqUA8IDKzMKpRNOuu8rp7
IPmCqnGE0AHYaHOTO88uKbhIiAzoTTXYbbxv7FGN+raZBuWaQDkS/0iiT7lj3gta
PEsvJZ4wP9DBrFAs0TPxmbsSqKcR1ZqbAFhxHQtyzQ22S4W+m9fMZc+mOIzDrm8J
QODOrb1dFHMR204WnTGCYPBB/5OSJ3IOfPJiwXYUU7P3C3FOShfGly+E2+GZBZmJ
MWeQZ+CItWWaQZHv5U0RWOBjqeEScNQKlwuyckLHSl+Wba62FVZaQ+7DydwGVqnM
jpGziMmWQpdCvtkQxw0iwqOAqxM4tTP42nhKjmMJxkdLA1q4UjknoG1ps8Uh/+j0
7BILGmXEzaYsWfuP1wGZox4MpqAtlmDkMbvE3a3dLZo=
`protect END_PROTECTED
