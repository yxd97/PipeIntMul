`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9ca8V1+zjiSZVXiPoJ4kpnVbkJIQHnMtWROlGCvRI2SS/p+Nq0cJllXdwiaRG/M
k1EK8vnZDghXdd5gVKdf2/9zigLyiAc1imZMe2Ej4vzBMUV/9L37ZtfbMmszirQK
PyUangb2ehXUco7TBfjap4lQHFX4pRhcpocgzZyJxmTisHE2serhQ4h/HWw4KgmQ
72GW6kzJSIRXTUZnJFbaQPDrN80aOR48IjFWe/o9hU8BIZtVscweyqYtUPLfvTwb
bZonEvOhI8yNbc7aTXOMXdYhMigi0c4TVSHHWE411M0cVU4xyMOkr9zPw2U8qgo4
dGYtC4pnjO6XrzH+ZSKZJWXSssySrqZguGQrFFw1f2AaSi2+HILDo2873EXvWAK3
ClpcNZLgyrsP+C8rghFfp7zPznfXNq5CyC0h062DH6262sg/qbYcH7kxLicntnY5
RzBG1Kb4mQjTM+Oo7XhFPG6Jx2sev83j5cRUWWb/2QoyJidDZksu3LzZgoDCF3zJ
SahDk6pxjSmP7EsnRsOS8tJ8s0vBqKdo8aTXz9mOxkg+LiuS0cm+uKlREuPlRe2d
wbtur+KgIA1vEimCTKS3niRd9bn1nEGF3CxZyVclt4RJVAAobwubgqTNagJtgic6
pMUw0KGrLukPBzlR+MP/XUzLsfOBGUToO6Ke7b/zbK4NO9CgPFoNpOuhCrtB8Gdz
D5n/zywpa8/Dhp/Vzm4tAZ48p7t+eTB5IUnbT+fTQzVZe2+Qg2NMowAbHXg69gfi
kQ2eQPWqc51owCcw8w61raLhh60VPD6DckW7jKQtGNtLgshuswG+tqeSXLBqX5IG
`protect END_PROTECTED
