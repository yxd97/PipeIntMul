`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrjE/arA1rThOPfQu7QLct+2qX+pJ2jxWMsGA1KF3xdvb1MHrR4V/L8RNlk+J1Ye
CGSvPEc32DRcohnjdIb4DNdMaXhK32dTqecnI1gdWlZLgf5Z2VS5diZ3Y8Nc1CLp
2u5VlRYtcII7P5z2B/4Sl/6I8aKZ8jzb7wuTkqVO8Pll1wjitKoQlmXG7IQeM6E5
wWmjknv3cWD+kiANaFYew1QIXMvclc6sJ3UDi6trCZkkruvAWmDZBHGHOjvitqKx
kRUHzIuaE6PNe6ABcckksDgV4ck23JcYhgS97fQYbckM7aEPoGN5+QlaeSLp+pO9
EcKWyTpfX291UH8ALezbhmUvtUrrVLVETumZAw0WnYLxyJJXFFOXGqS19yLoweX0
YUPtSJWRjYWV76vVrNO29yuapic2xXIr2FK9725lbNs=
`protect END_PROTECTED
