`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URKXcq4I6TvbfuFPHqo/vYg74dFemQOI/kS5MTStOi4nFzoWtA79SElUerR3eTw0
gHzjdarnv7OZwqkSznes9HbWkimlMaO38hYBkX1yPmx+ID9C3PmAKLrLGRGJ1YgV
or6VVpLNLvoIaUkgbzVF9yINZiXrUyYHG4OhYaatYPCVjQ6NdknkmUcxMHCp5Qri
qZtb5jie5B9ozwzKHSc1b6MXmRYRDP8WYdhgF5PD8z4raVbKrmDiCJPdUgcm3UbX
kzi1V4qYJdxz0ye34m4YmrLf+AIBIBlNOhAOIvH5XP9wNbQfWh0LbK4qSgpgxz2S
xsz37S+TFw5S2j+wUijKTyxiaKO+M5kpJJVsgGXVEEu+7iuUSrtl7DlLQIAk+KhT
cOK0tze5pPXLtCbxrDVXDner5QicwwBJV9MH3kGSyv0wR5APD0HXYshBmBUDdtDN
YjjmUljfIPV/sEddmuw6JrZNt+2cneHBGX6+HplNVo6nxZX4auBSJMOgeb+sJCWL
yJuO4hycp+JS4BP164N76QgWzG27xlR6Fr5qFhMPuQ/y/uy544gGWzz/X6PUT6KO
YoacJo/e5OjBeMF09o0h2pwwQIkTIHCGdhegONO82Kc=
`protect END_PROTECTED
