`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+x6Icxjx+E2VG9wjClgsu68SQa5WuQ/f9bt83/6R6T3UVNqP3clpS1CycWWW2Tz
oMCZziaTN0uq5mJRQdb2VSamLApYxsssX/HnWOO8zkBq/XCR83g5yN/nh6cX3FMD
ImVggTyUHdrSXThfeO9k2SzNzAAInwL76Vuj545c3xAdY6xAN6voaLyLExq7p294
tYG1wzlVfKWOpuGHGsKPHIjRJnUfOkqZ0uy124tPZfvfjxL86dMF5X/4QR5KANsz
wTmY1Dlu3bP5+cKz5WYdCgVvIYEQBOAwM0wtZ636jkjE+ROHAbwPQgm4Kt2GLInj
UAHR1Do5GvPer5zGg00tH05Uqt5oMwl+ZapuB3+Ne+wA/JmYJu2q/J/cpJJyvbv/
GNtICttnvm6m/Dfjl0i91oiEAZxaLJFleavG1uxsKyW1EOwZf7hXUsPO6ouSrAkQ
r2Olaf/giM0u1Iar6FOsOvcU8Grd+1t7Hg8En7csoByaGHnOLndg3Ttgxkydf0q8
6xKM4AeIxE+vnIMLnww54CVDX2K0ie2EJDynRadTLUQ+shsv+hw4twPTByjqVpM3
BNUIxhMX1e0YdxnalUmTLjv0xWgk1R6Hh/OQfy6lyMoAXU1PlpBpHZZpFDbvEdaj
8wqZ27njh5XfkXv2EoQLvAYBuaJSD9hpNMr+8F4odSG/3NTHXXUOgyKRoWXbJQvo
y2MgUf+IvdvAshu0vhT/sElfnnL7DCLtnvifbRj7MvMHjxTSZK//gQFlbE2voIH8
I8VfzfLsuxAobEtH0fJ20aQgpGy5mOuFS/ZEgQTgHMNWEOSeP8BoYXXzl4rKkpQt
DL14NC5Gts/eFtKq/C4w3+Vd3+DuHUlCWbjtTiAYa2E5mnt5nBI5t75qbTC7iTqE
YiSfdlCQiRqvC87pi/s/ZX8VDNMDmrCisYRuY2apw13AtaayTLUIN7uAVK/JUVCL
`protect END_PROTECTED
