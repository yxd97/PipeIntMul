`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1y1yE6FOBp3jdv6PvfCA7j/yTtBnbMTxhKH5gzOHnOJPLuR//NuZ25nJrAuSID0x
0pvSHhFOHyaTGUrcxgx0PAqmHYtCF480Y6WiY40OgCd3pnN7SwXE+PIn1j0IvF6a
xK8Vdt1gH2ROvLryg7H2epwtVsDNddF7srJ1WWje2St7a/bHsb7+k4kUvkc1J7/N
TMnkvAzz9bG3LocwzktnXfdvF4tB2RPWOhuUyhjb1Pm7m1pT0LTHaXdj+GsAO3n4
8bs2Tni6CN5lpcfDo7kUU2Q8ek1evYWk1jhFdw0MFbmpFVGiePZVIEdqX/LhCXVV
ONmnL5wA24fvt73fja4vFQ==
`protect END_PROTECTED
