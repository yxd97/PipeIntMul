`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X8n40mPYL9tCW7U+1kjq/fVCz4BjH/crruZIDmX0yJYiDBhb31eO+1/Pun4lS5Cj
uvNcf/EnLl2QMqT+I+bwDdpz7CzvZnzs5JuDjACCY5PytbQDSzOn9RZehgRznhsl
DbtDTqVWbI82QKKXxYcOcDUpk48jRuN7cIfKljsLlq9QSZxx0POO7LwRFdoPM2+Y
BBXI3Blk7w0B7Z6EV5NSYmER2uQo56mpfwF1NNohrSNEV1+jCK1s+KC2XMJ2hOGv
qGOyf5a+ol90ScA/i5TFM+xC5RivWB8cj+bKT6aU1ij/PmPEh2RwehMQVJrntezf
rU/2Q0Uy+/7teIZKroM5nA==
`protect END_PROTECTED
