`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UvVgHeXmmcOxoo9+sRsQVPh6LnlWNylChfRTLDdydJWqQSJsMh+WorSEglM2i0+g
er0JWpXxFMKHTauDnf9onr/4mQ7LxJ5B6TVa3kuBkwL098BjLP0rI2ATkR6rFDkR
jRrY9vEemBpIyG3hek7DpfO6UD4cGIGEjRdV0FF6sAEQESIOXyIYFEEMFZmg4409
mbpLBYoL7H9sMsNQA/QcO5wNZMOouknvb8dgowRs6NGZyOkvTuCHbeGqVRhAFXmv
b58oTFEg4Law/v2wFbMEFg5Zul4AOfRo1H6wv3ud4wb9jD4JmfjgCyPj0ts76KgH
wO1vlxUcBxnb2OR1qZUunzDquomXItuGEcbUGWpIxaQJRW0svBV2tX1k0pbFHz0z
yzRIJ5DhjoLTpKK3wEeCI9/33cQ6xsR7AXMKer7nKtY3m5CJVj/4Zi49ZnAlQ+SJ
gN6wOleDFfUCw6lqq85e0XFHx1Pq52HSXTkBM+XLY8ULjwWt0r8lzzjZ8+9O8PBn
JRfHXLcFe1O4zrpDyIsqWI774yMbMrpYm9qmTyxz/oxwuKVOAY7IU0NT0Cnb1yWI
EB9o59KixhvvhEWNmb2DZbnreBDp19Fv1sXriRbqRyB4uoSsq6tKvEsD4D89juQ8
7IzK0PoCppV4h9iXdQXte/I4rOBwhU9sn55EQMQaXuXQglxdgdcFrU9kH7I90/uC
t3NleNDJuZostKzJmDvc30b1ON0FCdM4YYeivIKi/U6m3SJdq/7Z6xzz6vFsWZ5r
noh4h4vQYvb1o/F2PPlg8viis1an87SRKCYpKaGuG10bFcjXPkQIPxvJBh5NGwKb
zgsKN3lQIZo8r8xXDTxv3NvOVMRLxeDsRWTZpoGgJqt0hckRdbvQ2cTf4vv8U0hH
TFEQatJoAlhkRqOAdiJ8nlM5AlUNwdbbMAGlJlpCxR0VkoEYoJOxXN7yw9gCRKB7
+i2PMRlCX6fREYEFiYkNv6SbPlAe0oXq9x+jlIvmdHlo16MgPkoRyvUwV7Xm5oSD
sO2Xym24/vokT0cngEwfxVAfyV/v+GEBiTSPnt0aXEsqXoJXH3BNsYdkerbBeB29
PLH0VqYFz5BvxmgAu9SZc2QfwhArgzCspP+xQm0oXLndUbIWvjVabP61od0z6Yq5
Sbwf9mHKbsHIL6aPOwNQmoym5mACUWNkX23GLCxDA05lS//QzvgmI9rAejSLlQ+G
WxH0CzdqQqO2QJB1an5zHs32qZQWd0d0QZhp9sUmZ+jbj6iTjpwNR5RjRaQsklne
+BgHUleVURDEDwK/Ab4vNdiotLt4UvtU5+GM2iz0w1Y7hjal1S979q1DEQFSUCU8
`protect END_PROTECTED
