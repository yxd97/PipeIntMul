`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cjjmpXxzPBo/KOBsYdu/AB6EefSrCMVsTE7+f1qls+CYq7BXG6D3QpayHdmnk729
IPcDEqLrYHu1sZabHT5Boh0iD6qsJe0L1O/dDySLRxWR0oYxbOaoNM80VZ60Aw3+
F3LVVp43meaCuwz/ixZ0+VTRpup6JhZq+exFqkQKT4FkZ8OY4jr0CNIP4EJHp2qm
6/2imHwHdrUL2dWHekYQkpBPr9mnP/SzMu7wDi1Xta8wixv5arRI90RW0PYzIpZ/
Gm4gxHPkEaXS93Gb4PgniSWdZgI2zUyQ/tJySqxBmppf5SprQ0UzJZGr20gnhCzK
QJH7+TLtHRivg2r1qcezMx+CPyaG1WL45NNHjAqqgXl4FvJRrmYbepNmQ7e5Sq6k
5ii0W7tVtMvTLipYFJq6QFT2XJb0evt8Yx8Ath6s2yw=
`protect END_PROTECTED
