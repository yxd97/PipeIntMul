`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/REfGGcA7FgDWAcSjCYSK9Zs9e+OFj7W7TjmZO548l+DeE0dp2nSvEKGSGYu0NBb
AK45hilJXNSTxwz/X+FGlUwHeuRd1nzV22zMpmGTyWLlVPuiUdKID/YB7EfV2sVy
YcDqH5dKe2bbbAsNR44dqJoGXfGp8sGTB68csK2WPWzxBMvfEwNt6S21zq/Cngow
LeM47dU6vItKPImB7ceUFvNTeqDg90EiAFEG+2yHULFr+4I1nCYoPQ/DgiGCuI4C
rJsR4Psblvkccs/hWkPMIKzcjkCMlkXa/sDSNE/Hg4NZb3y3B2pA8xAf+hT6u8U2
/+gGEld0iuXxfwaoHDCsa6yqcXxKz5Y8UjeaZNrs3zUHoYBDohtgXCKlE7QLhC7w
Gr4SO28nA3SXuGo2WxRTvmE60ZL4T8Fpl1kvMKuifC/m+ejBU/mnqBMShfiUGeER
hzkNPUy722HG1HXRkX0QUOPm+33rlU2KeNG3bgRdlYj5HcDE0P5Pwj6NQuV0lz6S
4ScGbLP7gYxOmcwnEhhcRcZdXP2+PM3XaIl51S3nA4iKTVh0LFJYnLv3mKfBQkPW
UQEfYBBpeg9R5qb8gI1RIrhxOQ8ZmmjC77vXZYnvA7YZjmLsdYJS+96XaWVjHCx0
d+c5xWMt5YZNYN52bLDOYSBTfTRPHl3lD3B96fTpB7CFnaBTjHp24XN8lyoPICtl
kpF90KApWncoFu/2bq7vJhjCKCBZC3/MH41F61CUa8mKBOQ4iQorc5ILBC5PZsU5
7Q7F9Ug2V59f5K9NlCSE+l2ohK2e3TSo72EmgHHBAr6rrasQvqGZc/rQxeqTPcy5
zeWrNNWM4Hrfu1EoxG3/kcpQaHijAtVnZIFVK9fmT8OvF9I3kxNDOlVs3CW/gN8J
iuYjE/1s77spYOVG6tqjSAfC4P9De3lt2kGXt2amZtR4QNBx5EafDHXzMPCNWEJF
W4LsmhpPHc4fcfXlDTkJ03eWLPdMN2o6D7l0G7JEDgr5WCwiyv+b6cY3Is8RGRmd
gO9enQGf+0sB8hTaQyNa2/+rYXdXbx70ZVigKjO6OBltldggHpKHEXRC9/35R6xs
ZL5IlHEhJoI4EgJ0vjp6D+qs7Ahd5jKXzUmNa0qsg260zEwoCGMtDyr0j9sJl3ix
c3eDsQ7xwW/FhtcGVaey+Wh6B4JX9FbUs0WBA6RBTsWLrhmK7lMoKT9Us6xGdijS
hnNKojhpv0G9lKO2tNG2XTeszy6Iwm3S6VJu750Vv4jAEVac3AuoXJYAh3n1FhdY
/wuVWru3a7kabMojeng6+tfNAyrU6oUjpXvW01rIKJ4GlCpjlqsVNVry69jqTrD0
KQgOnq7C7fPh2mvC6GBWrc6MfdCor2932wLNWQB6ZbsS3+clIQsL8qN5UFtNR0mE
DWAhiSicVkJYuySWFyroKfcqQidmQIzOXdqXNFnpxKaq/Wf62mMIw0bFTSu5+YKH
7om0ZE15KDlgc4H6vmO+lBHZvdhZJCGW4mXgSdHfvaMGp9+yABjdezC9afg9Ev9y
zUZ2ymDML6ulE/QhLqVkq+ysLk3qO44MpLXe0u4n+gIQnkSuri6PAJZ6eWiSlxJO
syPekqQmwjdLqMJDXtHo+Esilyl5qaAKNxb9tINc6P+k4jN1G4hy+OnbjX7MySR0
Jlpf1KaM6RsXW5fSBv3LFU5OZVwFPAyprY1VHqYWk7604YaQ+Q/kv1hBLPUlthR+
uBRvr+pOuX2gCeSZuUWK4pg0SFggWxw8Ls9POGL4W4stSY3iPbUa1JLT6FSmC37P
cLRjP6Q2skvlEJJYpdHZlUggH9z7PdZNxenpyaxjEBf8Mfs1H3phYgXTbD1+q863
7E9lim2BMvWd/G0ZjNhllzYopGu9orXkcJAfh0vC8s3O9FHWr+7jcx8qCxAksbS4
cXOFmRVOQ4VfZQCvwAZTbW0GJi4eGhoDzu9G9cgku4hlA8vKkPlOAh4lwU9DJx/j
teRYq51pOZ8Bv0SO34QwU8raR8b0RqXpW+AvpUwj9An8Goo96HyhOWoCxW0d4FCW
RJLAkYJNJTqlzq0YmuhUE4x3rtIzQqXtMnwrNWt1nXVxqELPWn4qdPIGUH4g2tWo
NQjhpPAPLnB/2SMcBx2xKBwzEAMVSWwQxFdWoG7PkRiQiMgYAPz1mua482y5uvKo
tM+tJOV/sfKksngBlj/6aw9rjcpVaG7B1Di11mZrTDaLdgYgbTwOC1rNPFfGnM0y
O4tjtB+lmCGLZE5ohjxzAu23iDMdbsbuO5clVLIkJ4356VNURMvqN9IpQztjsGbi
DN7kNM9HwQHBRYaKFY/9RnMTH1sqfNVih14kRRnnjg5ZQtbYmimtI/8KPOsh0tdz
fl5I0ApOyawQ7QLZYwgllPS1V2UqKEe1zW4JshNXfY4IHJWrMhgjVLbtdsAmK3d1
rvtnUS0MtbdvYskxiLOn2/kVyEb5RPretESuwzHu9mMImCzsHh27DTTLjWEGS86/
1JWQJa5NJwSUnydx5788TvkNe3NTZPXnvaIgXJBpNlj1T9ryitrikCB3rzY+s9XC
LnnI72AHf76G1W4dQNgExK919Wjftrx29j9CcZWtdNnXIadGKaAijUiVPBreFw2i
wlfasCh/TC5A6bdqG7nyd5C2OpliI7u6+kH7PdIE/CamDMoYIinN1FE/qcYpOenf
V7k7YwrqxwF6X2dRANhnpimaNRJHdcgSA99YaG9D/yTnaZN5W7kmYorP84J0W1b+
A3J8IN6p5+W21Q/LkZZvr/b6dGBCLSc0YBIhT7fRpN3V8M8K8WHi2juJZPDCppmn
PCvWgnWKYh5j2vSgJVQWZuKNIrTL/u2u3wuF/TML9z43Jyar1cbYGQ+Gv3qeDhQp
yRLMnILBGF1G49SKmQvdhwjfpBCcAEqMcbWLnTcyJI8ndNSxNx/7YnZGMCYFlsm6
zsqMwfgG+Bt3vzfHkbpHU9MEfweevjvZiq8Wv9UhozUqkRlsam/0ca40rnWpUqsn
jMOQbWYpzXJyvdDvYfrmKI3DXNn7uXFNCNkSyPogR7v1+NZJRza+gS5YKo3tDLfv
zws/8vG/Ehee1ugDVvjRHzQsQLx7o35ETYsrVIphO/h1uzco1dM4w3lTeW6TzsYl
KhREWYLfZknAe2gXkIPQjEx6ZTFKALd0ha4yK8rZ8zwcAAL2BK5mymb2Pt3KHS8D
xb/acn+i9j2ZBvhAAP8CP1Dx1/7DsvBuPwteOa1RFtx7rrGIeOiBkV7cUKA51Gxt
+2gmn/ttgIcQds0lo+D3R0ZSrrohSQYKFY6Lu5rYreWijHjLyzeev5PG/0s7+gHk
ocL8UaZ0F49tIkxaIOg9fFiWeokV21LwMwpIF1LrrHD2e7sLr1pD4GUmdNDGGX+F
IlGFYFG0rTMcjUxJW2aDL189MBuUtmKje++fKYnfT8gseE70KH0h1n0/T12kdLZ7
0gUsN4BdUDC7geT4mNto654V1ekgx1l6j7bRrDlL4XmBgEq/Zq/kvxXyYuf5yBvc
qcyXTDiWOSDV8ykHGGuKDg5s/wEm5Wd44etGfJDcrxWZUS86VQmIaHsPib1irvTs
bu/IE7Tzah37Hdff/H9gdRix8TKUIxcuZwQ9t7j1lSVnjxyVzQXKRkz7PWagm7w+
SF3l2+XfFoWShEF6nT2BBzunZk7I/Umte0atzY+MPravCogznWVUKEzyif/GvzDJ
bt8vfz2IKpvE1x7Vziek/FRhHHHALbHfdTEJMCXavmOVLuCw2dwg8JuxtMCalaQF
uqF3GklIyUfPy6rz0GFpaq9f/P7t3dz0FYQ6gf3jP3Gv/cM7ebS3BFrUSWyAoxsn
JjXzQoX9kj+ZtD5BhtaipZTjKaYVt/KBBp/k9Zq+qxNWHdBtNI+H6QazhFzXJ4xm
Jg8kr/mMggkV9nKADW6sJAFFyxN3quUwRrNJCqFnEUTPWYdKJ+tNDNng5O7nAR0a
Gh0LWBab9Ab4h9AOczyy/O/a0X85f3vxewBs0OdcFap9sLY0W4EgZ9UBDgarCaYY
2UWUgNqXwj/hYHwxuPZUH80zFIIQs5fNG/75GjgQEO0OA9Q0g6kOBeDaPaHtqrJX
aS/LzAXpJnF9H5c9c/9BkNtnGUdKPdnNgt87WFxVwNejzV9z9S918k7Ew019mIiq
QB8lCcbkwgRaqaIXrd67rcBvfR2dB2ra3MnK6bPfqeCweFz4ORAcwGztUnrT9VdN
CGR16WijI9mAUkjsja8X9hKtZ9vj/hnJ/Auucpj7UYE1CV59w8giVGpKvjG6Xns7
Vlyq5aK3qe1UQ7M29Z5l1Odk/205hhgM4tBVgyB7jbJetf4lqOagb59R+eyPfCZ6
Ao+VATDpylKuKQ+SkpmIZUR3mfvi03hHMGXDXIbwi2ygeGTQPpdVAs6F0nD9IWIF
Ad4iXmvZ41QahfVKztH0V+DoayLdOAaRf7vfn6ybDaT9bSE0jJe1f9h10ENESgzY
0FTYAbM6FigZegTGxdWSqtFMl20xGny6xqpeeq+kFpLPCp6vY893kdy1PFp1yr8N
yt/3C6Fhqf35NRr4qFnMmfD8vEXjtX+s/EMWftiHAT6Z3RGEoLoLiFE3fZ6Hr6HU
WcdRwEEJB73Da4EiUhQZhFQoC9lVsM10iNeBSs5KlwMUvc1cbF63s98i5RVciHGy
IHpHw7CEjyH1GrIqixnfAtuAOubWdzkDYkuhOAfpZlQiq1imO29wTunFqHJoPQl8
a9M5x7rqDBnBnpS1EsO7yF4Mo3St+ylZMrro1tTx3732HXLhT1frI4TCFcilkK7X
8BmC7edIVkH5ArP13r7arS2ZJMLnM/aZKj0LMoouGGBw/jwHnbVrkPFg5Gz5fHTG
UTum0PAALwkT76PDIpicr2KBIqydJxRsCpcWdg4X/73cOhdCBrYxPEsdYygFXiSc
8zJI7upi4r3TBBLje3cgf8mttt/p9gCLZVkayzlovILhxZtdbaaheshEPQqua0Rb
GSM7SXNjdUWMy3KBe52Xnmk2+Txh9SlUx8H4frY3dYh0A8hno7VJOCZl1Pvpsy3/
reOxsp/+bKD8/YQ3obQJC5Lf7QADeVPRe1KZY/fEiCc9NYXj4CzNQ6XFguQpuoAm
1DICbEi52RPiY87rsYGizbPlwIIqIltSSvzVZK3hIxb8yM/gqJPa9wxp1BTE7nrW
agpg/tiNa7kl1O+K6+C8K877W5C8WC2Yr/4vucdjPVHmSnzNKwsrGKypVU3v8IiR
YBS1DVUvaJnu7/WipRXjIP9sGCQ4OT2nCgs6aV/hBcT9cvEqQu3XazjK+QU+9Hw1
Qto+iYvElHT2XUUabHJhVBrTkoMPWSUxddTIUzGR7ByuoFvlKiXpPUaFlJ/RziFJ
HhZ5KBEeGp7yMPIIBv50n7ddybCvVaCfoQB6oOZKBR5ZX85NRgV7ltJGCZ5Jaoas
mwEVIFhhDXKJAWOWHXfcnMt3FS15NHCVLgdSrSK56oUE/eGYcsL57OKosdxwHscy
0+MMbXahQzsE9U7BuXSpYIP5jKrbdk2DcHm9jaCp03/qOBlzbacwiw9V0DSYrqAJ
BYUCZVom+jPcyU1kraSZGei6EhvRvmL0YTaigezboSOaZb88PLYeXcF1/TjDGkF+
4bdSQD88hWrshU6fFZGKUMGo3y8IS8vptZAopLmOxFxtuOy5HhVq98DRyoIa8jDp
`protect END_PROTECTED
