`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXFkNO9xI+vudmNaV/dOxwxu5xUH/KcNZ/vg2TKTk5K3UTrN+B3Dg5BYfnjh+Od5
zbqMXTAtxHBzOJrKC1sllfi2PvlHWf5cRqsKnUGNt1t9e8B5hFonaqbhlXFpr4wT
LpWu1i4YGM7eVYo9J5LrfnZlwHD0OGqvbGktxMCBYsEMPRYAP8Wh9uGEMobHSJD6
NSKBS20P5/cJhTdt3Vk/k+jjV6vhMXUm+N6IrFHtaAVujxXygOAm+k9LhAr7R3yB
6iowAvLuA96uOI7udOQzIOukrBLJqi03CkF0ySms1itMT0BNsaLtzgNiCQlwFBdr
/o1LkwRUceA3Vfx/3mo+hJEbBv7EMJ9hioqhR9rR2JObS1tDZKP/s+yWPJx9NuKC
zwQmKLS9wLWazZP83OpwTEWZ2yQAXsOZKU5cIswIIlMys7qD3aWnwm/uFa+PBQMh
7e2SOBucrKkgrkohXxRZk1/SoQabrEKmUo7ACRw48bv2fXCmuNgBHvI+WaL0YKSC
bBeSgstwpOKNdR5B+iwTbvUI58yeamv7uBjEU38olefxCKbfHhQo7FtbJxUwEmop
xvIsL++DspzIaPuRt6L9GYpUOGmYLkdIpc7StHVzSwQ=
`protect END_PROTECTED
