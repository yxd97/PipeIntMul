`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJVmlf/A656sP5UpI4K3Yh6pJIyvYczbN10nYHajX41xDJ/zi7Dgv+pJNRVjcGLj
Ft4bKkk25bb4rbxTMBfU3cSKV3kSSDBeC9HdmVmiZFhnGEc1moA6mGkrwedK5jan
LmJzNX4Y2jAInS7PJ2O378HBB1zEEiJX5g0TWCAF9OfgyXkgO47msuo0ouqjrIpV
fV/JyvtWFC9sj1djmqd+rRgrHM1ew+qB1+qkxTkxrFNHMkl7HkVB9t1+awbZY+Y7
hzSINROe6AAj9R78W23gW3QGeElXmf5rdMZ6HXdEpR/GNVseSMKtvqbTO2IX0BI4
RpHPQxV0DHwcJpdEfldOY3HQ+as8XSDbQ8sFu2wta/6iAzYRBpbgWrdDic4QxP1z
ggUfqtb87s/lq6wRiL2eARTAWn62ToVk67MB5gy78G4=
`protect END_PROTECTED
