`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxs9/zJ/iBl0u2r63Y/3Blgxsf5E/x3leAJxkAQFZC7fq/gFbs2X2psbh8vV9VwN
I365G8QLrI1Ne97RS5xONbuLvn2E322fcVG7o4SA/8vtN4g1EJZplbLpfluLHahf
ZaoDK6Vguz+FzUBoDipAl/yxx8DgJZKRFXDfKVwVPWjG4I4QxCYS9Yf7x0WzumKP
7PFyhVFXZC8Hkh/54ljsghsenzBDEfL1uQwWyu5CffHUF7KriiPiGTtfo+OK9ETG
kI3arh18Pv0l71xRtyw8dB3QRszEMLpWnV/Wj0gaUn7xCeF8aRAKUowGw9yY+7hs
7LNVKCOVTq5KZeEnQJI3TJrUdQeJ68XXeUvQpPbPATxY9R5kLf+UfFpWoY7Mz2Nd
Nor/g+OX1nAxpW3GjWGmZ0HH4L63jQQH8Ypfd3i+Ja4vyoF+NT0bsTGR/zMo4iF5
TOJxnSY1v5cO041oyGPebNZF72AdLPHJlqwsqYfP4+dR5zhrOy1/Fc/prxNbv4qm
`protect END_PROTECTED
