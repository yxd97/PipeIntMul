library verilog;
use verilog.vl_types.all;
entity x_dcm_sp_clock_divide_by_2 is
    port(
        clock           : in     vl_logic;
        clock_type      : in     vl_logic;
        clock_out       : out    vl_logic;
        rst             : in     vl_logic
    );
end x_dcm_sp_clock_divide_by_2;
