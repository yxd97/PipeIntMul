`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+JkwC89x1DIcexq15sIQOWWBpPP9vP2C/2X5eEC0Tu3TOKLHu8dlrg8wk2aIgwt
taKTm4dXEiCIYHNtIIC5t4brNEgltlTUzPHgJT5fXTapQDYElQRZMN53BOVLRSBv
wGdgzetGB/ycegtm8cQ0Sqo6WZUSEs2/CjAGHS2p+Y43AE3wDcb1n3SeN/wnIjLO
cHFjbUy085DAme70rCGeGi8f2EoKLrSIhIOx8iC/mPZ7BPM2pGEHF+1Tg5WmBXCS
9BHLG4Un5aeufHOQykUTJD/7mCNHSth5zW+Xb8wqqO+QtjOvuCpYRK6X1/txhvcI
0RPUx7SS0yxCv1CouECc5LZYD7cecVcWLfNiIVYFI+Mrqhcd+2TsEng4xlODzF4d
7MSAtaKm59QpE7gY1siphFy5BshoeHYEdSeqN31e06kw+scR68ckJtUY6FDWdX6r
plg7yC540qpPPPLjVQKjjIDGbOloK2YANGdVNxu1cZ2FOrOfKlWWY1aGB+WCYv6t
+SuHq55LxiBZtzecFBr/tsERWCyF87Vs1fuJa5tyaLpRsw0K4W8xmVhnjipTo9fv
rW++GkWe35k/QBeQr7ZlkjWN+pOLeW+QDP6KrINwNhB3sjvcMdRkdaOo+Dc8x5FN
H+NDWleBuRHVdPuDUgW3r+swdvxrNs+ASwVyj0lY0V4=
`protect END_PROTECTED
