`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdDKLTS+MOQLIZrHucclqb33cKjO8TTdhZwI/C9s0XoZp4z69U5ahjlPXbvI994z
zJbF/yiYzjsKPihSZLkvOB/Ask9V9DEVjbKsoTVqp1YBU57sTl2FMoAKi2IsYwl5
b5ss/lg+kKSSSHUm23/Wex0K1oUssKA4EQv1XKjTxFc7cnn3DN3OqdVt2yMZqF8i
dYeQyI8tSAegQnmNrlKCA95PEniF7YEIyJ44Ber9GArMcXiAX4ptUbibKVYrh44x
kwoL4VuAF52LKbU3TFLyFJk+gATfT+BKjbzLJ+4o/5OICjLaRmVVLVLZt9YTd6/K
xFbL9M0pg9pFVtZYm1pFt3K92EKm5nmagzUaHxXe8NCV76MLpcgeG57cLPuB9YIt
Gla6/GhWSmr1rTLJUNehQtwoi9jEiuVFXUWecHtOKfI=
`protect END_PROTECTED
