`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vUIwJrJr88PipRbna73BnOT8zey3ziH7wq984cja09bGAl34I0+50OkYlG+cdy1A
PKdt9MVmlOb54t0tSOnm7k3XnziiHn36Jc//nZWDmfuU+RxYk0UuwGqsu5hoHsfq
f/pU+X93bkO60/qgKXZ5xZUXGXMXpQYveoPKNkKgNPjTn8h30wK/mcvFQS4VFpiX
oZy9zIKVbnzJONWDk/zeSJwKk0h4dqyV+ij4e+XmNsKL4olV70VB+uXf9tH5ooka
K+PEvaMI3VwDM5oi1NYao5j/8Z82rlP/7X2qYz/dSW38gX9+a8YKF+1uhAoRtlTm
IXDqxwHJIhEwJ06/dJ9F36pqsNVromxZGCOZxGcvlpSgBw67USI2OaddvLHk61bQ
seJUXzztnA2pT+jP2KHOAwlYh6HHxXwOr11FqvruM0lq4qJXU5H4uLexqkklNMLn
5GrXNl6vKjCpwknweAi0Sriako79B46tthNHqAjBi17Czw4l1Lov8PFL+d3pydLf
WvGexlQDOPXFysHALnmUfYDeohUcaWUmjJhojxcQY1P05ymg31ZAtgV7Gr9MUUlF
S6gFwf6pw+loNpkNwoAPxCDfsI6xe1WYF7qmXAK2Ohw0215yqFgZQeGfiF77hNEc
jJJpIxaJSa287jEC7mJ7x9hMeG+LBV54YwOT8JOfHGPORlEOlb3rY1q+/yeHyi36
OES3fTSbfsW9uES3Wwe3TdJIWmsMw5rqA9oVPA4ss/FwvToeJOtDwjadr2y44Bh5
pXF2Yd3cdfuMdNrFQeKqMt5wlyHsSufHL2No0mPwMAlcFSIqE2DRuAiYLyHkxBs4
iGxLSx0tLchD40e2qD9oB2k4VnIoCc/L60XIUk70rTDFOnLykAbSc3LGs0vKTfSy
DbLDf2Yq3ZlM1MLfyaiNkH7UyP90MyxuN0alSxSRZDL0IR7DUYOejS31uv3VaRjI
eM3vkzmOIqLGohj8BnEokVSbS20Wc2WpoQi/Ee/Ca+5HE7zKe8J4dRO7weht6Nci
O0Bb3TS2gVf7x4kSz+gUQb2gIihutblaXT7q38pTQ7CnKF3sqCh/4D7Fi6AevJzw
WI9w3EroWUOYvFvmGtAss6uWxu4l3zl5II/2V5Hw3HfuIeYnAlhE6TROOS7KfBTK
X+Ife36pjSVOd9UM7TAKYwbSXaNKQ/0Z2qv0hOIf+1H5Wi3dkyBXF21ere2+KLVk
HYFNo9ehxuw0/Tz7JAaUiakZqBeyhXu+wdnpi3pvu7jNTEY/YF8h9RoVCr4IrLBo
ZprqYZiM9bZK3CCS4Xr2+g7VOveSTFReIHyzfTQ2H3uaMKaZjHaZMZLwQLmgZyTO
I9KX8cz1YZdsJHhWaJijS3YzBfnaLpkcztawXeb48XmsI7/k0FD9b2vZWMP5/N2W
O+9eYNkkgqHuYOwn59PY/Pl5LnDJpTYflOaPZtrKCOFIar0Y5qR9KmxHwnw8IZ8M
PpXql79m9gXuIcSaqOh8SfV8fJ825Jlg/pzRBLyW4zkXGbjQw2ON1TGen/o+AD75
eBCdkIh4oqbwvfnVsRVh8hxtQL4IYSTcY8K1R8c6c/gKeedn8Xf9fq5DUqrhQOFI
5KOT6uiglKYK8gjE8pDDPmHBZOhhNz7CwlsHhhCQCV4nb0hIgEF55aU8ui5ajouG
YRDiQ057oodwpbDybrkz9klpHHPl+734vghCOqs4YGumCNvO63PFeR4TGcuRd5MC
1NFXJWgkDrHYXdKMhplOU7QqOgwRKaFQxSt8avX/VDf88FCsXeiHjJB0X81VBSJN
ximBE4PEk2POvpGgWhD1T8NqWIKucq+shu00urgwkQTBjmEFZVC5z4EvjbUmME2N
B9WrZrMOZvH4kpUkDEEeVU82YEHGL8j+0Nbze00eH/HZSDgaBm5K1QJzNnT9yatR
gC3Aho1aEphR4NDteBK/VWSLU6WcEILfKoaovFH65tnTDAe4fKq8VHzQUo9hZ+G8
7w0errUkfPzHSma8ZRXCido6iWFdbsETBsEf4YIncb9j1kaXpUYksrCQdDxbggeF
OJgd55Zgkv6nWTBoGoIPDOLgidPVsR2GxXwCHGPRWD8d65H940GfeyfWn/ju7r/h
secNhHYxDRaSb/xtI9AgCeaYL6kT+7RZFimQ4L0fPZrB1b0tGUi6Mh/cQO1chSIl
DYaHq+kyV541tLdq4EEUFeSju6k5NNk1VZU4y9mnggbtcR8k0SzVCfJAV6cfWUwu
+xdDE965D3yPhJnXEk+HsDyQo2zzpJFKA473JNegGbnVn10BsksflyhDeSWqNcB2
9rlHP6hv1jIKFQY2r76xW3HsK4AWeLpnSuB0wZz5XVbGKitXTlTZlg1xzGXYg3UW
4VX+SYdEvQ6reLP5e35Z7DDP69sUVtCdtE/vlAliwpSinWpXbdCPQmC3kcpzg0L5
1Jn4DLCbD3UrN06xuRP1o++AqDnIjNyTJJ2wxgX0mm851XDd5XOYJbzjw3qJKqWU
6srS/jCb7Dzr+b97CLhj/oTrMIlLzIP54bmRJ0+77cUEmQXvtq1XlNesnZJ+LN4k
FTayk6GaQgELoVQuTugQfsXN3WlDCOzx8dSX1gTf44DaEHd392oV+YSsuPXDw2yv
HlQARmmQyb3EFIMR9XEXII4wsy7JV+FauJeiAkw9SBRQaG03UxUVfec0u+1hiezu
hLo0nAuGoixNbL9PFo+c264uNgx/kU9ITBQ96wYiTMTDnGBNMY5CGTbsZqdnpahf
WN/kvglPJRfXkS58UdCvIrxRGlwaG03u/caK0vXt+iDttE6zupFqf0DymaUryOSc
xqHP3LFjIBeTzZbvUvCJH90TjZS36jFsOJ5iDfbcaC7fQLJdanqiuj7LW8TNfk5a
EvKmx2TFZriauGu3Vg7A0l4K2IoVXKfSL6s5xG0/h2UJlm9b9saq0AP837Q3Jb3s
N8FDA5/JaQscCsn46u6n4oScE1B4deMrfNnvQ7ZBsl2EDeaAJO5TLR/xG5JlvHyJ
lC66pllOH9QmOYWHIya4QwxRskZj73dTLvgce1iP1Z3TJJ8ScDEU20N4pKMXvnnG
1M86O0gy5PgQM8P4psxzZ9GdrmbkzOWZrG2w0J3nWjCyd0ndcSXCTGNDlLx/FLiq
`protect END_PROTECTED
