`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0L95FPOmCNo8IUgedO2MYnY5gYpr806Bxxr6oobtUVExd1U0X3jLOuw/XC3s3yC
ATVEJdCDLXaCTMUUZNQn6BiYYpSImc471KP7lyXVCz/zm98IG3UOhEAJqfvxOiJp
nB/6n+W9a1A/LJhZiRx2z5cXf80sTGCwgMDumAyId9ZR3ck12x7CIIrxqD3/iKx6
cYw33wLH/c+3WDf7B7pVmyoZL4xxYm1oTvMCNoNyexT7j8Hvcm6APYDkQ5lcIULr
cH695p489EwjUH0+x1jGUCCwGdughqlOazmRLN5tw30zOwVr84rquks8S7u23q0X
jIH0VxdGdMcVeIy6oLrF7bpMHhTFGLvL4jxvOgzrwfZAqMPHmF9k67c8/mVkQRcX
`protect END_PROTECTED
