`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NLXElmb+zt6KvsqHa3nXnIxJLAKTDZABWuMz7Bxq4BwUrQjEdvsG/d86X/cL3Zcl
AwlUX0BpejxUW3eOVLaPTIpOy0LYQkSCtgj0p38LJVjW+jNCdrdoS/XWjS7IVl/8
pVhxl1Jw2mShaL3M+bMd/Gve4wYd0WPLcaekLX2pVLdMfLP7Any7IXcuIZCByhM9
CHeKebL3kocT/OZLLKZRvCmqVDGfVX7ResjtEGLlsEHKFf2Ea9zVYFLEzJvZr8Oz
7zKe1+tH3vb/Bz3TDqfPx4zcXQhfVKcboQoCR6RF8eqnc0x//8Bu+t1fMSlntAH8
CvhUFDIg8n8GEOD4KOr7u5AaoHT+QnpOjShFSH8txrECTbSxoiPdOx1I058+gUow
s8ldl5MQ3/pbQ7hi/7wju/SLGXde3k3L7EgWtLkilMp6hzjM4xjLKuQpFE+wGLnW
EuwZBEh+G4cEkGo99D0xtEBEqf/1FQGX6e6hui5MUi4civntF2runezS8iOpCAni
ttofFMRF2r0/9LU2a2uyujMwL5/smoOdlSNotRH7NNV4sOmW4P1TFF+25CBPLOqQ
Jxuey7yNWI4tGrFXhfeQmbgyW9nhR84kRFr9jMFV4yD91UT9ODbVhEqdYHwHK4DC
jAsmQPkEQFTFa1xkcuuZb4uLOuQFSfpe0YgBpdbx9N2L5KGG1pa5ZRPXd42TaZGn
xWwqWo3bEuVtCxcbL/gnG8av8rbREwBmm/NZFGMkXgqVpySVVJXwPRNTNRNePHnF
sz0+Fo3nVmy//5DS0X85+zMPZ5Q1GbXw9YLrUZ2T9bIGdAWNGvgODLBFnfxfBcB0
5DOZn7ELkws4B2ct7rZ9dw==
`protect END_PROTECTED
