`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5kExDMSRnGTZHTH60/GZzn+NHA1Xl4tatGI0vF1cVdOIDRnuqpRqude21KB0Ulx6
3XoqQkcYJBHgfjYW2evgII4AUlsHV6B/8rKTzHak/E3ALrXGtriMPt7mEAz8QDEg
oI5Sqk2rgQnXnmoktq/+KM2wIuJaP0HKMhU7PzmZhgV52TkScc83M48j8b777Ll7
CiZ9+eGQZiBDgNO0NecR03Ki9jVAbRygNbyfys5M3R1L97lLO8c+Vljivs1GcZY8
Ywkkjyn6W6akVUTEvswQhA==
`protect END_PROTECTED
