`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjtns+d+D/LbG/QxKGO/gN8uI/X8mQy17NPRdGGGAtChmS8C7Udz/DJGJzfZP3UN
/UiyD0TghEzYdXBb/dV4+cy7BNEE7IhPolwKX0lLl6KUvxGmza+hYKzEd50mc3vL
1GwiotA2UvQ6yLVllL8nXnUYiU11lQfcB6xnQhR0WJaWCEbW0unQ3TxB37hCnaRF
FQb7Omz7GyWqHniNHknyQdMt2Q5ByrGuu1wSp9TRbLDKJt1Ep+wzNVTjWf8ZREtJ
1ARguw/OgNGouYYuj5Uor2I3m8orT3WOl05eV1cEaOwCA+9+MR/0NfTelKeSuNmh
v2cSYVMxyEWxczvsr/FL3oZXqTg6+dLFZ9i/FLwoWdhF71YFK3hk9i7qItQ9Z0aR
231EyuyqSkPxAIsDYWTah+nzA7RBfArAZwd22bL1uT4hEAnmF/KricrEyKei5ZhB
H58Q4bpn7f4g/7fZiGUBvqyqIjOiaTa5i15AHGEbxxLiOE04qrcELF/eS5BZ2cEW
`protect END_PROTECTED
