`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJTb/2z89WYbyYj0yQFV3TJXRET56ckQ/hXyO6IzpR0DT+93FRKg3MmQh7zBO9ic
kKoLlbKLZzb4jy0wjJEsbRqx423Z3GK2ifilC4TDESp1d1CpcsCNa9Y/wM/eet5/
jtptUaEdnvHCgtLC1av6+631r97YPTfO1dOXbrwN15/ilWUMV7kzRjHAls4hgfzd
9a5pA5xXKKDDFGYMJlBtGSpL2tRfW1FEbfoSluRmpvUgIQjzHF/h/qCw95Kh8GgK
g1acrtGsalbQ7JHhtbgj1KngGEdXJ19moqp69ll98DQYfkYapfZhNAY0ORw00PNi
5l/aOfZTYnFQhiGc6f6q+thakx3csqFy8NbF2EvKP2A1T4V3hthZiqZi5k6KFAJX
Ip+k+lShPqge3tSgAuqJKg==
`protect END_PROTECTED
