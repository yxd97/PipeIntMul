`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P7cwpD3YjgC3ULWN4U0BXbig+ZSi+a8NSAkROMDtB0NSe76l7STg0Ow4zX4uyLTS
MIkJqUXBssTBrM/CFqeceQ/dH+mkPZe1UeJrjmrmkK9ww8C+fjsImuptLLIX5vPv
o2DLsMb/GK1qgPCxUDjLNBm8FpQO9lvkN6O2/LKHxN8p1YJppXFGJZeEnM+/6fL4
G/s7uRshtwQMsi0U1NH+4tGv4qEtj3lCs1NVjb6STzysLEsjidPkNPKfGw2jx5zz
IyswbVow7EwVfpI5sgjg+g==
`protect END_PROTECTED
