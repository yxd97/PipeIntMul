`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhfDMvZ1FCUSpS1dKx6GS8kHOLFZVlKvAMy/g2fZ8APnqOGY1uHPmGkk63FF7jCy
dHjfdR7zXInkznYIuEebSVt/zyDyZFaE+pXzpr0eUh+kRe5yrgt3So+WGPlTgdlV
QqHIPKpFVrwOmXn1RxdAmmFBrAOJ6xTUURVktSNHadvHnN5aeSW5AHnC6liN56/x
d7qLnfUA519Op7BHnqMbyOlCd2y0u6n1ytmsELG+C55bNNBx+/TzVnyKLonKr45t
0M9/qaWUR07S29oPtQy0UvvSl/4Mca85GnfX0+jhRZex11k9vaaLuqniAooo7584
2kZpy5WbkMHIGuXnQ2Jq9Zam31g6XSnqUD606w8otvYZKDyVILox8pMqVZzAdyCW
Upa/z93MiarlvQNXKzon5MPBZ/TuhlkxpLX0mIAbKysKxgF4YndLx9F4gjaKPgAw
t1fQMtF+5Rz8wqwfWPUhpTlYlcMrTNp5uGLBLI9Ko1x5e3AXAsmjLgn2J4lJSjl1
xXhPfaJG4qOMyc2ktq8J3Oxk3JnwqN1m8EDAaHG3xKf0xL3IkrGDKpyYpcPuPgd0
TNWxlyG/QQ7dpxMu/I8EbvStOeQ/J+KVY+92kWqV7pWTx/eDZIdsQkKzAHGft4YO
UQ0L6y7KWZL/pVkiyxihmJUpPG05SwRiBU5affF8WZhAh89DjjiNydrxc9I0Hrcy
49QZ0Sm6spDku76YREDbxw==
`protect END_PROTECTED
