`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvF5U3Xj+C3u77SUSfc2I899glSrl0nD+DEUs48MiqThP4GzKlA8PfWriQ1/+BnN
1LwQJw907kJ9XoG3NRoX62JlxZSlgEQhfa8lsoIMuJVEkbsr9YM2oab6Fne/3uVB
YCFq2dZZpSW/zUSJTuwceJu/kXNfB5XfFLR17/ILPhwi4eMF9g9nyatJgcUi0P0r
TgbVEEEZvcfKTGnL8xJs+3sxhyq6zaEzpW9PfXYoynk3hq0WetGzgS5dyu/967oM
1NkRC4P46Nju/ivDhh8krw==
`protect END_PROTECTED
