`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ACotatm7NxJ06C/AdMJUx41RHVdN0LNEtwKrhdf4FbmRV2GwNkfsSoEuG1DeXDLr
7nHjJrWRmJ492xEDf+/F37AteqF5/siKMGpXhHzTun7bya6Tr4n6m9ibgt12Q5Md
dHHvjcmLXVONF/an56jlxkqbnKdSQwtl9ftyo5Ar/DL9KSLTmfQC9ebcZ8JX/R6U
rmH6ByGaZjw98Ht+jL9CgKTUBr6nyVsnerTebsvon30UgYdEXRqExMQ9tEe459cY
ZwJYDCASZ0q7v+w+g8ygIUtSJcfxl3bLsHFnuNnsJoaaAQBiGM4uYUiZdYbUSGi/
b/M7+nfWXIIdBHzpYOQMJrSn4qWs7hM8iebzXosx6Mb7YceSkQXQkRW7AYOIIvVA
KTEwZyWh7fKg+l7cRjnQIWacBd3LxxxCMCsfAmV9I4Vg9oDnFtq8eC5uzkfkpAIt
dB7bxQKfU3nBzxsPnAkpOt8Mx5B+Y6s1AO7RccbCrKZPK314SVX/dqWjbuHAsI4c
uCZUWflYfMzcD9vRvW3My1/rpWUAlokrhb87c3XhdzvSwbQah5YT/p0eyCV1ps36
`protect END_PROTECTED
