`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VJ9SSSq44Q6Ftp6rNAyBg1Sxx14Ozb71z6iwBfGQt2xujMocatABpftt2Wqg6ceq
qKW/BujJQCa2oqQM2X57ThYMDk/EEc9L4jpsQnfPhvncVmaQETY95RGN1cd/dv07
lhx4mOhNqamRB46I8jNwJ0wxtGiQMmScMk4kP8Bvzm8BAB7LSz45rxXXQSCpsqDU
jBVo1Ct/xSV8Z7asJ1Kw5EkimMA0zTTX13SIZ0EMHP+UJNFbyOmYmDyitdV/LVN9
yLdr0PxP/ri6e864ENP1cLtMsdjPjGbQtsj4OsapC+lOB3wiEissJG7rUGWpjW6k
V6p2kb90Xd3e0JRCAye2PIEtugpFFau9bHVbXVXQNXQ566AcFVbxKQ/BXBhZxeoj
PjufkurZC2NQ5QHYdV/bRq51apyMCD+MYxR1+C+pPKfz09BE6jI2MTnWeTo8H09d
v2Ic+A1UQUW9EExbxuyux/r6oZEKzcxdldTendazJrY=
`protect END_PROTECTED
