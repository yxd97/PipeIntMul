`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PSsVf1xjAvTkwmrv45Oq6x5j/0G9PIdvjG9GwZYJLG07FK31vTIoO45ImIPYE2eR
9VuMqaDnK0ABdl4dKKN1HQgDaksCLzpRI7sioQ+rSJ2JZKWJDTCXBwYp1CHVJ2Th
syz11FLYB1Bfg2OmlnxVun1oTIx3CgDhcNexd0Fa49bddHap0fnlLuiLAtOPJcs3
MJmFTZ62Yp4li4SATLMaAH2NQ9C9qPLFjSbfrUwTtjp8hCrtUStLNpqpUeWn9xgO
VFl0Jun/ov8eWXJMY6RPe8uhoTnEAUTNjTGiEnBM2NPR7aJmoBq7kBlGDetv5WvV
SZQ4knfvYx4nBLVLEmp3vZjGNEn8UYDEWY0xtgICxYlZ//27lT+5JS6mpqhvE+p6
2QSJleUpZBsP1IRec6wWPLJvFkxIVocwMwjzZzPXfgTM8vFkrV+tqJMpaLhBbK6+
SzAz7o1LYTtB+B//kikmV7HII6hZw/Av2RXE1FxeyyLORmALGxwvpP5B6993c+Fe
qpvf9brB9ZwaspYQ36Kjce0yUv8BaTWCzeulKiMODraADhaoqCGsSVglVfUFA0zs
amwnrD9ZjRgAu9933yN7TQ==
`protect END_PROTECTED
