`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yGo7Je60TrP/pHKSMQ4qIQz/spzzHK3qcYv7PIeIByj1USosCr0E7qJD/qbaAwao
TRuPuNQglGyQIwPXOmhjbuxx2Wn/AthXxs/awRpGarDMt56jGW37yePs7y0Axx9l
GTKMIWI9H7xnVNYVsehs4LeK7mVlVyrg9e1Ufb5U6FflpItr0GQ9H+yQniYEAfKK
PXDE8oMnNFLnFzAv7ba3qZZ2mmRdLtjDnwOMJCdcuDlZfBDfvP+FLHu9yCDJykh8
VyuaPHMir9iB5wfwuysUGjc4N2/gavNgNQEjSdUp/FHhEcUhvhYu0biqL9crYIw5
G6rXLA4BDGWR3lvfJMbldwuviM560SuvZSzbi65FufM=
`protect END_PROTECTED
