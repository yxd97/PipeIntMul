`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3sBDCoKGyStaFWSRxLGmIjKjMpnBuGQ+CGnnbi67WLYqm9p4IrNiNI/VzlAZmUaZ
b2DLKCGF35+e27fR7vVVJpS7ncKCE2RmNhvtzbmlzFb8DFtsLNHYlE2nOoiCQspu
/+K1698kd1cUhhRUARTFtNKfd/YefEVjp8q1tEjzh1b43RilZjj72fiACD2br2NS
p4WsOTiZEu8MdBqy0IxN9L78Miy1Kwa59lvCqAVS0XqpkUhA9Fs0B+gqBARxAqfJ
ZXyxp0v3i5EVs/Ey2fbn9IcSKzcRXoJmX4bQQ1Ef5vHVW9kozFJ5e2y39m+IvBLm
fySdlYD02ImGlWss/pxWay11b05xf/jBtesR+qlqolWByfCIXkVIov9KOFyxnev9
v/T59nW0Pk8AW2xdbFR3lZyn8Lp5sIjVqVK/yBmKB/LqYcfdf9Pvw7ki1BWPuiZ9
bq47x2E5VwXwoXBqEwp79g/1AbdkQeR92cFjm6d/3m7S68Yg5odlvPsyqnhK/5iO
ANzTuDTlR63vaO7WIyVWGi3VasxOAAe/i4OlZZN6PEyB6yCwNc42vBs8wI5dwdZ/
lKl6r1C/CRWi9tBipzAZz3FqUQHJuvGsLHkgffnL1x+OMz5DR+v6tKcxGbVsIv1o
774e8+rRvGi9bmu520Wtiw==
`protect END_PROTECTED
