`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCJJ9EPK4YgpkA7yqzw/VrkueZZZXjX8HUELKV7fVu/ndriknJWGjbZzeOHYOy/y
aUMaWKsyRSiVC2NT22aRStzQiUMcngvy+97Z7sjrq/Ogyjz3uwQSxmxZU9YYGLUV
aleuwBLhj/J3zMXPuc5fJIVXo+R5XaFKcZkswVad2iEWjEzinNycQPuuAuG4thV6
OPQWcP1Dh7shRRJg8nExVNx5tvZfTe16RWb0MlG1QrIRxmdimZcDrbv+Kjw3jK3t
60i5m0aIAS9Tymk9GsrerfV5FTf5vxWEU0Mgezw/EPoNdlovRmRprMTWk4YMB71g
oPaq1Fe8dWuiDqb+p/JrINNQChPXyPb9hZXxw9UZoCE=
`protect END_PROTECTED
