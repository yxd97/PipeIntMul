`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yvHhmVoFCbBM4eDZKv4f9PeT3V9670W5VwWNy42vKKdB5s4mEhw5gtic05xGs5gw
D1bZVsWxgVjzK6mQKuF7fVZquTxPGyO6LL/hBqkLofolJrhwqyPyzeZKAWFYElq1
ue3yQArB2QSgDLzw5ROQ1xkgzTiPk32a2zKrkZlc9NiadOg3AefJrkl+GlWJjvbc
mSnLFzD12mCj2e8qk1CoLSR1KJ1KuQ/gJiWuiwgdfH/raMsOK0ameKqHwaxks8G/
8x6X+OoZBJQcRNYd1affc6KNMurn1/9Lp3DQsfUJuH5nAoyNs1GM2Z1QeYcJnNMz
lo92BJ/c0WAHlehjRLBbRF3wSyATHOb3Tor5BrdGifiT5MB6A1z6BPEzZNT7O9YI
yX5Wc3jBXZ9OsTQ5usX2OoT2k2CDUfoHvqtwCM3a4wNF7WCUxykrpgwvelm2P3g0
ucMZNmsc7OVxBvSjMMy5pfXXEVP2mUGX4yLwH51b7m9csoUW8mzP3idgjn6DBQuM
`protect END_PROTECTED
