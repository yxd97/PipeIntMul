`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TbtMDM/CjDMfOk2sxqVGZdu/O962WIeVf1SQDjee13FI17rBUx2QeqCHFvvgPTs8
+V1V80GOcNMM3vallOseK0hyMWYy8JXzBF1vGjT8DaCkwupmnwTwz6lDBekXZz4A
VA1JrN42/v7f5yO22Z7BuvQAsxYOm+JfUTZPGNKTchER0ToI/b2ezt34OrNogRUY
9OSNRP1c6n3KSjoonz4gnb+hvnf9Z/nkxmAylRmdloKzzsPq+MYnmqLSPw/wHWt5
3+Us+dn8AgmO/DJ62vuQpDNBwypHzix54X807X61579l4f3sZNZnQSfl1bwggvT9
e5Z+faEPQSFIce3dCsLpcHuONWoBQrYm24AgIx1+ViYVLULHDvNHD4RZVGAZK17S
nloIKbW53BXJf9pVNOg7BL04eB5TaAuM/ZSvI6SV+zRqu4hCZWel9/ncpi9t6ZQ0
7qJ0nGEVTmDfUfL4s2Q68xCFvopJXC7JiTwFmq/JJgLhyvKmB4MgKe0E7dAiO82a
`protect END_PROTECTED
