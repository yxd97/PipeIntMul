`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W74shfYaZS/pfZKoFdNyV1mlZcNgbrhf7toM0aa4k7QOojSNfvSznWjeBh3iv8cd
FAyheJLbQ56xLMzMPclXcMm6EzRjZyaDE5fNuyl2CwkQexWydHq4eE4XBFySFAlD
T9KiWpEYAMW5XEaSq14rVBeZSiBsGA+p7jPwmGTGD3Jhuxne99d8bSCSzlrNyUCq
BQan2KA8sUmNGVzDHK22989rzTM+AWKGwLhy4i3w5FJA1y7HHAJa2eCdT6cq9HYX
yr9nRogBG+/Gh2/RIdrt5XpGqg58oo+eemoSfq6UwaWfyChDeDkhiUTKevU4zcHR
yoL0BuM8eg9LXp66KeiuoogxAJ1lKGUkaHOCg5tdQECyC3uAnI7ykNlwdQs3g26Y
X4QPyEp+qaNZSb3IhwSS9BBJW9xVg/c23pLpO8Rwf4atKLoQc7UJL6qsjbY9g0aS
ofhlOeZ18HWkgRYch+8UDXOGL2cLL3iY0T4ObF758B9VTubse1sBmXlzZXjtr4Kb
AJyW5TLiCbaRhNreWTzVUA==
`protect END_PROTECTED
