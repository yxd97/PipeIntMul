`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MdNlSFcHecSAtRM8OtVpsr3Tr8Xjp7/9Cdf70Ksn5EKrDV/SbNGis4dTMG8TUx57
StRX51Zot96gm1buTZsUzdcTndxwhE42CODekVreGAV3pzQWwNrSEKh+5agdACXd
86WmKr8L6oKDDn2WiX9T9lHgKyGfRm0Js8YPe5Rjg2FM36HiCU6GkbGE8iYQbVtw
reF749yqZxTg7V8ip7dkKAtZ3ke5dN2JDPsuaopPDurmUmWhRRCeHIUPwdR2eDD5
irOURLIu4S2oIdvwGGAtEcX+kZMiOrNpZRXkFFPp19f9KuvvG0aLDmvAKdKPG3Sk
rZYFvNYlS+/i/DqpobVc6NdY8Phc0obSCFCERTpSOMUaHWFtnZeiMHrCp9Pr6IVh
CDmeHINOwRLPpOYtyCjFUUyLWRXWYjyFp/JGjU3tmsbCzHlOwuQu9NmxiBZuGg9A
nGXsLZpYnpFAZd0mZREzVShEPj+LvGyxPTmxm7VGaND0wsKW/hSj+w4rvnnXBo7R
pGkAnmIgPHMp3Mr/GEVMi3lT8abUY0FEm2ZX+NeCvIHAMeNJn8WDt2ZVQq/Fj40V
ZYKRCzHpa24OyCn47CpP/EXjnBZqJOU4RnVfEHPqrNCI2GVnlDek5r63T9b5o/K1
dHeDqGR+Xpz6ApMVOzfzRTXIUhgjxHMjyepKVlwHaMM=
`protect END_PROTECTED
