`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zms/f76jTuOXSLbJXdlokv7PFX53gbyURa+SfAO/LHUsbcMg4CZRzHIeFe6vVu9b
nTX+1rV21FsVYJdy1MZO0ov2s36744+otz+0Q7TJu3J88PMdtCN/VVYGczRMEjjE
4IgUDN/LYVKrHHoHWiAFZqMNpTnP0iEdILhymX3SKJUwMRXAHX05m8b/MPHtg5pu
tRt+Lo6M8Y5N61EehuNkM34fX68WK6cxJcvB0y4AlSqQS4xmEYpV5x+xbp0joC5v
XJ1xnNvHGUSMWD2qtk04/A==
`protect END_PROTECTED
