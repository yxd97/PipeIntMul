`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2yybYITTf+iJE6n2qq5IKADbH4dzr4Os3GxlJFDlNvQBNsI8sq7cCeuMZyqDebe
XnFjO6tFsa+9F1K4RlcwiwqQYoqJhSP0JHgk2pko72E3MylJRO9ol2LtTL0JxMgG
dL6nivRk2oc/KeNDnoC+8wJpJjo0yLjdWNFSIpEIMXH3FxAr5ne084Itf1BAqnL0
8M5MiYwYZOh2qykhlUtM3OplPm6lNhtdk4NtEyVkM0/PxCOfxxF5cRk6mCbLzRIA
wlA0cXtIznInRZJQWq3MBGZ9mxBguQ7FH53gc7ih2aA8CaP4UNgim+0/XzzQaiiO
gFyxJyBTgXHnFSWlLZwVEIlvQ5//c3iDdvc/irQKDIkkIN9mjZ/zY0L2ZSshzprG
6TbJ5VJ6yQkBPnEegIQeY4Z9DYvR7Hqkyl0i5BcCS2vkEUwZKD/0tGM2WgDrn45L
ducAAC2DkboVXzRUKL2/z1HKPT6SAL7VjHyrBs88k6Bjr2VgenYMcjhUYq7oNc50
Ox4x4VaQ/GzUPzWwCsh+A4JZmCjMWDPj3qDft7LFvFijLDnuiM1w2wavDHAvst1S
UXPhjCGcFJOLEvq+zR3dlTNENaRkWnDhriAwGFxEI9gT+Nr6sisx3QkiOGGoSI77
Zf5P/XrSvRRI0Ex8/3JXH3rQs/zAO0VtGMUvDs6XMw78Xha6fxr68Vd4OV2Uhrfy
20XSZtm65C/DngoCkQri+q+BJFhhE8puKqU34L7mYPnqt9r/ao38xqmq7Q7v+gBL
QA31LydyhWmCweAs5y/g2Q==
`protect END_PROTECTED
