`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c91YE3JpKMC9uOmNHH6cccpcBJlT+0UP/3BswkKetQQU54GwVRg/StrTcQVvV557
wfxZPk+3X9SY8ZtPCj4PhsjsmQRRavN6J2K8h9E9Y95FUSSqKuDbV8VCwBL39jNY
nrATltNGoF83JahHu9ObokxWvY7mehisAoaDtdlqrysT3YF55rsrco+otYsFcobO
uyLd9q3Lr3w2xh6CSaLFSVAJbTAQW9tROND6Qb3ZQX9z00jTiHptbu+Jl4EOqoz0
NbEpWGdqTnv4IjlRvdMa2925Vx0BMrP2/2dZ5IQ6Cgw67X75FNKaQv+zGN1TZXWp
WCuknIqeWeisf2k83ek2keauoMaAEN2E3Fo6xeeB29APT7xXnVTLWEyOVcOUqaU+
O/WysL/WhpMzNrJg2vMk9WqVnWwhajYW2LeRiCF3PEMXSNMuy3CuuKmwUSrZBvpL
WxgIPSn7kid4LjEcaxSXo8Q9uwdEj1aZMse+vCA/em86TQFy3kRdW6wqlD1nZyha
xj5Z2BMP/Kl1FOvgMl6HllZDoE7tnZ1tGWX85fMHm9GxxMZmHaGx98kZflp++cZ1
rrNuC8OGr768ge822geNXSZ0bKIUH+/SZtI28bUWTv5FvP5YzQM2WGlcbFQFgF3i
sR4QNTAQXC4MUFLqBqFv2iasUxuGNQ6Iv7/u8SBVMw8AQ/ipcImuTq/ODMF+VAc1
t4RsJziYmuoO5mtiHWWvuWx+YOT0uW4Os11Ua88vyQk=
`protect END_PROTECTED
