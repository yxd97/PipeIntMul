`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VSNpEklqpap/JoKFDs+SxiC82+Bx04ccjs/728kBYqTZXszghqgeTbv0I6qoJSQ
dT+Z/SVXHkyYoTkWU1DvcvuFmuN9uJXwH1qU1V3vwAcns7FDBvuNqif3cBFzFWcq
k+6UrzJxb7LP8LfMsa4kB5CdiKMAnYnho0FxfIYJxarhiLbFFSX1etKRJ9TRT+oP
6wtM21zwGdctF8sgX4h61/W/U6A9hE+88L5MeaxohZOQwnCo0/oBeeFa3g68M+QE
666tW7xEaumvChvfM9ZNvA==
`protect END_PROTECTED
