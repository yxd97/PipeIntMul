`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMt6lUepiTy1YqxKSckg7G4vVvltLFlA8bARjay0pcUI6cJ2evb5BvFk8qVmOvNC
bN46EhAxz1uwEtTJL8lnnHS0EeQHjS/JfXzg3dz7+DvrPymUDAiTOcV75JfIeAt6
bKwdIrTxA02/4DEXvmGvAe+pXP5MRMneL0vpIIWv33v7spq30PLZAlwndgTKPYHT
99v3X5fBRdxnnf5UMBvY0YvmAjLBQ0GZ2aRo4mwopISxqa40tdQqQRYJnxXvKTiX
DZRzDmZ1jbNeprOypw4tJh0vQ8D/hb1ix5XdVlKBut3wHlmvO9vY8nDifZr4XU/b
fOPLXD/rUH41ClyLNVLNX5QqvNDZthNpFtPenqUbx7sgKqCO5C70h2H/YS/1QMJo
aQNN+2lzVlr3H4DtwpN5ebHFXKqhExqwDjY4ZvIl1NRmseLQESadDjgpkx/DIOWz
`protect END_PROTECTED
