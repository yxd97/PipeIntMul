`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MlTjFTT2ChLIQDVjxuw3+LF8mNlBUNNGhF4EQoc20NxYQWMhvCF2d9oxmxG25VY7
t10MBhiP0XaRe4nEBvDnU0heqzLX2EBgreUVRHqmWecHJ1Gpy+51uyEl7CJ0/B16
FlWKl1v41pvrXPPvIeI4vkUKZ53641qrBhJ7fQHaWOUUBv7Cxia6WQmXQ1AiCfuN
OwFEToYz8MTorWrK1gfbPmN0xsfkcLIkfJtPSRUTOFuxsRU0DD10FGXe4lwu9dvz
kR6wWDw28pkPxGborAWPKacj9BRf4bJ8JdXhsXfQ9ZW5to9NOK616ZtbVCTpl3XY
`protect END_PROTECTED
