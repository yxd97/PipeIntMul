`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFiweLKhCm4Vlwbmu4fEfGK29gcu4XdHCY6vq+TXlJVFF9D6VBYzqX6RP7Q46gAr
wAWQpZoYAryW1Z1YET60CbjU2pgpnenigdqonENpx1mqd4j87RXRvAdVj8IrUZ4S
q8mKDAnYfoCay0zPuitzxHZ8S3rtGZfxhPSDmXOYsUbdFMueeebKTzOl+bGxHy+I
RR+g0RBkbVLzSFIpb5xkZz684JR+LTOEMxl2L2S9toDtgXJb/E0OFRA960ef8wRL
bNArrJ8UVeueLpgAKj2WyEFdut/V1KHVdu6y/R12M3qLvpDFTBQLL+jpyhX298cg
`protect END_PROTECTED
