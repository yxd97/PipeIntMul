`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
st/0fh/tLCFukCdlOcPzqoFPe7S+SotLLHYl/SgCh2duC8G/x1mlZHhJ/dJ/tYsG
Yv0jhjtUM6YIhGWDTrMGJP328ot//HM5PBXiQb/6w2r33W5Ys/9RAdSm845hnRaF
gHXOEww5Ia7ZeLwswD0d+lDihYXJJof90VvSk0jUIzXkzBqUeYlqChGmglyyGimP
vdO7pB/Nm73r+tjxsiz+l9TWiAQhCNznU6qSp01ndsIL1PJi/M4QroiWX4Wq1zBT
SIXkWyJEgnDji+kQpgZSHpWUDmf8Ex6uofbHU3mrv1iwY5wRAKnz4dxm/FuyOCf0
uWOAXN8ngIIO7fIeGL1kMuqsjxgtnAlxCGKOYrlL3ib0Dd8RCc9Fjw3iw5/Cv2Gl
QhRGizo36bJMr6xOfwiYI3XOsTWfIUlcYXW8/PKu9rSuChyPbHBV5XIC2Nw6pst+
wGhPRsDuYKqa9Ze+8zZNi2gFhL4SuwNSH2++PFREpF3DPJvXf7wiodRLsET7UcvN
KXnjCwDn+9TCKFS5c6CqAUsNaD2cIsCc8RqQN192vxHzhDiW7OTUm91Goaa6OPQv
zwnEk8FwFBz1sYqOSacyB6GEcz49dTtowbya68gAEEFXnu2ZkM8+CtZgKTblPXPF
7gyVScTgoU+V+eFJHfkmZA==
`protect END_PROTECTED
