`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
51g2XK95OV7r7cyxaFcuP3xao+fOrIR6UjDxlkqE5UpdKx9jxV0rBisqGi39A2n2
a1fwk2A7iOvIVXn+8qA/0zJb3rJD+ULpU5+/b8lpeLbPTjj4OhEx8nUfBD6jY+HA
YkYyWWTJpaXc1V0zjjAbAm8vHEDwieYBqheOheHf9TQBQJOCzSg0zFMDdsDfMvC2
k8PEKcVjc1Dcf0XAFC5+o6uSus4N3NKL7mtmghv4FlttqTjXfWncgC7w1qs73a3D
mFKC9U86e5i+dU7Af+a8iyIItpNPiIYZH4Wb8hpxYYqMKyY4uOD5rv01+nLsuTo3
vkxIXGsCKsbk0OBiy7vdMg==
`protect END_PROTECTED
