`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jfw17KmLP4ND2TbpBhqDbALXu7jbZ5qEo8zGUGFGqABx7k+sMVGP6EW7AyndQXRy
lgHKFl4SCwVcN2Tuj1w0CRvlSifvTqLvtuKwFrNoZIHO8DVAs2NCnkeFCKZFxMHq
urRB1Rz64dv/yYIA+/TplcpMFuOnVA+NBqyJFGwag9+1mRxIgt1qQA20qvAbPfql
44hhnH6Hp1/8lKI6nmM/GL16Snwfbo6RJJkNrJWhZhTwqKbzTY4nvk/tCqMMkYN4
Ehs88l0F/x4WMRaJGp6Y/teftMwcR/SXvRxFIBdFHgp+G8vHeR35bjt4vqz9RHwr
xUR/JsXKKFFs4teh0UovBK6uXZtXyH0yyD6+Jw3HXHW/JCCeZg2vfsXo9dKAgAz4
d8PjacaPDSqJ45cERdXI1gErZSpp3hTzBEV2GJcSWgdJ2XZpRRuDUh3ANDw42G0v
FeDP6lqLRgZWjn113z0zodeRyLi2z51lupCiLmXlyGkhpakqz94nzeHn6JOmMY9h
EMDq7oCsHWso8CpWHFY2QwwDqMaQjeQP95U7GX0jUaz6z8I9QS7cj3bfSB3x9YoW
uKwBomKGUAT1wkprRu4a68RG5KdTE2yqul3SuPc2Gr3DnFp3Y6Aluuc4lp29i39Z
cdcxTUT1Mze8ktPBO37/np74fLDOvwuqmXLxLWpPNVgE9+l9S3ZyoanY6deo17I0
qHf7lKHjW4yinGBJMcI+N7eTW3Xjm+sc/skmprrzQJIYZwFeuMJ/UUwnn9UTdWxB
TisD6j/66dtOokretGo9mg==
`protect END_PROTECTED
