`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0dLCHdhlNL0Ba4LwjWGLT3dtLnHE6NASxU4nxehO8BA7FclgPXg5fvTUxjmP7JT+
PFbpdmVuf6iYQAjraWHfbAFvyPaO81LzKwf5AoPak+tfugJUvyFlvoxHEuNYf72U
XEKzTbGLVMv/i7BJx9cfEbs8g+yCD7A6l5z5+F1O6vEsgxJ5NoMLeHCclCmUj9aI
baXpLQgrOnlG1DOJ96GyM3Mj2psw9u3ESBTWoQgZR0YNP+azeJz97/q8GlhNmuHc
406icPgtW63BWHqkJhSMLUelYa0XywcRfYHTjzdTZ7oxn+bqgyZKqlCJdsz4qi0U
yKTJM5kQUOi8SVgo6QA2aj0jaJ7qJOwPN0FWGF8iSBBjIDpigzy/UDWCNuPXx4fz
aWh3fSPsY47WW5No2jjJ1NN1KLWJHz0IjmVubKgocPCIHR3b1wwfeW+3afYquYxQ
Kka/1BevULco7iU7vRpoZkIumczAvcmlWMzG6jdBvGEQvCwohlWGbVoxBHmuHDdO
WKnY9YAIs1ulVZwF4rEprOTH7WW48ASSlwgQu8bSzo15AEEoa3jAEmQDrlLDXFq4
Ng7f2jSxiHXYLAcmg/PjaA==
`protect END_PROTECTED
