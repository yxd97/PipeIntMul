`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Qblnd4ZV7LGb9ABze5Pn4rIUa3dvLceYNHYXOFCAlquQuK5ddnQpMYTOUD+KpoT
cb6NFjEgrbYOD/SK/mHAJSGSKkwsqSiMOggYYavAmXWfNX6QoFwnEIXblThoNTWP
BndnW5avVEZTxrxU8nXCg6aM1dMcNNJeZw9BXKPU0FAkdhTx86pU0101iCWSApWj
H+n4F3kerPxEWK0GEwgpMCPJJ7TfVaMmmc0XrF64a7ODGB9gIwUWMNAUlt0LernF
EyL3YwBYd+9LUl2w3KMY0No8FruOM3LXca82luuU4wsTP8cuLtMcBl76BAd7RHI9
OTYrG06mQz55hu2uqr/8Q7t6IskQTt5h9d6Wny3cnAp1dIx7ZVluleCXmppuAVWu
FH602+hNQDQeCdB+mcNc/sYykWw1kNLIwjsCWTHq/vuyDFSo/ccyHE3JIc8+wgHJ
0OabKxzQ3sUqdKY3x+ZCbX4WI6Wlf2fffACTy4HhN4s9uhBT2U+vXaAoWOzAmjTD
Rw/iunVncEFIJVAHB7IPXAIFQQJmORho8tKCgB3MR9jeGwFdd1ZI9tLtLCuqkHTH
kEbVvh3zO+X21jMC5VdRfxSuLrtIO94B/qk0QSjocMfLp/TPA0dLJxOKUsH/Ve4T
`protect END_PROTECTED
