`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWq1wb+dBVOXkUSlZHDy/aIZum/rmGaxssCW3cr+YzHbJik/acmfCot26ua4CcbC
TBcPCNRgxcjRRFSgDVfFq+aF6VNnTH2dwtlVbAFvERoK0cO+aGYelsX3M+JQwIn+
6WJL34ubZy2MFLwCY5wTzM2EEke3aOp/2WzXVU2IZI0bmCsVOn23cw2flfNqajbs
fOnK4+oeMRnC72wN3wSPdAZFJ4wj/FjF3WzBultFu2Qj6XFGw2Y8hc8Pzd4fUs9u
FfLA62ZlORYLjkamOBvjLsYuXW1WyZoniu1A8MdvcHdKx6owDXbmNc0cv9r9Ulrj
X5lzhWXcTOeE34gNwFOBxMgUN32AKZR1TocPd7q//b5j9jgP9k47DsFY4UYK8l9y
uVG3D+e/dtbzmFzIKFWCDYCI4oHWg+epzeeusPtaZ5mBDPoIh+LpIHUftWIHdSod
yLkFTC7b1w2fibVqpumcHnvm5Yiz5EcX6j68nVXqx9ZJV/CBtbmwLn6zw0IqpDjC
CZUkDLDuXVcvXU4SSIwEBxyDYBa4ZIj/pl52V9zpBKDslBFpRPpOdSSaRp67AEzp
5RzqO4UMa9OvexEtzbGCRAM1uF6qyVe2DF9KKPowgg8CloMf44E9wFo8JrDiwZlz
hpnpmVgAP2hBnMoCPJ4nyMk9xxzEBeV6kSMLyVNGRnhpSymQswkio8NvOuybNiy4
kIjJMACgf9x7ueC5f64Ml633t0m1sZyw/UJI1XIdgW/aGVKgusSP/EkVg7TWSsl1
DjIwbAPgY0DiqdoJ/b7MXJ98LZzez/eglBtoDUB9Q18ZSu4j4NEDHJOfYTCIG5Im
7gDrpcjODVo6VTZp1XM7YCY9v7zK7dwgIHBOCVxUgfzbwGWVHNlTBwh7KvXnkFLD
xWIVF1sg+iYc8C7Hrhn6lliD2t70QmPphagNx4xrHJiGBB2usa+0VNGkYm+1UnQe
`protect END_PROTECTED
