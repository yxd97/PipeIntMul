`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCGGRBXJ2fs/ItjmKn28vdFlECHXjwUn6ikbgiPEjF9fZe7AP5LYCbT0zmrRJCQ8
ebXeSh/ALdFOt82vezHBSbOSnQd8AXynuVRIjQ9+JrWYORMjehNP4Dg+xDY93FPd
DbADlpbcRaOhCHZK/5sfwjSXyQ41hfcrN/KJyf/R6mBW38tJ7g7eWtOFXwMryNvl
G1kcNEGJ71MX/J1iPBfUGIP/7yxSCgrofLlu/ZDKs3Uv8wEYRtGCYwya5WXd2kYb
c1RO5UwWSnh91j4I7/BIo/ANpyRgpR7RQ90zkGjgVpUCfrV8UdmxKbhaDsulp4nA
HVL3EaZKqMRw2dN8HL9sId4VPxhFNUukkTrPnpKwBh1Ggx2bH8vdDFsvWfD4mQub
Fh5vfVRD51L0R3wiNInSqVQTUp0pRQgAxWZdVKoJI+FJWJxAmT+JjC7Zxp+e32d7
h8nLFN+JVTre5zK+CxsoANu8ArWD+Cyo6dANofWL4RI1L86edbBR9/Ac7M8prgC3
qpJq3OwQmbNOtwsLFoLqBH10cA065TOowaxJYZD7QpSSqCldvHdme8onWXkGBCmZ
huU/FwJ4qIzchb0R67IkWzsXkj1F3IJ2ots94lUnWWoHbE2wvOwJXGLh4t53FUUo
3PK2yNo0maqpZQDzqhQZ8XYZN7raVfnDHAj/maxHy1VZ29rzNc0eoRu5S2g1iVib
NnSeJpGPmf2qptwQ0nUpgcI6Xl2k7k9p1ric5skX0+y3WB1Z7hvSCwz5HtV1YgEk
wuMLCHYTCmQ3u5/kLWRJdeCWaMT9snTWhT9p3e5x6YxBQRU4wTfv5Z21yAfRjQbU
xd5UGwfTSWI7W6KyWbROgXZ3I8q6Sng5Lt+PQe9LvK9IwODnByoeSbE8nldRWnhp
SWt2pjhOoy1txkQFJYdH5fHuY6z9ldGMXnGN+e2M6R3Laf4SKw7uNZBRtieL9Pac
bqMC2oNdBbXhu5XARXFJf25ha7qRlmzsTAzj0LpQQDoa3H+XEWJy377NZCVVcNnA
NqWXUQQJJbmXLPfZfvsvOi0ZTvg8Lt6JU25sc5s9oJaHuiQYOl4dz5N32MBe0Br8
LUmTYDduSj0lfiDK1jb6x8voQYnOigjWDX5Tl9RhD15rhm7b+9bmjjTBv9F0mZha
cvg213BWgOP8IAPCj5Sr/e2HzDli8gftPdjSON3+3G2yHQJ3qY7ZcsY9VE+RkF6r
LR6o8JAH5pv4/xac1xCaQ60NtT6vAwDHKMLEvOkzzYJPMcXoUTJoZACxfjhnM09i
WdR+beDuONvP6KeALTCaq7sQfoXU51OZIVLxy+IIGhNV62iwCYmrzbVWNtijfVdU
jATpwwUmEMaVKI/C82xWSLf+JCfNsMp1+/2yPzKGf94iBkYetE04KkpGbj8gNAwa
km4jtyL2VXPE8pY2MD8CTnsYRWqbXdg+mWipDGv1ip45U/DQZzHeBIYybFn3vvXt
W6ZvzMKJi/neJPwEPOV7+Yamt6opazw3/boCvKF4CuZCNAsh6ggesW/HlLfVA8SN
YYf7f1VkRTWFnhLGtFYz4DXrZsDc6LcaWy+m27LzmuxEPQn+cyA7H8xfWjdVZ1Kh
Y8DCohSRuxCrzPAlaU4jUDaha8mPHymjRL9TEVpAmmXODvhMUfrw0S15mtK065dt
Ri5GITOjmDYAn6r9ayjkJ/sNjXUxwtsD2Gy8ilTjVj+KB+KjxJ9jQ9dxeZTXb7K1
4bxMEjw89ulKJdtbzha2zS/C1RbS9OpwDNZWR8e/ymup3PcUg2h/hMQ5Ywxe0umW
KWFXkzcAk3A9DItOw4pJVPQLQzfcSUIEkBSIpxWs6HLVmYHFgd/ptSYSLm8DPjKQ
W+IvW+VYutfDIxaAsOQchTgi0dKCKhVMUTaQxq7vjrhkTujFW9jo5+c2ReiRnmAI
lMFjvMY2sk4s5sHGlc5vKU93a6CduXZNoUw+qDSN+gGa96hcUP5zwCsgXYQifpOJ
wgA2MAwquiBrSVl2Tf8mml8zgsV4hZimExBQ2lkLyv28zGk1LphS+TRagGYA27kU
e5/pA36csmObd6nFVOljmHyosLLgUJW2HTMpbOJXsZ2AGQDF6cbPEoBSj4kQ82UW
nUsosbR4HzGK1lb+f56CdzMY1k4ATxbBz8n9rQrFK56CvM+yI3xt5Pade8IpIgCZ
yECTpKY0hN+VXqQ69zuvYB0j0ypNCyV6SUMyuf2gcTdqWhpHq4qymFY7FZmkZBx/
ZvkLD88dBQmdVD+SlzaraOeZl8ZBKfg+YuhXv1oHXkxMJuflyynGHYzuTi7yRUf5
lObiEs/CciFMHBZTJyehJiRuYqfP7r1yGtzKrwc2zzNmZ+s36XrI53Zco7XFzGu6
yT585srm2Yr+pUWuHnZS/xHETEcLTntF88pmYYt0d7FEwzyA82besX975qUrAirF
UfTU+DSFwPkmfVMtXKAewBAdn1Nc9ua9+pql09TeHw/erFM9lu+S1rBzmjDm0oso
GTZkJJKF9GKX+WsqqO/xySAB3DzO82Ql4Pgr9rO5c8D+C21vRvT/RWqIanZ4hdHU
wdhACxIRuyNRvA+oBsU6C06V6QZXMQYiAbg6GQgmq6gLbRJqXH0IP7ONMiHpARG2
reXK9wxU5LgbRiAlC9hiDZuhF8H2ajNooGKUvcWubNwF5TR8uc2ovIJNsTo+sPcl
2mWp95Hb5OBP1R3q9lrPrn5U+KVb0po2dkyhGtF503QwjN+DS/YrnvZ9jkvVkT5W
rC44DOn79Pd924bhcOOlH5pvabVTXNsV53756OkPiBcZRezPOaE5t26JeThO/9qc
iBV7ZqJMqg2wFRHw7nnkhQYfkeE+ee6lnQJI784rUmJrgtRRQOSoeqzV7USbUBlv
/LrKXeqoIK20LIkJh3HTxVTYnADmKH7gDIYKR1WkwOtlsxZHygI2P2YsDFtvAmOV
8dpZp4S4jCJLgoQTniybG1rH/b8nVKB19vTyByPPxmkqPPx90Oxvyxac7gt54SUY
pWipkEK91evS5ytlYPnxbDDjiQhNd/g0Q2wHtTdkL9dpWXCbl1YQvtu2xGobhFjA
YlQPQK+72ABCX834YXoVuV0tgQFSPd7vqAF5i1H7UC1SEb3IjxpRdEXXXLJ4KDpJ
BXaVqbBNpu7YA/2BpESy4RSX7+eB9RruK60PvDpexElwkiAXZiQmrybQMQMTfUEc
JFVYB2Y6SUl8tFctNj+Z3tBdiijCxpZYtCAPQm6nGsKI0Il7ob/9F8hS+7qQC9iw
WR6Sjc7lxaeyNOEhCwsbwiUsLh+jk8iN4e4pD5AyjLS3eUPm6X+32ZCyfLfH7DgP
zhJrzirJJELCw1qHYlc+N6EJoYVuRI38kJQ+2IBnrqmzUB9Vu0pfAzGAPDjujYzj
BIEMsnl52tWlZ9DxGM1b6WV1UCj05MYB//w/43gy+H0Dj6GPGluuhk4IeUXvZvH6
HZbwFHJi77rUvZkPBFaLdyyUSSOs8TcXf9iHaSH32yXBMWVRm5pSY6lje0+UQNsz
05fXGR81iuC97eShDSM/fsEtezPZyEhvcUIP4sEBw3pWrCBxGf3Zt1PUfSxZ60eq
llqhx/IKPGgQuYEzuYEFuhz45yJ5snUwaKP1w5OAn0IGOGIj1BFeFyJ+4Rm2zpqX
1FPB5EZq/lB6+k2mWik5lZZtXMKu575scZtiMhXrE4UYVQ83WMkXs4oy2Uau7JjG
44FQMC8CNJEaS8L0jRKix/DMAQ6TdfDXj/HkqcNnnDc8sLfmj/QSVT4jP5Rja0wB
Lb3oK3eAXGTkMCX1O9Ol+9eqiBSIqEqMeZLd94n/bky01NayGSRZ1NCn/0eLxjql
unBk4aBdfdJj7yS4Ol/2zAjz3o0EId57pmi87xK1O1looPw1Ydar4xqOd6pvfNOc
JRhXdfdMqXZe3rgJMJTlPIUZfYk1BpBtwh5jRHzda0fyVZw7nqXGc6aO19GxQEA4
5o0Pgv41Wzs5Rknk+1Gl64nihkYHiqcxLN945YMHD0Z2XGJeaKFOXkZuCNYnHTnq
mVTB6QjXbD86ldL8INagULZ2ocPLab1Oj+no9pGN6epGbzLFQgC+KplkXMZBSupH
2zZScz7dZjoWxyxfWU5DJwh8aXLtinPr/7dOtO7DUMWsQcuZFbSZZm+41YlE+5pf
frZGPFOyiuA3i6i6MYzclYaUxmZ/Z2aIZS/AjvuFQC76AwpWHcaRTmfwXuk/E4e1
/9FRZujESK0fiemC0oOV0GrxKgBBwjwbr64FB7eGlsFiCtfBU5FUFzk+fBfUpaN5
XppOMNB/X0gks06YEOQbTvniEOjTVIY28+JYYQWYsJzYk3MRKvqPxwhAIyB+YfHO
c7qlSgaFnMHdMceZ1oH4a4O+woUsf2ZQTATRO9gAgz0GpWYZUWmQKobdusy/f/C7
GxOG4x0atl0kc+PT41hFwBmUa8nYRvLdAru4iarR4+uJ5UFb6PvfTyT2/MsY3Joq
v3roCwcgIhxCkIDi3x82s91Eubj1hzESn8+6kDA87fR3zKB8O0G82eLAnxKSWG3d
6IYb3SztKq4/rEMdNjY2fopV2+R8eSdSJInnoFD7aCnc2ouXCG35PXWegs/cDUU8
66E+hEn+rZhBtz2IFxbJ+5gKqQo4x+tL5dmIP70XVXgq9TPgOKabcXl10Lm4Pb1R
ww6WseB5MK586zwZetrMGUo+rSjdb2blT1nirL5Plrl9QGts0+xu8tIsTJP1Blhb
dPRUEyHQCPa0KNj749oGlIjdA8pKu+uVXJ1zrfvc4/ERf1rTqYoDt9pSLDDB3iKF
2egNsN+mPt5L0/L77Qn94eokqMwirovOBNB5cF820psk5Pda5HQhz8DPxAk2AkiQ
evoKkQfjnN74RDxDc4p/OlYdNFnzWUBDJHNynDNyY1BkGCe6m487FWERtP8Iwu3j
ekGD5squBp/tclvvvIutEaBCb3QGKndYjoIuWAV/3PiXO2AFEnWSyO2bbVnDUAA2
hxdTJO3YQN5PRR82EVdp8Y6k4Hx79otkOqkPDV6qqFeOkWfJUWQ1NR3PZY1mHeIB
tk1ukRbF2haEA//2KksHTi33OKXt9JjcVIiSrOH2THC6uEl4GUxvM6M9p13ZQ1nE
ri9RHM0LTP4IbhtLioc3O0qDXcRy8G1qrMQlw1l6WmyaAdCsxuZqiJmr3/XPbnVv
7tsCRsle7TesoQ9R1dkWjHqyqp8gDGUCD3oTy92x9zmyUc6Ju7+zg6YdZOYv7Jc+
6I37SjD2iBAlMHZptrY9kqedq1YzlD1/aX4DpugEIZye+rtbwk+YiRAjCtC1bo3h
lj4Bk+oHxjJi6kUl7aXFCxY6LrpMWM7rdddwajYFYX1VDXntDdicDtxHiDCNm7lz
0vor1ReAek9HKMOFn/Rl0UgV1Ood81CVpUXGx2wVd/DSV0Z2XS7YrhYvNvqIfU5G
dEASkmZdanPtFMyV/FkSbIQYNU80fGCsITEj7hVOzyx85tpXJ1KZKF1ltarkYfCg
za76QWBvKKtF92BLwjbOBYCfzq9mYCApsS2fV4gjW5C1XwUecyllcMRHfbhQDhMr
t2s/c5KDzamsm6P0V70chyChiVnHPeWEoVWaZ8SD/Cwuv0aWMubLEa25J7+S0Rin
feTGLDQn+4ymolOpuruT2XvY0pVzTvCz6sCuUoKNiu8j6LJ8auC1A+9MyhGIOfb5
0oHCzo5TNcbqpX887uPQeAr4xB8QPnH16Td9OhRq98oPk5wEEcg11yuybGk4bZJZ
oV6T/UccdHEuIOW4pRy5wj17pyfOL9ErGxn+BnGB84G5x9YVoiFCTCSdmKU0J6Bn
jwmwKMJffsWcr6PwMZjnE+IQo2GO4YS98WDGV3gB28SbqcxwUTbpG9rMiS58YuQO
RSy1U/bWHa72R3t46AMrV3U686RrVGV3MWvnen2PiEJ+Q2dkW704mo+B9StePeld
9+Bw62o6js1uik7lNznTuJPuFth853UAqhaTlrfhQlxtKsSt8R80f2pV1vaMhEPC
gN/4fV35CKaqMiiTqUi2Qu8yoDuuo5sM7l+iNVr10MhCdm37PJf01GmZ102KMODi
pO/gRJ3Abp0iKPJYoPCnpwefM3sFc7kDT4f4mM0FAdiFcNCBlKcie+7QWl0gTRF8
HxfuGcxgVlwG31IjrgXXwW5OcFUAHLb8k7TovbPVq8cGvHtIc+ifrhEpUfNFYpPZ
QdwzAibuCn5Zh6sSwgVT4aXtlgbzt1vuLv9qfO+QaUkOT3RZlqv/sAjjbL/uKQ3T
OOLQ9Zb6RzdFp0EERAloeWjK8fbovTTP4t8BYw0/NLhJ+kkPdadx2Anl5b05oMXY
FUQS70lzZWKZomuKoi6U1XHro9Ksv3Mpu+m1yi0JVbe0E14D/AShPpXBgWDsRosr
BKvDI5JMwx/nsjPAqkD+QrJXueQoFM8Bj0GrwwDi6Mfn35Em5ydj+3ltK1XuHVGV
1Dm+10Z66wNNWDqBPSESsKDwSb8hc0Cn6WpLLKo/fxqozpFIVjKZzEKY+HRKxldl
YdOyw21iEeYj8TikTkyIIB+6gFxuZcCgmPcsxHcV6rYGgACFZdypxjLQcokPPRbH
9u7yMOKK+lCVtF07fhCrGNNVZjPHdCBE6lTTBS1iKKEyrjFYheNlyx752I+4JtUs
l1NlP6bZ1HUZ4E4XlPR+HPpd8kmzN9f8Huqv6kVkouTWh7q0QVd/4ZBKY1xf92M3
ePmtY6mp1KXXHb8+xay/uIkXPwrbF6ADYcx+e5mED1lP4SJm8/uW7EY9U3eX6QjV
h/0pqqoWvLN0vuF2JQELD+2W9d53IkvPqKfxIpxdyvL8gfdnLuRZfnP4egNb2uXB
btwsTe0+JWJy0p7oVNt/p05uuksP/kZ28YzllATQ4+jOLsykdxKnSdy+yURBWe+A
ky9qlE1z+YcYAyEQnjBcA6LMStY+PUJSX1cNRqnn5NN4waMz5QY416WjgExf8YFe
qQEYrbjdDNSxT+qokj6hRV8OufIOqBOrDo/Efkwr7ShpHrGfIeuW/t+mjptogdrU
LWcfwdJHUE/rht8q5gUxa/qygS/Ao6OtkfEHxd40DrFDtutngddqnYd4uEM2roAT
/zBNA5T13H3T9cwyzziRg9kBqDiMoHcu2QoVYbjFfkTP4m2yxD3FxPz8BTaFz9zX
AIP7ne7ZOdhSzHPXq6LrjaTpp0A32blRpgrEzI+UGTAWM4/Ei3heq5l3sZZbk0o4
qgHa39qmQRSoQyoA/2Kypc/Ui5pt67+H8+JMcB6tQeZ0OUFBLAgwvh0xJVv3AmSB
5SPGQinAePdoDl+GM0O27QdN+yssNeJPEsDPdDyEw4F6DXoVOpbTT7SmIIgv8IIa
LVv5I+ePFk5lCeCQ6esbbVvIVShek06u8HsH07ysa7IQEoK7n7CWBSg91tk3oZ4y
4CEav9Qi0G6/3u9fJgX5XFm1H8+N83fxVi/W1ObRt/hwirPiI660k91x9WvAlAmh
A9mJNB4jDDE2y5W9zIvgbHe6UVep0Jx5MS4lBHrWyJl5tPTXBhu7+/w5n5OjNovE
MsWQpihNZuwPvMJDHZ3Ge3CVhWAO/swnaJKo81ftivRb15JKwcclvKb/biX1x/tc
08DYQPNPlWYr1j0QNt3oXCBLSKOYoI5zbjSa8DAmgt0RxeBmdPhM+2sjNrAZpiJE
QXy8MkwZW50N7z7q2JGZY6RHt1fZU1pfobdIMtEVSbEx723FsQ8AGJ1OBD9jrTCs
1ShLOXkFz+Ei8c+r1GTxgrRuJjMkuJlkou9y/rInjk/sh/uI1adxMAIblC4tBRqS
9HY+sJgEsKtSeBK42PBCU4ld2/6nbx+Q3sBlPLNW0BWP+f7k4Z7du7qY7t+iv0lc
uTB8YbXsr8hi5UGNwMCwzlzk4YQ44cEDY4O6uNp54uHGIeBBm8kqjBaTy7FrrOzz
VWCn19zw584oZEPeP1B1U7QIv9tCuT3VtHuBgSI18AVsGrIswf6Uw9C5ZeD2gkeL
0BOCHu/27orpNj2WhyGjXwhLcandb09BILfuQqpmrvIWGdlMZolydLoBbSwhrIJ1
RjUkA+7IiW8aGAzAVhtU4AxvTWAQAv6wXq+R5EyOBhbHAfv1R7hgsTW3OLHbVdwG
3+OWQu+uRq0hbfSyDeYkuKy2nyd0mIpmVxMJ+kPY0mCqAUgQ3LKp/AkLpVQoriCl
P1ODudRNpxzYuqcUU/2dVOYcrJxKwViPP3lbrAsF4emoEO6hD3W2TY3AU9EdRZef
XgikBPzPRt5t0lBiiBbs1KAQdbn41PijLCOqyLn0EmHpu2UJRd3VYEfUuzItsAVg
Sa4LrEx2dS1WRfxikRdxYBaeQx+/abRlVbC8aQCQgGmdJtO0DduqQ7Nj6hnibo9u
IUWaIh/qo5mIEdcFFKj5Lr63JyNDLp1o5zXKJvW19nXJvzHAdCVo3n18CRIFtnYQ
o+oYM5AbHB8AG75cp1XYR3tb0OmHx2Xqe68Cdw7PZ/UT18qmTEMvBp7D2gMcyu9J
47aKFrnQj3wVKbrD10Vea2GaiCPZ+TV29UymsQQmP7cBDg2iQNkS7Xir1mMZ6Bec
OiZI6r2onEaoAeg7t3w+NxxwtZfgEKNDPEU8fo3+X0IO7fg0blluTlqjqDmWZcBZ
hD7tmi65gmFRzkfJ+xY534P6p4nrz9S6/tXOnCJy7hDGyS38MMMGbJNn8OKgeDiY
xn9ZvnETvCasUx0l9XRYesWJ576e/iw0rFsEUlOm3AyzS7H6eKCopIcx5RNDiWNJ
T7tHYJQhdaYtu2xDNs7xI+VMT5QziUG8YYDrCdadqBu70nnbjcuAY68kwbweeFyy
zTkXh5saT1hF2tWREsxi534dt/Inn20dhWVTwUNrgK4UObZ/NQRwwCl5KDxOmltl
A3IlL4KGJ3DS5tdAEBV56gk9sBqjUKa5VrXlkKCJoO6rbA1La1C8SgE3JybVSGeV
4D9yNh/jj/Evk7I31GM1Xca9PxnpDNq2L/ktWKXBOx6uhA6sRtI/RXZ3xkRZUVMF
S7JBx5JeoJJkIlt+BSMsxGqA1HHxsLLAZuZ4w92iXYuoSi783G2lCqQK9FU5c9Gt
f2iUz2rmwonWx8JEKHEB8G608rTEwPPcJpAkusr1LPlsLhMdXPdLblphTMahuojq
/BWeVdzxK952hO0q02THcJesDnGuRMbvr1KCvLivSKQqwlRgW3hTNo1Ho5W8cdR0
un83MmB0jvdRRHozfCzdT79wNcidbUGtnkNgMm+AEZpEunuZERaKphRoqi4/qNaN
VZXCFRH+mN+SpIxbPW1WXZdlQbT98WM1U03y0BXCYcLwumQkMa5oQnQAUt79VOVG
VoZ5AoSXxwpz0R7j3ovpPYpp1UZuW+SVVgiu73k2C22TR+QFC9kDANGXhsoHcMsF
YLY0YwYPLstCW92gN4Q43GDf1yJnlT41vGZpXcU7If5uAKaVeunzH73B5uhWicSj
qG7yYwvGJuNr2GaOMzTi00/zup3VYJscnFx8vKggzb/ify9n/vnPxQ9QXWooMOb2
QETL0iYKqQ86kUQ5iJ2PBaOcJNXrZ2mlcGEzSs/+C7IuGQsViiYRgC7RtzQ7epbl
FDAVFDJNxqbweYv4QZq9vJmKI21QUaLRv4EUkzoXyQUoSPTU1W2RcjQrkCK/JrLM
MNvdQcAZoAZc8HLMXVeSH8ITZ8E5fH2Tzyz/mSy28aaSK9utObOEkvFOrnPa+r6p
jxXEeQOZuA1BROfT17spSaKZzdrKSmfagCb/WGHymUY2R+fz3lU4uDLvr+zJ61+m
pJxhXd7n2rhxol9+Yt08ovovg1+kLrx2S6Iud4m5p7VL9/fLlgkurvlzOgbHIeal
Rqqp3uqJxzs7BIeeSi7PB+bYI3EuCgASsrGnPcvLFQq3w5QqwyDWJ3H4AkkkIJG1
cpU/MjrR8x8FvgcYsKL4mxpVsTD4wAPxG2YggudbfIZvqKLRlyZPJo2Kzh22iD0M
XGSMmVIPqWialr7Cje6+i5dKS3tSfEfe8Fz5IBysWz2w3xHHltBgOyJ9ezm599a3
QDJbGa5b1O3aPyMHTS+x+VNibyF7NzurOwmVteI6AnBVxt6jZVSQJgcij9dJeQnQ
7BUI//1LzDMy6y1Ic7v2pTvfSvO0m9bpObB99wqYv3JfdWR/Q9Yw1nSCulXZcsSp
nNuPZrSxH4nuw5oOy+MI7lPbtXfIwRDG07Gh5vBxHp+hWUkx2pNBcX13vCrHTagC
m1Dm2HZlqyeOQF0K7bjTlX1jLlCBwrXbP+LgF45P7V7+8mytPa3mNMeZshf76hq4
EVvv1JkzXtNr0bFl2hCl7ctnQV3tZTlh9WdN8ukacShDMaNSD7tvPeNuYkFaaDoD
rBhPNVrr5fvJaB4PlYpV2XPafxGWCSvl3ppLdxLVwUHFCfzXncBgbcHKlJOCqk6a
6MyUyM0rknvj4mr3iTZlVDIux7BUU5cK7OikB/gtwqO9jHjUAzAHARxEwdIPDyAB
06FA7M+8zQnGu6DZiwlIm95JTlMihPGE9gTVjkZFQ2lWny5QUrWCKFnIiof5YbXw
0zsMSudQ4C+bAvTBdyltdWVJOGAASbdG3VKYdcckM2z1iuP8AooenoAGk9I1JA3Z
iEi93292XlvbVaw7aKKNwFv3F+c69hBmdwGVkQA52XAZOfjpdMygPFj+wXeSdKYw
QEx7rIoehIOBn6PUCNk1q7iUTpan3Lr+BbI739/I5iZQxEK4TSN1HjE43kNBHCq/
pyHZyfSExzTKsmZRj2Ht7u2g0j4KX+PUCPtpw+ZVCq19mC0pZlY0yKxl6XQAQ2Za
B0mDJmyVGe2mGpiVpFirrIf2Cz5fMLr8v4dowXg9FBvUxGnN9C+iyOgXPd+TYTUo
BKieT0tzm/I98j+Dcrfpam9PsoY1JuLTojWLtF5DzoI6nQxjSFZWJ9cyR6PJVwR3
YZua5yu/5+WwiJONtL5vAnHZw+TsqV3io1X8B9K1hXug7cywXgKdzUqUHTZz2ODH
uCIUPtl3YB7b+6DolJIZaXibB0gWTRLhtNELIDG9CM3PUSg7dGGigTPsfCklvLZp
bNClpTUXwi2uCvGzaNadwFxScX+7Uu7+iliq2ZeSxNdSdf6GcAschO+hH9I5JxhU
oocL/SYhbPuVHMSGPiW7klwmEnDttCuzhfdekvV72yXT+inQm3sxENdXbwz5oWyV
TMOfY2NeV0t+kTLu1bOE75OR8dJOj+WD9jMi2HFQedqP6JsZzbg4JBoAx6mQ7IAz
/KFKGHGwLtWUJx1ME2q6JLzpNwhvdaSjdNLKJM83UkPl58KKJovkVFDukZdS28CP
WoxVYR6LyXPVnD1UqEKLmklMA5c2uIv/M4wHf8RFhIQOTVGGwOXNJSNq2iX4U4s+
tt4l0OUILCsfd4nZHvtLlClFfmcw559rh6BlBNarPWA8vlWNU6LDe4jQB+W+4ABF
qpP4YNrMi3pA19w6HPa5qVWHJBzNbmJ1qxgePry+nTb8/N4whAvGNE12YpUYtD02
fzU2z6vOZUxyIvxhkWWz4hf/+rMAC4Bmp3r9y5eCYETNIcG1xC3FADeYKO+mFvzH
fQi+DgR0c6wdqwTV9KvReRKKgZDD+tGBb18+XbZB8gMZQ2KE/WIJ4xzIVtSAu/yr
cUVhsJtaBQ6nppgLO3F8Cfi6JCULG1wtymKtjMaYKjeu26ulnGOPOaYd3uZKfCsu
xAmLbsom4/bvtokFfXmgtYi6/2YtCnIDQC1+38fTCbm58IfPPD8eJ9YXyaAOeSNL
UOnZLfI8w5Fi4/6Mjg9OmQXs9If9i2/iqJbQOP4s9hrxk6dC2kkckWgNngDuej5P
/z2FmbLiCJe1v7xTAN+/ZL9Lj/ZuGauw7GtGouCKXID4TXDXAgp0u24b9yi5wSaV
uoI1orQSxoMBDEf8uP6vFc+pEUOsXFnbLjrsVUZB16bD75+X0LFxA+6Q4KAJecB1
jNVH6zPwobWZY7aS3TQPZZI2GkbFLzF2mgpdtHVxlXfX+wxVIHufjV8hZYo31sN7
rgacOnUbLExVBaM7QACmAgz+2CBydAZan57u8KSLBiv0kZn1LzMsKWKYjzlPdW+n
4f//1dwIAZ039inH7dQ3A7DTnV39+unuO3sxxCVYspi31Y9expdZhSgxEzQvvdF6
whPIx6w70Jl16Zu2xVvU/UOMG/7YJYij2grDtyBrAqgsIkbEuA/hqruhEgnclkF7
ayeTnUYJjIhY8Be2mk8wsjOxcR+89L6bgGHUoQQLGLV1SoTLjsZEG6BrdufVU23/
6YNmnpptV9E0uoBBzP2viT4aUUg1o5lDFC+VTe5Xg1wJFeExvz59axhk6p7guUyT
0Uy0WvcLH7G4/lPcwdV1N6WcmhbKQJk2xI22gsQo06Ek16BHcn5WNnh4eXESXT14
s7TP1Kx5IF/tTOGO5R/gRpmmbaXvjvDTh4SEC5NMB2R15fbvULrQpIXY0i9UMjDu
LaY2tgR0jm9UkjKXYBXfKBOepZqxk27MSpMfg4bIzzRiwu9xzxedQz3tEV2GjyDj
8GenDWsEXRw3jfpwERkWIiXbVD7K5k0FPqERwDCzIf5NiaddS0Lnk0eGVgZKMZym
He5jMax/KSfK1cbFH9m5ilQFy3peW4sg0kuX3j8B+FVc9RB/0qzGkB+nv9vKWF1m
dS5ExNrZW8yy4nwXzdPaPA7wZ3DExpOJcF52zvf2mxgbl5ZvTkySK2KClgz9vi2j
jbfwEi1L3xcEnnt2vm/iZREBZgCJiEn4VMYD0ZcsJ+mBqUm+XRPe8VlPsLxvysh4
15xA2JiHLD76/E2UaQXMFfw13IGbyK0XeLMxHJoxJEb6OiuK6nKRQcYpKShYF1Nw
O2ONnsqOEfzU3scgojHDCF9iOJ9xG14F3elf15IWLyKBTzkC9vUtuZMLcumx4taR
iJe6P1Yok+ZYzWF37mbK3qvhumsYPlxBWUyf1PFfxlj8jJP2hjWr0j4NnA0dhRO8
6dJzzsDkuR3D/lJjqiE8JAQ93nJzZfjJnYY4/QDVW4Cokvc/JGO8j+JsKff/pJRz
3STHPriC6fqFfWbxsXW1feuvpk3bIKuVjIkEx6UFnY4fI+AJkPXEuhqFaIh0BuM9
/FO6cXDsE+0ugw9ehykPtTA89K7pIZR0g4ENqbjg/c0EP/hRktUJ6r0iBz4kVPjR
5hijY/7GjQnGEiLnRZyT2X8o24BQTThJsAskBVOpc+372RSKEcRCPIZEi3G7E/oP
kd8Bi6H1UIf9Xuk0bvLKfiryyJ7MYvLhk+c4b/OiAXOyvmtXG4OIsEg76m8er8IQ
1MmYoztJjI/dmlkOW9aBsd6Q9dTdKqFe63MHFQD+aN3yzDXfBVn1IOXcWisGpl+O
qzIaCIAm91EcvqwIDSxnQuhJ4gskSD4XvKdkOOu8WLpXVsAaUbro9ivscMT6w2Hz
KQe0M9qMUb2o6twjaf15YB3toSG1nMQPR+BOpSZQD4NKcEZ33Vp4IyOQ1VT21IUV
cH52IHxbK2bkKaW4ot25doPSrnC9jb0NNBYsFFehUoxJ/R2BSqHmGZ1GlkvCTrTE
pX4kACgzyyPTZAH/lktE8I+vSfVgJctgBCePABGio43oZmv3kQHc0sYSsXO6oCiG
dpKrSVabacZiVv3wzTmQh2r4Mxe2xzmI2NPVrJ/g4k/F++osUhVpOtSs3h/fylN6
Ku8Na8eB0udcabh4VSmk1plLUcPYLmX1DLmh07vr4M4D+0yBnIac+lTpwLqRfRlZ
TfxAuJikrL+IJdlSwf/kge78dUTDXWxp3+KbzPoCWsEXZir20vcgfdel4dn7TdnP
NHVzJWxnKOPdyOTAyNrl/Wd9r5fPelCdopORRue1n7S65/FHSnBwYfCwpy6UHV1e
F6N9jxYu1PEOoM6kk2jEdYf+Wuda4/dhT/HG2D52RjX56I3pwDYHgqEm1c0x30Az
xkMiE3zNSpWIpnPJ7hPuHaQY4Dd+jJdZ/m9/gGqxDamyccRrk9by0GKJy7O3P0cw
LOl9gKIhhnsY6O/TghkZ+0cmQ1gb8pJv2M+fk7GT2G6YGch9jeywf+wKZlQJZGHR
7XP1UcEB/9pZkaXWCbbrIT+iWjAFuc2lQvmLGV0Ynw8EBpGj4DtkE26p0oUmmvih
mO1cSUezVhEFDueu9gFTdGq1XeBm/LH/98LWSuAQLpEBJwLNK2IX7Z9Ay1aY2HL1
4eG2uHaB2I1N57WAoHXuQC0meJIQ9Mz0tKJUEqg4Rplw9pRp4EtPEOo2PEzqChU/
5z4cywo0Vj+wuqwJ+RgKlc/78GZSYqFREkxeWT0Tee6gUMf4ezqlFxiA970wpcIN
BHtIIbTZlHfXb28pes8RoSuZfpiLIYD4Grf4pUGmNTBWAOyNuDYyklvFh73ZUnrR
xrPkL2h11zrRkMpNR6o+ZiclS1Ynh9vnXWii/z1jVDkpfMr0SZRzR1pDM4lrEu8H
n+KaRVaIeSG8l0EEpqr9pxGcToHzgTHtrbk1a4y64mhTPilEsOqRAZdbJMG4YdAx
H6YWuv2U2OrSzYAdBtGYhknGg+vn4cNLc6VTVBhPtIgR+KuSKVBQvd3ggk6ibYPL
n97ntP6ycxVdr3fxswrLkVNzca4dOzs9hElqguRjl/45/3esH0D8v3+YJ8Kha4OG
TWUymQ7EWnp516qsHzWI0+BCM7NEyz8YV3zaJRHb/NehTNl+gfpdYDLRsvUDD9mD
iM/efDTX3zaIh8ZPw3yKeQorkSo4uWgVw8Fou5ZcX9BOdGaMJS9AFHfVikz2CwLf
I3CfjK0W2wgAr8eHNhMj8ngc31tIZcTkffJSxNy6+NAHxTiWsAIpVi8GfkrfoIxk
KRBYKPY6XlRswMtSaxPwb24UrRijS6A2mNN12hYx62Gay4EqB342MU47uttFb5vj
t8ximM/WtC2hgko+ujrQU/TSxrII2az8zvSPkQs/+7snfVXD6svpJqlvqzsiUOVu
MkG5QV5tHL+ywR/7OGTyDrzlGP7EgPY+wXXx0aJPJkuTc+Cbh2sTp37mrCJq82VJ
sn3HlTsKrtLHPGm1GW8Nrr8jHzIcn/Mvvphgse+MnKTjbj3B1FLrZ0DsM3cjI4lQ
KDMoE8iopyzNav4owjOpcDGOko7NrTg+akO3x2vCD1Cr5jq9m9A3AIxIO0EZcaHW
`protect END_PROTECTED
