`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UsuJQ0pEjOSZ+aKEzL2FRpPBlVmC1QwSqG9hqGXxnPhKP2yU1tG4YgEzp992PqX1
BLHEMN2yXktbk1Tj2AnqkwisemaWEuOgmDfU5EpVBWATvhN5/0Cn6i2WSHvGerBB
cuGlmagAWB4kxOK01QaanjvOfKtpxsUzqkLUTSonoJEbGOpZQgxNvvGN99S6wR/F
HcMXqBDkSBgiN5GjdUxFY0glit0W9U/R7Twb2ePdsYWJQlZku2M7RAcA4Z8LJikQ
VkwemStxN40ioViP49DJGdnLEsgA4LMoBcvZx+rmlclCqlBMMJImW6GShxtKyT+s
vD/FF15zd/oYL7zNYqbv4cRgQLq6US3gXrycXVtttFkh0yQ4qZlvhpeyqNJApWZ0
OdxkMMRge9rDDNmihjj9fA==
`protect END_PROTECTED
