`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3EQ/S8Oz8t2scDozNbpXtNRdBwM7Y0EK/Lds7DuA4TyIuVyxI7J/mQxH8Yndl3GB
/Za6y6627qYin/Iu1tpMd1/ielKqrQ8dmeKj513cYLGcYtuE5Y6SymiUs7vPzV7M
RfAKA5bDP7SzkCjosfpvd1Bh+kP2tbwUSx5F5uHA7GMs8JBQPVnAJiXeKf9Xta6o
giTeOl0iUR2ey2Ye3XB6f0C9hE9k6vfjl3a7x07kx6TYOjT08RQTp4Ug8Nfwp6po
vuXbRaUx2WutghJzXLVi0Ubf4imCzG7SK9HIDtVoANc=
`protect END_PROTECTED
