`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hg8YxGfWMlsMbNVSBVSGI5wWh4ECDprxjwBfB3kwIxpsVAhgjVlvo8HZ5NK6/p4k
syfKdUJuYropk4++y9BfM3GXhyCunrtXOzrDgbI05aSHYHeHNn8+t0tsuHUJsYa4
fOrKqcfHh0QvSGCuMgc67XQ4IVSlzzSF7IiWOSaYc4tIt1dq1CNZnLa5MzHJiWW7
aXVrLpgPmuKYAFO75khfPYlrg7xkuktpULCqrvJh905jGKUz8eFEzpYrNXmszHpY
gNsSHuaK35b0U0jQztKxtidyLKAsbHKWQq9oWugM30KLK2boAUDYI8ez55/KdUYX
v6+jJwZzQ6w4kPjRdHuizrq22WfJrEgK+4QzHT6wG14WToQ0DZwN3Dg/KZXuOin4
8HTPG4oFSyzaXFh28xAN938ov2f7n8JP4WJBnx2Gs85rqAJkyty5YTl581ziuV8D
G3olTDpqzNagPnOA8q++V4kUuRdSAU63T6rOpKRGtPqA51AF3xxt9tjl98H+xRBH
gqnRlVulSkRacSmCJU3z5OUjMG1q4JuDlVaL8ncgMuE=
`protect END_PROTECTED
