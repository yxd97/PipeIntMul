`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bhEGpnunB77/YCHNdUuKBdaKDpLyo6EJEF3RDYCt0BxGy+PGryY6Bt93Nq8ErGvz
2tr0i+V3FO7LAmOXUA1kE1qDd7YsUvX2enpyTYrHVfF3JPvZTj/3bEOh04EtfJV0
vCFJ0rbDDNFlzmABlNMrq5md57aEuJ9g07o8NlqCSRFUTshNtm+nSp7cZb1Gx3J4
001+dwma33zY84vCQfy481cqaQDZpvHzb6yYGHfFNbpQ4QKS7bIDZslOW9zdHmbk
X9CKzmtzrM+Vn5vg0nbdi0UOnkdocbSnAEt1vMwFx2Eds05Go1rtxeDFKsSH4cnX
EfottD+Gfm9GZT9nq7hQp8YN8ltmptWUvC9eKtaFNw7ShMO9AiLC3S9AJaZAFYNx
1r7VA1uqmm5hsI9V+BWIHxPinYbtEa3WM0edfFHIDkfyOBWetWz2j2CD7qKwtK4s
wUW0FgZzqM7+6uwj86pwew2x2WzDASgl4SmAsnjBrxf0ugbd4wDxVuP8P1zD2P1w
H+sS306/PUvA4mV+K3Z9rLEbJMasZOpVoAIvVnJ3+Yk=
`protect END_PROTECTED
