`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
svM5XcW58EPfr7wB+jqN7rvWB+xt5wjpjfbmZYu+yEiZ1OzQ86saiUbwmG1oqhNW
qfC6isbnd6CoPkP2WmZ0KeBynesCm1Kj8HnaXMsKl1YDotyl40aLfPN6a0JWBfjb
clALmYB/Wj66G8amkDXcEtrJ5n0WNlz0+C0649rJ2LZ0kSTmwtxKVdYc6Rgpb7yy
jiEGugXdDB2OP1iTvOolVCldjp6HXctGBjy9wcZ3aCzUNl1l5JbC3Cx4iNJ351Qa
Uf+g85+C4bs1v3ZGNRWfe8hJ/HQllLxWc0XT9SqSsC5ji5GOJ2A4mVv7VWkAYK4v
ZyNoyzXfSnot2sumhxvLh2IZahGsz2qDXRGrFLmtjGSvaPa7xcDhjiLyrxRKSxpM
abmgq76SyLTY7TcVkjcwh3ym979RSDSPgHYBqj1JOHqAPR2uETF8aO3GTRnViXW4
GeSn+DQWaRP80mK5wrAEXsDZFL8zuq7t4sSTVYAGlqFpjzg8UaqrTckHamBhzYnB
hAfqo7AXDLafK8TxGWsRqMXw0GEhXWvqARYT93dPkEW8ge5EvlBcgUEqhAdQWGtf
Et89GwmTYAm0z65vZOJGZJgHHbEH31yJKEtWfZ8LwWaLyRcJEKpbqJas5fsr/PkF
406tSXH23kgwPduTV+cEuaZVgZ3d0CzI1jDEQkranlczUnzQgVZ4YcQcBrmpsfwJ
cmrDIawx8RL+lWNTUPPlFflzqzIz2Bly7S5kQJuNL/fGVd7TNO7vzV7yeg6Z5PMt
zRalZrpYY9sZj2I3YfjQ7I/t7UIZvoEMc9O7ispix+z+FTImNzIyN+f1183TjBjB
iRen4rBCY5NfZHztnRCEs/fOiFIxQVbRQn6LTj3XBiA9zU+U2aNKAWky7oC58BkS
EhmNkVVg6nAM+ca+5vNyNchVhzZ38nWGjQ1RjocvL8uI2Yrc08ISDY0VW93ZQ4HU
LJ1GD7BHUgX6RnnQmApw3PPQWCND7vEO3d0KimASUqNmwSN47P70dQa3YYydyO0t
5rFCaiLLboh/UL4G6bN/yU8eWuYPHM7egRzXXuSMfgemT1xxbiJMv/TKpddGQrsb
2xEv7Vx9XCTP6G90H/tLqy11n4IRhr9SnBN6WVfCwOom98oEmq9uuvbQ2hrH3j8x
/dQ4JG6hO+7zUXruB9/6bROcFxSmdVPP/92y6BaXjsBSkkSC8SCHDgmT6HXA9PNZ
uqm53yw0m9PseeQHeXvqNOB0pgG/n8J6/oEyt7tRAmknRluNPfKbX5Gk8heJj7tb
EvoIwzY4dpcIQOsRFHXx3cmAVA9o+FHW1dpmWQXdckLQRY3POPQLkQ7UuBEP9JN0
4oHBbqJKt6EihQYsGncB4k7Kqq5TbBG0vXhL/nMnhFCMPIf1N0q/2hwD1RmsZ8XX
mQRFDDRTXSUSvm4yAJzOb/ahYKoC03UJWNHXFqEsCZhbbcV9kPhbQeSiqBTTbqJa
67YO0cVm9q9lGDmpu7Y0L17lmXa6CLm9surMUNIqiwIyg7nmLcOQBH3HBCKPKsPY
lRVWvZLCVIp2kjX7Nds1uluq/BZfHFcHQdo3iKjEUdgZMxLSrDniN2ADekyFkj0E
8SQblNlnSqJ3zSEAjt0k0xKhCNXtutBfnpI8Yd+wdfJCaZ9iQgvxrDnyGAIamIFw
RDWWNx0bfBigvD7hoebusZGODH35kCQdaTNudslCbpETKVfjdnf7gk8VUykq1YOh
epqPClUr+fTIRxcXJUnVKvMbKK63Y4sJKv6BtvkAsJ6HGc/mxTnyjANxh3c4INZL
b9AJrlmtKjz94T2BPAZMSmScEUYDyPpjmoCRN3m4JuOrw/rRIHcQo98dHYfYWXFZ
ikLFrjEOBPKhwskYs42MO97J6OIp/yRYrxjINeJDQZY85B1KtrHI13z5VbuTp7Z1
JHXtzHIp+UjeZGzlgJxKDfdqEdWyG3IW/oM030Rq2SznTsJOGjSlRVOVI22Z7bgv
vx+7+Sd/4h/vuM4piA4gq8x8R3oWhRk2z1NviLIVzgUTQOKlcEz17ga/dc2QldE7
6jNaDzIH32H/NLYjdakQX59KNCnKRRdggo+vJoQQ0i16MRvZTaRMm2NkWmysDk2B
ImWqXXN5+XInw+cOUFlqgKpru4sFYFa6WJ9PfhsL0Cg25wIVugytKSVzY0hkWhiK
e2hIa1PgxsVwclMIEEA/e+HmKN3ZjvTPohiLNj9DSRNltmrFpN5jpoB4TrMui9kX
2vXE9s5gTSgLcSEqzYGA1LFg9xogDE9qkxLjo7CyZoLS+2LRiFYmHknwcTZoDlWn
EJAn1qlUP1+kY+RdkUagle1DxI09K54wXOrNqClLN0Bfz9C5qBi6lpmCPX/Z4oXP
VBRQK8p8Wl9kQSuIyz5M7njSb4x7Jmg8kzuDG6sQ/jzC78IKmepCAUgp2udbB0+H
7AHebtfdNUaXll9FvDa4cqfEkAnFj+puzFszHeZyPF9fhGMVsyfquqr1ntacajWJ
8hbcoIToKBpmzYqfKJuoSgutJGN1Qb6B27dRVeZttAthAZIdGCuOe5NWMiVxbO2p
rlGQ3F1zUasjg90oVvOGX0Ydeiq9IYmE8D8LM75HUu7ufuNXDWoirvSgQ6/iTJDG
L8eD/z/VLQ5TkVnxUD++8J4MdoaYwIB3JDFj7d/06fAcF8Dh60eeMZy6xRW3bLXO
+AQ7khTgZ8smnb52p5gZIHr6hEUBXJC0G5x6akcZsYXnGD9qRUe/z6qBC4zV0kNU
JrPZrRD9q/C2VJTqmv3Az4DtN045oK0qNRCi2rMLef9zWIucOi1fGU31tzpeSS0Q
rnJNI8y+o5onvuwELKsZKsDLGelJhbvkKArdosXRjSyjP9q7Q3xoUcSdIzhYVnK1
uFy17VGWN7GNsInF5KPOBiLaIR4dmVQ5Fmq9R2ZywZPsvjsYkupQH0zYyd0GsKaV
I8UReyYNaS7Qd2ZNWf1UWD4X3GKwF38Jmejk1zBur3HQ+N99ulaBd9NgfVCWY8q9
FWpAAnxzc0t0qgnwJr/Vjn7pTHZtNNQT5WMrkyPxnQcUFxgNxJyyDLzaYAQggG8K
2R9GmJZVS1BBCGPoe2Y+U1JrHX+YPkIGNbLA7ek3ZzwoQho4Rs6vCzYmvBfbka5I
oawcDWiwDjzrSXWxG80zq26emlapA2ZWCtPtcAV72BKwzcfY6BbIes2C1yNEUyb8
A9V4PAubzQkmNGfo607ZBBLroEgkTZDEI0GBi296m6bdOcnwbyAfwCHuTB3rPNu0
vTGJg7J/PkXa7gjRRmTQk9sq+YpCAW73CFi7ETne5N3SPEZaLtf7m5xY6kqoHaTH
6cM/MyV2VUhS0Yx29O5C35Sx4rZw1R9DOwF7pPx3vEKJlGHEPIMuQQksfzQYgPLL
psiYHxfLg9nk3AhSUGqGamaPgJ3GtHdN9r3EF2nCMw/yXpCdlcS/NcY08rsYnriU
bw6X9L9750BK9yuNBpnNFLaNHi1s2IoAfHis5+jVM2op0ihUEPU8wEfOsRR2CmXb
HspBck2UUx94uf9FemBydSFfEFxj/KwIGgHIbXjc1sZKQt8kwXkBQJvf0hwmTKJY
DorMwtusVX8vmiqLmGny13dlWyf+2C6DZruSIPsiMPkAR2ReFBG1g3p0OzKDA/HD
miY0XIPO1o3zbotT2FCO59Of2I2FaZ61d7ACuebBM5BliWCuoS4gKpWZ0cQzNMS4
ZIcr2yQ8W9wdShYfHWX5rUP+HZYLFZXNEBMsh8T9/9cfVfg7aN8k62QGx6284Q3q
VRUunjDwIEZIqojHQWs8fynKoAOsTkC1gBnKnmtGYPgAKR4KcXO5psJ7ypmHoNEg
SwROYuF2mrFt6EnF8HLam65bzr24HyMXHjGdOC9GPYQ/uHnxq8xsD3cSwPqLoDBi
BR+A7QCOTt0vAUnUDt/dcDJ+lk+MntbOODPSnV0eA2OvTdrSVkZofQzx+9jpclSd
xrx4TnqiYTjskdYrGwmX6SQs2Pjz6BVRBbv5bC4sVqXONlhf7vp5weasgMJJLw2F
QJv5ehjFhACt3mdW+A2MLu2W0LNy2k+wkZxc7j2MnV8iHBSkW+9555D5y07+z0sb
EkEXHArdei4wuK3VMw75ERe9hgOJAPT4qGqXcQFlHBKw7BWOhlXFOYGrsL3xd6OZ
jDOHfun23H6+UCMPo+rluTiwXbKPRBbObA6kM41/igI4oJDH/dpkRqJo5xY9jonK
IdfVrEfFLJhTSGlmZDxd0ktFHp+b7rInEwHgzPr3XXpm7SOoIpXal8RgVoMcAqAw
wQ7VZBx5LbzJu3diEhZv4OWhwCNsZNLvcvcd3pMQSPlBYNRUQ0HpcmdnUU4y2snd
0LiXIHz2EVUueISgyRB5xiq7XWpBjIdtrEHfiLpOVm5Zoc+pK0+JD/R/D3rV//1V
+Znf33YwMATIz2NOx9QSr1SY2fGtfnUxNDAhlXzjh7/UTPFOgvPmgvokNRIk23Sd
DOREImMCsy6SQRYlbVmsj/GSNpKDH6QwFnkiBSHvzL4bXU4c4h4Phf8RMKAOjR5w
Fm3Wud80T1IjwR1E1nNgeR1VJtkkh5+grWDJh7cwdPlGDf854I5hLRvmKS1fDhYm
SvxO2ZvFXHQQsdl4t01ugeeR5R4GlI+cEKWyY+8f7ITN3Xkw2MfYEgOH0eAkH/0W
sGII2fhMdP5kpbym4YQ1ikfGA2rp4bLtAO6MLU1FTQst6daQyF+IP6CDSBFmM47H
FFvHx5hIFQkw9a8RomXIIXlAYOvozYWJ3xh5Vt5RZ7I/nUn9FkNEflcfbECYPEkE
nDIOid03/UA1cF5TNtf4fvmvwuoryjcsI8zkQm8pXD8Rn0CwvnEM0B8/sUoFW0Jm
FOzEgc+Xrf0hWW0CyT/Aq06IZ9F68okHGu3kNjwDB/c/MwuoZFcsxTDTyYvpR37g
UkyZ+ycv1OzI4Z8s6OC28R/T9Cwtk14dRT6rWJ/RTPtzSj44BQHGGSRhYHgGGH0d
gAaDstCfJj7NyC4hJNg9VbAvv9CvrV3qgciQHi27vwpoahMA/1T1AXAJPWVooi+A
QA/lKqXfWLk0iyVZWEzAUMvHU6LZy8gNIGOgRHN5q+wp+PS/rKuv7vy0fVB91Zty
+U3SwtFEEeNabLzK+lWfB4dqSZZj9IOqmrVAU/3HqsnpwnNOIB65X+Gyba8b6q5l
eeCnOxvZh+wmrGJTe7utqfEsXRqHb4bHDjQbK/ZXIp9t9Cf9j3/ndDIr72+Z1r+i
OBFdTgP4MTu3xCw7kQmdfhQR+XuxG7zOVcBP1FcbkQA/YnToMKoScd+8u6I8jggR
N2ugPmRSK80ikYxqCCxJGA7jtnF9VOe66Qc3f+t3i1STWmQeokJDw2Bw0XGHSfme
Sbyla84i0L1Yg0xy0uYwYvdof+gZ49mFxGpoidB2UA513KmzFcLqqT7YEqY5Q7MM
BhdBieSK0vgjifhKTgc8y7oYE7apGqu/Tje/TaC7pVV4U8ikaRYYHN5PUVY5csDF
Chd2REDwmVHrgV326NQWbObkfZJWmLBnh0ap5SKhZWBSF42IdzEskoYBffSvqUJd
6dL6RAG45QmUuvvUJNl3mQ3z7xo50RHz1JmqDSwimdup27AtC8s7Zbm6E9MSRw1M
0VGtSxacMg8LJccPUA6nNg1xx+wp8qpZFlfK2CJcwCBgJZ+rFFiAJIU7Ll+x8NyI
ObxckKwRVydjKBYO1CS78XVJa9IOLsu9/IaOVHJGPyzR8FvNBQ+z4TXOvJN1u2ct
unqyqrO1rJi7aTqFZaJ68Ul2iXhvYeJaveRxuDbj4XM8TIqFoLNi3u3osH3K7vs2
PFX0udQTnI9vzW/XDISNUMHUBoN9T2P6iCC5pWpckItETrH6bra9H0hH6bElSTuF
14TTz7uTAuRnuzR3JbHzM0sEP5rcynvkIVSDPE/sNChtdXofG66emqsrQ6ZNZ4BY
nPvfypUMxOau8g7rKV8BjNLhv7eSffOxEbtEoL1VDkAmwtsVBQHxf4HQx5RWJCqP
O8VSBujeUac+2Wlrgr7HcQNKNGJododtjnITyEF8qcdH2s6HVsZaxg7oQCtTM50k
p8SjN11Oqr5L57WGRTEqGrg84y62KQoSawO4NMz66ID1rXzRfGDrP/htdGBi/usQ
0oyIa71JAmAwWBs5lYUS/5VUpZSN/3gzn+FBpwNL926hyFCsNFbG0cBYpP2Q2YKI
OZGe6Gx0AFxb8l3UTmVgfuDxpHxoCsYyqngNpgLF+LPOB02IapLufyxYQrPGe+/g
WY3w6l7u9ZsqgTdFOKasjKXCOnY48SeTCr9ZNWbAqJGLQLG3+zc8Y6zb6aF4rPxL
XaCkj6touVWnY68nsjpd0tjnHlpq7aQ0awybZPQuii1jqVDAM/Wbba39A0r8inTC
fP+M78DHkGdWcn5oeD2IyFpfufAuklKLE7N2ClK9NivqJ6yHrhzyRyrN4r//Eq1v
XOrdehHqklc2lKVvaIJz+Rlz/jqn4tBKwNzvlDRUmsMZJeiDXqtxP85gzCEaYLg0
ILvgdjNrYps+1ICUersj6RBr2L1x8+KNUSS/EN3o5ZlU9mVKkN/tGCJioiJtY/bB
oqiSvNmrka/f0owRDlmVKUA8s0ZDAgC+QXGac4G1iEVa00lJdT0dBRc6K1zWEJBO
Jpl00hCozqGUn0MT3xiJ5/4Fw+wQGMvpWDu+HgI8MU2Lqnl/TR2Ar2Z9Ebzkpmwj
AsQ7tcDhfhtjbsM9zUu9Ol7NcYk+v6bcbU+zhEdrPVNl9+wn7k425v3BLLNK8Vzs
9fJOjIPFJc307UQNwzE+ojbf15bJbI6xi+vqCtJyq8jYaV4wsnAzVEdnj2gQAA5E
Jx1tWwUwP8XFNKK06PbvX3WIVjLSgtQBGPvsYg7FHMQxLtR1SmXKyVDppL3Lfq+F
/2OFX0I7thFlNGvtzXi07V4RzV9QPuuQd+4RsR9ngJOrLVvNyWCrFABRuTeQvDFX
KA5jMC+txwHQQn+iJgb9D7rpBAPnobUSEpHHIN2L5BKMHpKBJg4RjTnRFGFfjziy
hY8ClMFDllPSzc0NZlGpx3YLclyYSBf9CeCkox/nEvYq4Xjr+ChZW7YRW3lqKsJH
n+rYeM0ZL9ywJ8Rhk/i2zx43ifkKeWfqwWbOQ9r1q750Dgo8jxWTzUFqWNs661nN
XMcnnQEdcjfSmnErhvs6fBhjmqE/nqdsHUBsP8mpvgJYo8v/PJnM0OMrUg5GT+sg
uQNnA3zChzTgzX4sySW/09luYHCKeZO8qFhXQ2exYetj35bnysWHo+eMw9FvInKK
4ZVCXrtLZK5pAo+1egcf1lz80S2d5EhaDPo8oRESNw3sU37xU1cyLIUdrmp4N+YB
wJl9AkOHxUEBXn52pqlQiKHyCpVl6cEo9QuBh9+JxJ0C/tik4R98UGUMrYYysnDu
U6LLaBsk/y4tEQJR7ky8vJ7cNaEs4IgGh4uhfPqfAgYba1MvEjP572tUF2vBvtYR
zTOcqb+HBuy4potOoxXFWkv27a5w7SVWTI35Yoic1hcQ6Nr5F0gQ80Hj7l66k5rH
JHRVz0ikaRH0GoBCAwv05Mg6PQ6DLR8yBdc4/544bUmeZ6fNtGapg38q4trovowh
p+jFTAUmlY03lxk+c91RwyA5+HLDLuuV9lQFrSvL29tsGdbAbHw6XEJNjw+XdOUQ
0mWV1G3MRJELQ7EODPDioDdqC0eIYULQyTx/zi+GiFlWxPRp2PmOEgbI0MhrOlNn
1cazGABT7FpYv9AHAhGaxVAeuoWcTHwwXMZ3UfZl+evpeeJtcsafGdd8uTrDmXjR
A3r7L74O7wX0TEOf5XzCsDiULzIqG5aWq1ke+IJPg5Rs9ZUuhYYpraEhN5MajYwa
+Ecs95vfR+cv4K7xr8Wl5gM2f+yrW69xpDR3mCbSIIBN+TjtfaUTAMHx2/mPuKQ3
gBLhHlaERKlXpuvdhStOxy0NsPt9+XNtcTSeIZIXisgA/eiUrdlpWRJ3ErzCQzBO
lIno2+F0duFjBEz2ysYFJ719w/Mi83FSAyBebbSSppcOgV5ipofAiaahg6NcYQFC
MSDuNZguCUxEYUpjB/OyCs8kIpeVV5FRZHMP15ifBTfPhfYGEOaoDaV7ZBFLP1dx
/otCmw92PoL8yM7JjcIzfBO39D+/OWDVNqRu6mf3YlXXAgrEvoXr5PF52SBF06Mw
UsECCjHZ/o8Y/PpWlTWBKKRhFS1WC4PLM6i25JQGKRwvsz9brbzBVAkPCATFDzlb
Iikwnu3Lhbuo2IaC9/9IO9Y9bTyG8n7kUirgHl+HgFThhzWuT+YnZs2RdpW5jlY9
3YkG9sXWTwnFb4TTWeLPkN4jb1WdjWDcM7AadBDRtpSGCnJwO8iNdpy5AlnQXY9V
XSk+xJcaEHeoQqOPwQ22anCT4vpq3rXb7syEaU0RcbP42HIf7v18QIjITB1ZejUT
Jls+LwpUfYZlokQ0NIjP1N3HUG2mK3yNxOPlXjNTk9hg1naoWMkuyic0iVC7QxZJ
jmcTHaHXUM2eBbpL1oYnVsCkQuvaFHh9Onz4i6jp2GiQ5DJIhvvdI58YNm3wYgbz
GBUwwpF21vJQMTRA6OuUlfuQGFFnPpFYLE7Jct59GwZZ2Z8bSJ2qaCV+1wLGLSp5
lNvnWC1FR15geA7hrE2L6ZJuycLMipEJwd+s4ckIksvjPCty47crFiorCqhB0RYq
jnvDxwAs7SYhdgTU+Bi9S0egiXDh09n/5Zi7dx/YXLfLRyHhwQ7puoGNF/97uCYI
tMLZj1sqjdCfLUFKMwDzVCxPqFOxHzMR+btn43q6Cz/1NCZRJyS4/d2jaT7nAy6r
+VIlbtlxU9FJIPFL0Pn+ikZBwppukgUzaEhzCAIC0VVt8vgtooX2A73PNztrr9Hx
Uh1kr8+nJCuQfjIzs7o6uFyeb4pSh0YHK49CgaI5EFUrMYuwcuDqrxKqcgMfbUoe
8PJbR++AEnFwrQHPMB9QLQt4Bdt9XobEFfMM5Hc23P/Q4d9hPGGY4DTKvSaql9ns
6K+fOLLJtb5Hjg5hmKbaFWRLSIGG1QCnpkKkK/u5/VT2PxVZCHD/+CPGtjblF1O2
mbzcCw+NFBsPbihPxZRt0HPwSWZhsa5wWXjNU0yg8yf0YfIBqYP79mIT6uZc5RxT
9cxKLP+mew/EkiC5V8U4Wa05Stzs04rph+2WfMAzRbTmcgY924qKJC3Af2ECf0KZ
KZazHfFDyC9/KEknBDzDyi/7b5RTA8ndblaaqpjwgrbKxoJB/MhNaKUguRyBoYuw
iqAMps5rhCbDVeR++JOJLmk0Q/wssPpeNKK4Aj6NjDVOAi/t/eZeFWZxFIWgXdVL
odHmTs17RmXu3CH5y1ovFksFeADW9j7pSHSJLjxVWC0FekTO20xTxk/fBoxJO9rY
YAA1DBsxt/7JDJJpvjWBer2keHo8ABOg4R9khZxNV71OMh3L0prHHlUxazEyJe4d
Xvk5c1Vtfma12xnvj1G0/xuYQ32ykYLJYtmqiJP5cMtF7JZqWpxHKnoQHdf6yYoH
+NvfKNUe11nOPO8GS0nYBzY5UtjwtW05Hjwesj/Zp54+H1eAWpWpD3c+4+0LN4Ye
gr2uWSPGLgRHdreG9rk0pYkgiPGXQ+Dp3txUoe87NbTVD5T84g/IJM2eZq77GtP1
M1COZyGN1BkveCHoWuxEeoqBj1NPxZC+/AjgNddl10LyhdsvTVAw4sr/81M8CsgL
de4N9QgosTE+ga63go27h6yOpvQ3usN9er2D27Wk6ZcQi9LofoTso2XegUD4S0v7
EEWVgEnU4OIfTOrgGDRuOBT1//UbhkWQuhYQJbvqlyWG01/yj35qlhqDaDcpSwNb
AEdOSoGxy4vU9oqsaqt5Ol65gWMG8rBHetMjLV2KP3CNKw+WMUEQu9KZKqm+E8yS
DiVWFpM9YH+c0j3zlFe+PK8X48se+TbcZ4xfzmPp5887qRgSW/5HFsuP2uKECqoz
T58m65UBgCKOAsD2/LEAGFB/WTYyU4GWt/4uMbkelIqXfv0j1xfIqtp0zTRTooYW
ueC3JXJw4JHGrvMxHrPbPWecwW4x//rRJG1nhFCxWqx66zpaIJoKf57qUB7rMOO2
RRrXRRT1W+unpWUcHoWKJMWhTZdMpuNSEV9IaSKLXNFfEgOPAZoV9aAyy3+UhDpZ
MLzNJreeTSXTYI2wMqXDqdWJAgywAsLirwJTQnI76CYixaTIqTwDVZJ0x9Nl19sb
GkhUxVzeOT786oqbwKC/xyqGwPEp1G4Y5nSejL8ME7Z6UTtjJUmQTRAzN4iSvPZf
nLtOe1PZhvrS8ll+2UuZ4UrncSWvsLuXJvFUMfy2BCQ2WYDUGg092saZvz6qAt2W
01J0QgBXVFQJpjTeXAwMzMhQ3KqRdV8F3vQ4xVXqT44LghadiVaju1zbCqXLfEza
cJWib3LnvGCPgPY5ykk6GMXl252v81HO3br9QvK5rt91VqoEIqiuGe4VP7vbUnKN
SiwZhlXFFD+MSfgPTC4RIgyl3kaOFCnqYhStHQyZXWZriqrdwm+BAl3TTkLDEady
fX+7Y5zJbToiZheUW2ibRqlJHsvVnUbw9WSy5yY9JZspBhpZhPqnfHzrvp0QiKm4
z/7C//UMsUvf31kkfHI9WA+7su0y7rVMXDDM9hkV81+a3SAU79UGDzeQBo+9rkMw
djGOL8IEaOg1QV7wQX9UAKOgkUHIuXH0vtYdOPeYu7e/8Jf6a1xQGhMnFgKPxrMn
4A6WGPUf7mk4R1Yab0Oq+frr/cpFIl/KEjpmP17ZXuG81WTB9IKtKDe7QlOlG1Bg
F1h6+TTnBE4q4TPgd7vFPJExIEyGYnaN/L0S27caofMi4a7/rZlh/6CxSdehebEp
Aw3Sp1vDB9zSPJPiVIKWmISRljWKjFOJh5VrSv5342ifwATThDaESXp3CFPVBwJU
odLz7icicO2Zn9rGAJi83y/a5CISvMqL1DvIMKLbL1ObN5FlI5ATJyJYqXEH87kS
v3srpo+hzq9Aj4urCRTgosJVct01zeokmIHgCMWfO2TLwgQ8psweE7JmRerhCR1X
IMRAElnHFntznZSIEnpxsHfS84H+LCj6DohnYBMdLWgGiVVvdxV4Kb+fDLKJHSaL
H/vR2HDbYmQw7KFLhYh2PwqKVbeLkrvwjE8H5birtOL6/iGIT3f/+JO8ni8reLom
CwDxNVlHckBfTsDwisdVm04oJBqApdspxPsib0r8s72YIB1GVG5u+aDHlqn7ed9H
`protect END_PROTECTED
