`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6MtCENSaXscZIBxyfKENqUdkKNQOFZ+8cFMO3im5HO/1g6+YeLZIT4jdG7gvjVc7
G7cN0RFMJ2qmX+C6Xxo57En/hrz6NaV3gcjV4CJU9Wcnf/vOCge3gXntBrZ6d/5K
XothNQZIqNn5tIq5Vu4nR8zq0BiLXhcguz7B9ebui8VBRacy1//ZIt/e3ES2MxwD
GbY1fDViUe4dkE4y2W8JIv8pmOM3rXJm0Q6EPNq6Xszhm3E946/RDUoFDGLHflw5
nc7J4V34GoC8BtwNoAwHGrpWBR5Y49nMO7wzseumlDDP1iHCUhqFv89g/wRTJgFF
8jkgCp8E1otfwR8xgsK0nDz+Na9N7GK+2KJO13p/QtDgpUNdzzgxr7IyTKCPeeX2
CkFZThmpF/DY4YZEqmXk8/RFekDyqocVrwEylL1A/ulLvdaSgO8ATwmTCDUeoqok
kAbtutvx/4zy71F0DzUEITYtFxYtB+RCH2Ry0bwts3upeg0D++HLGap8eK8OiIjQ
4DViIbeTSTc9nsap/UhX2WkxYEqozuLF6GZxv7cL91zoSwloPLbxqYfIiJrYcNuH
7QecapqcXlrkFZnrxjCn5Z6uCehJj3Km/LTp8RMyvjhnkukiR7y0XXvErKKwSQWD
qh3gNtpCNlhGBpLyqDTzMElO6gl4JGcffHdeumu1mHm7RKLqflzDrUGQDzKR8/wi
TyqKiZ/7eYT3AaJhyp+JBwODOncxgavG/aTy89npOKy0POoJYBtvVynGyaQFP8Wb
AbfeQ1b7vMJkGOq8i70KACXm0h45GabXoyke93iLSfQ8c3MM/DLDNDC/EI+XGDeA
9Iu8ozu9w+gT4Bln63KFku86T8Vy6KrzgRH0rmAD9YmvUXfxqV4/HWEzaIP72ld5
couzyxi0400qQqanUqZ40hw13KbDbVCg6VdCtPm/NkhcF7oT0WgdlhdVI4qnaoD2
93DoywungStT8jMP2wdjZj3MAJaHxBj1H6xBzdO+WIW0gimlkslnKvIYyqqbopsw
VfbuXTKqFuMUUqM6uxB67Hy2DeM31nVAJlxlVjHG1g/zHCQ9OD5dvZcJ76ynjRpm
4QmfBI+Pv27VOjqO26YjDxmy3zvACkWLW/eqccBWKP5QL4gfkpKoht7PnVSgLFW5
srPKKT7SJM3sOwTwPiwHsqNytRZcqS1mieyBT0SLZssocKOs05eoUGHm7begI3ta
LrxMjzeq00/POkXPMi8oLb3Dnr8KIcp/UiZ21bwxK+HKLObSt/rAFOYzHDwObqGR
`protect END_PROTECTED
