`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g/LlHCVzmRSx3meS2Mu4+5CUmK0vvWgWxJ3jN4q56mUsyefQOue7SUtlwRvmqWcH
TXg4BW54OX4FoEZBt8JHDO27yW796uz99+b2OnrYfu3I0xZLwhUV1GT4jgL0xnId
ISK71zEItdVvNuVPkMjXhNMDYMAno6jFgc7xT5PGXhMlwyTu53ftowIUYja/6c3a
YfegOsKkJfaCzuo0Qh/51nhC6g0fd9i9NFfwNFp7zVtrxYHCoSMMJuH6TLoywKAg
xbJtc0L5JFR7t0mbdLOEnkGEzFjR33Y0+JFQBnlmvbSgIPXy9vzDCCC1XpY3opfV
wZXrunqhzG+SbTWI3gwpiBZ6+Sex0qaADOkSQYUk+eCFBr/e5QKY5d7U9gqWxBgp
zpZrWvAzme3VyT4Kt+3YJ13MxAxqOK/cFt7j3CA2SzQ5JtyhBhhVunyBkyjJRDxG
KXYbKeBORFObmi0auAbN6W7f2C0pcUFjc9mOfn6JCMJMIvSdHNkqh7gnxYKqLXPx
92xvJydV4tOMbjOl737fNcy4GsReT1Z+R0vF0V4ozR3FMFwfB5Z4/rGC9LqTPkEu
KNCt4uzfUEF2tXx9zJp2hBcmY/IuF4rATTcjJn3KQo/Mq9WMrEIGvgAnVV+VKFIb
SaetvFjWgw+x+syWT8qkyrUzpfz4PbIrhFcXqraHXCzXkVMuZ8go7GKZmLZwKIVF
oYbb6WSH7Ew1dDnH5JWEi+/XpmixbChpRZgOZO9+V8aMIE1PJp+P28FdGf1+ijrk
NkZ/RkbXi2qUc7zZAQGzQLPObaex4FyO1+a+gq7ROZHoJVj3E7J4WFwUAXODycHq
ZTlD3VC+pnWO9e1GMcPqvQKM2y2PRPnp6mt6jsDyyKL4PtEFxrLP+yP7Qa88IQsR
6TfDqt8P9lAtcqBACHd2fcpwX1Bctdze1cMhDVRGyd3vDBCZgyHd7WE1axUR1Xgp
G3mXfJ9fcPvJ6Jxkk9Q7kYXqWDs0C8HJtC2s7S42AcXh+0G7ETqOA9RS8BRb3Z2e
LgP3BOES+olvKPrPnjPP1ryOwhdGukHlbg56SyH0C8dAeLQtQj6I8mdbhqbbmzys
xMwGegK4N6+R2uKGCkUbGDSZuxlKcdNoZY39JHDV5Sf2ehB8UytDgAbkw9SAHt86
bY33OEl/k9LsH4oibUKczKf3yaUwNYgW2trm840PV8aww3Y3ngu53bIncj30liDO
4BnGOxqACOJvcIhN5Amgd1lihSQQ5AyIg7QxMR/iqHPussAgZNBU0ZXul9+WQ2I6
GcjnZRgyhsSYDhbxeXXOgil09LyF1nS+xp8heV67rojan4mxhcE0+GxjZz+cw/un
tenufIYwBNA72gm/BtiWPVRs+NMqgWs1AGRY0yAFJ0rZ6noAc4xeHT3lhQIz1Jox
M9ndhK/id17zkOObnX4BJeUuEmFa+468fnHJbEACwrv++lS71kIn+1b//HtT8jZ1
KMC/zPXywcatXcZnls4deqkDeSgKFXCIHWf+mfXCg9XOJZuBLNdm3cxIEhH6iK8z
OsSZKMFBvuc5lcztOZ+DeboZg/IlfbaKix4RCsTRqJpnb2V7GjGtL0+vGm5NqRjf
mvEmj//F271CPXIZZsksSrDqDZFpGEpASYvInyTmt0PpnpB3PcRW9r/lk7NErd6Y
iByg5JqBx1qOIn3bK5Knnwrxs5/+RThOTdr4dWbUtALEdlwJ6Y1rNPy582zLsZsz
zPi9O5DVWQYxmEBl1v3+e3O1pyopj23OxFOpTShgRxQ0HI7xnZUD8/ag8fGiVeyW
KYXsxX6nhzIIksIJhS7O+/fxD/fAiF/j0dfnQnI5jmaI3wH1nXF0JSMf+5M7Bcme
dXo6LK1plnK8ya85p7x5PTqRESy0LcU1AoMT6ndwXFKc6ReLzqaQtOAoMI2kIqaC
qwoy3GDqcyB3GtVF4fGOYneURXXu+cSWkiAtHWASytTrtBFNvO0Gyn92brWtKMXk
NjsTKY3x5N+Y/kEUk5P787kQYh+578GjiMC7EiAZQrrilqt4riJxsAeQ/5BrPmpv
ot6rYpo0pxcO194u0ZtKoLYFClj4+yoUdtPhAie5dq0=
`protect END_PROTECTED
