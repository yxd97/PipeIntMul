`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4iHYa68Aor/FeGN5I8xrp2pL5wK065B+x59gLJUi+e+LhUaFXzQ4uYYG2ECySTXh
LraPgf9NPzJ9sDcLs9PINHT8HPTjJN0wfAWO0GlkKCGAZ4xTbxtamQP0Xj5lWpVw
Jg1sINbY60erBD493irU9w0a5S+Sc8jRa9mOJtuEOlSMNOLDpk3mGryM0bcZdCv8
ZYvlUbnj2tsEFzWpUqTrSX/lBF6nLo1KHBhN5TsSqGkq4/FD5w54VerncF70/LjE
2wMuPV8WgKte63QVWgsOemXUdXlyJMX+ICjA6RHw540ZPBHVMbebWGZSy/ulhcAv
kGJ+1+JEHOD+9EDj/PpW7oo6vHkSzcweMPN7rFavTG3k++J4QsZd0fb3HKAozfDg
IPHWloaQtE/MbsYOJjaZ0w2MRjSTiOsq3UdMKKpvpOC11skC3mbpIk4HZdCrWMM8
5h/mtTqvQISMoOJcRRvhChwsHE8bbdK3Pfv0/3VVCjI=
`protect END_PROTECTED
