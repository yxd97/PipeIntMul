`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6uUW5a4om9FC10K2SquAHBDDUXl5Rt5IQ8i1lcQItctSoFPfxv+rRFB9QECRbBQN
ntnCiedfrZ40nNx+tKkaWOi3Rw4g7a50qsp2BPQpkObThgfd7FlJJp20FQl1lQwf
aTmKXkYMxyzz5o+4NOzpTvHcCDhmvDh4mFW4ala+SV+BWjOLdoBFM/C+hyrHnGrS
Fn2+NPAfHD8tPvos2m63YdvlkqdxAf+JNpCzH5zV3364Rx5PrYdGYARzEQ9dx6jW
OYtSQojiSBnUzuCm/wliBGXvz78bRc5GR4pZ0+0/7u43H7DwtocZATYS5Nmms5qm
BZHb5ozUF4Wc9pP5m4xsIcakb6QJEzDk23yMA+k4Picth8lPWHobB30DtS7XNtib
t095XQwdsIf5ypqehNsKItxGKOx/15Dfz3GQNUcKRxRpTyhjB0Ntm7mwYLzppSQa
qguYxQcfrN+1lrC3srwz1Jnrr77TTi4SgPDjQ0ZeFDbnptu+CSmhz1S45ihC2fcv
apLLMqcgkovF0tweGsgDbzQnvzMSVkIb1I91t4S/OVr9wdi7VV9q1TM1RDM/XFyJ
qaAB+Rbed4bmK2KPFOKs2CNH8DEVsCsebycDJACLcjUWBi0JJBrsBCt8/NyVC7Zo
5K3wooh8sXgTIChwpi+TvBvJ3iAdOB1IOOmxqZFzsJWnEq0wdBNphdZqLVrH5W7Z
nZ5Io+Ty7yWeivcBY2xZ4T4nzuBiz2zZ8AEP9CqSUXe6m97fW1Dh8rjty7YB7aTV
CSuNyMNdkCNvBm20Ctiimw==
`protect END_PROTECTED
