`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NpZAiAiFcPuFHDFCgl3qC6cEdbJK6zm4W4LY357kFw3psUR3SWw2hpXjAqHD+gDO
XWdNhCQmObybzvqn3afxDlP9Wa0hin2pXFPmMHC8nWdb+N2nXxQGCUeEfLbJzpSk
QTgA5T/Y3YalWpFeVDZKrNF1xxOP9IP/Kl+FSOOk20tThFs3/T32oBxzTXNsZkEO
i/JM8ArXM2Lt+GHwSZkjWm4TbGb+Ddzn0Q6n/edo79MtcyEqk2wUYFy/BZg+11t+
d3VVpimAyNtney3bgYX4h3/UKLYMphEpRIBZr41OCHhv1A4nibiyWUif1eItzA6a
1J0oDmK33rLAXPmO65rjaBTkXT0dC91evmuw8EDhGbfk00CyfZLiSd5hIDFOzgck
e4Tod50Ax3pQW0MMMfRKytRz9Lk2oppUXnVowuOZoeTxoCQ8KfgQGeeocc9qtoFK
mD04rnq3iYHC0O1pMy31lGgcxmWrcuJNrG+xvudzXBJ5BnzGIDXETMlDsoKt0Rmo
wj8il1SSgsn1zHUnfXOCqpXzwhgP+4uZF94C5flSjoBAi8tpmW+qWyP5izdmXV6c
xvIGWynY1kF164VQwPeHRhO91xpc4zPQQSDvmP0G0pz/80xpI17lDRQ5hsn98ESr
RnKY7w9U5QrRl3IkXloKqreAOpIL22H+mcwwGNlMt3wVNe9itUD31E4/Rey9dD6S
Ha9zD13HSsnZAVTgA75D0HGOhWW8PBlrmlPi2OrXUToQGc9cDV1bp4sp2g4OLDvl
dSxTqiMcCI9vqFEys3lKDQ==
`protect END_PROTECTED
