`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L9XdKpNxOrTBsnxR9VYdcl4tlAoC4evadErO91Kcx6Yt5TKNCTV+LxJs2mn+3xJ0
kQsa1DJY6tBcXfiPaMc+wL3LjJzKtAHW5t4Q2iSIZivpFDkQqDTndp1dbL7NqvT4
4gnRlqv2KCd9d3h66K1VxIadb2mWXdB5ebqybOy9MHVZ3uF/0TpAcwaviakVI1Gw
e2pNehIlSfR+2ajx2uevawOTeN3sxEpC/oQInypfSbbyEgDCpLX9O5O820KjdvVn
Y2aq3HXGKULd3mapfCGT22IWcBf1WiXq4m0Iix+Uw+R3ZvlUH0PNz+PQAthBBlhK
irPg5ZKuuGqYkrwB4rzlTEp9yadDuUKqb3tn8UrYrlp2VWnk0Rm4dh6otvQXJZqd
mO/x97HGX78gq9Vmp9lziQczBcm1J+C3YcU7DyOpog/zcHTQ904SndQl4HcT2euv
uxotrgwfGDsS8UH4IaeLYMjET/lgY74oeCV/U40qHVvpEu792Su5oVE/qHqp0nGe
Q91LBljvmlD1YdGyHpU3/PCHctsUjt017k1LsKIqervmhCcoBk3qStXwNHhqaC7L
`protect END_PROTECTED
