`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jX4YYMdFwKPE7x7FuFnA1GNGJW7LwodJvBKB9Aw2QNdFlD+J6wr+8LSKHOGTPgnb
N2yZEXoBL00hWYCM38pibZUQWm1QeCUmkp/AHacw9UrebBiZNlyVW4A9rKD7ZBN3
hnw31jK9mygkueYTxgWCqioyHxoVE7h2a2ym//emkJT83X6OKun8bdLoOu7qQnNM
1Bb+WIxj9Ox9OmdWb/4TfvpmQ9YV+oQqmcTFRBukgsgxs9shODGot6ZpsDieL4RS
kLQ++qbH7hkeubMkRz5wRdQgWWgiZRDhkOh5knocfU67vXY52bLoWoJNPSTQXy17
zp9JNtSCub44ycM6FFmDMvHBPUnJC4GHAyADJkYtojrEqJRQJw/6WdyMyrtSP9n0
QTPp82E1+lOgrKDXWmnmRATTrNzT1dnoQ7U6BfqQzy3ejIpHLHMgrI5CcJLfb069
briJLo78VcrYXoyEH/4kvc5/4Du5CNLpy17oDm2+G3LrXEXtbt5sAUV3tmCVx4U4
za9b9w06uqkcaSI72KP9Ol7/4PNfuQ/0cbPXn6DEdfYtkmLrnSPBYJsuANWL8k/Q
3wqgdl6swmHzGtjj1QSQ0Y6Xq0ucb5ipQ6Z9iBYVoDGw147Pz7KakDchzfMce349
qqU8iWBcUYTxxVfZw4yrb+tQRczReoCz6gJtzCQZYGZIeaehmbyOh4aM5Q8KFmtx
ems2XuSBrhYPMN1WIdjea0lPbPox2Nvo3J6zZqvU9PG9BTL+iaNmPIftcfDGGkqP
bVYbZZ4eRWm/jQvWhLodtw==
`protect END_PROTECTED
