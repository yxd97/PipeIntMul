`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tnlcckYA5mPA/8YEA1LTk7COG5I30ws/+Zwc6wVN5bbixC3LAHSa4Uw17dzzcvKk
sj++bBWdM/cBEQJ8wrsrzj3aRFJFILXus8dpQFutXIWMEKTeKTFloPD3/ly/vXuS
Dbb2Is3pvKzGudkPIeOnmOOyHL7MOSI+dm02yfsCSMcvEi/Nue4q7X5yAyh+SiOy
11HyoLAhLT/9Gd2Q1EFJfCRwnPzgW+8ULSAur37chMI5rLS1Rzdd9TbSku0xnc+8
ARSm98TAxSv/0EI7jEC3DHn+N4D12rpsSAKU4NV5CPZQcQerMfKuT1nT8E5B5LUg
d4tW8NywoMHYgQIrNBMAfLpoFh9EgpF7IbpKXYLOQs+iU4N7/I5yo6RB1KZEpp7A
FBDdM+QFVSk7ym0Pu7WXIJnBGLbcQlPzHgp2Exdk6ZY4cxUpqjOv4v4hlQkpkAjw
`protect END_PROTECTED
