`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GO9I0ACgaMxhwxyIEKBV7PiLrNocepSu46WAu9K/80CquMV5Ct4VP9TPfCu51QzM
YFr4GAqSjCPabFA2WHfKO1dfuW89t3lxbsJN3fhCj8GJtCZKILWxw4rHVS00cyF/
fB5fI2hO4c7+sZxINNzsb0O0ugOk9WGkDZZM1EEwVfkL3w3yVfu3a4nd/0HdxWcF
2fA+QnjMu8fHI79iwXBom3t6obRCkvjy7/7Kqurxyv8ZIU5bpgx9+FhtqDbWa7FH
9SiaiZotkcqW97qXWD1dBZhwrNzln3rXZ2VMdaUCGb+dN5o3VV/vwjmL4/NQuM1n
dEij3PfFSaUnY1/6Rtg8og==
`protect END_PROTECTED
