`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BJ4FDJ/E+q23bAUSY76wTvH0HSNUYyeXT8Dgq+tI224NPl//He7GLA9q5xG0dD3H
jy6mXGqU3ujlQeVcVNMbRuxWbw1ilxaWl4LnZtkdJOIcNkh/WDB03zMG3DGq+9xN
162zqRz2Q5pnVb98EU739LyZum5Pmc4mx7b61Sobz2lLvEHPuaW7aVt+iQU17qP/
H0oiA6+usWfU6kxj97E/aA1dfvwrPibigtigJ8LjcqpQB3vomgvrS5tGWnK+aKbc
vUno7ISmjaph7oY2tGh0FvuGkY/jIB7WLeVVsIJkSSsmH4sm8rW+vxKW9nw988Em
NvDdlJSYhy1AoCeacmo4AvKabXpW0Ia/t+Lj5blfsBiP7BweVAKL9QxNRD7I2W8L
Tl158kESTJmdkSFYD/DyKF5/GAv9afbl/kszwor77r4=
`protect END_PROTECTED
