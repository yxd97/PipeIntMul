`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lsMBHEqAZVNzX/+9x3LgHDL1RTeP832AGAB6eo2gVOt+9LqVHg0DpMWZjDUmhvnm
eku01N6b7A5mfaJTMLTNx+Q8ULqZ3ZpzNS014T8Jf1OJa87bcgVEnOHoFAT/t7S5
+7kF8Da1d72bXOUpxGhQzzxQEG0UXZWxib4oZlcUo7wvFNXFIIg0cR4Gq01yfIal
qysUhJrqOJpxf+/rUEe1vsLe0Ze06OUZWdpGFzLes+UR4/SjgQG/Jn8hcC0TlEfY
fHVXB9ve+Am38MLOuy7U3vCpxWQhvUWxJCotefYBGeVhhpo1SZT9pJ4Px5y+U16S
XReTvhSlrpmGAUpo67nePI8aptD77+6SvqPAI3XGpUQhPzbKSrEaIGGzOXZXV8bk
rpinhZY6dI+CJQMDVMjdKUXpwSxaovGSGVLbVYAonp8Etrqd2I5mYOUFtk9YP7R+
84G9EUKSGYQcDVD1OUkFHK5yNOTbgfqtvOxIIu+qJNg5gZBWoiQay/eGrMXofEqN
LBEyLu+G+lhwH0iQae3QnqsoMhuW2+yj58M1PgostEo2LtTG4sdFl5T+lPqVpWUe
EhHW7ZKlQe4dGrNZ/nq0mwI2gYgnS4lLuR3dS0t6ACQ=
`protect END_PROTECTED
