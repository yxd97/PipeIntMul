`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67hZQMW+q4+w0/XzPmf8JWp++FxW/F/iZDwgtDy5NCjntM3d/EeYlJg1sd+WxWkn
6NbyDp2mXkt/YdWehCPlPgFOg2G3Fauv/hIAxceXCSvAQtkUhBUTznQuOuP6Dx5O
4wliVZhu38xQSUoqkLhjN9Hekv8ODDIt0O0XgMvB+BiBk+q8GZ8NHlhK5FBFrWG7
lqPG7uV69OQmImJetFNgu8lA8wAu5AE0DbhAsob8PWim4h0rycXueWSwAelm4rhZ
0cM11/oGm/+4aahHL7CHvH8kedO5i8E0J3BZH5VSIqyPianBWe3ZQyg1Ao7HcuMB
OycJaqVugkNZDmSNK1UTpU3RIUFsIkRFvbBA6IEo3YiQK9CFuZK1tmaTLJZhHCyl
7Pux+EgrcHTd6mr7+Tsw24qwXkuNS+D2pjpnR++6S3YXATHLRI4KPKm66RO313wa
Wzms15jt0J4KHGP9qyNK1k4K651IBn/fL7K8KYNZ3+l+h+2tWlBtx8upUp0jBn4+
94R9V4/XF6CQ5D1HbwbuniZrj8MhM1qCh9uMAh0wcZGTEUvGMXKIIhRJ5w3qnsam
`protect END_PROTECTED
