`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6EhjJ7fWpLQZM+xKe/RgYHYh6J/sn36RozfgPa7iJHNR+mzADf9LOWMx+mj1KP6O
l9J1Fpx+ENYWmDHq9xyCPqxFVrorldlm9h4zIcHbayj0M4D0WUBAw0qaiuPU4suX
dCJS8oE5dbtudIHGusgBDmp5/LTjuGXSzOKzVbIYqYa+Ija0FU2UFMbowbxpKGG7
oL4Q4QZX744kU9h0y0N9m0Ey4UNPtNqMLj2Tb2sSukgGXIHX0fC3o0gyg2YYjEUH
Hq/Cqu9+JhpO0ZtodafCBZcJRZNhRBtAWvx29Czt87gcTRz/8N5UTyG0Tn6DU2g1
UBejmInMMq5FYUtP7BWsQwUTHvUVk5yxKTWhNNv1J/RnnYLJROGiudIS76JB7zb/
lMBxl/QrZZeqzRxCY9MPJNm1ekt+tDWI1Txyy/hy4fcFcVMdTvjb+7SXo+yl9wNE
srRdFk3MehmBiruT9ZaY0ZumzLB6zXsPcgOLSLh1akpXLOqfs+R3Ku8ZIuL///X+
AMUQ3cE/tB2OE9vkPE8806ECw3FNP0qb7lo4o8cKk4Rzi+KH6MPhaGhpNV33wC6r
p04uxPwJMwLcIvik+6NGbA4LenSDrlXlcF0/ttElQsy6nKCKvz9avnBfP5rpnp11
8kPYLVdeR5s6fzC8dYtqNlc9XAnpj4kwvN/B1gY3+JjyuhK7P1ujkchQ+US75i+X
hDCJSxtOkRgFpxDaXWrTop7NDOMh5uBNIJLkO1PzswJO+JR9u9qyz2c6OGYFVTK9
o8B2/JY7VZ9YNk/BVdX++KCbXcimhtfb8DMu3Xq04O+Dgdhdmn+Ym+K7gFvDzaqv
cz8R4YszRWnKqx9qqXjnJoxXUnJockSYRLOpPm3I42mER8DFRGDkYavcvkI7/1Ro
Bs6cKt7DeBUR2ZT59fGCjKi4MmPpE5NpyIQiXCoc/fZpvfrUp46v4TQPOzI7YSrA
a4s3QFoHHlXN1dNat6V2u5LAo31ndjizZAiNxa2Cgh1uJ1Ws3sOo7WpBJN63ZA7V
IKYdw0buKfBG6OKHkdWsHediBYvrSlBvFnhoAW3afy55xQ/+FN5FnJE/YkslGdKT
8hvLgYit467ysYQ6V/grWhjeyRtT9m7CiQot1LgAr6ohmUQErwvek7wlCujdRPfu
qy0UoYi5hUYwsJBUNerx9OzwjE2sj40KAAbRBwpyso8AmFzz/uM+lQzIp0v2P3gR
c77mgEtCKs/xTKuqasoUpSU9L3IXF9k5kBVpQ0Cd9EkPxi7cF0ckQ+3Rnr7WX/iZ
LIIIlXGe/D77Z2QB0DM0xdN7DPXGoULAKhK+G8io2X4ipzgNi2SDKVZw3Q/wv52f
YtGBuWJd68AEiAbBYj4xYgSf0JLx99gsBKJc4GCZ8+a6zfbBRnZyuKQuXxLMxB9q
Bi9z1eKeLg8GXL6/Ggb2VSDfXc9dQwl+q2Bmu537jMN451xAlqYzEbaNc+yWNhqH
ELIBXY0giF9LJV9nXH3KVkQk1Z75FWksi2aORuZu63jfM99bxbrl/4gTyco3ijj8
kTNTvPCeEELGMb/BpszK43V8ZXzsAM2jDluYo+fmchuHJyKiPKii6ncS6T4XY9PD
pH2XM535xWIJVSMimF7kZb0MGdGl7ZPsS1qAaZq4aS56EjIb5qdbReTGw88Bja3v
0O6euVh/2H5Owibt4CGgUyKHp0md+uvTQAcSfG3PAgBty6JlZfPC+EZismVj9z4q
zOqZoQ0XSt1if9TPq2Ig3B/C0zoJtJlL+HO/Q91gXkruDlwcjiGlRK6LMiMIjfYt
tZiItqPdF1VOKZswc4Oj18cBG/Oo1vBvBA50t6P9qeZHVFTRbG98Dz1yNx+bUAGS
IFcgt5ZHZ/FEktrVlUAbpf7eAwQmESl4hiHEtkkrVAJDb6DYX4VBe3xNBUfs69HM
w8/uO/+Tw3P3xETYaJ7KZ+tFmMZEQZNWyJDekqx4hQJiQiuC+FLe+49Ur7k6S9lF
En13ZN31FO+WIwy8xX/Uz+jLQ/KNoKiUM6+7mbOqtNg6CQIXw16sTwhGcwHbaCbx
YZQ5TOxm6Oo9JQA25vlSI+MCiKYvlnSwvZboCVYt/+xeXuKwZC3RL6vH/N72tRgJ
LT85gC1/3qjyL6d+iaNWeMdNmePrqHqONDKiOGemqTbexb1+N8i4rkA88oRTFY5G
bTp/CU1ecLA5444HH0LgVb+8T88zqbrMWf9CorH+fpUJjUbWdSa90KUu/k/3Fhb2
g5X51fEkFPGWbBUcGKrb7WuiSaNuADdk8BP34uj7hCJVERRh0VCiLAnkpL5Ie5p4
p0CQomwdMwZZH7SX0clCTDXIZdSwqq1LfJHCy4sLtMlHE+KNOl9bRQKIZXpPzNK1
bwm48NnTgjA2VFFnLpwxIk/RpCyMyBxRn9AFBGnhu1cH2vNnaU+EPQylkVQC3mds
DnSbFE4ZrxRYarHBtJ9fEkm/r12ty78CKGRkKiAhL095W75AWO7p85wnHUIK4ueb
enEgDEbsywPLNUng25C8DYCv5CxWMnYWu/f4nccPm0ksbYG++bkg+Fwpmb4Lwt7w
C9tM1rczsvFsLOxsTnxClOu+vS5SxZLfqv4kyGLERGJd6P173Q5yG2OTNuttQGmm
juFiMJXgVsIBmklGeVc8gW28VjEw0yJg/usGU/A2DmhTs8xF3cpe7y6BTnJrkJRA
taaE3TFGKi+XK3dmLm0QTU2LRA9H4k/d1k1ScDw0V6gc78hkE+N7oaZEZq1m8gSt
Mv4c7dbgQl8gZz+jGCl3wEbrANE9IU8LiyqDZ5+cOGVNPuLsfqlrHk1fm7vhmsRQ
BxClbVPobzF38vpsCILL1/tw0dSp2bTdZbCi6ST97xY2XmcvN5r8MOa/AI0c6ucy
A4oFZ8wql6kPNqUO/C/PaU7/OGVk/2TKog5doSrF3utM9RxtGqI2VQh/iOizzJml
PSdPqk1O3Kmh8ZamdZLT6E9Lq3htV+GTtVAF/n9RaozrWLa9To2M4OsWZVnexeXS
HAEktuu9b3K02F+tEyMJyTWwuqWNMdgV1OVjInAFlSdfmttdFULrDv1NzFqqfbD+
4PniY6bG+PpH7UXOUDKoGtGw77Uv1RzvQWPXTWIIBRP4ZGzbrZxPaMAo80Q4gGU7
DXrX8vmkdos1EnlwmVy3hUeoq9ONhLZ5utZdVimRdxo8TE86oSNSKF+ydpTnrr9X
4qZOy6YVH68dZUz0O2CbiNTDrPLuRVjY407xy9056pQMQ9T3qk4nSll7zSROinNa
HMxpZsH/yJwQ6xkSi3Asiy1yl1yB1+gMAUPnJXa/BzLpMM5CgEqUMtzyUci82mTy
TvIRGPukDj1riEOnPDfa1gQ4EoUekDGCclIrfpgg3SYVX3Nst3eFkVpX98ZTGaee
Pdoct7O1CGqMp9hDeX8NNpQaTG8pK6JqnlYVnBOnudo7W8bAhnIn+am0T5pXqqEK
dyQSnosBasyhitd35T+mq/GxjAQARo44yy4vGnV6mERXpMwK2+N17AowuFRf7l6u
WoBkssEWYxoMVyOF09oZJ6RJDiAD00HGp2xLMI9jaOaN5/2cnpc/u1GzGHP3lupc
2Cf4OVKmfupyPfYTBJWJlekCLPq/Wez5F52ZZC9tiMGUKLO8jvSgAECcHTCVHvuz
3FABH3S5HJbHFqKCi8QObaGK+AcWs8jiS0TKzZ3X+xL68xaqO2HP7wQK3Dqv7NWP
QH5kc+qNyPdQAAjtfNIGjeoXo9SsF5bs1uiGq9I3fUfEAcYn4FgbPwh1erf4j9ES
vdEoWwuaG+u6nYfYgD5/iHV8xH8uZXuNCgfhClb34wnJdvuivjbBGcinA8Cgw7Sx
RThh5LC0UTkCoUUxQShUrnq5wT5VSQ6rYiiXG/tu8YusqN/L0OJX4cBaqwjCdpgW
b/7SYRbmzUf6CCHs1KAZtgF+78nVxzRSDtrTMV2zCXz79LgQTWe2EjdH1Udp8ONl
iEFIsR3556XMX4PbYFkdU/aM9D4188ClaHUrZQW/x4Yzf1R4gE5LY/5hCCj+gDps
pyq3JfQPWTIhh1EAnuuWQy2sqN5p1TeccVBNiPvuU4wHXjlZ5U48Un77xcc+fLbU
4ZQ5vXCiRhJY11Ngrvw7HEU329cWBuLC0IC0ldCwQFHyBbmgfcKAWEQQQp7QhUcG
HTJHMJ22x9DtWAvup65K7sLMJl2zD5gOI/3nCxuT7/LvNzujgVJwaBlNFHSiSYmG
eBocHvStS/Ace3H8dUxcPaU6/g+2SLhBukBPZRDPr0Ja9NaUGumoFxLNW2gEPPRR
I27YRtLfaDXpuvPbkrMAS+Q9icRSj4wKdl3me2X0nYUjFwxRgx4QUt0CN3yzLqL4
gCo4/Ds5XdjiG4VJHF8YxNnXlCkkEytR60ZErZMDhIAZhDwe3sSOsYX6h06dz1s2
aOK+QFf5qs06NnAWAtk48tK1arq4HSr67weU8iZlfms8zOH2THuKWNT8Zzn9faQx
cO74NGxgpcAg1XdyOOU3/ZrS+gEerYAZnVG3antszEjsmwcrj1oktJ+RQ2Kp9DJ6
toKKOIXt89Kud0znFkUlOcpXmlkcfAbHyrQPEHAXUgTKkMtRMUnfLJIwfS5PUkzI
vXVmlxXdFMgnGC+gXSqBGNzqmfmFcN/zf8p7MvoHEZmqfzEccqgajvrJyxYmzSLg
cweEIDF/Yprt3VoiqcNulWhop/Ej+uLwodHxea1ukaxWlz9W+P39SCMJmdhxg8Gk
qVBlip2j3IM5FLgQVSBniRcvEbP0yas2ToidAl435gb5c2jELBGFR9CHKFf4aQli
SVGjl9p0shXaz6GpLJyg56nSsFkAvf1YeBLrPhQU93DbizMZIZTaTPLqFuouioE5
kwbvFCfpb1kmtV4BxCikBqyoqU3k6N09CxMskccYAK8BXzTvR/qdlhGTrPphnjg8
KTluu7/SdmtOKkhhVI7wQVnzS2AuWIpb+TcV1nt/Y9tXmJ9/g+UfxE9omTamw9R8
XUODg7tjcDPW4NSOMZfb8zt7z1sjXtYMD6/U7g6AR2VrZ5XxVuUH7iM9okHTxfj0
xv/aUcA+kaA+0wZfdDEvn4VdujZVWSlLOo2FHiSkSVgcKns60KT9yBsMA409RcIv
YjsLInryT3kXg9KYpONAC42977CKZpnVn3Dma2eqB1+1kkTVKboggr7UnSYBOCSH
99hSPKB5GWSJAfWGnmuUcK6leN8GNt0y0dAv9ENf3ZQYgjhnyFk9Dj4nrBGmsOSa
BEAAPkduhsW7Ih+L3mMYK8ZPr4DYhAd7FnS6webIkJ1Kzb8qLRkPgiu0OtLerqdg
ltVWIy9wsJgniwOR8Af7b7crGJ8JmajaSxM+Fs2DuioThHmB2WQXw+yKZ11lSaeW
5ogr+zfXF+7ykAZhX6n3CHKPJEIKng+e+r/qIyDIiSt7UufZlAYPl+M19FX97Xhn
sJTs7yASkfMtNL6QPka5WhsFHYoc/t9IUJE1nEnm9x0nRqK9IdKLIacQePybUz8l
ssp0HA3bTswKsgvWDbBQVdSKruSkCt11kL0rMjcI7GuwHVkjSMcq2ZlIo0xMeI11
DIldIdq64dt3oeAkWfokIuWPyG1KI+qL/KI4CI1O3dS4ozJU1+qkmJIfkoD0Akxl
UZJpjd0qEvK1Oew1A9fU+d0I5xq61ao1eBoQE4Z5S0GYltpufzGzsxIxCwr237Mf
Aor7IkVhemqwDTkCM5AwhKwQ6KTozf8Knp5e3TTJb4ayFr6BGEUW9NC5OIJhZy8v
1ohbbZ2t1+q5ZDUYA8oatPP99fGbusjvJFXVhTUbLsoYeJFiYFq4Gj8qXbK8gdS9
dE/viu3MMHZds1I+7zg7OwyslKUHsk0aGPhB7R7e3HWU5HtMMbkC/Qm0cCgke8FB
ojF84V89OXutwRtDYoNnjKYAcHuy6FkuNCsp7oomUIjh5E8ueeI40PhD9+fy3uJl
EH3f/ZiBULVXf5rYjODJLkKuXrccNm7MdZRsYZBjYnpyiusqi2ptYQUWRftcd176
sPxTLaaff+YajZ1kLv8p9HCYGiHeNMalFeuL/zZB7SK4Z44eG9oFLi7ZE+Wbiy34
1Ztu5QID6jVj5ymmi8e1otVFJI2NHOfsBb7TWfHGXfbRGDw/vHP+f0Yqt2EQDkg2
7ycYE+ZFheS2PuPEOAEniqHDNb8R10y3sp43PAxSzyAnYs158hrTgVeAVgOIBVdb
heZM+ngf3l1nDMFG4nd6qLqmXhfbZzodyY+vkr26ULZRGoD1PuH43Cgx7PMmxKiz
1bA53cU7bzJIPCDbZh61ks3PjsGeNH3pKAQHQJLfz8GMwZCXoJYw6xymaTdipuOg
QQu6u4TLvCGlCSUK734W8Mnny+3m2RrLFMztB+wP2ZwB7OEZMMagDtjsfRTFBhJ/
V5cqgnZ0z4oMj3W6nIqAT/aRZ7PrHhgQNGaupOzWmU/qRnwZ4sWyYEiudluIUxW/
bgqIxc/4Xaq5jw9RH7IM8AOJMCx3G7NXiNjsYZ1/amz2nwAdWLmhOEb0L2O4VhNG
mx4NV1ptnozYXFKsVQLk2qSXynclgsThV1055tJnPUzclf0BqS37zShFxoQ7QXq2
dqqxRDf2SbHI+tg49vyLPQ9AKLnGmAniPS7zWgpy1npTDCGSXlW8mda/byYG1BlE
F7SkEqaJWeWkTKBY2jXkH8WW6Z+boXPUGKoaTmwLSjqWjpDgyBtly7OA1af1jULU
P0XEie4o+uk5fNvGns4tOiUdMt8mc5EpgLUwj05El1D1BASNliGBRC3tzxlFTwew
sXwQIS9ETjP0Y/wPFscM0+rWuWcDzTQpAogqonLZEHJ3V4RDnvuqEhOpjkc5Wzjx
RtSvuqvsZAL19NLuw+0IjCoY3gn/frj2/XlB77R3WpFXfyoNSbClYWui3o4KXKI5
zbcdcLxCytVUkSS9AKgMmeTXR2hwLQIOoqISBxePB5fLdHNbCS6l8F1CYf8HWqMA
N8u92Vf19SZU5YAsNMMoPPy+FvxY4nmRUImV41b2TQx3dArixBZoA6eB/OHkC90+
VIui+924d6OIWjl3swNeNzQBzoOVMlb1PvHo/GA+jspRJfBGNHpmPN2bJSFBWH3l
G27MHNkDKw8+08sOzGVDNaH5mAxzZphjy3Veg63Hv4FDCuYg2EPx20hdmEsLSM1s
F7c6vRJCGRqfoJz5lj+or6fYIRgUhVw6949HNASkBSrRNBREoDdcZydXSrHhYk24
3ZlaMIdIGo0HxOVG4NnAHiiIiENRHhHsPCg9uDmwsLrXlLAFt1nKFNCB90zvQC0y
3hRZCqIB675QK3OyslqIZOh+44nl+ldZU5NMOYVcQnV39D5f8AhcApMT/Sg6dA6c
vIxloNyUKpz4fsf4m99/gAf6uJbj8wMsSDXAZUGjagq9+uwCTBoUWpSebuhOW9x6
iBqmTRjjGxqIQgBeUaKYPfBOx92zywTIc8y9xHvpaIq33R7m/UpnOE+C8Txo7cSj
KeGKtzpe+Y3C5swhBwPJ7dgldh3kBaWtKcqjM8lJDI2Fsguy2zpGV81w+zbGwnRO
e4uyK20ZjJCWgbC8u/E4oQFurIFudkEm2P6n9VWKH/aEGjCF+zLjO+Q75kOIC8QL
ak51VQ/gZdMywLcFCUxycMrO0Ep4aSly37YqUSVS3cSwvNGv2ovUeErfE/X54bZF
ILjvFBTmikJPsuSFb2KNkM0BM8KpdMqsXWLAXmLfBL9JpHWEqa2NU6Vcap84zLqD
y1lREJRh1/P8vCMVk4u8TO7oVUS1a4THg6+NXFiIxTqxbeJzUs4tDb57Aniwmo3y
0Gv1ooj8nLOKERHNgxh328qcNFxsCxsRCl/YoqFTGUf9Yd8QeNK7xiIiObUx1qCV
ba+iuy/pciDQIyhBKj9ZpPOd00Kn6rPHxE8l8J/dva71gTA3q+2pzT6qIOiRiTv6
BmOJoJiI/LRmztQTgAN3YnQ+e6McxiBaCk8f80G0njSklKEThkZs0azDpwIatHh9
Xyfmcf/+QAxFSmnn+ZCPf4PfZO4A/h0LPGMjaTlMJ3np3rOCZybV3r/EdthX9WqZ
5pHQsVYu2gM1BBuGPEUjaIcQ81HjRbc/RQlYK/itLSAyuUo1oOLQ27SzQPJ9bh3m
AuK+PMLhAgjCoyIs+YfNQZSY7Cx6blLayqPW5Lw+nEWvf3gP5EgbhZNghlznwgq5
C7QSAB+o5lhTMja2XsA68QP4NvB2vdRx7wHe0kttbwWqr4tQwLaIVC6wPCDQ37LB
gqGkuXOg8CLgEKytM/NUCoT1Q1+xQfu3PUEy7G5j4AQWyjeTLEyH2DzC0bsAwuiG
FPVjE2Dz2K0slgYnZPHNqZb1Qru3NJ40UkH6ANWjRTS3fw6k/h5vx+dRRZWny49k
ch6K335Wf9vHqpR8olAR4uMtBr5F4w9Xe4HFRZ7RLib8yeTVOshOi5Dm4a1vzTUT
3/ore+elnoPWt4biVaBE2ab8tu9l8CnrJyP2uBuT037xrXxksVZOk311+S9d0Mh2
C6LX49otYAUc/GfK+XcnyhaLw5grBZx3RNuC0jzCzCR532S8bwuOL5N0mmM80O6q
slQbai4mWt9vxI7LGjrkzeYxu9R4NNJbHYeDrz4CbRsL5ODOQNCX3ZT0dWoIRwDV
Uybhj6CCc9sEgs7lBXiVPnZmarSr4nLdt/JFyCZ9qzH+V1pfF5rYX3o3cpQZ04Fh
H3yiWyZNf2LXWW7HyCaPHw==
`protect END_PROTECTED
