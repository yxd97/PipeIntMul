`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vurz17T5WzMS7GOJWRrL/JmJ48av5MEleJkQZKS1G7Y85t26oORsepw0dfgR0jql
6GcRuTtf2SOtV4nGkyJmu4YLGUx09s9vJ0Gcbjzy57I4JLA0t08okOFFscYJFKPC
LquUrnoa/her35zFfYnAm0DF6rGXb8mwiMw/MwLGID65G34mAQJWVCqdaTgUZA+X
PMwKHB5zyLKTnNaa4Nvd9aA2Ct+DuIR9QzoM5NbAXFewMevAGEbK04pnEzU/zJDN
3maTq2irGiwxDVw5WoIN7AIYsb7+e09igk5iN27j+3owbTCN5o11f6A53FnMLAv5
rj9NPk+x4dd8aof4H4Y1Pg==
`protect END_PROTECTED
