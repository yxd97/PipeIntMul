`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5CqcgHPWo/XYTzTypHO4VMHeg2uSoAsvg1Sj+hw8/k3mMYAmdZFKz30aT8iAXvWu
95owIqjnaqI0/zPCKBJMxCqoN9FaQvSKqPfAWzTARYxbtSf6rk/RfBOYYCzs9GVS
PrsjGAIIRSI80BMAmHtUH3NwL6diZk3Iq317cGKBRIhkvfxVxnQZW1GBMorpHpnc
0YnKpRClij3Cf/DszV0C3+Z977acNSacz8GVN7XAy5k3XFd3bHa11ctsG9tUVtXd
rirIXIjfr0Io/R0RSSVuQ4yrx1vgBTG/Le1pZZRQ6Adt3+T6/nQ6AvGAq4dpC6n6
vyxyKP0YaNBPdxw40W0I2K/nk4JVfRPE1c/GB3+Eq+YZcohf3AnMoLW6m+Ro4ZaQ
fUvyf52JZS0JeVQ+bDqX7t4BL0OOfGiZdiX7q0IQAGvLYW6YVNs9PnFgqWRlksRx
VTLznrPsq5tuJw59OgzC4sClj+8zVnuNFw0sqyweDgTHBJcSMX/pMwIi2K92ldUN
K2V2I2VLsCw5Jjypl3dhjael4B1DPeIbrBGADF4vJ1j5jVk/kS5On+/m4kLA2EKh
2uHNPLrCV7Jc3SCubIVNEFTgYcS2yRQTegaouXvdQYATDDAFxer/VFyT889FJNN3
DIxAbhjp3Y0I60CpzXljVQv4CFY+xUTtLq+/TRiWRSuFwg7wP3dH78SKzaUv2rRb
NpNji2u9GZNdkv+7ymyqEFv2/BJrrh+v4ZdRdmMaeJk90lqY26WSNxNf6S8JyPwJ
iqhLC+3rqmfuyPcUpoPifIt3ax3iD/4bhUzfarH++iQN9FZdsK3G+E6fDlK7hOSm
tnzgSj28F/MtdpGPwYC9OLtIAj1sXMmUlTowS8T+8ji6G0yaBZ9S4AqsHcy3huvS
UtnfDMb7CGl85rbNMrAHwoXrmnN8IVr5ZYxt2viHPRVkXVVsYqqbluhCYh9gPBum
H+k11AxzC//7BGK92Bw+tV/jD9GUbvXxEBhl802wP/njPYEnzguqNqXW5LmWbLPz
/4vHBtW8i0HaMnoNWXv47ympaPqbbTWGWcMiKvPOP1gESIxxGtFbqOm1xzVJhmUQ
hx4cfaPKRA6UVAYv26Tl4YNWxSuX+Ik8jzmVSJ7bU1YfYmc1+uf+VgsDG5dn6qlo
rT8p73oWxmGXuIzjIrFgkv2erQGpQJNK/nifv5lYN+uhcQVvBI0uDqssLfcsOdxe
9DKKdG3hz+coxCOtJ75AYRtXJHOR9s63szLSEmVvR89Smcg16rL9IaHUHCX+mRwd
avabJyCMf/OADtTBIkCKSuVUNxmEdNr1u97D1xObsijdeiFilB0BzVwhrpMhxnZc
Ht2no+YcaC3Tbvm33F3cCnDXbRmZ0dUS0fVpOt1pfrivdksiIfETLknQdC3WRobG
LmTeBB7/IZ/T1Yt8cWI5Iu9t1hbrFWB8ttspPCNpKY+6oSQWjSxni/p77bOQlVPo
DbPmdiZ3s+41bDnOZeEuzD0LfxBvX9tIU2gt2lE62xduroCzACHrRQZGLN5+daIo
wRhQO1bECOKVYK6w2m7Rw5RmLGwTCStk8o7V1MsS2kX9e9B0SzcswiZlL6GMfwwd
LzMno+4Q3cU5sQRpcAjZzPgdIvhx5GZc9TzO78GrnX/Wl66k8dtCmSPFaxNrOGjr
GmDoX4X9asr9Sxql8kd5wpRcOsEuf2L3ggVePEGzwyGsecgIFybMM3hERqpqh9K7
oNpoKs4Hd3tNT1eEmbiBOSPVYPYpH1ppNvPdgxqWIMO0btXtfATXUNRrxq54bETd
vpjQYqjIMMEw7YzXwlt9mNbgdxvyYvlrHO8GmRFio1SsLATwUu7lG/I8fpfyVQQt
X6c1wzOnun3+kGSX0Frf1KxAcvf8+GS5z7gImPQ47m5iSS4W/icgww5IPFnGsDjk
jaUC4UUD4uJmqime9WUWXbwV4X9cTO8dF6k6k8X/wfWoURsZWH3rwME6GC+RQ/a+
pX0WoBWjAYmEfYJP0rT8x2dDxRE8AZ3pg8I7wYLAx88wslxgWdcuT8TBfeF+vE2/
+tjFlG6PhGNVjOAsyEY62YwSgBUKaUnEXndpJrHiEDih12uXOaQLZP2asv4W1MV1
JZnuP+zEgDHbl+Jn987F984mSg9IoAcbHxEclpjqM0QyXTQxJUEnqKy1pZi4F3Gc
rJGWt3hvrCOv2ldqNr/eVJtxnYiWWp2n6EHLskTvRzGG2++hlTL1Dxbyr2ZoMJ13
Yb6Zy7VfGHJ1exyfJ27XrHWWBWLGzwTmI9Z1XckxU60pq6OIJt5fVbLIAgCy2KNv
s/XY4eggbWOgzR18zLBX+JKAGjRUmkYCH7kPVVO6GVk+QbhZKm6TYnw6sdV4kObj
na0YFmbNpqY/Vjeog1bbuQWXShXvx8pgOZ/yJTGzEJP05fev/rXo4DbgowPTACfV
gpxhgBQGEzTk3GlHSKMyTpis4B6lmSzIvL4uZnVEqFQGkrKgKmlYWgHFCsA7SHMc
ViBaOXIYKImtGzA4z6KsC3aNXcO2eBEmH46VWhahO0ZpoMZvtPwIKX7nIj46TZvQ
Xv5wFPcW8Ynim+HPH35pSA0TuUi+MwNXGxszKGpX+3laom5/4+ECAmpmRVUo/qXJ
2Bu96cwkXChFaiXb41sT8OTG42n569GSoiAEi7r3HB670rHE02rQTYf5ygTnuRln
RuFjGVzVy6Np0paORRNP9G+NaKv/0uqIZauqPzRmQy1lUebckOdzKZ3vdEOfkuRl
tco1VAEvB/izuV/AH9OLm8ThSZ9rOP8u5v1Eg3vI8r7LzvMMpDEtLoeJ9reOiXKF
QyfZGhRdHW8W8GzfYCYPpcLonyyx7OLCLwT5rdMYJhdrWKgdetMMUkeNcW2QqsHR
r6eJyg9wmqqoHwDHIw2KzfG49zV+bEMmLarXDe3cRUkDe0r1+iBtwen6P6CtPeRb
jZ23N7Rwye05Q6CCzJ9E9JIeOJeMDPHiYAdpZ5mwlVZyqaCxwBL0Ikk+PHFWW3iG
XAfwA0DLziR37BQalYtyBD+0a6dNt5VpnPK5FS41S1TRd4I+pT2GXAT9M4ZeH6ec
1smwj1StfTMhbv3T6Mcx5DY8/xNfkCX0pMuWmz+/0tywXymYCKjE7jgzhwW+dvau
XQ2uhQuV4Sl0L4Pose/OlxOO9Ew0p8wsqUJnm7El9v753pq5zdpcImLPBtWgL49E
pl2XeexMJaMvBsE73XfSrocnVk0mpeJS58ksH5Y5huM5Quj8JuyJi785VCqX/vjd
NB9cB0VeGUkuwpJpWb9zPL0JiM7GnGTrBPo5zqoKo5cJwa1bmctkPgtBIe2sCVs+
UaKL4V9L/FEK7jqvWyLVpOHivX9g2ZQh9/C9xKZCYGCFWty54Q19DZjFlG5EC/MV
Z4p0MaNZR8FMhylkrVIa2h3PN1iGUl6brLNHliVXEAD09qqmkLlqIUAgCO7NF8g8
4Yi9E6tL2v11bOwLvfliahZF6Nk/EfW9bvxjGhx8q3kSf3oNWTnDCfkvQxa/gr5u
YdSHRrOaa0w7XWzm7eDUHi6zFaN1wfbdkRBQltpuo5cmJm1xsXyOdkTFBHij9GX3
bJ1+cOiRamNYV7RZWXup1VUiSPsiMgXeJSI477aKep98QpBRKzuyhRn5b6JhZcsV
QsHLVPJQqxwWBGQHArPLBQOn5bsfT1HMa3pqYF2Z05m77Fa3Hdunu3CPsjzlCMOW
0UrMoI9VvszkD54anx1hcyCTimfVeWDWVIykRILKecpqFvBzYhBFz3AZyxRzkXx6
3a+r7H5rpJRY1xqQ7eAHbMVTj73uBsifgACX7tNHadw5deHsewglxNWz0GrrSmma
SjRg8RRdBngLtvqVYznSsjdUbkTw34nCRMR6lWE6C3JHktcP0OTVBSQb8JTcdyDL
2SPXI1GljB/fwTcGOXHAALEC9sLseZ6fRx4q+BXneuINO7QOHx/qORtvYMPIEA5d
+firWPhK40awFDPv00qiOJrir4AoB7QE/BSMQmYgbxs/DW9wxJahiyI5gM6D3qMR
73MByAUn+/xrQmmBuATnSq2W2MjknMYFLX2BDUmqX/q7k5DASPBhxyjtUc3E1UnU
RfSr3pRbV+YeuXz66HQausX/mcmZWPxfJ8N3rx1+j/9Kxp6awHKXty+FWa+5Vv3f
acZHJbWxIlSe0wFDuh2h/cXdBmcXqQk9to9UrizOQFgenaKfzW2tIrAgt/sJtgye
JtaSxWSxELs3bZULV3kQDLnZKC+vL7MiaKOX/flFSAY01qYZ1tLudOcj+Csg9jLf
+pBD5n0UMxRr8ilrdBz3hgN94pZ57AukkEqjstX5AZil/zGF7xTJjOMoV6JXuvbn
diIORVUPzA5GfJTWA/r/rq5yH8nlqMenFGDpOx0dpCgUxLleET7ZCIpZQlGtW8ev
Q491+xy2BBvsALiglIQT1iDd/0v0esqzMtKnTFgrOCSaSVusO+e8IqBTe4q17XOh
WJLH2Ti+BWTTvPpacRARc51qTX1TaFsc+mubKWYRXXWha1xFaDnOx2mZ3JiTT6BB
hmZBv0sfYg2Deo4KdGprrP34ICAEQZBS6aX0QlJYRpqA6AesHJOoxIb9Qu5DDMo4
y55+SOF+4+6CGV/JaCYiuUNi+myp1yWoaQvUGJPMYHS96WU1/I3/KpUi70La3VvJ
a+IAKDGfVy+KN/9ol+Yc+65Ezpm6MFXc1KXMm0UwG7knpI9VKhoZWENimN+MGrFb
RUmLvBXRnrVaO5dAAsrVs7TgfXDjaUrw9iss1mGGeOHXVoLQzkuAmx9FDHyvw6nS
p2VSeiIOKf12xto6URct8kklwhJl+sn2LVbVAIooVJqae4DfWUnjfLXowu/Yqfgj
ZQGE5n1yPop5FP+X7fhO1nJ2GIOgpKrV+SukaAnYm4W9nBZqosg1m5CnQR6cejKo
aaU4/PZKgOSUbsIFLwc1+GedkGylvh368YryNoBJ7Kq1PvKP5Dys0R7lYih7CUyD
rDVTwdKEyri/tSo4jXHd+feWqyC7gKS1rsnWSYHP6cZIN1PD8vlC4aEB9jU7zkNC
ZR6wyoy06u+qSkVicHwpx3UnfTGJ72pK0KfQSorZCOfEBT5vLEHqLw5t8Rkj+lL9
fggMmPW0VLmpkLsNlbYp1KmQUbDcsYdGJzilgC/d6p8vtq2up5yVt8fBhwXgb0/q
fp+3ioYiyS68rJ/bX/uI6PvVhDXFCj2JRrm8CRSOwJGwA1kvaKq2pu5C7ynSmwAo
Ke8S+Xe1C6PNr+9azJq4WhFMw7jE/YPlIJEdYVV5nwWxJXqQMJLbQPSz3i6WHbvg
HBA9a61iRr1BbccB7JOonbX5egwB4lsZzj0q58qi1VHBIiEBIhDyMUkBv9kRTZPu
wPgPetgksHCVvAT6NiNegzCLg0qZZUaFLtkJcPdZCULMYTT8/HS4O1Ogx+caQRkD
qJ/6H3HkViFG3Mjgd4kULNpSyuwJSykh97F5ewLULomYp3Y8XqZbgkiQfDKmkihu
6UE9pHxnES//wLJcZyBxtQSR60ObYa4a9rwJ8ohSwYioL6ffFPZ/L1JTbChKFJjq
D16qoO/4/JcNt8J7N8wVJCMSpv8D8rX1lPkTwTELsv/xFW2o2np1ASqc2uvZsgnV
4ZLNu6Oiojg7HO60VkytShVOQwzbp91J3NQDE7vXrW3cAcmvb/8hszsPXZB4+KFE
vCqnBbs8jZ7dNe/GmczQv612f2BtnGl1IgW/sksHUsK04k89iX9y5rmgRTUDubsI
3yw1rl4JxJxgt1Ed0PVIVcX5PKiGJcXyDTYSo5qWhZTs7pQHLdlq7QAQOhx8pGVm
AIZdHBXLI5Szfxyf8humYsY7ExEhEbWDo40NXBfoPHYbWba90+gengoSAEevpvpB
x2qloM+p+9LEeXg9WMg1sCtcQD8At+lU67jzI/wcWuMCU3MuiCdUEmTziSC/BErF
10uhJn5THXaqm9+c1ICuX4Wrjhn1+FA2PmWWP+LqPvrR5rjdJHHeEXLZvBzwONzQ
qb1YFDvtb6t5a0cjZHleihQUdOewSU6HClhBqZyL+beBHjmTrxYUETG28gMGtxHY
Ga2jClxpvkdIGYy+dk/XbVmEFvYNdR5Lk4/QFfdaw/EjlQJix2gppLN2QdjMEmZ5
Q3ldqdi8jEjOWttSTGPeP14c7QNxMxImCxSV6yVSFsCbTh6xVBJsFQtoDG2+Ii6T
Z4kbfNPYuC4Y0H0w4mb1N0RpqpX0Icftqq5SssopxSpd0PrXqM7LDj/5wsYjqLKC
FnEvN9/rpawStxmbQ+ZZkFv+FXP/kQSv2KPtjQk0mOUuSo7J1bK+yPwi0LdBpbft
LyQYj+G42drOT/tCOIwRDvgFEiPR9nZQO62URSx3+53kr4xdt8dVY5+uY8ZYXD3O
1oQcjD21nGorRFXH1TkTMZen9ZiafdhxlJtpWeM0tQbMrZQ9MtqJ85LcLuXMON2X
enVEjtrBAkhd7H54uqbt7DBFfTe/z7QE4VhAQrsqd4wiyICs+1kW/7mIInqtmGaS
dgbVzMSxp0HpZvFFTTPTpib7SoSv11CdzKFlYi4GVfIJo5QamjiQCKJg11whgqRo
NH0X29O0jSdQVJ6vA2Vl/R9HiGBBJN9Mp5A4+aRSJv0x3ejift70s/867UJHeg96
FIrg+N0kNGiF+gAj1mD2JV/p+5O0aIJIEADmlYMoxB2OkUgE8X+qUIprp3aOTMOZ
kE8SxHNi3Hr3+hqa5LrhC68cD/EazSVf4+LX0FMRRsmUhTo357s/leIPoshPXBgf
uilf/hFYrHQBQQgOKmWLtJUOpPAxy6RkMFDcFcRP4N3Zt1AtnMFZYcHvsMT6Vkrt
1URvz3E48trg/lpFcAvQ2juCN3Y6HoeRB28d7NBGl9v5gufbyYP4Rg4t2X+zNdbS
Kzg+QaEzC76RnuK58oplqrxKB/4FRryNb/i+obNfS3N4xcPRcm/dNWWqnS8gzJxb
iMEQPdvewEJuyxsd9yN6mWZDoKeRXYbyyDmygeOMhumJjHVmw/Z9OklGZzNNhSQg
qywtGcfT83U6K/8SWKk5VIomGG+5e0IVM03dVJsdfML4pEhB5a1CRf4f8d9nnhpy
OQM5wZ7t/4Glb+90GnzX1y9TUA+JQbH+7lY5ziJSEtZW4DyK09iGNZXU9OilPFs/
nCcHypse4IhIW6zPeTWjsnAICvGokmEBQf4xqae3h3D6Hspy04UnOHCdPgdt977y
fgrfN0ZbBKUkhUc0+RsdCICAB/NeP/rhHqwz9duIrTnXlYu44iZt60wFkoRvYd1x
ni6XvoOtW1/zg4DMOi/eZ9E8jVuZolzf+2LGzC5m6qtd/rOY1C+ZDgG+U2qGNq2c
zsrtQnRMdN0qbR6ne16kmOtCTO2NLWpY6aHReiMu++J+qgo5OnPGw+/CH+cW7V0E
69/pGrSlnSvTNR6tp2j8zqa2qoMc2j4j1tAfxsLe0Qf9kic84ITieU4S8lYYoRM2
gFFi6OsQ2xkqwahOi9AiOzlv1HirVwjQFNTTJwuu4fke0BlOO3Gvdies2j4GnuyW
NkSrLoGt2UABMaaa9HDPDNqmv8elIsCOiFphROan7vxO6JqqQfrx0bNFxE930xKR
mMInhupjV5Q5YDGZEIq0BPYu50fVLmdnxQ0fRnJSDtgHW9ig3MJKB4k0eYo+vkq1
qclYiyNOPCzCfarNmtUws6KZt1rCr43iL3RomlQ+pIxh/8xL82dJotvmwqQady77
vS9mhXmr0OWywHUXVwj9Inlq17JHR/fAxwV0pXKoSY42AEeix0hjLBjbXuheNjpk
iT0mWTkOKPxGQQp2LS6uyjYx0EO7YPRjEZZV8w1Up1WGSFySDvDGogu81GUAuHyQ
F2a0IPortVIzyHCR7QthxfVYhaVwtvyiv641i28CbRvgYDMiLsxrxKuTq+Pd/OKq
9BNaQq0AADR2v7Hfsf8g4pt+1DIGxkKQOIbQGzAyu1m7oJS+iknKLSzYc2lntgaQ
VLc4dTEtIdIHV2dBob8HYaBk8NJeW3hmtsXnYd4e5kluo+2pLrTq9WEjUUnhSDoC
+NA1YhNqQiZNmBSQwh6biYizAzNSjvBeguktpx1Bd2jAzFl/dYA9YVgyTVrcgdv/
ZT/lprYWfs0846CL0K4sUyU217sCHDh9Wy9akFEcbTCdQvgyU7cQkzpfgfIbGvuK
AS1eqRLU/wM81QUZX2V4R7/OAtHrMHV2qNbo7sOD+UUCLM8DDVtH4BrgFk0CqTl2
5RXUGnoBn2oFfmKzRPG9Nl4bL5WoYeFZ60pWOQTg7KIJUGA5hRSXPuoOLpiPkGTJ
4VDliyahAMo7RL4gvWwnyyRkKZW0K8xrZeyuGWKVLoJY2kV/wDo7Qg6tkIZ9m/V8
cF/spreGYA1r+9C/GCe8aR2kdlTYVmWMu3Y8tywwyWGpjpV3l+cluR0eRMYCW26k
4ivb3yUZVSC7ly6GsQHdFOfhdQS1ajV4nmufSrpGcq/48euHFk4BT7bl5kHxtN3U
LI4lD/1t9jK/82QXB+rvOZvutEyKb5DgSMmvXm/9DPIw/+1aZtgdxdPVxczInp8m
SWgGQqUNtsRqY7Q7gWu9//FFGFaRp5FYyJHjVlsJ+HjnpkPl/cVoDxvqQnYvtyKp
K4+c7K8RzOlw0mSFIv0RSN6J8GfamU0Jvm1kzKCdPdPGdztN6cr4jZwDnzEg6Aqe
AgaDRWAyxxWskzMkLOmk7lqE64pjfVxacQU+LYWTG0KFBTSrDTHTypJDHMa48szb
rI8HBt45lKEYHwwb7Z0XHFWsvku68ykL+eAC+jNGn8R5+ms6YE+qAf/UOVxjEI4a
r3sMvEyUos8Oxe0BieJ3b4oON4N7th9YUEe1wcHRNHgmTy/JYvgtJf2g2bSQ5seY
wzcgdFu75EmBkjLWV/t7j9y/nU9S5MNUQsHs9yx2GfyeIlwi9dIS/lUfy1aPJCac
cuY+z4/ogZDZHhwgpwOp+FS+ouRjYCeIfbqp2Ami1WyvytrpgJT38CMpG8pCleUw
GakhYGdm+O/R3TwrQ34CiHue8cYIX5VxdbziZm5SIK5cZjSZZwk7KD0EK9M2Ns8C
qKNUbYj1A65veTX977mpY5WpWIgFMA3DY++vYxIlWWQS2+4peXaQcAoCo1v0VP57
8lbf1/A1zRRibnNKKZvXi5X7F/D0gyLIqPBmd0GER/84lv78Td8/F/XjVqEfaiTx
gbbeRCPNf16GFKs10ro9leoThDCmNgQ1+FkoJchEOeuaNNqPN1bgL8MWXYA9EKsZ
hKljQHx2iVRz6r16wBLcgD8/Jz2lOusTWJAfoPepvPGCA//Jdi6pqBdVGKaW7wD+
LtBA1xPXNUjF+uf27ZBLEL76j6WLHC6D8U4tYAWUBW211a2XNLdizrZxyEQf0ZdP
YrHORtwNEYIE3w3/CDIgYdOWcuZOjMTMTh6+vxsQEj0Tkh9rFVNN+EJ0m2S6ENPr
+JypfMWHihR2C9dKhTcUtD2nOJpuxvjWISKT6NigJNZecjRuZGcScmRWqHw66v9T
6OhxC+vbWPPk8AMdbcPo03wcjxreUCSTbl/HvDZu9x4KkRp6G92JfDVcDWEiUP2I
Y984ghR6Kpa6Tc6B7vExXmxCTMigYRw2ko89Ejx1n72XkIirq/UDnGLsxAmEJliH
OxVJ4w+70WJKIbW90DX9DEWNW5jrnyc2yqauL/tNdqeqDZSJ3KAttuP8LhZWxnOD
mpXeq/LBfGSEz8eR/pdSF7byYKtGLqmxz4jK7bOUJgwB0NMue19pJJBBHiJ72Jvx
VsTbCTIWtuNgdRq8cPiSzKkxxkKwPqMfr2/m3KZQSnoQJ9ykd3weiGgNk8HFfOAz
iwlAIxCwWpCEKX0mFkNrvgffWIuNIprj6M+eZA4ReOYYvKUhCxRGf00l5nskFKvy
xs74hMZVjZc8qgupl8hQs+AnQ4gJobte7EnGqglBEfuVwDskzJnPCM55VGTHhkYs
9IZmIMyhzZcP1Euoh7pz2jx5Hfd3pmQ2zZ4fbLzyikygkYXrjLZxuyO5OWNH49rR
QDlRycE29CEN3zcq4zgYBfzoedMdd0C/z2yOsGVTq5htjBxcpwsO+GDe7D73tbrK
3rtj5/aq3VUglv/iUSclAxH/fFWYvCRXguthQNI+IuFOQDIGP28zHG0+ZS+bL2ch
hzDUFBOjVDj/UThc6p/d1vNrfMvh+jVaZT0LV4S5IT9zC3zeLftt85gu46Qp/cix
vccs8m2d2MQ5Bq3TpuCit8VT7DPcksfkRWlS5ysBnIpmqLP1HYFVnXx0rexwvmjo
abuK/NaC8D/eccl+MplUjUhqKKNdzTBTWOIiCfuBsLEIXzFKJZHia27rnehCfPo8
K8s/1A92pXblKGO7Pg1VvXElDbwdiqZHXADbzE5hoHdbBDQGZd7m+Z3bTh7Fa1J4
o3a725gmP+jOKzZsmhDc+Fbi9npTF7ccLlA+Y5ITV0zTdhjbo6QvPOscsUZqxpTG
6qU8REdtb6/lslusmm9447iw+FZpVRXUZv6pRcYWKaoi/mKukPKlo77fusTDf6Xn
nlXJZuC8pkgjBUMopQnWYvU/LxD0rjIhnP8Le3Zeh/Pc3HUvT2apW0Lysa6YfhMG
lAF3stzLcmhJFEbzmZ+HTu5Pf+W6+BGRpBZm9jhE36eDDeq0llN9XJvdYydX8BQu
zBY54F/BfwD9sBh9FSro8DNjPd1hpu6467hJC9wNITgL4wRN+R8xkE6PDoudZmDN
xn+KUOaQrUVGjqIz46SOkShFHm+lWN0+uCLaFPaDR66j26BxAV8OrhjPi7Jci5Bv
gw8dGzmS+BpST1Y+AxrIzI3QBCzV+X7hSEVuYXSTi/dIOTZZHcc/hQ8A9NuVembp
ZYFymcn1Op0GmuxgwvnzVcbzvJ7ejCFwrRnLN2T01w/yWrAKJScU64qmdXokQBlY
MoJJ7gZX54dJEDXfvEQLv3olhbG83XM8hB3EM9O3XR5gSOHwKW2viFvmD/Xn4cZS
zP12u1vPejn3CiB9RzBLeQoSFxapjc5cp2tpJtLCpFWMu8ACMp9Lud1JYNWIP+qj
Hk0TJqS1eYLQY8Xt0khYjH/4dcFlPaW+Z2dF5DkGNHbsaon2mqU/rVJ8lIMOcKj1
G/BJLezphQ072ffAkGT5omKrUABbuURQcZMyX0QCIbACvGd6f3M0/q2kOxeG8taX
0dBSYFeBNWNqnstdY5zxNYTlS4buVuJdOgQp0oggaAYLXcsok4CUA5YulKDeTCI6
Vn6YhsW8CISjMU8iyeGQVDPtPm4+BH67MROn4h7SndWvG/icmboRhbC76TgNMu2y
nyU7kpTMmGE75FxrTEES7qbP35gI2+vxSYZHnKq3G14DavJeE4MjLCWZQJDzv1tx
/IUVVq8z5tDXGaXMspWZCChyp8YU/o9foPstaDYrerCbZIkXey9vPaO90XaZkeg0
MKjajd1B1ekGJgra6THhJlACQSKbverl6xxgdURotAEBP0NbBlUPEdwgghSc9jMP
mm3dQ2RHmL5v91Vt/cvhuYSMf7dIPB5a4tNxpnlkBc+T4YQRZZhSzce1evZ8oPpg
ZUasfH6QR3l+YqVqaGnsp4cYN/oqGUmtXjdiZYyO+8bJ61cfZrZa4oUx9fqKaa7c
az9TcBWVEonJqXy/g7aMRCAaXUjC8mjETulWV/jei+KbPOI+drLPikgk8gOGaEAl
QuQTF+5dhkhGZCVh6SSbSmFEMGcQt/eo/8NJHSbTHPyZmN3n6TGMh5oTNiU+96de
lA+wWa7wvTcNSUcJJw9NBHDdh8csnv+yLfz6yKExdlV64B9OyUy/1i7WpPtHNUkH
k1uLw5MdmpZjlrCsfKZ5HFwDyOp9UMf6vy52Lv1Q/CE7y7yNYTrouAIXj8xnsy19
boBn5WI+y+kHO8hohRs6KPFb9xjvT9wrJRGedKvAGyVLgIVUcnL8KLqUnRQ8aOQD
vdq5y5sRLNces9mfrzeSxRaLSjNm2aZ3szlb6gpe7HXHRXt1mnPxuTnL0JtlA1ZW
MUrS0P40DKmxeXDAOTqRIumlB/B2pNtLBueg5Xa0c7h8TVGplBj4knGdfquJ74zK
oLT6SGy/ePowGossHzkwEYN33m26RoJu0g0Tg9BH372EI1dPgNjAszCKpuYH0RM/
zdmQWAgrPmtsRo9XXCQ+YDC4X9LZ6gIVqQh0MZp5LEsdWs8S2W0qAXuS6JYSGRS2
NCxHjAje5Ynr+DR0YtDR51GrgCVmpF96QV11yJQWkMnTHdVIE3SkQO5EX9afHiia
56P/FRV4jErdnGJJcnl8euwMSBEyoVmlbPMMf0b49oE1kkyHitI3cp/OLnt3fMgx
rP/mNhRZVFEIwKR4Z4+YiubRtTvlmbJs4jVDZyBsjIHfXmFHYVSI8DoOsmw2HPbf
n+wy0aI+5mP+L6HkNZ/kwrZ5NFTVVpG/r2JEB0YxwkXJzWsNVRAS2egQEdgWFEbJ
9djV5Uqs6D0ZPCs3HgsnKmvQs0LPUElplzK1xovoHhdWWaOxdRYb/nxUs6CfCMz3
3wxrfSObqzPGFabZYkaL83FtIW8h130ixI/lBEFt2OUY3MRj99vgQS61kWN04Dlw
AgA1YrcTYi9hH4yUkWHbMlCqAKgwiVGhJQ2Dx+ggdgwUnG4VQIu/5+svUGG0Yvbk
2DxHAXDkVeCTh8zC5nHSpXJqf+QmxtF3nAArkup0gmDdlw+kiUej8Y653kYjubZj
ag/byELpQOAomkI+o0qLwiXI1oDDUYpLGNyRRSf+I/mtjlmcnzN8Kjh4h3KmksIp
FeHUCCse6DmSpQRQfJepyJb8SuElaLduEARHo6R27njvjHcK00qteYw/6zqPw7xX
KT96JNttr2ljQQcPLfAmPMg0tWWlU++n09UBmjLwXYn8t8Hazr1JV5CN1KImxhqA
2WbEy3zdglbQSzVpOAgxaW94lA2iUHV8+H+eL39hpxzKl+5y/jqsCgvpLLit24AE
OkWZ1m74PYsfq98v6wDnPfdfj5y1ke7m5hh5TiPFE7B1lI8lao+6VdvV5ZLTk9iA
o3cOsxJo35zpvXZNRKrEFm0+TIIZ1uYMaeWpQXiy6jpYmCzjKmXUa+FCFPDeRkFa
f4bNIsYKwyqbjZCv5hNbx1CsHgkDTWPpD4JyZjlcpU7DO0chvd0uFEGaBcZynVPS
ijov/upCd9j4LbRZAjYohvj00ExqdGJTcvyb9z5dbXJ9a5KJQhoI3y/G0bskFdPP
vOo+qsIDKHsd9lkU6nsTcGPWRWwhT86u4dA9vTsVC9pRCMZTL/7Aa5paAgccJ/9v
biIoDjxpeSU6yVDyjwRS7rSjd0trylV1BXGNiIqKTFOgTfCmMlLh4IXSQk6ILpP6
lpBoNaE6vKej93hieO0jFlbzHTL7chc3qvI22GSf3rxFB4VYRHAYPPd0lewy2t8j
VyDGNmbqsCVng+yKlMYn16QY+pf5alvzj4itsoJ4sppy4HTcfmj/k1clkVEjYX3c
Bmqj7WHx6WW3b2edZwPvltEvYnSP5085UX84o9LV2foLTkma1B0GRuSR69oOB/qo
fMDjo//4xiQ8gbT00dhVnv9Ve5ao6gXmn2ipINjCa8GzyHLeedccgf7bgYfUUSJY
/byYHi+TjkZo8cb//15TYjHlckLK3yV8R+/dxGzcyqePUKy+FHcnJ4DfOpqyJ4WX
/oBPmhIhm1GwDbjD87c0G4uq5BxPc1dczpl3+F8zfL2g02oLYn/iSY2/5GloxWy9
HOQyyFiWlq22C3rrj3fh/MP4UszT03pNFZZEx63aOD+PfhvSbDKOz00lSWRfJYyh
0tlCFlGxjwV8SBrI20g3vN2uHItFkbTOqTELRGtrSVSPpF8nmpXBIQDLf9wnFrLl
qvVLR08Xl/oqHQKJJi+Fna1KCzHp2pFU5keVE/xoWe0FXHL7XusRjr6CoSLuCvvE
U5IglDVxIktiKQ+vJ4pxLH7tXVRUjqddKik0RO1ClsN0/M9DU5O7ZHjK29UGf8fL
JcjLqBymdZWdx/YiTMtHmMIxmBzh7/tZ0EWR5Lo9ZKRv51u7fYKA54XZ64nitKBa
SjEoMwjMMMW5sA7Ujui8xMYkp4Uw6cMxRDbRIyGXtyhf7JyOgxJSN42P4N30QHc1
Y1Y5UqwVTwH8SiRBF1XfzEJhXMDr+Zn1vW952FbJ+m0foKDuyHjnQ7TX/Kj3fANp
lamx3fybMJZCmfcvIhrGMQUykSaWs+KJtm2EyIjqK5bgoZU2ic4n60ovVxlb9MQu
3M21v0xgMFoqovacBWCJkGiJLpEa33s4YUDBXSocpYat0QnlZn387HdWOryBRVwI
sDtU6V/3j/fGFfslbEz39a4T0Yc9CE1OKcPpFUItlJhThYhV8DQ0Huho8Cwsdy3P
v+cPKl0cdwMX6PalgziF9NnflJnaJX6PSVtLPY1xXunTPl3Lu7b07rY2GWgeMgEG
jUWyqQPB40sXsr5GRgzNSW8w9LYlgbGIEDBR0fdDE8H4WrVsmUZnj/lqDu71xRIT
CSpXAGQd3arLXxArGTwWfNsKEPp6odReL1rC4anA1tmZJW53yfTCMF0YIQgiZCYI
JnSQsidH8W17UHTa0k65sOiXVt4HsZn50BkGEIAZ3mvPJUNVhoJBKv/K8enfxWTZ
QqDtYAIIDZeFat6HyyD32vfpv4fa9p4B3dMUycS2VQwun9wY4jRpCeHVrS9b7KSm
JtItKB3SCsoJQnwuyIrwFsAMvY+Yi+p8bl58eW5RFZSRbP/QXek9aFCdAonTZwc1
zJlnBDriLV9VfGDeJyRQA11SvCSLT8bbs49JdjZhnlgJDxJy2a8cKP8rLLbpUqcz
PGgYXtTM0tA7CDzSRbtXpbu2FT7JaeY2/C/4MGmmPbufW1Dyri276cpYa2mLrKrk
MYWmVam9ejcvwDBcFQxMhm0lti/Tj4vkBXn+7pQULVtFB15mGvcpy/oSskFHr0d5
ZYH/G6AY2yY+UxF+WYkBj6Tf4vHKAe5ix4TKZPzTvqdXsH+gQLmcZ5KENNG2CfZY
YEnzY6S88R1pa10n+1QXa6ZQKX5clDlZZ2vDQlQc++uEJdotbOJwwTYmtlDdf6SD
PwBRg7wN7Y4FeNp6P20w7DB5zNZ4i6Y9UROVHN+zynakUPXQpHXw9OCoCOXFYNLb
XAGlWXicbHLqqFLxOHG8Arnf0yeB90kMS74xU1w+r+G2odN5cY2b19BAF1AP+VGb
JDMhmH6eTH94eWAWDkoV1iCj3iKGx5bpWDQyioJVId+TKZTM29vxTNRl7oYjtWIc
GiN+XNNGsafS88FwuFQLFB9ls54BacKeIn12N15NI+m7Jeo5oWbupWXLjnlW5CPI
CS84HaBQOmk8qJ6bytCdr08zmiipfAK/SOqAmJSvjRKH3f9eIlYg608fK1KZ1CSx
GnQSfkIGDoLxeBfrPdF+xSyU7l5NQivVp8fSipvaPbn+2WnLzaDg7CbsIUoCLWKb
ZedkK1/4HUt/C+LUuAHVXP1+uCEYVDMB/MsR7/d7LH21Nn9yhSQSlb+JmDH/AAtX
gBy8jgqsJX53GGHsCRNLm3NCZ5AkmOVszY4xc/s5MaF8lTIfOFYfVU4hgIyYiZjl
NrdrsYadOiGrwoOvFnfrDSkPD6H+yH+rnGzD1hJMkLv+nNyzjCTqIkYDFvdbz8Fl
GlzddLXfYTT/CnynpMbxOaY4Ut65y7oZd5HRITJtX5KuCrNv61cYRViIoWl68I99
ydyVhXoWSh9qA/k6MGUbS6l+N4jyLwbPfqKJIDr5ppE6vHBDkkOISG/w1GcKj/uL
ECZ67c8NESUKTfoxz9T93VCAQ9c/DU+3HfvLrMPh0XFOgXoz1QkHmv8I0YPvo9RW
Rq+QdU6M9reZfxoQaiyF9Rny1kNSs9uRObGHsEKkGZYCAmhnJ1kZOG+43+DcQWaP
g86mHzos89OKwxh837XT+/3fOHKqkfwV8ZdHf0LdG+ESPIMUWq3Q0qdOzRmdjmDh
lUPTYlyxlKr2RzMIKGPMfin4TPxQKF9E1JG89MjAyBhp6nSpiGMLi2gIy7g46FdH
t/VqhsfBK3TaotCSFHD039mHOkF3XdA3srzniP9XADwpRR4cTVa9MwGh5AXpRjgp
ySs9SUPu44o7eMg9cf+T8D3h0qu9CxRnPFBk8ZvXZJahAwiz+CPYzAozMjmNkxx4
+uX+aerquUcaxeWkMu8kwmXe85qV2NgNopPJZ+vnwnUjzwAI6MzYuuB8m2C5z8TU
mxZhc3muSFWIDj0fIOXCRZbaL8nMEmnUGz270Tzpn2YlcrYv1v1j28ZTuOZ4FcQi
5FBFeo8+pNt0OsXTLq9h65BD8ZL7tZ2VU0M3Lq0/SBe/hiU+QeAcX+1ylMq1YOmD
P/kXwWPzWdtEsnBdbeje82TZHX2DVCbfEsBtlCm1kfRqkziqL1bIKwrdZfKIvzUZ
AngA/35Kio5aDV27B4vrLf6m7Etr97rvHRrcZmVGMc3YxBPQOexs+OjBUsXRC9Kc
jZ5wHis3x1oTSOxFLOOmvnUcJl/AqPf3Q8UCc2u9Tee/4zqRRxS31JNvCEMI3hkP
+tlwvhuOH0rTFL1icJTGKCFIbu4DKkfVXUwbwqJpDAypFU+wq4d3dL1a5FfPxZ2/
FNwu8DEfMJqyWToqBKZ4QoLBMjekooQ+iRJELTp35NR6cFbVr9pMq48NSLRCG4Z3
Mxh+M6lQj8EmWC/hacYFOKyoJUTek/NIB83/6xH2W7EkMUBPn9Au29k0SSULfv7U
uGNhXaxY1/RpA5bnouNJy/cUN6w42nKqiJQqUrKNtGWA+ZnA1NljX/b8O3Mt0ukR
YCmCwQLw4udiBwcpJbxHRxL5WPvlPhyyxs6WW8BQU2nyv4CX/wnVMkDkctZLJqtI
mWduYMIZiM19x98SjFFn8W3o6R5Ze+fwbLoATWPKrOqvJZAjdtKppY5jImI6kqul
ulQKT7UnpaCLcEyvtMennNoKnV0wFmOPevEpr9b7cMPvHwcF84R8deVTME9QCzHH
BqNAyTFOWVliyc6hvW2NRVkdVKqKBPgWOfDziAesuhV4NLGRnFTT3nWuy4omXEmi
nV+LwUSLt9SM+3HeoQz9O0qyNjERSWnidwAYEBSRCwa6PhhqP7JKE0d/wtOLSA8L
VCJ/ojhpzggx0IAjcSo/nzWmea5wZ1vRcWao5AALGUDrU6TedSuDCiCaToU0H4FO
btW1KVvX5SdrLh6ajMKqwiNiYw3JKyY07DHdHz/4QkCw5Cns1xFxOV2/Vh0mgoQ7
whHd46RYeHT/wdCpa+3564WeQkf/rYU4qyeYrywyqnWJdio4/5CPP+edVKiIWutM
7JFuB76c8aBT6BQlr0JTcFMksFnTnNZjXY9cGlFXkBYTGI+2PbzLJYpzXV9WlzF4
yE3/chSs9BABDU2jsnULkvudYvNkj4D9nEP3H1YVBEnDPfSDbRuVqPDOK8OAbFbc
q8ARLbZNHpwsvnvOhcIfJ/Kke1u2LnacRIOFJMfj4ie2FoWHuwIjdfN7A6y97RLO
mp0yAeXZtQmaIpqpTBI0NdL2yN0QWhTAaFtcOQJvdtsKgrKF+Pgs+drzt7+a+aKU
VUp8J4va4/JoPvvf2ar74rRrJFdUsD9pqx9dS0aPcYwBAFkoNpaEgri97TH044uS
T5oEtW8DzmcpzLNIonQDiUeVI0vo5acNEZxSS3kiberjEhlGqP5PYo5yDQnbsaW+
t4dt7Z/IBTR7R/0HOGEM2XDiHbrCTX/CgRWaXinJ0Z5oMTDTxGJvCdsrpEj7VTj9
p6HQF249qDpSL5aWfgxUj/UF9kRdcEUYPlg8xKn7f7PbBsRTI6GQOQqlgzGXv5EK
+TQCe1p/PoOHXrSeqEQ2HjyljjHK4pEyvMu9NyAlTEbxZeSA0PcwFafp6ZbQq8Jo
1pYAuChG9RgjrBoQsH3d8VJl7FZm5Ks3SbAVouGRdXrctMFoplhu/vQpCP0QZ0J4
ADFGUSyOsHCzLQWE6Q//GH/Lx1DhONXcxPaqSOZnHDFDdaGr2S4JrdFFye0FKQhA
gJR1svWFUvdMP3FSsllwXEuWDoAk+TLYOOtOTwRRwUTeD73WAb1/znrOZsjZ2dx2
iNnRSV6cDdOLyw0FGhFwDv+oOV301mwLAfzuZMKfCANJcRfYRpw7E0tEGLWbRgQs
4qmEtT/bB0JnrKyqOnAp15n9nhJQtnesKrHukONuv2dF0YuW6nxCBcQKOC00sRaF
dArjkrUTlh2XjfeHLUxsrx/0OkLN1LKsd1ZTNYZjFJDGTLafUatXJQa3jPRTW7vc
XMhck2UnFlGQvPrM9vWokla2YtK/JTOuuXihTSGqUuvE4vmayHF9qfpxSK9RHd+B
gZDX6IdFd2vEzNpydFLL9RCSkOuAbUFd6vcxR2fcWE6GkYMAMmhac2tmiwe/gzCK
9DRA8I0ysBha0S6e7EotfKo3ycL3h+ybmVRtPbU+gOVUCSBv8C76JwSS5tj03Rbc
79GVJnvXNhrJZORQqLCq7W18G+68F3wVzbY4N4WhdgiKvK0dajVvdHZ1SHDBKOnQ
Bwg+8LFxp/I1C1IFgJwyWDI9oaYZo+eTUYyIKF+6RT/Ao6KPyfDtFuLMfgWa6Qjz
CNpaU8lZmtFDb3OrK8Xd+rAnQNdYBeoEGKhW0PRJXj01N6+aUnNaxwPVmNCVouCu
IR/JIqF1G8MGes7jn0+Tr2q7pbZFdlHZiLuXVkQ1Oif/7ma/YHvZXJiRmVi6n1+2
IvAScntuAldHCcJWGIFgHwjnjR5U/eXgmW55ngkXwHWKTLbWaZcQx4Cx9WAUKOYt
9uhFQsVVl8cdcmX3Lw1bs50Jzcu6fm5oV8EnUKgKbPTlsFDzFIaCR+MS15bAPiEs
CRpXQ7oSw3lgxdtdU30mLyvVUHARDp0/HKKA95mA4T66FNlZXnrtjUE7uDcmZ4yb
RfmVF3HxPvSwtO8LjF/zdHdnfXVUDPRdMccQZIt10sMoegGkYBf4hYXR/UX6p9qS
8Rx3WKt0VWA0gjQzexuIZeZWrtEUvkP9PhVs44qBLZnzOCoEfJlKOL/l1zJKfBao
LXofB8EiEEscpIVH3kozFJnxxn5uosSG+UfBwVP96/1pzvk91z6XC+W1238sXQ8G
m0U88qaMiQDMinpA6PcsjOOU4Vv5QXK6PxJGHUKNS8DHAu/7gPY+zS37XO8Z2CVw
nQI78Hkoq5x7DgNRTjBkEXsYlO3Ar8OGHvsvm5CIzNjR/TRbXppXho1ZRxjsM1W+
I90EEPRwA4V8JQ5hCF5KNaRBXQ2qDdIkIJELFzQGhDtHLlc8sgx1+QT/FiohCiqT
On2zSx35xBCOkQOkIZsa/nhKSodHvbiaRRo5Twbc/aw2cBtj4Pl/AOsrA6nEPG2N
unQYQ3CeqlomHXnuSbLCaVe6P/43T+MfLbizOH9usbPByxKLnsGoiFiq/osefM31
D38096ZNM2k+cLyPj4hofo81UZSWprY94AoxiT67sbeqSLyOnEubVS3zkqbdnzR5
7C1ZWR1JN33hoCvWiHhRb/BsyeQjRjgidW8Z9N7sUCChVSWIw9OsYekCb0wF4ziO
UsBjNezwvpZX2AIsMh3sBFELMly0EsjosbyiZx1rwWcOg6oYNLgUzDK59rHMwhGO
QYiZEPSqCvavNQf5AITO2HcvsY1XT8bw64caCeKmvsbtnPnfRA+mw0H1mbdPdCZi
I8blGq7O4z3z52dOy/BV8V6pXI88vKnTwtQSLiOZBHZffGvuYSvI1XsEXAQBY6Jj
j8uc+LxWA30B07V3dhUTlp4cnY7Eu3zJsxzMNd82L9Yi8yL0CHJTpObWdkK9UH7S
bmJwud6Y7GmV9hKTdE0My/YhpZ/7sJkhPUgZwHKDwxXIm5cAHEKGVUXEgtJwNTHC
RSe6v5Yd0laNagLOlzk6FBDuqEBW3ACb8IaYMYxb6BiVJdH709edujyiyUSY2pOx
hwpZrqT2hqRQBX2vGZFBM8sXEfgzJ1V1Y6XWpvIq+52+2EpRrqbLmz76W4MJ0PIT
NY653T4N/hCE7MXjSmB1+/8NIbLJUt5/yGBYNVWeP3UOcGdJa2hi9Rc94YyWK+XE
oslL6F+fKYE3mbXEcuyzcfjEGAsoddGafzSs8pZcC6VnQwP1fbK7YNmaoAxu5oL/
obv7mOTC6Kr+xSBEStOD/MH4pXUlFQIitbFTwPI+Vz/Domg9EeWEHPPokFIxq1tn
aB11aG2+FUerQr+ZFEKs6E5oKbD/kvopgeviAko8p/e36G4liy15wY2yfvbj2efD
DxRJm99dKv0kf4iBeEOv1XTq6qzNmiOAkULhKxUpuRrNUQG2toeCp6GQi2AOHYTS
j0ip+c6v+nzmAJzM20y6PGLuecZmccGna0tPPKkUkPX9AOEBc8KTgSJkZLBXKAM6
+yn5RPS1EpcUyVhoVGN93DisfMWo7oWJW0b28tv/yggQnHblxgboIuLWU4iaVc1Y
03RvvfVbW4TFPapxUDrNIfViT/ilMqT8d95TrxDsOqAEq0C95opfo1ZuXfM6c3EH
oKp5TVsOuWjaIVgaGdx1+UpQrpoIELwi+pvkiKHDK8+MTXbupWhimMZF/SoTWK1i
T043NqFkcJagRZV60fB+FWx8pEqAc8PuW6VKa3oeo/qFF/jXc3csP9jAgsAoPCfC
H/t1x18XqOPi7RQsUdve+IVyKuM89eJrVyoJcBH93B1paNwDkiB0qo4J6T2uIvYw
42gvlIlu3O4o3bc4X8+KtT3Xv57YG7t10YlLox6FTFIjT1dtSat2Nv4fFV5sk+SH
IGHyJ+BKHFp9H9W4RDj/kNOB1SY7Rwx0pauEtPRNbTYTlX931zgTLqVyixILPBfD
a1Yp96txzdPdz8B/cHr4H7QJ735mGQns+q6Jq6R2e4zdRh/v1m1QIMltJ9uo6Nj1
Em4zEuBY7mb5j7xCUijK7bj3Xzt6NNi8zOmH0yvK4IW41T2SyQ7+/i+klWzwNMq0
+ju7Kyz0Lw4pXP1aolqKGJsCNInuOblXZFkJ2EWC4zrmCpFRSwloL9ynExK6NTBP
qG02ADl6i11FS4ua6+VqVWmp+f7TtiAECL2aPARaS9KA/DIw22B+qYxF0YchyXlu
B+pLmpZbn3udZmn7Ywcc3fDxtS5LXM/GDFnO3Z8AOZe0uGB9+iSWfdcyULBRZ5rL
FYkS2nXTYliCA/uM4AsTCjh3+zF8TI71eZGCwFBwQ6bBBwAZmV9ZDTmL2+lD6pwH
tTvE7drZv9U2gkdKzq2/2jYYW8vE8Gn7PuvCWNkmvmAuasg2azBTXgCBU128wu+j
i1VkiYClViuxjm5sTdLQLkh2Zv0lAJEVnC8h09nF2NyjxPB4LDEf/c3CidVGQ57a
MsEvMnYEdRvoD1kJbX1QhRSVIOq7MRKoxV1lwonlwAb0vmrBTvBJcjZd4c+bGURH
7esoIBNkAdEoBwlKNq6Q1mWjNuSpTI3vzpxT5B5zLvp1Op+EQdSfAxmhAKxXS0S3
OVbrINgCkeY2q/FvB/VAg/lXoFgE5uFwhumCNx2KgkwconIwxO3YKpkN9HAXnzvM
BuxHhEuT6IvK9VwOMC9Uz3B182Of1xJltpP/OkmYX9QlzeR05EF1eF7u3khCrXmB
jYShFiWKif96JPesCHiragilYDyBSN9f08hI/WOxTWe5T4fSBMumrJFaGGNYaEQU
fJ/f/8UqwTIdXkIJlqD05gwQReTkLaJ1VwuppTTcy7RZ00itEKhhOHY4yCqqH7QH
pzeRXRAfF11WDj6Jvv8EYyXTru9dC2vVKoBvr2GaxzUCf4CCdQ/sYRJjaYltQQdl
0ueF4+v5zGwV8DTcd94FSPuKKHnAfgnYOG2Q8v7yWa53oVKasvyAM9yUTjH+OdVt
scZ5RjO1nWNr/SWd9Okgx/rvPnxSAWQuzQW2m0hXUkvcIXB5D09Jk0KOT8KfASL/
vHyQdhN/+vZ9oHMbskv1ccrVGoaRKajYRI7q6n9AnazkABWSK5+yvHJt3keuv0mL
1lzXj6vv79DrwWX2k7TpsPcE9hwnWvObxW32h/0PxbKeZTgzBM8ZLo1HfiuhBnqH
zmhp+VTn34LUvILGTkAvJARUMGcisgB2NiJSwPNzTrlCqU9wnmmiZqeFv/UzJx0z
lpGh0oZ+SVrfd/ketRDLV97lohPOcNEEptUFOK6oodF1RWnIdXDiyPCsFHAWzKp/
DVaV8XhnhSZm4NZMMX+FDCpW4UuSGhXKXEB9JnPRLH63Zo4xZfce/yxid8uM+Nxg
gmR2I+scfJL1I2XcSxECVQUuHQ2jEJa21vwHXsOELxAJPKo0YOKZ1Vxp++ejQLSf
1DTml/cyUcMXpwFom4aUv42GDa8xZ2v9vW+xGBsr+qp6/0xXOaN/7+7veFGavNnY
bDU0tvdqukp2z6zsdcSZrg9TjejjlTRTb038U9oWmPWFPgv/6FRC0Unky8X7Ph8Y
0Int9oCmup7AUZc9jJhNa1Ecald69Aj1JUJUVXta9X8FXPStSG4YoUS2O7jHMOUW
9lbFxz6yZHWYpaNeofgdkuwKt4QkCaUR1ySsFpYYL/L6W0QTYMDFUcqb2L6uQ5ER
5bHcy0aCWtDln1crtk5Z8tl2FuzNa1zTtzQJmVgYAN6YkCbMHXpvgS3sHhGiLmfJ
xkBafgo5bZBNQPHlmlbFWpcHQnD/Xvq3CdOQGR6FAT6Dp6WSCqbvOrVtrcGqhbu/
y8yg2WxeY/fR6VYhZuAi9guT+g6nZqBD/ODObfPW2hhwYTCif2MH3I+AI8ISXOrN
r9NxAzvpFxjEOtwAbAmvknuDmn1T6/G9q2HTnVYoeRcKbEPpuYZO7byz7pDl8Z+G
egveMqOXZ7gF1wOfjzA3XhXDuFMX5SoDCME3lPbBB6+E5R08nwK0cHueKoaA16GM
xzjrB9GBPWOr6HOMa+tdyd6ioeGJddAVdZJM4oJzW8qzMybz3PcCiSg8X0xF1wEk
LfAsLN1Mu7RSyaCCe4CCGLkpBxu5xgRtXY08uVKTG790D4X74vDlonEk40dFB6ZP
uQlT5XRy2bCG81+r7tMYi4h/BJe9HM6d53c8q02HHzU8ywQHemv2ezzyMgskuKxH
vr1ayL3ZROOB7YHYYg8uO/rtkHE1TAS8VmM/CjmS6BIkPhcu8DSNaiFNtOTxn7xU
vqQ6xglz6qCfI2KfhBO/H/42Mw0fHIVyYniMeS/M5nKfUYm371c62CMB0myWI5S9
4LXZOkc5lhR+E2bqwjRAeOjLEScHm9izzNmIR/IE4DLKL9M9mbzZjR+58vsSepXm
Y5LRQDBzswQ/99ZVLEwag0k4F4wkDalNl/LY5ul4RTLa536orUcWk0dsIuB/sit9
/rCGu9uks3uOWn3FRrSt/vk6NdIRpahMgKEcKsm3GKShwGK4uoXl7OsUMaPpzkul
Vils2mlvWGqL0dN6tdlOkQPQvfBX3s7u/IdB1ymmDTOkEzDpOgYKAo24gD0zlMkx
cA/1lg08wAhlQNlzh4Ggk5uaMADX1ua55gORnFBRkNrMkmeTqg11eQrxSJtniXlK
Y+VW7tGACoEMNbYffLks4p5JNcuOaH8nKHuAJKprl+d8Ki2kLVHYnfjzqK0T65F8
CQ/56CK0/XBdisEFM4JkNllEs0CdhtizOypuSBnL9dSxYEamE41cEojnfqk7f3v3
gHgO55bGZ1HT0S0n5yXMURGgIuCDds6j6sAcsa4AIISeVu/11/IdH6EAGnQXbMPN
6nDbTwTyJGBoYGSJAd2Fd5GQma0z9MuJCelMH+GwR1lHj9WwECnz/+xX04s0IwJI
l1byV4/q3k1LDlHuSVPBEd/+BVeymsIYKO8gyU67amh+QUsngF+gEbypKXHUNIt/
IxKa7eUV+l97TgwAbzl1NJOz+2ExAoSa5wD3dClWBqbdClpRjjNXXPhBRsmAaayc
fNice3jFTUPIfQFEF03PImJDfrmjfe0t59dGqxcFq3XftOBnpny5EdOCPIi3/anv
VCUELSyMm+hW5QXFc37GANLwotFOKFCn5BWD7VCiKM6SsiRnxoLDJGmy2IYC4nDP
mPEKvoSbOjE4FwmUSJYXYhaPFnzUXFGgXZO8OM8kpwr7ZdAxUSjEqt1bG6Inq4Ey
0RaWWu9gvVLQO4WE9YsmaUv8LG5SBE3AdPj8Vto667PkEtJHiOU4NkjiAjuOc93b
TwFKfYMEkiW3IeNUsMkpiM1FAgvRZSzO/weubgcxW44I6A9YcTIrWsmX8RwpX/I0
9bRgU7R8sWBgbog1R83+LaX1MMNhCN05jPiu0xD5Cnct4ZcAFwEY/N2kSe82PnVH
VC1PBLkGMaOtk4+GHadeE8NbyEfPQTMhcUlgvCWWlWWkc7OQmodXQ3sc/o8a5nia
oqFlkjH3U7gxnqQnJoq75IKXEFZhBnkIasyvhuNNv6yxoaSWBB9q5kcfuRlj5oma
fCer0dADSuIyhDMnIuEpyL5MIk9ao4U9aobpnOB1tDfWWNU3tOffgmvZOCNOFYHy
rYdBHK63qns6lWErcTWEzKWhW1SB/1iJBStw8sE+Nc9GC96jWS/8tE9VKog/nvza
FYSvty2mXVhsNqHc0PsOxDy27gvMFs1Mk07ho0PR3CRe5DjRwyhmmCLAhSq0J8QB
w4KtpV91QV/5fktPrvzEa238wZazKxTbM1D6+GQ/InC6ZIeggUJSuMz616x8f402
9pN4sechjqeHKMVK5d7ehi/D6OgzfMWiItydzi1SKjAssUB+uIhCb6BMFXfi+wqT
a0zIwAZzTYksZCMxbWciK8/cC2y/J2mVuVadk32tuuOQ2gZhYvCQ9gKoJQaM+lcP
HcZrJMdVjddso6BDxqgG8wZZoYwhzwj8aedgObVVuIa2k+kM6daF4P5YembDMYdx
CUdL6Xv4koLj4K5Eiv3n8hhp8uN8/eb69Toi8KncTZA33ln4G3TJfi3S+9Stw+4h
A0mVKGuKOBFsd+KfKBsYT6xrLi91t1zEZKmvHyElHMcixo/2m/1jbqtCwV2PQh3z
Q7O2tGk4OoLr9ab0RzwPagvvykGeyZ6mMbUQSLFAwcMHI6RiLQ7BLhyp1Qo0RGhN
dY6i4MdJJt0tmtqTHn5262oloBz5RQmuH2F3ddgKodtW3AXEivHhOrI1HVQAUX2x
th/+NG5vwiCpVXdKnM2Jyw1EKZ7sHwvlMeXw/O//aruu37RS9UY+4NBZW8xDB7ID
Hl7s5kh/b04DxmUU6+DOvDz1zAf6ChgI8awMHG0LujIyVbPV/PhFssuN9cXbQ97o
CaG5mrwxnMPUwZqRUpzCjZeI5mDhzENBtyHruaxS+BeheLVNMfIg2NZLs372h3RQ
fTCtaIiW3gLVu9r0IHmP3NWem866ZW91a4yQ+Gt99cg0GF/pTXUBptGvX0IUT9AF
izCEaZiGcASTl4E2qve2Ygs7nXh3ee7KO+1AnMu0m4XOxq7CUTJaqbdZcR5rTNpK
qSFICtcomIEnqaHglzh/9jfq3XS/W/FvfNT/vWp0UPk857utr+uMRbYpUzAutKx8
lJ1pvTylCW2mdsHe9gZn9XRfMgyQufZd0qpjjsBK3DEUEo7+/Y4xQitVyL51hIY/
kHkRNEhV6VqHbXakMxfbvEZISA0X6A7FkfDsPhmrIfOIW/dc2AZSBS+MkO9mJfMK
OZwgacovyzYO9U7Fk/I7h038UuYY/P0HYzW170dDxJsgkmrj2w+gICwDhNShlYi/
vVzFMGFXlEw8Bq16qiEfAs+ZOAGmWSSASyqTnVp6Zb/9bjTb2J9tH1kDGEWZjYEW
C1az463FVnyzNrEY8icUspUvsA42LICgCe+i+xlUYvB5Ne9wT6Ro5A9o0vun1kdK
zWsIGH3kdkKbRld8iWhMOaz5pwqK1d6i1TpcgU2TtUaBYfwfnEy1CeJkLjyCDar6
HbqR6CuAFpnsilEs+SLCYbd/irInEkDLWNkC64VqbLU/bo+ZIMdjwNoP8TfW/yP9
RmOBZyUyH/AQNL9LQ1kDWSHjl35WQHbyrlTxC/I+9vblpKiwRKf72sRysmKe11Gp
PFqvD7X0ZcTDIpb3FtY4MfXnvNsAQ32fvSwyJDiYSB5kthh2CxdiFDLpKWyITIgB
wKyzl1wSyLlG1op0StLaFQbuum0p+FKZ1D4S0Bn/G5T0UPpWM1urDgVmPdaaO8uw
8AHZZSkXHLgS+RyYiL0NhTY63sFWPH9I+9uqDJWPkHqGka8WXe4F9Fb9skQeTKTu
RaESFJEschIQ6lYtJNPz/3LnKaaQUf6fK0B8M1EgThY7BEQVXx1SiDv6eK5Czldo
aYVZwC46r0gswmM6GeFE7TBNKj2fTCldEQAtifCAIGgPkD/L4VvOEXKWc75oy7Re
5TVLvQh8v3RB74EzTm1cDfwhOnqVzQvtGM58mL9UbLI4aesxdyhkdyXqWD1RJknm
TBBwOk2+r9v5sV+/RPlS/jmH38fcrqz21pEbHN8bD4GnWUthZid15gKWe7SFWYfF
ZcP1PhdyisBktTuKnKnoDwb4yA0UGTtnMHVqGcux376AODrjnv1ZVdY8Idkrn2e2
kD9zsyENeWRdGEBjcRNrB6LgXCi6x2A/qna0IHz8XxYld34/P9FWZxkKEqhlDvxA
cszDUNTwNvzW+0jnowwBlng7a+cCJ9zu75XRJBTUmKwQbDp+thMchAp6Ah+gJ6lx
ADrOKZvzAKxcPfUkmWuXoHP6DtcEuLMjX6klSzvQ8n0LWvsVNaAMi6xzXzKg24xE
RqxOuDYRU/tlTF/Uy5tIeyad6o8CPmXAMqPj9pHA2zG0FxTfR5FVF9JiYZ6cE9rt
d0fi4MTldqy6FVjb4aDZC/4eSwHPj7YmDXkfDe9SRw1Lukw06UVQAuui88u7tJ+5
KQbC/lx/5wvLO3yUkuQfFtqMgjfz0aO/PNPyCA+cZCy7m0hJbtV7bv4Rkfe5kp+x
fcZUdL7xtcO+OvepMdB19Z3VUG2d8U//OXNxrr94jYupVw4w7ddNJaoqWjU0RoCQ
X3Y8elZE+Jof7FclNpmU0wZp/RqE5WuAIEtJNmB1wiPCX/f9GDphn2I9HtUAAqx5
UqRAWG6aAbtLo0H2EM0PfUGG/JV/QSjSy331nAkRFlipZMVtimH2n0DmE709A5yo
mfDkWH3wFo+UIWCUHTHqEPtIVDERXvdg7mubnK+yCdK33hUMjYtK9363HskAzb1J
Zo76JrHL+PqFbkCfaVS17EqoZ1Wu1VX03eW0TZymZtOV0jkAPZT9t3ozZ1o7PXCc
Ei6fPkKYDvyG5bGHHZvCiIc/rXCO6kRwKE57Y7jP2i0YGth3yxkvt7gA0zhXfBp7
YISqNIw/YeOC89JwqNLvG2ITtlPgeBAz0myxta2sfQo85cUVMEYlOAGIsygFbUDm
TJSDpvdJzQmgZVlVLj2ertR9y8U5pSuiOZMyUQf7STZhC4XyAuSxAL4vidn4o75J
ih5gUNvPRu0Nb6sVVVdXBAiAmQBnzgwrXULvRDSl3XtKA/w1FLloLkUJRFlRYAJi
9Wms3p9DeAOsHsfEbsapaFeljTuEjW+f+o7BM1kNCsM7WdU7jgo951Wo/4/W0jg5
TIoziEmtXHK0MP3NBr12mC+JePHiFMg7KEG4Pv2m5a0njwYLBIuxQus3sfbf2sN/
trXw6/LnDGgpVhWRoUmNuWi9LZh4N/vD+DNcGw/L1qKyHN04Q8x1nah8iGu9hP1z
kAGowRQi6LC7VLFhY7qJE1/75Yn6zCe9srROBMMXu/XhEWfukz61RKZokuGH3zQ/
iBIVXl44Vab5Zh//62zHPogFm5Gr+lW9yLrrSBdBHBn2JaSfQHKy9WCJFcbnTwo8
OUjFJoYh/b0ZKmjA9E38Yd1PCZXu4qX5ZLB187HioAfPiM+42vPkFzecbfRYXp7A
oqKZNfWIjH9SHmdfLynKL2rMGd5HdRbfM4AFGvzZgAmbXPsCbjqH8q9KQrOvZvhk
Yw6bCKCR9oweHUYx37Bk5FpPqsprbIfhMgDLeV8PE6NywsT4pnNyG0V9fLLejQ/z
EMXPMvPVIzLnGcwLmzheXUqYOiSwbRFqDt90ioH9MeSDHxq2rdpgMokzEEEJLeMA
WQDlhAi1HJBgDCFlVn99KlPoFr0314jSXnDJNf+TrRQ1RvFxn0sIEB+NIxfno48k
Drnyv0lsOHkjh+9dL4iKwTWd94X0F/5fJ4bIgrItUKvf/Tk5eFvHCUgS5jFaicAc
UE3Zw8hOErKG/V8K67Gjmzl7c7RevIcugeLmIZ8kc+VZBjQLWH8hROPpVlSLQjkH
cpqeQ00vC8wla6pKhrXj677aBZZEdQLbwFSmcU90mf4FR4gP4UqvVk9ySmXMBAQR
dN6yrnw0poMPwueb3QX9aIL0fYKPLMAFt6jsXnvyXhzVe4TmcRsnr4fOA2mW29U2
CXMTG1g7Xi5CMJsaKtgpfgxIR42xgHOc4WBkM+GykDOC8Vdr3KuJkAHs+dq4Hd/W
wXIVME/SLZpclvTjhjJx5lsykatYqOIpvQvKCftENG7gWW8+TTrXfycpzvu6D3io
QTA9CYzPINdn/PuX46hrNKEmCrZwx4BpYiTwHq7L3frJP1mdGM02I9KqSXvEtEjp
j0+BpzYPTZQfNN4RxI9csbdKMmJjaJK8+JJH+2BZZFGgEidAuOPbaXTe3n8gJpLD
8sqwHmUiDQ6K3Bd3kbMHuDhGxdKx4f/WULdDA69EEEQDMBoIQzeyCxHZBZaHcZQS
aY8+3WuzIpoUy71xV+UOe0HEUdsZQjr4J6Rea1plLLf8rkDg9FDhtATs7r8ZKozZ
OyUxGgQobVnLuuLKM6nobhbEcS5B4NzJ2LYq8Oa4jmXUI0n8xFkPJ9ZYmrfdCdAc
TfS6p1zotLms20++XvYbgiKbAhKGt1hCTDI17flh5BrUZtCtD/VYIvCaW55rYVYg
33yRY3G5gXXmbvI/BEQv/yyIvnFTjNMlHKktzVWrMt0MY55ljvod3/sXzuoa04N7
ZdtyLX4TBz5LuYsBSEgzzy5E/I3wbkNEAaioju0biiE67B2sfOJkuwjTRCT5dl7A
iTZSzF9myRUNhkFIe+0uQwVrcZIr+EzIWL3KBpfXrAM7OhN422yhgBeZvsWmraO9
UreOAeQJflxeheijRCfskrviRUFiUWp6+2sRGaWOxfQZjuenAFfZIc0gnUQTUQRm
ABZXzqhK+zulBUnGtSrupQHsWyS4lPe2/QkJ8Wf5tKroJrj5wFL87ige5WN+GmxR
cBimE0vOS5QKgHavypJ8kahCE235QMJOifzeF8B0BO2i6ou2s0qwepbFb3+eeNln
Q3814JDCsbfbait0JxfgK4I0LwNxldplZv71G5hcREeOTN+hLoxYlxhHhPFMxxDt
sQXJxBUQLSd6qWTqAsSWHweroAJ+z0FZ/hT96mSSgfOJMXGWAn9JRYcDtSKC/zZj
ovE67GDLWYQ4Wwf926+M54ulZPyGDzT02o69s1dpi0IQucq97xSpvC7PFzF9vaJY
e/G9+EbKrWViOxSt0LYaNtF57LrESRmh5EXUymEWdCwkSRy9enbbk53JsH+wR5qW
rWIfkj2KFNwGtSNUmi6egVUGMQ8kHYZ2oMW1FM7iV6QyUwlt61QA5aTqiKxHPCtp
UDIVfmEGmJJDNI+4nOl49xfwq/pweP8qOPSNgzVjuXEyf7Svh6MEgotZlfjZjDMw
W5MVW7yk/wUnz9U4gcU3kBINWKwD3CJjdZXzCUe5HEWnktx9rDxXRDwCbdf6Jb4b
UIGQGsueRziImJuErSXYAa6YZQ42k88k856lYo8EbaJk8xGiL7fX9E7CFKCHpwTQ
KnSKCsht4qWrSeisLAPFdRiTJuH4pMrdxKtxTipOuENiT/I79s6Bpd9FHgJ0wFW9
eq1viFV8NlNjHbQ3zncILMo+M1RLLB25x4/Zrr4P3e2FgsSL8eCUAlYHvQ6i6kQx
22V6gzxU3Pk4WoZB8DlzUy3RAiYk3qEihy2lxm/Q7FpguAoEcf8LiLT3ZxfE/qHu
c9bMVjG+5vF1eUhwjFmBGcUADbnhmhbCLdBHSgGBOsJXGFEsa8da4M+FX/cNGSCQ
GPSroqWmNMJEFIHE377toM9E5yhkB37KVRy7WEkg7j+I8Wk6dDHJQ5GaYUxpBRj8
y/tbj1HFr6vJ1RNB8PN8HeJ+RBrUzfPYtyuVAPIcvHQMcIvrDSohgvDhvErMXu+Q
0M825iM/AImtIs0lStsaJsEbF0YrbkjRhrFQrR1c2BZoB0IR/e/qm3KK8xA9O5Ng
JKgZbv0NXsnV6+Y14ey5HTWMIw5497U+ftG2IYDXm3G3Q0QYnGS+/Pxn4qJRK+o0
dYjhBBBOurZvPyqAXDJ68jAHHE0gxtQuVKQLHycuDMnCA45Gk/USaAtXWTQSqpIb
CZbYEEnseY/pLqLHTygQr8PIZ6YGllDD6kfxiyRrUP7KdcyZJIrn8akJ/N2Bkd7+
FkfmVO7Qxa5TqcljWBtgfMZXQ0ZjT4pJz6sztW8PWsdMoF6RjDSQhGkU8Tjgqwix
5kf+Ede0MEfl3Xry/wOiQ03PdIadUSBqvBFa2VYoDwVeFLgGGVH6UqjRdGXW2BiZ
eB9pryTkjfek48hfM+YMSHb62Zjwy/Z8KG0u8zmWhVBL4r0ihZvH/J9SLJ4HhXY8
6YfH7xIxVoM0Lm/HcI9P/8MZ0Hd7OAnF/NwMiexZo4szqeMcE2f4gjJHozaA2/kc
56b29SoKpzLvxlQ45xec7B451BKegHoCWmYrP9zotPyCCay1xMiXMdnuT0NNh0p3
MBcv8yVLlU1PSpZerkjWLIHbfwfQIVEqtb6ZCKDdgT4ZGRcJSrOmx6mfixJ0vPAd
klHw4fJErP/om1E8x11agXmU0YBdvza+0tC7/m+xAv72DOwvEEaX78VrmwlVFPWB
o/uxxY8WuA+GEBleHzIz0ELSUO1jMecWXCQZGOie94QsiMWZ9CjzO6/U9NzMHvly
hpN+7C3zTd4hAvoMooGkwJAfcvAwrYK5O9zQmVPijAwe6dgv5BTV42JiWx1W6kLA
ESSOhGwBjDEv7jU+twBsjy+imlqEnOJ1tzBOvBZIzVzDbGu6L5Q/Zhs1AIWca97c
oquSzcDUQA2JCuVaOj06qkUmLA5WU/vsG1pZ7IBgAOIKSSNeDaiBrVR55LlaUbl6
cZehF3CXg3ANSYJcpo3wQPChwIx/VJWnyBA1e5f9wJIirbyvsWBGY7QIgZuHPV24
qKwv3hh2JgtKmXNbwhem9wcTHcirui+iPYw6hL1GDtW78AhpzczaBIRdRis44XjS
nY8yBBPz/REJzx6RUIbwq0koD1bHzZZtcm5umYZlK7uk6LpVZTB6++5rVEVaTOot
JrRs3m07gIjYR50R1tRKNWiSkEb2iK8WNjips4Gkn+GV/F811+svGYE+s3U/pfwO
LtUjvL0NMb87sZrEON+23dhIjX4KWb0vve9lSZ00GoFaymXLPbgcbw4b6X1U79JP
C5n5QOzBF5ww7pkVG3INiSW5KSvOPYHX+cUS7i7exupmW9F9dA4Ft7lwaBLkjHeY
kfaiN4/7cyNTQmny+lJJB7kAMWAe7rdHr2g2tpQd1td05jeDdkF8znEg0kmbXa3C
L6bvB4CfEpTzjaP7+wbngBJXNdk91co+3sX2h4coH4hSJTWNOF3luTah2ADqDdfO
Hd8DGHRkwd/9KrSo3ChliGuvDWRrgVhGy8U6DDO4IbaLPSPKQc/x6sFc7JwqJY74
+7zdyUFsAZFTGSErD6AyoFSEhNYZ2uZFqVgzozG2dDYkXZUz0+MCzJ1Rgp5uF3+N
8BhlgGpBwllIf3U1GWhDXz4Giogl/vb+oWEWVWODATbdf7eox+6xp3YbC+pEAwYv
oM69ngPzKXj7nbgrX1L/xhe+I3ZbAKLCEs+0HRv1k/rtSJ/TezjNo2O+jjTdX+Sy
VFE+UD2MX0DhDQLJ4AW/mPavTwzP4JP7g8COkfOkUjEb8jmZ5Tq7sFT7L7mBfxw3
zAjrBX4dve1k6l5Bfvs1/lf0/K723A66TrtuvB/a1tG7pTAwM4kBQI5nlzmX4JG1
HC30AfvmUjcSp7DA8yBR8ddYiOxG8MOb91a0sha3Qo/1/K20Sq3NAYd5w579+ONe
uxzApAx3tLjOQKA/5xS0XPE+HLfB6a64Wg0xtMO1wj6OQF4KU8M/g8kmEMx7BD3O
ya2cCr5DusnLexBORzUIvZ0Z2mr1MNfIIQcuOu/woSWJfPu2qsw3YaXfSAbtQ17d
rhkLI6m5tBdQQ+CCpnEcFxpue+XjaTdL4A4MwtuwnYcrkJhAVy3m3VfHOB2vkKRe
4C1JIazy5lmbqShh5cY2PdcWtlO76KoSBrtRilwRRREMITjcr5DC6eKZseijhjRn
m2gOkU6DlqWzrJh8Kn26rKJJrtsDhIUr4/lSMN67c8/bMzyTCcRO82JN7XYbvlyu
mS+nT6Ldrxz09NH1OnyGsYBD6GhPT194QIKnCCI3PA110Yrx8/HXTbFXL0Qa/zal
E8RQK5YuZvaYESxf+sTFaSZPlc7OagntfGYiacQzBKipVn0w+kNUjbcqxgGGSr21
NIP57JIO1jdkUwElL0lMCPSqTErXTv4igb/gcNe71ZUpGUzkvD9/tA1VtN6X9Vbe
5pct/lkmAJa+k52ie+HGeOfVBlUwv2g3OlB6FlrDggJ7YXGBh6VDa7yU5ZAbQpIo
qZFE+UNvryob1ymsVusHnNgjppZTTkh28n1ze1hJZLjJrhvAjgY6qMLfz6xQG/wa
7xvcBooL8X5jCCI0UFuTnxwTIu1mRXUpwT0XdFjCHZ7hos4ZVDJasU/8UXKJ+pLi
yoJxM1g0xWT873lFDmoutmYwqq1UIyRKBALqCgYIL1y0CyzZGj5iPIoxT9Fl0V8c
CZSiesQfP5bZip1K9/rBn9ZkEOwL8E2oioP2b/tmUPXfoIxK+mC6hXnQkJT+TnuZ
jUOGephoYlIZDlVI2u7ahklkh8B+S+rALa9rSVEP0KxUA/dI2gHIwL9V45zPI0Tt
zG1C3vhKeZp88q/F5kF6AHvLqgrwV1A8BUotyRWqdNYhqAO4294bj1Pjfe7e7QC0
svYhJBOHSSHGgj5Lv1p5CJ7V91svsl3NI2cvkIBTui/jQV77KmRf6riDP0tjg95J
M/NdPb/coapmIOMo8x+1SEltUH9ennsrUdwRj9mN8XGvRAQ1eGcFxaVPEyO8RBKb
+4vvzu2B+B4m/xdL96owHNrvUrUEZjdAodVsmty4izM4nQoClS8knii60A2H4bLy
lvVJsKYBh39orA2HKjZkX0njcPXG2xchFPhvVBM//iq526dFuGGcItmUBR9iyQg3
qecTQZbjKD0EpTikAtFqDtEZBeJfielpSo2AuhOVPL41mOVVPgWxpgGj8bnS974z
QjrjQhQvHLIL7PCQSr0DynojPnlDeKX2o3JkhAqCEasDooR8ypKuTRMlEYUTRC2X
HB6KuUL0AddBCBvbBTa/9397hce0pyD2CfYrubzOQX4tA6EisFaDIRpuZCpFEHzd
k7N4RphjnqJOafbkmw/7Q14c4tPYXOo95hYhwuZeK1JV6KCVdaxDeFcj8NuG+XnM
5vaUtRyqKNFn22SJ16OTg5iiFhTsG77v35lEHNANuo5XvG+LauRvF1ac0cMIJU1H
ZhLO/H8B8gjW1ISGlBVIBzUXVkuiwkakT3fqecRf2MJ2GTr9Z+qQxVe/BzATP5fk
aU+K7UVs0lqc6t4fwhEXtpxFslxJv++nRcSZZ0kSCMC6NROWor5fvzAzPIXDh4F3
VEaZfy++saH51Z9eCpChnNamTT9NgjBI8qb0yN8+w/NXWbmWPTjCgBPLqWbLS1jm
2sEhJIkplfpKklGSoGFBiij28vymw8j4J12Ubdysgjh+6+XMWa8iDNZ8076Mh2v8
KjrLW5Dq5Q3/GBCucyXWVCdCVNjuW1CuUnNYD6mdv+vHoY6qe6gtE2ctSgEEEYz3
lisowc/qkk+rr1ub43CqT+biBQOk02qx63nPpX/sDbC0vSgsfPTQzYsErcQe9snz
GhDzzm+CSh6lUiYvQ9n2pJHSvLVJmvGdBnGICfHyXwzw7xwBPUI4YQrZnS8HL84d
j9au7ymuvKvl+fAdpIEk/Kf3IHFAjx1aRoGOOs97LV0vyp9hovC4C1yVlh+MVZEq
ZHtBR+pLxBA5U1bPnBPUM20jdKJig9anm/Y5n2vCl/4IDK+ySTiiwZcuTXKtIAPx
ws7OfOSw2PKon0A8bgJgC4kSvvP/lCeFY7v9tgVK2nKFGqMEI7rI6D4fG5IHU5hl
B9bqhQ7N+cCJgWJFehQQt3Rj1+dIOKMdgLpG280gCcv7D29d3FQ0KFLb1gmk7lnE
SgyiBb5LqiW8n4974I3EYPYrZB2cQvNM+W3jYGpE3XI4jg1bpn0ytUVn0ka1y6L+
xQVYva3oqDYR4tIh2RRHoOwIwOqHVgu23YNcKlaPe2paKZP57vNg3kl60elktWuG
EGXbATk+OcUG97InGOnsAGe1g4wA5KANCBqxJQ2E0BCv9iI8FekIxYk8WqR20V40
Yx9C2OC/snnpZWeklaYSlQJVAeYEfDkAFRYyA5Dhi7Bd+EBv0bKgo4x5Ir4oQ0ro
GWrpwwk5OQooFiwtAOE+/3kFii7JbQaapGYumwDG6yrE0VDZhckzei7qLoYtDuWd
SRb7vUWn7g/VUg4yrj+PIojJRBLXw1Ma3RcrWDmSYZMLlzDUX5K+mljrqHyhIudO
9aBYbVR47625PRMQiuWTs2jMeKTORW+7ODmQIq9n2BlfagWjgE16/tyHqgvflpbo
DFLafJk6V2Se33+iLFM5SLcyaRuRnr9Ux5NOO8ZSVMvT3lmfNofNe4QjmlW3leci
0DElpM3MTYKyKY9Oxwz1p57PQfPhZWwzBC7DXBNII3qdKa1y4l1tPVV97WFhtxH3
W05cL1B7oo2Nc55yA6VeiUufoN82zCj/ozgPKSgG7yUzWnIKwNCv35/sQmjB9PeG
yMcQJ8BoqJAGRo9AgJE5OQ0ia+sDkzQDX9IIr4CMQ3fAhaFjtVhH1r//cIFeEAEr
EiBJMX/gWEbwW1G7zPXWr28jcmd1Mpn/8AvpqQub4lhvpTu/JEsCHcEI8AbkWwTp
4UUAZ329HxUAfTFKh+harnmndO65Jog/kb/vi+G9huXFPIScKxg1+BuWF9jfbWvi
VsHNTfdXa0zj8VGCZ22TBq5ifmamRFAbz4VIKtJtGw0wnIN4poCL9bfbm+ZM62y6
pZZOki4DtpY9O1Iz5VGO6VbWYK30JgByWENkT8eAHwnjT5iFPhsLX/O8s8OovsIO
YZBVxIP7KhWGqZK44m5J1TTh1D+napE1WBfb/6GxflLYO8h62eAsgMCrF/PztgFa
kUmR+mhWS7nzt8KHreg5K8zdT1Lv9k6DxqllbbBZIraWWDQRlNb7fK8w6CItzIn5
m8UA6G58aze9KE9gt3+W8s3LVI9wSA89UAHzRqBlne3KyuH1JISp97cju7+ZLb/z
13s6V8XbghVfBcQvejuczOhJpNdAA+LWa6JNSybTXKIWSBYDxAgN5BHxWX6YKTPk
TbRpcrEuU6ZzkI3Gr+zUIImdpsrfdn8tmBJ5AV056vf6op+S4hk6e+6CxIWBTGKs
8NPPMvyS7WVFva26/FN7Xe2G8E7W3pHlyFEFrJ7OOmsQGIZkETS19JvLqsbSpw3b
1UTefZ/j3ht8vO4JYmjr5ZswScMeYnzj0xWUXU5xZ7FIiUzPajjBDIBqi0r08xiL
vBCENmY3ZpRce8vwkJN0Sp7ltIMiw5EMsdPfoitHD3PSq60CVl1z5k6iiJZ4G9Q0
ZRb2oU66RxsszPhLtIADTBUCTtc3rClqIdL/i2StFTRGGzXg8O7ZoCJaDUchzSLt
yO2VyFcJO+LQQRTcNTsbS08MDo5JWRXRlcJg3znpo/7t0Tzd+2beKWMPz0wSvmlD
1CqsQGOOyGbQN9X+bGkFhyvzAKv8YT885XjYORQqGnZRakOsPtIoiataiJ/t+sX4
IjkF7hnNnRyPZzawfXkLFM9IboIhhN5PE6iGZmroSp8fRCSlM4wgzife/rYa8IiS
JIYbZFUuBAsQNdnpMaFyHCEIYO/5SEdqFqpSPcLyuxcuEu5ryZMY6FVj3AHyZdby
NzeLLdMedYlGCGMbJBRrIsQ3wfgQBMYm77EASLVwJ+UJL9UvSYqUTIFHWwtcAQ1d
H/CDQeA3SgMXzCTsOogBJN4aGtXE+ddtt+o8FPNbhvxe8t9tG3VhU7wq1Yw1fEud
+UfoCsXri5tYBahf07DM6XS6qjKROyJcRyG7nScMit5guPTvH7Lh9YKSI2QZg+IW
VMC29czIgvS/DI4p4wEH+cq7Y+p/atRpKfec2WVfjfwlVrHnFkg2JKloetcHjLoq
coMWCbc3mjCeRYBaaoHpWDqAQ2B4u9MVnpl7aQ2ZWDIWqzsb0DO71k/sznaqmKR0
8KEFF8VV87i/GMvfTv0RQQQ3uetrGN6kwctCPXpRuUn3P9w+mHzL01Lo/rLI59bB
EreiaCPn9c5CGC0jm2/aFAm7MMTMzE0zX8yIXvR22imKund2q/HAL93sJAbLWlWk
r7cE3RAd9oOPrlMDDR5lRtGXf6UPpf1AIaaeeWyXPRJv600Ydt+iio/v9a8pDyxk
0rmWCkPEDFmOOOl3Dm6DfG2uvFhnr2nBxlMVfhc8kzsByiyW3wb0vJaPv0sQb7l4
RkDGZEp8wzaGvG+uvIru3rcARe9Y6UUznMhzbx4EvvjH4QHEu/3UaIA89xsoRRX9
X4PF+XPkj194GCz5NNYZuq1QaMjZDRoElM8FzxLvIn+AQOxrAA1dF0Qo8MfZhX73
IJmv+1SqMC5f4XPTti8YlgYYh2AYHJiBMGuE6RVY02TMYaosxgKcsMz9Rlm5XZ63
S/0ut7KVdJF684WDHBqQtS5QhieTmCFTrkG4rwD+jtGC3rBQteDxeKMtsSX0iPqC
YzFI+ds4yHUjepXP+22Bz/UXNLmIS9ADfHZDfaGcgmUI6QhzY+dB+pkhzQUyPsUB
V3wUrka0k/qQLYPXczZRQi39CxN/0qjVW6bf1GInRtGgqGgUMg9HPvL4d6fpn7GD
UXnM/qaxPKkJaTyFtYDPuAHat5fIiQCys7mZN0yL9YO44vxKbsNth46cdA4fDGAl
L40ZQCUw9IrIp0/7hlXDIYz0Z8aJnLcEdIDUzLFpSkYxa626XvtRQGjvtiIt/U+X
qN5rWz8kfEvYDdA9k79U9eQLygbGKn9y/IIOmzCSbPJke+4VH91lgq9Wbh2zpyGb
vXVeeuU3w2dYvak7T3Ck7uoW8a9X/DMZIb07qsb2sj4fV1O1xMc4zSNxDhHck6qN
bggHGTE/eP9FeoBmvU9PkUMCPkNd9Uz3ZWefutAoAZqaO6Nba7CXzgcQbcQsnp8c
ix+h83DYCBCiJ/e8i+5OGw5eB2cNH5enbKd0t76mM8TkG0ZY+1IAC2lmiLmUd7H8
ZOVBMbFSMWdh5zKBL5TP3hWj1t/iSJCESXXAIXw8vsRoIcEu6l47mzZtnSB/Jq6C
qX4pHcIK7rqe2/8pBdLc6CkMiNbHUp8ApezQNrIbED+VWYZQc+uQQ84w+dhMEKsC
VYCJMY2la39o5IaLFq+eQNAWDOqpCiKS/c+lJsWVZM6/sb+VyAgqoUyhtfgmW6gr
dY4+gQoT+VGfL2WTHKNuY30xLrEl5mDJ406e/g6XXsOBpzTTiqRwdQifpfAxMxfu
DNYbutPp9YtXipMfOvTSr0jc8PuBcVuZnTykFQtgHHkuPp4auXEaKflVL+5/6sdg
9LUpRIRVjR3Tpkup5r5b7y+RrU6NvCZImnPgO16yxklk5Iv9hvjenwZQi7M2JPxc
C8x1KFK9p7ziYwircJotSIaIheaOQBrqqkcG05p4Fvo2dOPGZsLPuMTaI9Z/jpr+
1vxG+95zsQQjtcfYMMtw1giV3uJAi+XVwQJaYCW3G+lCMujHRUTJhLeXWUAVwSZO
qTR04Ca0IjuqOqs7hrW+StLDpemfp0/pjQRthr20hgsThhJQFz5HnfLGZb/MoxMA
x3BnO7zxHYyu4AvT0hZP9g3CU+LOv/lutpewQlHAbkz8VMK4ZubTLBLu4W2Y0yrF
cyantX/eh/uYfrFVsTF35aIhWlyRBdtH63Zi28w7GzFfzBFRu+Zka+vZuMY4Q/Kg
YnhW2FccS5XwqJNqICx01miNj9mHT2VWi3JvdYHGWEHwUriACWoeIk+hm1vEIiHY
zcgQMBhv7WUUzjUH/1mwKZlD/7Ay0oFM/FB5ZrowEVacNFsr4B23ZFK2cmPBjEPi
CgF3HQcTxwYuC+d4BT2ZKPaXaOGIS3jGwZH6GuJXpPf9iKwmbpvB0fC7U3u3mtCi
LTbc/WUHljyzJEBMK6QBewk/7+rzu/Sn31m4qxJtGEn3bDmd8tyU6lPnDKLPDFFP
suj53T2KLJfcc6YaNjq3Z50c7iNsze6WOCfrEIBlGV3e+G0NQhqjQ9RJGLii7hus
02ZSqkTkfglgFMTSi4iqEIikXeDAL6RaScyWpfOu88/sw0sv6wZZEdnvzVMrdGwN
Hn4rpmwBztYw1FrkRsDzG5ZfVMdafNoaeJvfrOyUNX2d3ZG9xEoNa51ASzOR9AOK
/jsGuDfEoxY+YaTUri/XVxeuag+Ea85ojLeZAOcyyVLIiUNFZDEDmF6sc8o/81L5
BsTToYkCQFwzjReS1SRVIwCxmzl9tkn9ElxNiTIYBC2hQEaZhp48tIbmEAe1oJCQ
9c+x70sGotx1lJlWum39TxO8F8j+UAhxJOsZbUhbmM0/cnMhM91Ga3mH+mhmjwLK
WysY/KKWvbz9KW2qC0cZWgSQfyAWRtT/YzffcZ0mrLDxFR71MLYTzPds+2SH3lxE
mzP9cM2jXX81jA2sEqfZoodZmmXQ9LjDDcYslJBO/+imL5tK0yxpu9yCYRtskwne
j9TGiI40HxrS2x8BDqZoxNkl0GtdP6COGmrWpKgTUDAgY4fWTaaBtPTG38b9ZTST
2/VDvKuxL3zz8KMBS6iHyKbh9hN2Z/4Ck4Zt9bbgjRjAB3L/7c3vsSu5qcZsx0eW
bq7dVs+wqmUVya/9yPDuvLm2xbiLSAUNYKzG47TKTUT+MBCcAnLQmvRWoTIZHSch
7N5mVBlrscDQw6wg316XF3rWIeTXm5nyNp70upeS13mDjhmzQPYRRezSewbyC5Ry
pkrj2xg6RfR54r1ECZM5xQI1Hj15TBdmh7Q99fBOiyffJIk/c6CNj+viG9bk1kYC
z/+FUNHw+7VQ5bPu8G/RSzdERiAcZ4p1T+o8i6nXqVD4XqhjDDlSRAyi5mgr9xOD
QoMrraJJrkPiij3Mwv+Mom1jsBGnP9xnz9mM2GLSCqzm8iK/y9OK+4u8tGBJJWZb
QKjdX+R45pwNYKlC0EQc/HhHKwn+BRcybgcYUaLTPD/oo6mg7r0QNi4kViIXjgWO
xqzo6RJAMehsHllJhzMxEdCbgQJ8HDhNFDHs1loJgsTUZVzcaO/zpfDwmQSZjARA
GDNY2adUNRAAp2ib+CzpIu2Om61Ia1o9wqByxnx1XBbNmgXSELsG1NSVelMSLjnS
hwRU47CSxLbv2SO8myz3nCtDdjQFap/cpwzCDhtQGjUjTxN7or9S1RE54lvsifZe
0JgYyoKw7QWqGGhwNHkoaxJJ4M9AwSTphDoJj8GS9xT0frYjw5LG7gbZk4fasj4t
PDuHNqumhAM4E0+6DX9r68vAAmQD2CFjEVKibtOtwxm4uF6/286XYgfJNLsUSFVz
o1CchTknMjOg4hc4i+Tq9/7vU66qqag9+PKFIJ9NCCOdHXIbpXLuoKkyQBjgrMO1
z0WkXlCjLXi5TcZW3SP5DAVtl9Oo6OWz3QwHVt+fD+4rYg/JfqB+AKsqXj7r/lLV
Ex/OnclXD+LFywaR0gnalrfSIS4MQqyK3J2Wgy73uiKqwNVeKyALbaoByjIMdsJU
N13zwvrZxcmov/tyl2Q5XSQaOD67JCaVedv78hV+z62GsyRXci0Xgp6+YxjkA+J+
D4uyJAuDmbvaVOXBS9MQllv6Y0Jkw4iPmiAKFsQy75m1EvQl9B4a0lnbsEluqC5S
1F4w70LEFFieu66EmKo4q/tlHQTkSsWD8tSU2FFWfmYCgkXEVKEFoUxSrT0sb+Sh
TEfeWcz39Mc3fbZohrvHnXCDKN4W0z1MY//+ZA8fbSr6KIeE7yKSsfquLKqltQpb
kkRpUgRZugKp75/a1XrmjyJjvDTQqWu3vxZAHRMgE6VR9CZAgk6lwZ1DkkBUHHL1
p0AZLQxWv3homKhO1O/j0SznWi036c91aLdn4F5KLtsiDtIyPqu5PnUwLzIt6KQ0
steomcng+2SYtc8tiOH76FWimg/KY7g+vRFUxqupfeASD21DT4foeCWcUx9ZRlZu
wIBu3JVGYBZwALS+ViPEvoyLSCIvBm7e/eqEDZXPrZ1/ATqH590KGufO4hGydO6N
rZ9zaOjwmr+g3dtCX827Agf0cns4LdYMXjKb2f5sKfah6oxxhKvmdyi3bn2GVKpM
iI+E7zOw8TJuli5VHg52b/fVCaD8MZY4NGwqXIxJA+H8Kcn4wIaUz9UPJMwcO5Bk
m/mIYXjnf+6JnlEhqepZeQREfWOyXg1FFO1wr/33HutuMDRocTzmWOIR4N8GWkL2
Bi5OTlZz2x3aD141EOIrfpWel9LifxdXod7h05q+WQrk8jr/EecyH1+zU7+TrZSS
wMgLCLLnVbKAAe0/ELJ3IPkQ74+KBtKgyGLhlYLlowOnBpAB1Yf8H5yPq15gRCaR
f0hqlAIcoQz4lhCdxXL01p4F5Lep5IyN2Yaa7a+o6DVXHzpUWJrMY4n0pNvYHXpa
2ukH22dZUPzdeYMnU9RIN4jbu07Pshjp/Vqk+Apu97xBC5JSYtfDqahGKkTe61hK
qV0eSPcDbajuBl7kwN2C0OH/AddVRWM4haXBpRcuq20PVU4sh9T2dnDJnGHcIrr/
9CqUCIkjSeLva7uyW3VSBY1Aor0tLGRWQTALa9MsjX85q4rOwl18qmnl5lrQm9I5
9NV5pne9uPxtE3WxP6Hr9Zp7hKSy3Xt+/V77BcJ+natoiD8oOKsQGWhMTyojosfR
QtbBQK8aPP6Wcg9oeCWM2vxXunt3iJIlF7ZSHlkSgw+xTv7XQg6QsJVK1dAwjCdi
VFe5VTeapTD5EF/BHcIzGWpmfpzM71x6fCiiIZHRUVke1BP7k9DHk3JmdZBpDUXp
i1ER07JCT3Fv5Twlxi4EySd47R4gh5XdoyDW5DV9/cbmlWTKQODpc/8sK/H40/4R
IOlnnBtesPDDTXXSAXEcFke2CRGrE6qKIOfFG4vMEXem/BiR+yJuCtItyzN2b9fC
mwfWV7hV3uKXnspgx2aOM6NJEODXvQZONUXOwWmZmcftJij2vUsxLgiLAvwXCVy3
pw68whj/nS5tlDyJogmPL5YyJZIkFhTXENA+gbppV67N3CYE9+IETO9HMKe+A9u6
EVSn9+zUgz7NagNAEfieuOOLakrjbqpIHLfmNl3gocLdr5wqmq4CfhlMvKQtHJcp
BwbVyLe0i6iJvKWKtdrBk0mSp95E2XaZ9+y86fvQwTdjUSy7NFfTWNTb7kyB2Bbo
4824WWXK3bT2RGPeN8YIuBxXlQBoXm31JB370P4+O0y0Px3LISdjj0SJEJBej1UC
MCQ1VFeo+1n3jyTq6h8CkxGv/5cdKaArj/cUqZvOPgK///9d2Ey3U3mgIXwfxMbt
2jYNysWK++w9hOWK18d1Sl9aB983TW6H1OWWnJYIPZ372kgEOQFsUhcu0ZbeQukg
gsRRKaLef5EOKuiRIBsxuOqrixwMJ3C8vxejM++aU24glwModTc3Fxl3UTLRuiNu
bdzAvfEk2UxxKlThjTqkX702qmatIVgcGaThYK3JAhf7jlgnO+Yc/IhI54pyV8WR
xD2/wqoTKPzANJM7NwwDMccIrjjoSQLkcseKNLZn67q3ARnTeaPWFqzVHyuG+lXo
vH5rbzJntouMqKC+/tXBBwm+WdTBSCwf1zGTaaEoWbrRcuN5LEeFhc1v6a1S8BkR
QY5AgRyJRv+7SBxATvCdSZ/l0uXoznMnCIF1omkQ8du/eSogj57MEJ9gn0HaIENg
O/v9zKn9D1qLxPiEbAYazYGRnS5V+Tljv7C/0CokWYQUK9Yulzfmg6mG/19cTUZx
fd64EH0O0XOTtqqaUiqtRPG8j3nqg1Lvza/nOVeYVZBcho/+qfljmkHWyCbPY4BV
R9/F0XWgqml9eS/x/fz5WqnPJ3SzT06ej+ITzndubZmrkhYbbPT1LdLVSYKxAH4Z
jTYub4dRd/dbJPaHXhsn0m++zkKh97h8/4lYlc8i9Zk09lZK7WyPMrmBpTcCPWYZ
t6c6tHJSyomWkuG9alI/ZyGHVLQwjk5ogvzEoRubMzPpTecQS/RsyATPq8zXHLW0
/hWrKcs8AESyU9KYl9eUR8da/XMWV+AquYR2+MDNqIUtmvre154PWhEY9iPQ/nY8
3UVdgEHUZPEetS8xIVo67IrbjsI8QlI7gDQPB2Jj0SWuiw6S6VJo6yPLIMG8rtKa
eYQymktgT6qbWHrPfl6KHfiQrOf+XJRK5833CnTu4/+fAvTkZj7zYzEt9iZgcEsm
WHDUzxy517lU3VDOthsu0sNYY0BDCwS73xvVChMrAzg5vCNRzQkm4xGIaxRUu75U
Mle80bEkWSv8xJJ+DBtbZsVw9Z42zCEizJb7tFEP0E7g9fjW+suTf6lBaG+p8FyA
1woV5M0FLuUWJNy3bg0TfjOluSumNoBDy1BKqVxaN+J5DGYIV2jhojSqFeSJ5KI7
+7ESSxhBRHtqONVk/bXG4mIVeEfyYmljsKTV0u8jQY9D5glHzH2mSWeEitiQK5cM
qOvGJtI+ZYfkKXwy3BvfNq/bhaQy8tebSdk+XU65VUjXGEt8GKPEK58LJV/7IBwM
xwdnudVrzlGx8g9KYggpiFDb6sI756rF3+au1PPZIYUATgADTe2EZEoaD889i7rW
rK0dokS/7fgzBlbmT46Bg+7sN+Qje7qS0nCRVwI/m/bQ62mDz6FkJGPdnr4TEkpg
5FGYbWnppLaQilPXxTi7qMjRYuwnr9u9isWENpj5pigBClQgF5GBD8leLvY84lNb
Fk1lyNLZDuw++k0oOUBS4llNBmOdIsCmHwCxnl392VuywNSW0l+8gQHXTrXpd6jo
qWvZlwfI3whhiPkrSKQ1arkTNGazeArdk5JiAWp5T1zCRCAfdhSiFy8IXKfDQ8mv
vZGdilxSNl1BUigvLC5/f8lp8l9MQzDQtxIkwSGmrRxkYalWXO5Eq68j+tjZc8Jv
rfb0KqelqVvf6t5rJlT7hU3L4B/ePM94bben3SOGjtx6QGw8PT540Ueo2PoMzVcL
jJn8hMUf/fUYchLqXlxVy1jSBZeXXyJGJ/uGbLw5DSi0EuB33XCZtQ7rkjizzHIw
05B3OVarxa6jUgW1OEInJiW22IZcMfUKl7ozZuwC0az5mmUelVytUO7MKMIOuxYr
9jMVpi+66E2phCo+BYLxX0CBOdZ1h6aotdA1KYbeSYa5f56rcQKRiTuGBTwkmg3F
iwEl/S3/zTynLx1HggBXu+SxDus9nwbHMrGMsBvUCyseD+t0cM3dzz1hYQJ/y4Os
CWuBoQEjQmZ/FPf18aN2MD/9hjfcoP11Gd+DukMKTOEcsaAIuuDLG7jNXK7gKZi8
p85+XWcSkLiO9lSTodo9yUUsl3UEIKuAlNh29vryZ8jQfG2k6Ndy129JniHFQUnJ
E3Tqd5H7udNapS95/NgSwaSQJxKlZugd1dIa+hX3GVo5kJWOtA6vaQlvL/fGzujc
9/o6lXUPw3AhrMwZPthyukLE1wSUsWIXg6Fpn74fuGMDmzaIN96GH+6NJ2+oIXTg
ua2LX/fqmeJG8Kwq7MYBkIAx4sN3Uz1Zx1dceTqqak8DjJmaTeVGPZV90/fTUo3Y
XuzpLxogW2loeL8IM4TR9KaIU0VEnf/Ouq1gqeR/y6HS+LlM6rlpC9c9OCPrgxzg
vA4gtFenY2o3/nEg2icVWVnGuIr058oiXyAc3sAwhM/Y4XxUMi/d05G4pnP4GxCz
z97aJRMIM14FvxwYgB3wSSFO0y1rC/pheBfb/I1LM630n+qBTj+pT72JmOTRsBq8
bvZXftUEIw7hixaFqxhbbs15uTXzEAkiuFb7KXE94GHEZ3L1mQhaIuzeFUskEpjw
xKUnwVAHY+bWfN92+PnAZrAs1IExqj6EDqWdagiUaS79GXfap1P/WK6CLO2jF0h9
+ciWs22HUJWyO3HvBoRC4EqHVn3u9KXvL+EX7ue7MN49USrCqoUvdISp/hcauCYU
1KU9qkhpd662U9Muhh4Hk1iTRW3Asoc5MOO4LVzVhnDB5AlMjUmR7CYNCDdw/jYk
2Vgu+F5Ro/f33o5c8xlhEvJeQKjgF0l5HIdeu9ccc7MOBC+HCKBV0/+kuqsx7bGP
+3P6D16+QEgVwzSEC92EeF9042wyotOtdDB9bSVDpUlVB7UkRcJWXHgklJmNiMW0
+C+940wvT+ueuU1p4Cs0dpxcOETn/oKUIywPdpHUJDbTp+88epZxDijSY25KNlQD
rkNFChefqB6u6hvBFka5tbmUgQuXPPEmfSVDLFpeI+ZOZopoCV43j8Xvo9XyzF7r
lESZ1SI5Vsu4p0p2puKZ0jnThYe9ZImcXK+OmTRQbKsm2+LiDYCLpF54IX4sU/6i
KiASINNf8gHSxY7b1pxMNhyMgBIo4ghMBWK9blWEEKIF3pRR3M7s90QD3CeZSh50
V9khQ0vOp5larCk10zJHhfYozKUV+UcbRymgJCJYpbpIPFgszNWiEsCGDYHsaq5b
b4EF5/1/+bZnOGIVa040a3Ien88dS0jpUOuft/H8nlu1tintbgFf2sUpQwU4vRAf
mpmYmVRHd5esOalQTbTwTmyaxEe8dfrlyotccLbqrZgd2oNiBk1l/6N9YjuUAlke
Y8cht/J2sLA2gyn19OimbQcmzimOQ57BEpGC24xLj6IJaYmRyLQxRuH9BUPPyOzH
O8eE40WDFPbjwZRWlloIkmetVsf+S32wFDoIHz5aOn0eJ4G1qAYFiNZpnlP9jnnF
lwFcGtRLz7Qyc1JxC/SQ/Oz3zram2LaOzWBsf9/GcHgK4D/eHX02NrCGiAzwPLmz
Vjr6QDVx3K55aOtZsW1/9dJ4HeULAw0a/hEeUnXxi61GQXHNEzqSwo5TRCkm9PVF
diIxf2HaqVepL//U0A38MhndB8HY2B6fefFZIOIxfTFaFY39L7BzsMOEbXU4yUhz
iUydbSzcUVMlBQ9OujSoFin0R50O55kzfg4TGAKo5+YslvxMh6L7/IvvOFHi/Uk9
G5JXT4pSLpDqmIgNC/DCLADypCJGHX8awyGdMd4GjRtA09+oaDP1yTyYuYAMiuaN
XrN2L879bACoI5qMkjOrFU34gJGzdikKUvyWyciChCaUU/BgKqTnzWu7Bq1cA/TN
G6YIw4XLQa+aeBp7TH4/X4jLjyYgjyx9W6hD2G6t/gWXhx32xAkJ7W0VoHzQKs2N
fQRdnKTMqbC5hb9ISzTZlq0WMZPhM46V1Iu9XPO72oY7AqePbKatmT0jaD5150wv
p/SY+/ZDmoI8xsjjoA7dc4YPZNG6TNRw7i08BZgklPiRU0e3BKF3Z5vWoTHajCkQ
sXyyFA1XRQvItzXMV45AfuJWiQI6HiC2tsVmeWue7wEfCnOnVDNCQggwj21velTg
Y81nvdPH309YEIKW8gUzjQH1/kUrbliijgSDSKo7dmzPVs19YDi8h5dSjmMWCMMT
qf7d36Wvgjc7FP3AkBfACfjxCdJgTUn65ap4w6K6v/e6ESTWpXYUvdYXNKu+6qEI
/93vg+WKlMwfMeQwENBWm2fkR5rJ8GOD10hEyW2Y/RHT1zaegmJXB0HU10/+mgpm
zo05KWiPAl/ycP2uXXTmkA3HgOB7GulSwwIMfJARpDbK5msobX0J6z96ex07T+Yg
SjKKlRCyagKpFZVnCc6L8+/NySpHz5GvPu0MU2FJ28huTtDSLXQ4gT0rJlOQZb2/
y0XMjksDDOrMchDCdgAG7BNTF3oU4yMfr0aQT0jrHSZXLvTT1vEkEvwHLqwTRWmg
LRJPWYl8JOB6Wol+PRPCcGpJoL/gfhVoqcYLfwtZ56PR/z68S5Irsz3H34wIZOE7
c/VDqiyss40qe+RB+9yXFwf/dsiqTIKoQ8dzurOtz9DCBmvQWMzwM9bs37gikMwb
KA5EGYe5sYQ/EX5lKifcNbh7I+0JnoE2nwPoCI4cDYQ49u+7k1B0iIb3D17Z+Olz
4xmG60YEEhHcXUkIgu2aI8f7dRpgPertC09Dx5TXLyhn2Ll30gj1YCEPCu8GagjE
2NRwWAfs9xeBOPpK4u91/5nedSoT637AUbhPogWWcOfchnC+Cb/+/vnIsnAO4RsW
gze65AP1JQiH99lysmSvuCNUJCQP+PLynGIRAktUVZ/Hfk394kaOxi+pY7OPr1Qa
xiAHG7Z1jWXlqOhcbImBhVxQbwmsqCPaz/vIY/7UN9W2BwboAQXGFEBTO42kpkjx
OvdS8MviXnADLrKtgEiOz4E3CQb/v8p77q9AAEkpr05C4nfTElAM9n53Z3Wk/LEW
HrhLJo0pcgkxGEHtLf82RGyUCZxzwwByqhiKnsa1q935uWshsBSK+/dY/5hhomXt
XLcMTuPp1tlmMdAeDnzIodPykir4Me1eTx9ZzNIw3DjTYGK8wurrk6MLBHXUR/PL
J7L3Ey7JQ6MzLeiYxWSPFLz4ppVYZTiZT8HmFU0+3QqG/N3Eqm5Hry+9FhGmGYbK
RetsCo/1darquX6jDHyxsYIFhy/InhiYj6t6dBkf2RqtfKt6AdnDrX8TicJ0XS/1
v9IgyTjMO9/ZGzV7klTbQPfG88sKd+oMmQbyaeynsuIqEQ76UY7H3wqe1eSGRxA4
k2rxk3QY4bvbl/+zD57dIslWoLBIwMB299Jeh+ARzEqAE/1eywkFNpdDnOB8DfOp
E0trzdL4E4t/KlsPuoKE4RnI0aBkxM030KPhqgn9ErUtHhIzLDD0tHbPats6yZMj
QEH4UtUOnQuXRHPc0P6ina0QP5l00EvKHpy1vg21bAj9lTjHrWwklkBRlOsouFS+
f8ipv5DAFD3t0E9T75kPqAR0/bC/9LdOqgP7K6Mk6laKtwaEqnPAfivAgjQ5rhgB
dqfiULlGEB2uD1b8rNReRR7s4//ZWWDg2syIJaaWrPG+hjbbWUJpOJ6XfasEKjvT
3D/HEIWKysDH57d1Lk2PNGeuCoGSBz8HkV4PRSMY4nvRm8r7vRa5dEmjrEjaksnI
eYzH7RxQv8m0ME2njcR7evBs4YrLeUcdHzzdCkmQ51Wnur/7lPANQslOyVqDSBG5
AbuMMI315BZK2mPU/Ow58F2OwK2tngEI4knL4HM/T5vhcTN4Z+BjbrGnIH0MvUUz
hAieRTk+4TMe5YElKJsprHFm87FnuyzwwBEsjH8u4wVRMR8BLCMeWqzFHOXhyK7c
KFrs9ePWwXjGeT8HBLVsFmOoXfQtSthZN37mpFBloTO3ZwDysYfjjDms8T4ncY81
68UnGLboayEeegOgMpK/V85gTjPiaL384BSmCktH7PaBt8yPbuK4YAAx3lAgFO08
gVrNr/QazPvuy/YB3ECoSrkuDcO/B2twCXbI3791OnXuD+XzPHW4lw+amNPcCMN+
RXaWx4t6+xkKs4kIzwfJZz6HgFqkicBUkFNKZaxjRJrvMsF6bbDOk6sxpyvS1jMB
x83mOzPqkoVTUD0wpT2QyJ/i3p3Pr5WiA6o1mcaPvnAEeN+DjoSeMV2dC/met6Ze
8CwWRR7sj4emKRJtN2QQZpXG2EmLxirQhe7Savq3J8PQKpFHLk4vMQ4k5IHoSU/N
YdQWFmTB9/cJ+m5AmkXttWIhYQkHLaPAVDcZtN7Tkvlbc0tnteqi2R0/dtYMPgRY
/E7GsEii5mM9cvZJ+k3ZChV8o1Gr5kXXJGBkWPce9YlTUzAWPk9MxONzsmoCbYel
+X5pKcgkEB470S2O4UZ2BsHRJiuPdo4VNiYRskyWMJa0gwe4/piUWipsfLrNcNTS
Cm8ehhkKgw+KP3aN443bT7Bf7JAoufBc1lmylJVa5XpQmgJCJEq4AbFMMU5+29X/
esAo1faA5Mpv0A/3FtKQcTObZSpzCWxf28GH5Cer0nRbPIEvtu7QHc2+yTd2zK8x
Mk0A6oNc3Mq0x/Yk/hnEYONhGABId0A9SB75WBx7hE87eoBSxV3qMP8bMswb+WXy
Gun/zRPfiov7ZzWDbBTKY5XxG5lKS5c9klqf5IDH/cGAvcpq15AtoCl2Add7pycX
sYOzwOLtyhng660CEu6CoZ1PZJRLPEggfl2hdmv0jKlGPSmjFC3dyHmLZHdk4q7S
3YPrUzQBbKl7l8tILyfu54zB+M2Ap1YPcMj7qhp3i7l6KjVPdR0eZY69CNAtNZ+c
8lygSf0TRiU5WZ1uaU5/cVNg2HWgXxwXMUr7fG9JHYhQBZr+hnSHWMWZQcwXCVe3
/74eNRACuYUQ7s51asCZCIBg4GP+Qww4evYGCO2KuPVDVVvMmGglTSl4AoAj5r+g
vxELbxTW/4EFSRmzMfb0OKrTkJm1gpD0yuP3ZsF7n92A1XjZ0Nj3b4d4TanOCOkl
5SWGvOtdDZC9Iu4l5UQxO6ZGnScDsI5/ru6zmMfEky0IDJDD7n8C5cVTXZyk8WhI
LBC3vc+Fsn81sfjK/wYq70CGQxCIQNXRZjm2UgEvEUZiQDesYkIUsGYoXOEyT8/H
ovGB7O5iOba1iKkI18quUCWgBA3Pl2Q/YrDB9wDAv7JQztqMkVYx1J/RmLEPRwCb
XbrEhWuoKBuyEy1JDc+csvQxbN7/iG9MSfFSavTczt1QjqxSiJIw0J03HOj3A4xe
fAb8GkNUx/sao5dK0zM6EVUn+A9xmJB4RQjrpJGzSr3Q5tUAz9V9PR1uKgAJCKsJ
WSuHMXcgEoQIkAjElViHuyWM3AI2DVugmn7IulwZJ2F8l5x8cEBlQqdBx8ifZurP
f8Lo3gEKIQvzT7cmLHusBSIksS5H2kWcbeTJyREJBf6V8OVJTTRNqbCVEEg55lao
x7RDdG+ytxTu0BO2lgdYDs332/19ws/Uc2ZbJYHa7x3Q9dYy1aILKUiUzPzkKU4o
KPJgYr6Rx8q+fg29yNc+pR2z1UK6bSKRK6vC4UfaDzF3YYAspNrC7TIaHLgatDvS
jVfmDsFxwRKL02+Cw+Cj2iksAoOfl+Vlcb0o1gyAAFou0jB6fp9ZILsrWZD4p5Oa
GwjlFa/wbVoi3LINz7CgzT5XXIylC2jJtxx/A1+hAI5JinNIlD73Op0kVTB0V9xt
lvKxIn/bx1ltIjaIud+nLbkP44iqZUMpiDdQA6MS7VGPkjFJuCjoJXtuzMDUsbB0
Oa3+a+UBzO/Hz9smyjqyrLQbjEq3GqlIj48VK76nTtYGXtZbFNBOH2GWvNmC0uBM
7CEibu4JMdEALq8PVTjQ9exXfNmsAX+DPcUxphfCg1mCEgzyLTpRunHC6FPXsbH7
JMk3qCxQKu0yKiFZTK2wRc+j9f0SWH8hrVzaPClC3AJslMKU86hktN4c0l4trfKR
A5+yRxWTsEOb3AXHoUKR9OqDV7pxOi9COA3m2+SRbDSqM6XQfLqMXk7qxmHf4iiJ
La/Jp1xp3G7WyfWpNdY/hyE1S2mcxdsE7BQsjsH1b1KsuJaja7pegXMZQcMTBdjU
VvMSPq/n0n/RvZaG4x9Hh46ikvNIRVSubDnLfA+eMOu0lVhZmZCz0W1PoxGQhtcB
f4WkCdDcLXDivnbgU1XjMhdBNBgtp5fU1MRnSdppDW8IcZfdu8IYxzt1B/LHuxCf
4UBRQMIF61EYiqgSurX6Ju7CxJh9VAMpFhbyu4BSjlHBDFzaa5APjelUIB16YeHH
dXVs9uCKoUWRrjtBIqhRFVHgdgcBQ4YBSdiR5F2LNnAqxzZB0mk+ofTc2q9bIhYz
mXCNLjHs5MuGoEfDBdpNX51WyhrXa6VMT2RXW48icaJIReAs0Yc8jtDP7kOlpxtZ
gCAm5Q/6FqlzFCv6fcBUnEfF7o2bGXR04bK1nauhyzeK94dPzGJg3P2ZlBXY5hkN
hzWrhPCO5B1pIDZd22sd6v8niw/sDKCio6nqz3WVP7QKdVbHY4OLet+Jd1Q4sQY7
ntFAFcqTTc0zyImhZ9IB4yCUMfpx1Y+WompnG4IiB7jXqZwtsdLEuL2eMXYLYxl3
D4ZsBFeK8Vt3NnGwUUWJ2OFNnOHC9X6X5YEBmozlMRTa7y/+LNoFymGfCV6zN4Q7
2as+ylDUxvFPPUYx0PT3ZLPSNapYIW7+qDTQb744EJDIwF1+WNgzSjkTp38W8FCP
bZ80i7btD8ktYVT4uGHHkB168ISRQBjN75fsAX//YWrPqbWEPdilcj5zg7vQhGdC
D5axobiwJw3WRmjNVjyheHOgrk6TwoCEyV2TvjH0P830nWG3PnVSecvUXCbCalQO
Xs+SdkVRUy5FHMdeM7PmoQ5LQlbi5psbdDYOpZ1FhuFckMzn91tgX91GaVgn3ob1
ExVDkbzzufRqha5Rkan0M/HUxnGDIYwiszOICSR8s3JTG9pxh7BPgKvjojM+uz+U
IsVXUUSmFdRQXur/Gywx15chFRRlPUq6HyDqqmD02I4smPeONF5I5wVtaZfKE5Vz
uhFwCGDxB2cNaOWqdDOcB80FMOQDsysP94SXxy8eGZUWq/1H1eGxC0O3ltVC8bgM
eQTO1zeUPO59wJw68rUs2SICju1dfrVyFxdsqe7HYc/YIn0mKI8LI8TBwYyAlzGG
OjPb/t+opcbsTtlBYrGaBvBxgqby9p+F1NvMEqqx5MxJnZNMPtTU76H7w9W8YOWq
/7TF6828ww/o0Y83mKEKpgmqome1nITZAPjHEpqTtKJUsCpEJCe3Yno4+LOfz+yu
6DpJJI8flPgHNGq4ktHJGZAdZYXkQV3Y+sbxJXqzDdl/8KjpXQhJOVJRl9Vbi3vp
aZDk1v4u1B9N93N4kvo5jDuZkg7Zmu+WcMjRiQ8sOCkFDyEQA4ybgux/eGrR7uIU
mL4mzdoVyv0qTEK7HkWmYn68eZKKovQsmTj7RkBjby/F8W0Ylhr8YxM9dnz5wDu5
8niGxqexFBJjowKhDqxE4GAyesrF+vUOL82Xs2aIjE/83HkcoKkhX1/4TkOJXgsa
gSBTzt9Or3Dh+GUj6RhyrqmOi3tX0+QpMlJ1n/LjXztW+4f0q95O02o30cInlgDz
h1biSGwUbh8AJSkiSI1c2MuZtRiUOX+dxb27cksohbpLMV452RlbEUiQZofNMicW
DsMlWSZpXGHPtPlOLLHoZQmW6SkWzeMQhOcgLKixNGOt6gbC8aHAxU+ouViaK0dO
atr8DvIxyClDFLL6eQ0xKw==
`protect END_PROTECTED
