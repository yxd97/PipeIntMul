`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMnZTWu8QZ5+BvLkqQMkKx9F0plQ77//YgHBEhhGx/83yyzZZzy7KyxJgKkurFgm
eGXUCdVlONinfsn2L6zYjVh7JmxeuJagPiyZ+VDfVfsF+7EVDLeT/g1U2rJp6Hgb
qwxun8zcqn/QgDjIS25ccdej5GpRjNjvsbTnPzWm319byM+amCH0qBkXyybWmAIk
KS8B1oYC02v+ZEYxgkydIdeZ/m7tlGvpoeb/YHTlv/bDzjIEdHNqtIYC07DnOHEf
WOLwB9gAnJgOCVK9lS6DWXgHKP0mhDV5pvvLgqqh+Bugd9ST7pZ412UHkM+6DGze
ZPChaBSZr7uz9i7u0Jt30Jr4VBvkLkUBdvnxcB+zYziJaP0+ddZDe8QvkTFZdHT2
DtBTR2ajN254Lvk+5+NeN/uUovID4pJK+7IlVNErmZNNXolPKdXo/PUdS/9gEJkK
/CFdi2KiZdOLBceOavMzzP+4OTbVHNQUFrmOV9utN9oBv6y4hBBfmlQuNGJDG+fG
K0Q2GI3dNFA5rDxQBKM//pwAYA+qs+HtuVMpN/gx1gtGXQ7hGi/RM/QAqQiUNIhI
YYwMcZiwX3x98wPHetePqGx3xt7Vl6aPbxiYL9QwqC8hpM537orHD6qQLVYPjSuS
INHb+DPBarHsnDfX+Gs5kEcwRDNl7KvDFtWvOnZDre4tXeiah0RIh5q0UDP33aRF
ScweOS/dh4fF0eW44ZcMD0/s/L+W3W6h4/S9Dg02fdgQ0yAtKeuoWXHobJEEQ935
Bd02rVgOnaP5ri6utSzSLt35HuC0TlyDpkXcviSMUu0Zlb5k96FpZGgiyKnEnffO
aSJxw1jTKNhE0QV69yUZO95sPqUyh8LyRjLTA9oa1+0zXHq5eIIx6A5dzWD8znlH
vMVJqmVueB6BO1iAKxz19O4e3v3JklOJkmVTJomcJpiuXt/rg9FvbYqTx7hv3TcD
jux5OCeoeE26JINF9Hmz0tvmc1ierYXbUuQs/FR+6ufXynLGF6wxmFtTtF4kQhiK
OawSLM5EaJjYDz/Wlu098P5UlltWvuk1Mamrth/pmDhu1kV5B5BhYL/UXagjsS1x
ZhmXdVvmr8v4l3i2zlWyVMN0/hiZcyT3lTu2Wm1DIbKSW2MDN2bPBO4FKJCQjBwl
jWNdBf7AUSZD/STVALL0BmPTDZprxtVt7lnS66MQBm0=
`protect END_PROTECTED
