`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CbfGvLmssz7/BShe7CTXvzgXpC+VDgww7uiIuEceco3KXfuv/0ffuPz1aEu5Q521
cSX6sn3cY51VzCcrWusRHTkYqtyz3tPjtGzRtg1EPGtlWe67ubVt0H0zoNvxD2OW
l0fle44XS8mqLPRv+1UYkKqd1zbE4BxucA8TndIhL9Kh+/IPtNCT5+jmEnFWfpAr
J4CdFWrMeuF7m1j9dXZkh2+HT2lC0a2HdSSPBRHVetHlv+nIWcFM0usRzHE1Bgrc
/AzYfSFa0j5+1U49eE32LA==
`protect END_PROTECTED
