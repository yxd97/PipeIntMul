`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qPkHfOVq2cv5M6ZmaVJ5PbvsOZpsCPZOk0ZVYBPr5EbvCOBKVb0tP3DHt8fabCkC
M2AYtS4cyUDLsVv0xQ08hc6VnSu6U7K2HvzNrJhqev2aEzx5tOBeeLBmTVfuh0Mg
rNEk12QqD06xA0/jV2hT7VE34ZTeca9Fo3cMmjR98piNwsTlrd1SPAZZTXF/ItlX
gTytiz1bKxac1Z8oAMjnquNSQh6pEZHREFtl/HTrBgwDNSFh4IA6ZrqCbDhPxteW
OJ4IhY6U+z8QLnjzYDgMx4vdpCn1ilV8BJ2cuE1Fb4g2j8k7gKRe6xKo43nIjM2d
+6J0iEJDXYcgWtX+ybCMMg6duCIuhpu4Kpet9QJio+jZhmApTQbgI51C3Nq1uLQ0
0Z10o8JxHBrXvl2NYnGHcIPZZqNEnxPyeBUUT3Kb2PlzC03UYsaXsDp3HEPYUMzi
OTRUY7ruOPdkH6Fb02WxIF5gyxsn2LTyWGhGY6BXmow3o99WX6JWuVZR6yE6nC58
obaY+/vkvNaXbFUJgGNu320mM/TYZz3Tnak4GK7ISp8yZJqhajxZiE86lOBFSE0X
1heQmx+VpSz6FdDzqJuTKOm1B2MrIupvyEs1/5B62l5FPpqR2u+uJ3xKetXLd/JS
GhI+ZFG1YIeCReYEWS0CP1PsKxZfusWgf/4yAmMQeweHrZCrZAcG7q4apFNN490N
9xHA22INfwcVYzfNTM/ZpKCtye6ugZICWaI4Fz9++ILiCzOhFmJJHOkPdUJnBvkC
7nWowPDrdLRhX6na5nWE4kyDE9rAkqhTlOREwibarW0DtzKo2OpedcHjMReGPTGR
lny2CrO5yhCj5NCl7cWuX6xo1EKGU+NUKcqS8LwAFGYOM5u10tExh2aYp+7SyX/w
npWct+2PnKVSdcPdwCaXfW86377vxI4b0fEW59Z8gTJ3ctnbRQJly4wZ+276NnsQ
NtONknC7J1FYJcGVDunQIF13t+fDYsAHcpF653Bf9m/qyOT3gvw9EECDXMY1cbRE
+jlb9pha9rAvRqGyaR/a/dS3LvxK3viAhMx9Ofd/nvI8YyWvWvxFHW+so/E2rHH4
sPUgTtB5CrHUmcjKCFXlzN/jxbONZt16VV5JbThbW+KRBV43Ij8bDBX2Cn6L8BTx
AiXxkO4kXAP2VRMTBvEvuElPFPstEPLOQszE38NYAA8jGlkEUByaaj3aTJzX0Qqc
Kx8Vk/zC/4hu0+iLnA/+uS0OCBYJtmGJb99kvuZvvt+7y0Vai1wJT3LaYpgcfBRb
X7CT/nvr/L2ZiDkQoHSIDJo1ZhT3UZbz5+DTmabZKmu++aOWr8FFyt3hN6Xa0CT2
HqaA3EN276lI8rox6GL9rsVMo9BN0w6vtx+U0pif6uyAcPgI/ql9O+xEKhd2oPkl
/Ta/wDQkzAetlzt8SmmEnOhgk6/aSYEDautKgZ9dAkN9sDoDDx051SFeeK/NqYOa
WbT8EZAxQaMXTvwzOt/ToNFkSx6FpB5+bM38S7ySYbLJM1lx8bMHm/7C48ukJFNj
qn7vWxqRmWVfKTf2D+dEIqteHvswXhM2ScrMtl8wLiGmsrE/B5FBK9tAGV7gDHfH
s3qVcjUjPHBWRYNJ92ESZofe7qTiqjpbaZzkRoL87bDSaoPpAx8D7mpS/ubRjOgV
+i7TJ7eW964yLJPTPd89KV/RNKbxDp95deuoDt9kIGqKIhcHpM61O/btybFnnWPF
EdeRh0gLpO+z9dMjw1ccLuCbHOgKae3APhiMgodXH9IyL2RRyK18ESxYYspwjtdH
F1w7Tc5ZJirwhjV5LQaRtqCSWO+J6/59SH59qNnZcwDGxqF1+vIpO/OiKzYAq64S
fEa/nT7V05xntM81trl84g==
`protect END_PROTECTED
