`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yhfqTN4qW755Nv8jTrFskrIW6UgRm9Yl5lWUBfB7WgfcaBhrEaBXfaQvh5ZJbNKd
M8JejZsO5gSKrzCjFAnqp2qjutLxTVITsatyoUUcK9ia+oolh3hwtapINJUKf7qo
JKKqL+S8ZKzDx/9bOP5RONYURaSqZ++QFtDEe2TvJt+AjV1O0bX/+tBOWwihoFN8
h9Ankdy9yLi7CV2EMW4omKDseR9qN8ZKGTx18xVKv91c51qDxOCU0qQRM567YA+0
ZlHvyseseArWrBJ+jEWiYNXxIsK0bm8Up0OYkQeEAz5Qg6+PhGR1Ex9ZlngVoV8u
1jtl6jMLPiTShj5Azzb8ovKn69KnfAsxecRpZvtQUhUqr8y50VvHFI3VqYd0BgbY
WtRb67QvZSRKOs8BVyPq2P1IqJJGV1+B4hOcjviLpiFFag2KWmRTDIVm/4ncWhvE
cWXAu10Q0NoTGdgAMODTrD7ZqN3BYlrqKeysekmakQk=
`protect END_PROTECTED
