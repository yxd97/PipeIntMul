`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXSX1ygw1mrehWa2ahDfMDCLfTi4nE/slyfZhn9zl4GVhcpJ0rY7bH5LbAdxEV03
8exkEFNaWOoYmIV+J4m+yubPkvaL0dKFvtSPsx/SvDLMabYeXVKY/ZrsWpQLlGfQ
siEzHhmcNAUEJBvw9uolYmTU4BoZc6Q+ix31tgMOuFxfOIpHRope5AjAEaxMlB/0
YraaNfvXE5kIC69hb3p8Wbf2UfsjKv/NDIaUOCzx5QOUCsjX59PQxk7FQbEgkszI
GkTGdxX/YVT61nGXIPAWD8m0vryw7Dly4n+X0KI6s8Un9MV/Cgjo1YEY+Sopc+EK
0e1izRZgHFL9y4A7MOu3+gFGSOJ0XwTjaqtaDZ5ChjLLexuTKWt66Rf+oZejbJnf
SmHMqjgAWsoWA3Os6CebIjb6OcSwkKsQX3c1Jru45fpuEC1yEPrOBGn8R41+2mT+
bXzb4we8vVGsLXb8aCii8Etd8gZZtTwKWJ+R8AfKLh0CLKRy6MrigUUP8Mc7cy+Q
1agAjSdMP4k8n6k3MZMYByVTsW4YStW/pHiuJF6QFUXpHyHLnSP9cEsackjfjr8Y
KWLXg8N/YgIk/3IDLO9AQGG3EwF+fEiZK2ICoDUfK/qD/9mIbKLanwYV/9pg7nqN
AjXkoW4/S3122+8rt1OGnY6lVyFaMkGslal6VdqI+CE8RpryPTpl90QpFTyPZhcm
pGaGmJJepmFtWK6otoAqWQ==
`protect END_PROTECTED
