`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DrC/1qgx78bzuFRaDalgmNn4vLW1jT+8nhqamPP9CHo6XAjOGxaFVmkxjqCqshtV
tIMP6BpyRVkw/RiLU72WCWyvewq4FQPD8z9xBAexGfDC42z6lKgUWja4s/fx7TeR
vdWFmf0Fnpwd4vU4Cp/xM0LF/v1zxiQCALO2a4qaRX3rN6wHii8lTXKpVs8KfOlT
g53W2J0Gan1DIjlFAVUjhP7xyCre+UgIPzVXIYYemzxBIejfdkEcyTZvg1mE87Qx
str6BbS4tteKMqYDKflHek/LRgqTOsCrVvhOh2RkXLe34YApgAdLhqvIWklc67tD
iP/qHgw3LureTJ36CEcphh0fPJ+82+BrpXqm4a9zioyulbqm/IrGLv2odJzrp8Sg
mTW5f9Hk+A/t8YkIqcfOakSLkh4gIDNKchzQKR/TuBNUQwTPxBVWn35hEZs16KtN
gondhq/uc3Rwmi4l8mSNIYw2/p6muUk8aHIRLQLPZwc4LBAcMvEXJCr0bnkKe0Wi
pMJR20tKl7xUxq6nf0ebMcfCHPuHIqW6IrPDyr/tGTSeDsddGOYgBEgxGfAaEI0I
0mIxViRHpm0x9llnRe1fa9QMoqxnrF5VCNtCShnXTAxE7CEU7b+EkoQfjyZlpwJE
4PAKE7d7h4f3CexE3i4Yv7JtKFPuxzOc0HAz4c+RjXmj9Y5rjIv+MDBRlzp///sf
b6HxACypiHmtLBEIADDxc3nFbE2peaezg8G0GpLqf5Ut7OSqPrm/c5oHLdehgtID
0MC68sspX8lzKdfZohfAVzv+7WvjHmIZTu7sNcoimC1ePQpVnz/Ccd8rBktCh7kJ
0sSbNn681S52e6Wk+ucxu/I9MFgiTzBXvjSM7bycKf04yNfW2Qq10UhhQCOEFchq
LcYv6CDU8blBtG0QhhFzUtc1rvA7DihuphkFotAjvGi7CBq+8hi9CW/h8B4o06pv
HEmUBH/d4lV8IetlYHpv8w755ZbVXIBPWXtX3Gxl/zqXub3sBWm1FttZnqM9y3hj
zOT7Z6fzdSr6MpkJB57LoSXxs6kGI4Ge9Dd2TOGfBaOsG1TQ80cHVLjk1kxpqjIG
z4i325ppucL+n45kl+jPFc4VUhaqzPzwUw13tP7zR9i/jaWZCuk5uKrRfUZdtcku
G/BLwyXaxy0iV2iteHhh1/c6C/jxUxV5FTI3scfDuvGd/Swrj2U9Ji7MfEU9gZPp
7wJ+Omf2BSb2650NNtYyfaiZ1LEabpmIVSJke+3YVh6/Hp2DOF3Q7A5vTFghyTGW
ERxX3Im12RCBuBGofk0cPDOmNC41wgL5fLlsyaTQb6716t2KGr7++kHtLa/jTh/J
6Ld7DP49Sfs57AgAwADMQ4uYKa1P2LzQEvKs7AttEyixi3GHOQXshN64q9IXfXGk
K1LvfzngdaeFkgns8uyh2GPhlTMf1J4P3nl3kCwfEq7AYTIIaYFbrPPp2PgrIYZD
ZKWNkGkSgqTvYFX4ZwacV6lNwobt/p28yKEqMyVMbqkzvc0B0RcDY30C5NR9pJgm
hMC3kX+pS/52rb1iTcWTpmpyV9G68FOgGiZuCKbcj/hSD+Rvsg0dAzRctQtrT26g
byKx/2PwclV+C649k/r9lVEN+g0rlS509wEiNJs4yquOCvaXuj/PyoYEhYt4g5X8
GZdmYebi3j32lgZBAtFLC/4hShxA8/Pu8TK/s3xDyhqQur9XsZ7Vth8E7cGy6l6q
unJyKF0x8s2nzY6v+NcKhhY5dluB5kwOppKa/Yl4FiS6L4M6MITNWnuAde9pw+KF
jYQYh3oYd34Shrult5tHVVRUYyCKg1OR5hKgMSZ29XxjZFnm20IpQQvEvezK5mqu
xTZan9r0Oh3pYLxifTlJBWdrZX1Nm8RSlA1til5tIsP0yg1ezcHUVyKLDgTSunLY
3IZwR0SXmsPtsNsL+KDFH8/WS/nLGTysEN2KN9i+PTA9tOhU9F7fWSlmpuCg1ZUZ
TIbWE45Bv4Fr9OH94lAZ583hHs+Vnsjw5BwjPGJGLJN/ATWh3MsOuCglPykaubLh
`protect END_PROTECTED
