`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Pd3EzZ0mn50jE/T+vcDcGCViAXIC0SPgp0aTwyrhV/nkBajzyskcF+OPwfYenaC
D0vl+xEPKz/evoWmZrFl7iN5sjyqHalfwWR6091QY4ST+hpshyB9ve27xu2q7yCJ
MRBUDcsvNQkY0IUbzgNJMdRlKpY/lsPyzBy9B3PdBzL1PINNpxLdnFRG5xtgWigK
+0pOWKHUONt4uB0LTLlXG17r6jrO+GScZ5ohCq0wXuRKD2rQBWH1sMvuI0H9HZmX
YT67yCklhCCcZiizTw7T1s+zrGGFLQ3Ou+wBRzDDd5e6CcPdUtfPyDQ2A+gIVITc
KyevEhMUesm8YeQwUNLSw0Z6YGO9xfMY8dWYcT+f176ygrvZSXWtWusgSZhCiTny
bPdc/gmDftebx58I3oaRiQ==
`protect END_PROTECTED
