`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nhrq/FiRUN+Ex4Voz4tPUS+E1AnbKFwaTzsMMgVkHOm2sM/3v66UosQfU381hBLI
uNAdac2fo+FiVdR9YMyQ1MWmOIwfVq+OD/plckKzmQatcPkj2mVhCNrlwuEs8bVR
O/yER5DN1bI8zNmRp2mQuBacj4AAAlxgSMQ3GSdXoNEoUx0kHcOeiPb3AAl/LBBp
sQ1Le+0Nb6qYMo05QkbLM42ALcG3c/+Sy4v2doj+opNkDMpEw8Ys70BoQbU3qrGL
v6Spkaf1Go321b0LEPvzJu+DrIzdDj5dFKB4f4K8bmdzEUh6wpBC6sio3LglmdDX
MDc4INCeSWTfYGcJO3f/xtQfoBD3Y87RMMXNMgTTI5e1teSTMDrPGGSuF2G1w2Zu
`protect END_PROTECTED
