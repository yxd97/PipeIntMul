`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pxfNmQ+Ei5dJcTWro9X69YsxNlYSUTcFwbIoMZ6FRMvqLgdgBFBzcEJqm8w4R8pp
gVsLMNt5zr0AbUPgh0wFT1d112aXGb0qQ11jXLJp3BeEgjTbtT8fjqwiyGinsUVF
BeXXFQwvRu3Yux02eJrlQC/JKCk1YhxabGoXWqG9Lk24iOHGDuNo9E7bQoOEo7iQ
0F3IQc+XE0vcTuFyHVbhXk8SwYRHcP9upiEk1CEJAFib33Da95BBPPMOGr7PXkkl
QLVs+JPvCtonA2oX6CBhjvBksqLRE/nebnEbrdBkTMWRMtX1jizCPapMGBop7cnr
hjJAfcoTtV4zGse3tLosWMUhxm4numN6IphIAfuCjnNypbQfeTSi0h3qMc8K3mWG
VwK5PZiy3nrgqcmCdHw6vXsQ/HiGtwb0p5c0iY72uBg8za2L4RQ1HL7W+pncSux1
jvtWdQ2MMTEMQndo+bV0gZxp3Qpn4diR5TnVeg0MJPZ5rL/+84ps/SZ5ZUHrO2QM
5gEpZl9IVEelEEdRPR6h7f3lkFt6G76vYkV7jwwQasx2JJlWlvIP6en6PbBr3vqw
jo+qqszIlFHhDZm4aMwAMN26gFj43tGfR5ynZ3kbGk3FgPFhMtKF8Uk2U7mk0S+7
BjcxgLT24ylz9j/CUYHwnXCEA+mMg/1/UvWEfWPb5i2JjkKACO853otlXPTYUw4a
gVsgFF8V+jfCKxINDcqkOR0ENQboy72zxdYysocvDVpMbnsvYEerP8oLyEJKWM2h
AsjdJXqHOQmLwQ7/Y1TO5w==
`protect END_PROTECTED
