`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgQWd1hP3RHwbZrQE57/ie6DZBjTKWUYF87l5JVLdG7xKw7JBPoD7gsyNaivNunC
yx6iVTx7v5chfeJTOuflLd67yUlQ40PDz9pOTPJ+I/w0Atb9+aeNbgxmm632PQNM
E7FeW9EIPDH7gTyUuI12QGqhFEua9UDtfX/smBDA0O5GEC6nObWZmJzq5KZr9DmS
2OMVcuwqJDxbNdcg61oYv/osKsWHtBIivg3Hd+j9e07pcLq0peXh3YLVhm81ShF1
Qih2W1CJ7YlOoMb1t06duA==
`protect END_PROTECTED
