`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0d3CD69IPzUuSfi32rHil9YFdF+X6C65pO751aFECJUZ5VK92BPmCWuX8Jbdvav
pRfzGseNMcuWqvG86gqnMaKDZA8kzZMLJtQZYEowetK7lwtePY1i8dQ4OFubjC2q
ppQJCxx+DjWyBukz3SCSeVNjYEHd0+l2sdwjx1h9wi3/y5sbYdMevGQXSoFqOSgL
iWhCNc/3ZTjj5Iio2CpI71KjLWXy3gUC1JXIDPjIupE6mMeuyox7xLyln7DUa9sS
Ij0RdbkgrC1/fuBA8/S27eJ/N8Pb7QRYIX8SPoA0xKL9ymg3s2iBLa2ikyccoQnS
xTy2VY/SDp8Is+vlTU74rPn/Pim/dmkoYM/D5QN78fjDrAkhmwGu12X155JXWMNL
qTNY/UFJOIS6YzU7gAC7CyM8FNSZfnoGn187hyuXJfE=
`protect END_PROTECTED
