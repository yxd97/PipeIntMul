`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fm7tjaTeMdimpQ+C9OyHLUpxvtsfCtdr4HwtwqdTTxtsAF/3esO6ZWfNsNcuCkFS
NYq63P6RZu0NQ/Vm7O17AjPVSbMupulbF9MsjpCHaliERobFI7n0tMrjtxdJjw+i
q85Tgkg/KdM1T9/5Yvdmrp2jRTLADfxeidJoSBMGNvLZ6xxz702uJ1vPBcZ6s3rL
97/Dbx6WCqA5Br3mRd0K27eIGznKBqg5hQ5cxlMUcPICajA3hYHtVeUKpUKVxdzr
mB54RJHAB41JbN6JfFITgoZR5eE+r8QLARGuz6n8tYXOT98lK0RqGOSCEaKBWoGL
PGn0byOFVWi+zotLFfWQT2KLhWBX1NT01OrDIQYjVwQAKCmQt7C5pWgGv/Reejds
g0MWQ33UnPFCXNFkYczwlaUj74LGHt4SsVe8qvqSbnhQPIQz/Z3/tO1DvGlt+QYR
`protect END_PROTECTED
