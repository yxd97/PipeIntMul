`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7PsvMzrozN/FxqNoYPC9y+zO+VOB+o43YGkpTdyQI9wsWave931iiwbsmOokjB3K
2gkaMVAFjPeNbnRr41pygnUss/3Tb9sKV5x7E2a6XIGXu5swPg1KfGc1oTnTP1T7
tuF+LfkFVfi0VVqlqAi0JohwXrcDBgRbjc96afwL5KWcf+6mDulYirEXFoJQoVGT
t77DFU2opc4w9Gteeu3uVvNXdKYIGval1sqVt+YixQDMkQo6TmuS6C876CvSBGlj
MLnK2iqAHnjVrAyYrIoyGYTeMNKQP6vF3GDOrymWXQTAfugSEug8ZMN+bPS0YXUd
m+kyQCyLVf4j8MjasK5KV9YrQFo3irr+usDHcMSqGWvt4FmJfCvGQel2dCuU3ZDT
1EI1VqE0YnBVT8bj99XX830Rf4IDNKBZgTRDdTMO6yEJzN8+YqJhQN0K1tCCPAvC
Rgi4H/QeT9nLemzziTkXwwmK/sxeDLKjjGhylywcXFyVgHHunVvlXarAhBVPyrPF
Ic21HxpVwm5hJXjQiBz87hn0waJCVJk6QJN4CQIw3TU+2mGNXySW9EvHgcBI3kmX
zVi9ww658gmYjcLKo0Sv6Ju+cDPVQfiS598eOaRXNVleyVZbjurbd4L64E8IzPNo
Km3ilekIbXcC/KFBf/dZzqSEY4zBnF8PALGsWrBS9u8yLgN08Ev3kTtTDuWzBB+p
RLGJCJwl7CNU4e7sig5V60fhVDRWJpRaWN1FzeMeeWXN2hv5wk74YuekertZ1V7D
S7GLfgj02hWNGPEhKSx5NtuwxUFdYDF6tkthablVK/C93PRSRlZJjdu5N0d0+lSc
Fm4Nb1TOp4xiY8C7Hxexs/CZfp+JqeJYzPoX9BogL9WR8AnOLUx0XrUwLf3kbp3L
`protect END_PROTECTED
