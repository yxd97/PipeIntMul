`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZUEExetQCvpx9sCVJ3hrbfopAqrOlZpN7QpgqrxdmU5ykxf7/00mTTHG1SxXNTlt
6z8wg7+eNAxQdJEZxpZW32IsdH69u8rzp6Tv31zlrGP4dMcDW7wv9yJjDc/HRyuF
UZMHb0STDAGWLcjiALXxKgs1fl0dNY+E/YY1ANQ7CotcHldt+b8w6kiPgSvRiu7M
e4lzw4RTaaz0yIBarDl4z8KugTdpcbZScsHQN4UAKFzBnEKdgcmkUnjYOX3tRT3A
b5ze22rwb1HPt0Q1YuB4Yw==
`protect END_PROTECTED
