`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gIEf17BdwEtoyRN/oNJpxDnslf5ySxhszuaxPY6Cj0WG8wOG06HJsgTW2sUaCtDq
/D7mlWwJVVRJ5mDK9svBi6tUAaERbIoD9K20ebwsEkylENXMVN2XSsEuVUqONgzU
+vCjIWdq4kOg8lXfxDuqrfHWSEAZV4nAQSdckYtkULWH/brlTbpwJllJ1TYLFGY2
IJPuEsRWekDkG82jSwQnc91Er3EKb8SGRbSlEgooH6zjTyNXiVE8en+Dso1/M01s
gtgTbduIBhXDtWGuXRSjcHLZAYNnzdMEHI5zgrqWfU0p1v796DUJ+rkfDbu+CsxI
YTlZEoHEQ15G0Boa4f8Vo2DrtpbvW52Bwl//U7YCEYhLVerMLUt0jEdG9txXIjIY
LKvrQpD99+uNROwGbKnIbpBhhVxWZydyFmsax1tEt16oPPFqhgCiipapZTm5/WNU
d1zUJ5Cyd3RFzhie/nabPAyUhP0WSUP5sjd4SOWdqgeCK8c+tfG8izICTya5BXRU
Qeu90gz4OBbieWejI/yUFOeF9SWR0abcHndwRpl4FbYKtaXsjyhKfOMBatApR1ZK
LJewmTtnNkD0Q4mdd83K+5vVDk26HEpzq7D2luKU4+gbOvCHRNGYeiKz7JG7GJ54
zQzn9Z+yYHNmSoACOHA/zcaBPZOWSJ/4WLKjjKivge9eJ+j4y5RX4BRCnuNOqXIZ
k/56kza3G3S+mB/0femHF5BEEs8v7FMo9IltP8si9voh8jB0zxVM/fn/roYiBo4p
1E8l4zaxcX06V8ks/2k381Qu3Ct0Wbh44yFZ/gjdH5EIZrADEYyEpAm74N2EZlJe
C7LjhqEq3zPwOghoFizyLOf/bn+DYW9rscC/PrG94doQq+uwbhoK3+6An8vSzl0W
2cinq3U+iyyMFQOmtvF52MxZq/ovgf6XG3CS83Z9CVl3Oa/MBmJLdEM8mNb06uoP
86rBXT36NRknRhZHyg7SMfzgSU+4nGlJ/1q4pIx/qD55jzlNaBJMoKQPfeNy5zbP
k8c1GrYWDIn6LesB2+Jj08sf105gM6ITnc0+fjp1BZi8RwiINLIR9Y9wqZI05s4D
qPP9eru2XyVlXgEM429sA9nE7vgVFjwBhvWKoPcsTLOcsjilK97bQ0OBVte1zOdQ
3aTOwOrtTab8T3QOmbmlNwKn74+y5E4BitolqYQo4c7H6SRMfVsR0lSF2jveJ/Fr
4pTb9MEZ3wj6GZS/+K7064+qGjIvTh8nuN0D1/7Mc80bB4J6dnDbDO0rSQ0Ql+5g
lAhfgGXcgtpfQJty0z64JqSr95e0nSe66g0Qtga18vygCj/ScOpI9SK77Wp2M+T/
fcFivuQ1EIPgAOXmsUJbxr7bB9K5o8S14MWSNVP4G4w5DJX+RXrgArt3wXj4Uf9t
ETSnyY9lMrtG5lUjw1rmzQIVbioVnnWf8ip0P8PDWVmGZ5eeSLmyD26pw+zhs/hL
l0pEjZpDfEykBwye/IcKXJHAqQtxEUMPlm/lFmNfOy75Dqt96utmDZfOoINOiFhK
1i/Kw0sVPoR/I+F+Ib/l9J9c2E4FfgX5LS5MY6hQ5k8AGv7qqKPtYVD9z1E5A92X
0cvqnfNzbNSZbvxrtxNw90iH2BALYxTxTx1tv2vOHT5A1kfn2n9On29Z4mY9fVNs
QLA68MwKrmI5mdQAY7J2JxByhUgky14jAGdqjXe405pgAHQl+pzAkRlo4HRNvVzH
zUG4lrlIwP+XeDsRZc42owlM9lsxzWEtA9ZOdeDzHM9GlS5DTYjLbbVgCCTP5ubM
Pxo94JtfX6FKTtxYBzOoe/m9k5DP98xCJTeNyMEIi8Zp15HrS4zhwh5MlW+oKw1+
QtctuKZ9QgXA8jBggTdw/rSuXncsZUxn96CzM0i6CHfH7aA9WxiRDR8i68kvMQ3Y
NUCviq6sXTKA2YaLneKqvFvQK3ANCO+dyNBSltOwPOX4XrkQ7W/tp+c07DXFlRw1
78117AZpanammE436dGDVpcOLINWiRleqykaFWioWDnlOgdrEEu4X4ulvxvVrfOk
Bs5PEJA41DuGrjUkWRzOyg+ttbtvsLfqzsa9ysBdvLY4L9bOxvzTqeaApuZxOc8B
Txp0ZE5DrFN1/RfvoMYKvk9/pSa7UPzD6SdjbESsZ5VE1y+uiljwjB9iSB7rVMer
`protect END_PROTECTED
