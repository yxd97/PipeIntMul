`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQMlAohfVEf9izmwuAFTfFj6aWfhWCNiAaSr3ux0TiDhcj5zAYoGiMc9J8RTxN4v
moK0Li41NrW0BQVJ3mNHuyzTs7anhNsSE7o5G26Bfiipbn0xNYG5bkT0CoG7ybwd
ZReEZSuwTtuUdRrRfMxrHf/oNPZrB7D6J6gMKxPLDj6EcE9tGYObd8hDxzmTNs0B
pcueqiLxwy8HzvBVxjj2gci2OhQMoF77Y28oyWXrIjjDZivJYVf7D6XgGa2aB/Hi
ZbFcriU9wX27tNbGdYw1fjImy5iZhB+asHbwkEx/X9xf2U0z8c6SbLxRffW3aSKa
tsU4hZKAHH8cPGFelQUaTpT1iKgiUlbBO/Esc7lPbBZe0E8ayJIMXWaxLLeGKzzi
nPLf1W61MZxbuie+Cx6yDVSgMLak0NLL8O6RzLGjS/yK9HWxzLoKAvzNYjPFR5ou
bOadho1CfW0cHAjum94QYFIayG8DXQ7bV9puRJtzF6w4liscuCox1SAs6pY2xdgz
PkSARB3AtrXsQ6rgAJn+5voQUQzhSRkutyc56DrkdMgv2WOi18SQJTo2QrnV83ks
GxCTWnJAOXeZazF6fGsSuoB+O7JzjOmMKnsYe5bdqUU=
`protect END_PROTECTED
