`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
imMBvRz9VqDtj3Gpe0E9t9Hx9lwlmXxa5On+94sW0J69cJqAdPWb34G1qV6aGzOg
4RSyEbL9X3ntf9LtLgOrC2s3fqiy59r87GzPCnPj2KK2jdkkoZgdONSyMsDgZyTp
DfAHSePnAoc7zkhqhL50grFU2i876bzSTvB6daeRYrQkXZK55j3kc+BwjHgCEOhL
W1DzFZEJQh6xqwVOYxCjzLeVSCPH5BBsYj+sVzw60NxqW3yHmmueBImJeKl+k9Te
0KqP+xq83M5Vb+FATXM4dr93GUnwVszMUdO2UnoaJHnOW9/8ZglKdUt3Ys3OiJof
l7SgEub+pcaB2b8vv+opdCHhCx/6CPUgNuQBV3/kCv6LHChVyb68KEvpl9XZVE0x
cmj/jNFjn0YN0OuTw90ASMqJGw0g+DLtJz+rfb+ZWvrsbM/fVv0uWmkbsyd3W/uq
xi4PhSE3mFGPYDkHVS/SAqk1/DCwCLIrgL6Qi/tYZZI=
`protect END_PROTECTED
