`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R3hcypP4S8aiJjsVrnmOamEZT5Aif1uSijLEqQ6O2tWzTWq5VPuuLZWvKFcTqhpV
yF0ywQO3C/X7+uo2s6WfHeInZivWoYYpyKGVSxsilT9FrBfWd8uVlUvhf+Wm8ynD
N79uRz0i+h9g9uQ65uVz+VbW/olg3v4HpJYuE7x+rEh5GjWcuxFvuGgSLT2rbVNn
vNpAkUbEIjYJc7YXzyAz+/7hJnJ5+WLXjBMBxQb1/HBQkwVJBawFePM6I0MLQ/lq
bd2qHw0rWbsfGnQ0GLHbQfIGFnvadIqB32Ca+yT3QnRayHq9m7sl63sJ9MuVczKA
52SIZMeh9fmy8qNsMDHSbAoAfSmf+12bDSM2ZFFDbIrv6MbaHsVGCw6T/XH8JAEK
LEnbXdOU4mjKSCdPEalf803d8ZVUjVaNFytTQ0ktObzkMwzGu77EN0mU4yihXh3s
oCL0+rvw10LwycMsfh6dnKgKsYv+oPtcSlI/eVKhmrm3ve5BumTPIUAOMZ0wjNWW
Zj2f10YdMQwrZe8qSv8I+9P3mARUqQ/ZZ1/5WJn2p4O+XqG0hK8QByfNW7UJ8Clg
U68YXPB8daVjdrPzaIxZ1GiwnskIsxZFo7NuOxCHYvUV+wYtPvWtQXy9gXYcJeUh
5rWj6xIoSTCRVmrQ97+yalLtTdCcipqUsvJWd1vE2U7Xd9ZsEBDSVvJ+cTfcmgaQ
HNTJJvgJPH2le3WYMhntCQrR2xDleZvg7etjOLLbZDn5CZBbRfmead2IpCNw6N+5
H5yBkbR0N/59Xyv5VNAiNlYNwijnyz3Siak+LR+rwW7uoCbyhvw5q/eEthSOP2Oz
KY9PGSE8/RVhEXaIFirS6RVbqS0rTZ3KrxCNoujnWZRUV2+I0xBkoyhECniCHjZk
CTWRZZawueSvSdbE7MiKfLFWUABkLLeqghX5fax61ohqmqhEi4M4XsC9KGmTF1HO
NOwb1eK9+Me15XeQ6KwzlLfgkIPXqGD7lEvLh8NWTTOl+FMxkPWcXH5lk/NTIENQ
H1M/7dR+U3VMe3i4m3MBRV3pims+0z8m8fJplgLcru+dCv6pJ0m8/eMpVki0HM/x
x9nBrb2UB05RtOF36UEKEyxJ4Pv7GfEOAA8/EJqjK8GRk8dH38jeUQYKa4JMyu42
8QwaspDTiFTjOG4QGFcQ1h9WGqiYnyvsXHcXbKBXDapHP26svWaxEhSUmQHVWeGR
mp3qL1ayb/2BTKltrtfQJqjmQJ8QhF68O9VTpgiZ4pQz3YCqlOkurGH/Sm8KQ73g
EhueSE8MeVH8mq0KXzsPHM2qL3OBGBuc+MVCmq/JLauJL3AiDbAtLFUc3bBwbGMq
O1J07hvtcklAnK3weiuVd5fSnD+wcl+60byt9lMnOMOJ73CpEWela2GlYp+F76Vw
wDdX+AimCma+PW8ycWtmG93jQfiafD+TsIRpWhYVjvIbc1ZLFLQF7OZXp5OT7poE
nUbsflSLYVpZVsW529jRgHnxLcVPPK/zEDxzYV6EzXsF/JTK0zw84kQXjz+RUdQl
Cwv5QUFXmSQ5B6QSjueG7y4HiAZEYSYcaviPpZIxwFvbhDaJc6r/vraGw3wUXZJr
1Z4nwSi5BmfbIANIx82qgMK48+2Sdg8PpWO9K32EPldxbd3wcjVWKWFjRQ98NIP7
tEkRyUE3Q+jpeF6P+y5gbieHzUKqoY0zz1wYGpDcSX6MLoc2Znn7CRwFfDRZkGlc
IWJ4O+ANbqEJSH2Byr1ueETeIW4LlLn2zamMTb5Ah4Me6XXC1LtIeT9cVCwoKrEK
dVAIjkSwaJJ5LOAwzQCTdGvWM0FRmlgy1V0ujr5pfFsaRm82Q5WOcJnHoZKmtz4K
lvFxiQPC2jvrbBu6ywOaHRN2KQUfpRDDj2zzKorMRkjhDp46u0/TbZSCVqa93wmk
3wXwp8liABoyAitVlMl0o+RHiLLkoTzCtnOA54ZkUfvpiOnoREcUg6qDyy9pkqsA
SLkicQw+s/7/Zt7TRhWKesQXpaLLm1u8z6bF36JeAUfuqBmm3vSMLNPpc2C4d+J4
8udKMT0tSujiG90AfuhPe1gAPiBlv3rkwFQOXWSJnL1p8xc32qFMMeEqlYsZ4EEo
YmsPP0sqHc9s2lQXIhNGbUCcYoRHLTKQ7GhQVGs0xHE7jrJ1UftbS+tYyiqdSgs+
5ogpJjd0ebEd2ZN+1JpoQ0u62tQpxBrlL+uIW5xMaftEPVRaSt3iAJFNu4khM0P1
E+ptV51SgC0IDlnqw0DVQQ+PJsePLCL4g80UIHE40eqMuuvXCYzLRn9ZgUar6H0j
8yiw0MwH70b5sC4iZcvOI+BQcOLY0HrdEV5okH5ekR8UjrHd1tKnYTomSLa5uFEw
1xeTBEUE3yWL6n1c9BQ8KObf3H7O5OyzEgqBc3owAF+FsvWMHul5VRvIcS9fIZpe
lxyVWhg8amVWydteO4zcwuL9PCK5WnecLSlK2uUioAQS09aCq/TCRcbutgjsENxk
eUYKN7viHAPb0wRp21475NLusUj5Rjv9TxK4RovRJhfpD5wsTgRW/6iaGN2aDeYA
UWcUrKlIdHQqWtP/SbxmoRzryA/NKIn6FNItyO4KT6i32id5+Yt+I6l/NuD9G8nS
AIWzdjNE7pj1q2lRlTZlYYPRG3mlA92+m7ZAs8BWEOzouVC4ba+T1Kmi9m1zMZyJ
M6FiEZILZ+7LB49ZEHacJ9aeKzf4H0eqC6BlHRdKQ8AOEqAc/9unhjP++JIh4XKZ
+9xjH4SFRP0IxLE6rczeR8e+uoIdL1QCMKMRZWsCH68cXNshdiv/bDzC+7S2e/NN
6mnSn27AzPlrxcqK8qr4l4/jrZg45FONHub3S9q0v7GMxphsGhBd7AgqpgGu6G40
fYgf1ZZj4ocIlk/Q75PqEQRp1RMhFvWZMKFYWxLHM1Y0tPDt0N4hxe8z1tD1JOO7
nMuUXZYcJQeAeuTXM+N5QlOnF6RhVjP33GySA83oCmWtmJuaZvPplXXdAS70EQHW
moYVwt79lzFmbWo4OPlKwlfCv730n0hssyHQdbbpeJkEjZ1Z2bep5PTYE0ULhi4C
JLP3X6A8yeZmDW2kPYa++IIgb87w26B7dgQqhZPqx4ddjLsEF3HeDLEi4o/Ei6Ww
wdS90uo7t1wMH0dABj3sAfYcyvwiceGDbEVmnRgT+QqpBDB7VuCAwxBd07CGDj0Q
HUugeYK4nboGmIoTWUzca16yMWEihXoxGrwCYOC78z72FhBmWXgRC3VHJKGuf3bi
JGOFGh6diXVQgirUxJQCTKFibEBNsP/4qHPDnYGPbjXN7CHjqS9fkHc78UELbcrU
Qu8OXRnFSYRMIA0GxhmtjFrBnEtJYutw5YpmFSJGlg+cLxxBh6Cu0g2qOEwtSKFt
3qvTsCYje4TxfCfr7215nAaEIIpIu3djurc8jof4qWWj9cHRbY3s8zFFGsGYI72J
ZbFil4ktW/OI4dbrXcJZCD3aSSWU+YHjbGR/0r5/YORqW6fL2TCOTuBge4VzUhLf
VuF4YxD5+niCsfGafNLgmdUzxtVnHRozyEch/57fNy2XxHwCx8xW4BBF83vfXqHf
L3h3lGsBzpZvg1Zn9tveExtSI6+DekeT6upScdboN8PbBjrBwBbKjpGwzRetkK/Z
XVRVS6jmympKYTys4ybsFQgsS44XD6J6lZCu9wUiudlvwByXsYOrnH7V2aaeKJj8
oE+A59WQW24bPomhtQTZEUF0dZIYNyc+9T4VatTd1CHphcM1oyGvbQIeSuh7slvU
B5lz8pRIb7Qx/3gLSkmn3Qe/3JlfgVNivTSxKU0jcOG5s9lK5jlLh+IEbmRZBWGD
MswYzEfHw6z0mten3mpc/QNtBxApusSNHQDuOx2yOFf65K52OelKGthKOMcj0UY5
HJhkyW0OUFBbnBteNCWhnEy8cC+xVPcLP5nCTG/x0Rdzg5V+TPVMWbYmRW1Mvp6q
Ql0PSXN/cvrgF4o8idPZFHyB8V6ZVUV+YaCVnyOw91zgPGvn3SODttoEj+C3Djhz
bGfIxpRoYqQv/WlXbnJqK5tu9aE9E+Usrj5fouh9W6uWGph3QvajtnEhvCF9vvIZ
xoNlbv5e3Y2i72UcMWcpTfDOVVgEZTGKCOnyUaQVDt0U7UZI28aSOg19W6cSmjph
psY74b6F606hBhBdF+Yb9YFksc6iRuY5DQX6Bv69XP626XJ23jyFK0MynEf7SQxj
9f/B8FGoQZpDkpFCfLByl3XmzrzKmgeLISRTHOr/b526QTAXCLvxRHp/jULD9kXJ
awZVat2a5nWR54nt3v8/0bWVJLkE2CpFrEAK6b2saZPZAOjDK8ceiWJ5vA80ZR8m
MAah49MBO4kwW0YAtJMBoJKIxvgLMXVZBqFkxlgljDEmNNbM31uB6tMdVfO/6Wzh
RBNaNEkpdoBpSh2RpIo9oNIr2b2gYBV+oCeKI68xGcu5eqepEHlXdXZ8k1OBn+yf
caG/6O1yZ+/M6gJy7GnpGJ09LeIE7rxnrlpxElWKKe8460u2bjtTKCFVxHt7ENsX
UpZYUD5IeD14hHB4/31G0dd2zGNYR2yKVaa7I3m8tMlOso+7viKBxmNjmcRJciw/
fg9Hwb5O5yCfE1M/egUVXc38X2hIUfdvPnANKujRYeu1EN58vQywH5BPx+qG5A9q
HAwLjoaqr7poQMup2yF4kC1Mh8H7e79SNzbzuMTBQxvwGT/LojFW2akoQgTlZZ9c
wvKDTR5bQGGChoyID0S73VaKeT8YdmpvUUD4n2RThFrhu+Jj5u93TJv3fhjILuNr
wrwBzVnmOt56WuI0NGvH3XdC6ufj7E2qmWCVSHbV2oQmd6hV+exJ5o+02peGWCgr
Yat9EwmYklbCnS66fHCHH9OVa+oNM0bw5oQF8fy30wc=
`protect END_PROTECTED
