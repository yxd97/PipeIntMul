`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZmLj72cHLHt2g1SnxP05aHcretgcMh5vsT9JJyvEp1qRsoqCQ+6IIc0MfE5iEsDp
qazQtDzbiRzHOmw+SdrimlV/JlhbXIF7rafX1OXaI/xRsFAkZ9JBnElMllW+DooK
Uq9GZASeMgLDAXw682l3pb4rfUZffKcGKD2yrt2sAs+LOabEKMh6rMBIvaX7SN9T
wn/UqewFGEx7nsolH2gjUN34DIpBjLiLHmLwhwGCBQptD2sgn81gfYdD88VrgKEV
PJhb/4TqmCPQVWiE4s5N99ZWfOzgVi9L5ej481NCvXcrQG/SHV3GlrdVAzocc2SE
t5HEOEfb6S4U7Z/k4/Yl0UX3YN6UUrKqOa32wvh32Zsj4661ea6fSgZeFWN6pOOG
ZvHm9TAP8eXbTqq5yxkTh3Ewy3/ZRg07UAuy1kuyAj+B3iz7RwjyTtXRcjCl4JKm
IGnbw4/yq8RnpnKpwK7ouyaPYeBDva1YLkdVflp+Ju/f0ZehVzkL+qZX/m/1aTCa
`protect END_PROTECTED
