`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vZU4W2M6AO58fyoRDmJmmFgaDxkI5fkH2KrmAuFBSMzOWYthSchlyICRNLQGmNMf
911H5nrB9x6Hm8D6oQH3/VXfTi9DcaR4uYSvo2wD9TAaCoC3Cjh0oi0xK23vElUW
TZr8jzBdKtSoHZ9c1Q+Zn/mJFCsYDFcOjiwspmds3CuIp4JC2DAdeRw3mhJ5RCxp
MfQoGjX9Q2QyMPfSvb9VOFnfw5jqxxCC3tN55THlmV2Zza6ddMM1AXynXPalJf6l
wQIpN5Cjpma/hvOBvPcc4sEw7u2x5AOxX3E0Mp/xSLcmfmybAgYxDciVqlgCl/By
sI+GayyUwxlbxgoaweuiPbTCdGZ//kHnsAARVWJxIKopRzC4zIxnkaqC5GAoswTM
B9BZge/wI9i9E6DMrkI2PC96qWLxAHEQSUQ4qOttm9s1YUipax/BAy7hjeUVGTwD
b+Vbb2GFP8trV34aDWpa+aOY+rds9AEEP1eE7vk+FpKG09isXIirFUSBrlnVnZO4
z1Q0X0h0sfjJ2IQi7+V/F1JymS5KFoaSxh2hnyy/TbI=
`protect END_PROTECTED
