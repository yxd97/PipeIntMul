`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXFdvr9G+uswOaw29IT8T2NOToZMBpHwuUOXwD9LoRlUnzMHBu2pwltDk9838l94
PCmBXTiIPSgLZq/MhRTlkA4yAaFjwRivJSmTkT/mggmwOK0lw0gKWiOAjJt361bH
N2zrJtCkeahfvkrQagc5r5I/C2qMHXVvrTGkfndGivN/oVPnacm+vOz47ymgFgeD
ogXFseGOzyzUHLR7JRgVEI9GRUqTrado05KBPnrs9EG3cpKe49UxiISPg7iBALJ1
u9TMI8RUxZn9ZZHcYVAVrvlv05eEnks8sHJy8/XOn3oQv0HY+cqlEsP5/FZCb1Os
1aUEY68HF5bKDjJOLfQUslu91SK4kSXHCDwLqU1CwIQ+bCG7owrBYQp2kq0doWuP
pnEo3six90r0zWTb+hznvS7fJe+JMBrX7Svx9HudFLEKSW0hLBIOUhwP9sUtwIMx
jDGUtEXWOGtzX5zjxpIZ1bjbRO3K/1EPu9LGkbcEMsumypOZoBymnZJNRkho6tuv
Ft6sPEjui05XW6IpcrUkZxkvplkxr0A8Z3LupF+8VpIIdn/EOoJbE68REhryEf0M
LanXUIgiZnWgyswMhgCeDEe9UVcaxC8MghLC/ObDXdTOo/RAspnRPsO3iUUy9+SK
hydNf9CTzfOOkfFcBGk21S7atXxcqfyEDOZaDCCVX42ucuY9xNjuT3EOA4D8ih83
QbcETRvUXQxGycnM3Egf+ISlydcZbw1rM9lUsfvaKL1fx9T94GxeOvyMEMsJG+Ev
0s3huDXc0kOkwGpeA0lDq0CV6aoSx6Vx5JCCKG2irt9Kyq/aa5J66YJFp6Vbap47
IWYCIKoBhSNDYJs2tscQFioDlwzrpNow3vJJgK+7USren4Ig46mvX4yCgi1CiZUd
bHyBDDBSrdC6ObKi1M0sPD7/2+ns/iTxFwwXa08OTw4yM//naVrzAUiMOVghU2oi
6ZSLMF1AWIr2DXBLefb2gq7q/15U6E0nvFiYasDM/J9EFabn7ihglhDCOkzR0Rru
IsTNEbfWw9vZQta/1dt3tQbf0YpuVAM9GOGdijxwTo/2jnWOd6SI3EqYHZG19fK0
2cuUdWcZso42lHgobw+TJGibWX/JY9rY9g7IozgLfq1vMZyK8WCuIXhukFsXX7z2
SW7MhB2wZKterTRNAomQI70+mdnqeotkn2h1Su/+dclHsp5a63945GEze4AppZ7Q
KlTH/wjBdgH/EMzoNxFqQg==
`protect END_PROTECTED
