`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zv8sm1rwGJjdlXiXJBAZs+SiiwlZlc9en7LLq7YdJsp0RLDU37GGecoMu+o8bBav
xGUmW54qrjWBqyCr6lSQ/7tqWxgX/9TFLv13WpcVkZSxED0+ObT2Q6kC4UEUE0oq
psdQ6vxhlz8DPZ0thR4ZpEGrS5EI/2U2Vpef2Je0hHY8eYG2UOBfP2GSmQ7mcoNm
IqfzYbxURoX4Z1StAJ1Hm00wn/YoR3HwFQdKmDyJMbN6N428AYMmEpI4sKO1hh4U
hrLtYeOeNYb4Q/krcnrcBSesnzX3Tr3+8KDMxMDvWVx8v8UYliXaN+ijPQ7BPN+J
S84HWIaCrPqS4BZHrs7YJg==
`protect END_PROTECTED
