`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLUbLmfe2pzNG42cGwU4dNYUxCfcTpOVxOOMIuz7fdzn9raGmz+ReW9cDOl1VeH5
zXz0tLHVYUXJ/Ky2dqi9JErdRJmlMVuXCFEnn9Mqca9JSZ2v7V34m89oFI7rkYGa
N1NfmqcY/CYQFB+ekSkLtCW1jXbryTbg1UsN/LN2kmMPQHee6/ofH+p7wXqidCSJ
xTztWAjgmOExR1erbB95HL13fR747MM67VqKfjKSVZvDIYkLPiZChWaAY479WpZR
F3AXpDVqlO9SktGWerSnHcaLcgNQ2K0ooOJR/k3EoBbpFAgc5dbjQzfhje4IIE5u
alM/aXuuiqkp1pt1jGFtzGjla5krdE9I2LGENdfHnDx+sDf2lTJmgQMPHh9pnl6i
BiSzaqRR1ivLjwNOMMtrsK9BNtHe8oDQx5zghQXm4yXBAar3tzXa7dyvKaJ6AFaL
jreyMxD3mxxhp7Jn47n4xtxusDtO8s7QV3I2N04qE6NGK4y1/HbVYAIrGnHpQnOd
HE7xE28fntRwkzumQA/1T8zDNpm6q/oY4pen7H9n0zTMeLRCDweCngQFTNL9VYVF
VCfdsE67xEN4szeL4+DHRuUDx0Z0W/OM137Zp+IkQHXMbRwAkavpE9YCYmxeWSKa
CkTRGD3zlYDZeYShLqXn91Jv4ITtPjpcAzLI31XzHuz/8AXH8AXGk7iNE6R9iFJv
BvSVUxeo/8ngN2e411cVUIKWgciYC30TGLOXCz6dCmTCK3JxSX1n06GiWOslDyH3
IfihBMLmfqS2hhuUQ64nQcnSGU7VDUDKXz1WI7W438KBpc6gU0qUctibJQHI7zF+
dSaOByTlHxCT1EQ5+A+llDmHVKAUkgH8Lhrb1A7/6o3ya+EWt0XQLSzrnApOkjis
aImma6CDwIui6NanD0CUZrwXDu1oKXrJZ0THbUGZtnLi6EL8UavJ+YTocI9i14T+
uZYjRu9i8QwpNj+KppTj8LNxqTfygvraVDI8E6j3Husvcf8e2nIUKk+051PhAP3u
n0TtPgQGxpkLLQaHQn6hhT4tgiVeZaInAcLY8kROSi7yCrBCynExpFdJExog062c
YVRkGJTYvY3qPijcWuZxZSCCdPaR164rWaA12NDVqIbNO68eTkSAwIwojumMMOY6
S7xH65q6QAO31zYYFZWvG5HCw4XmbAWO5zoM1VWtVPyPTAA/X1pGOxmYKj52sOd3
QvVbnN4Gp8Vw9oyiDuirKO5VjZxP5PBH51igm41nua44oB+CYbukRHQbxWwIZz4n
b6E9jRaN/rNLngZRhpTe80FoAY8w328ha+TX4ZwP0ro=
`protect END_PROTECTED
