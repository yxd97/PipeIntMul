`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KW8//qA4yaZSmgdXGEMRkIMm9SGTvd9HJUNzLFbOSNQvT/23UmgAuXI9OI1hM7om
qpAe4xCfxs5DDkuE7j6CVIxfMa5k39MHmz9X3/6L964YSQ/qLjt9RN9U5VK0/bZD
H5M3m964/Kfluo4TowDsDXXVHsmPmjweYVQcYZku682GHJrciP/gELWbxAtcJogy
IP60KDsyKWBIZhakCsFmhBticTJg4RRwHcg+64ECCwsv3qAn1CgAmVgn+Ap71/tl
GHFZgZrJk16xP+q5O1wE95AG6JAqZcbhP0wihDqkfz8whG3Gwe27BYRqezYTkIVu
4AEVMp1NIdH3NSvZp5JVyCndf2hfOIEVakbxVeiwngaevla4yDMxs4PAQSanz4al
pcYnOHpdIB+K/igC+J3uHc8ZqDCMvFKSZNs23n8utnYRe70tsK4Yg4hIJG2vEmkA
WvWG5I1DvX7W/hykBCvBbPB6+r2ORgYQqdZKfIgWdynNKE9X5XuRglWi048orltT
/7sWivyvIE+QPmfi8Aaq0zoEwZetAiuBQUzC/0APA30TQHcKEHvepp7WrEpfxHML
`protect END_PROTECTED
