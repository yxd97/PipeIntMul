`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sx9QipssdKcoL2pFyhQ16XXaDeNKIIz6eWD+CmNmss9SVUHK2up9iYopY/PQ19Jf
MHo9TBiuDUlE10+YW0fKH1T9aejSYuOgrR/tf+SZcuIpvy+WwdVEFtOINLWHOmyx
cJqbPRpSKvL+fqfLRI/krqn4LEpHLr3zNuUdxhr/9zx9u/66yfntksDkRjrawO08
TvX7E+bsCjthj6gSd6IcbK6inY4RRFWEil5s5PRL6k7/hLdRDA1iSSqXdOQaWWKI
cGJ9LQs5KBxgXcVV3kzaa9sVEr7/+JBV6pR2pXoXfMzIs7SBIVSF3RMuWrJm4pnc
STuYUsV2z52CII/dX48dxEdYZ31NusjC3/zpGSrFimF/SJUfobrl8UphTS5YCupZ
tRj32HvgsT2S5q+mP3LbScKaFH+q3DxQbKfvdqtVRXs=
`protect END_PROTECTED
