`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+Dohvls3XqY6/CZzX/eGvZx7506tLDrghEVw0MS0qaIo64WWUk241+6fOvqPoBU
RsUSEtAygwki3dyE05GJf8PV/ayjh+jKTtpQBGhGwPrD2sol7iIC4Fap5FJU/l3I
LjPNpprIDN5eInMY/Omp5UlH6wlwgP3IutsGNXodWt+dUQORJQpGpJs4Yy43GcQL
XXtloSzFCNRMDJS3gE/U/9q3uBlB7gAT43bSveCNshrzyVZxP8cHmug4yEeMqZN3
VHicp+9g/2XZjOE0dP64l0d4xDi40640AFTF9eU/9H3soeKEfcPue9Xqi0IkhQ8I
zc3/Oer28nI/8lVSelgDZ9NrXyhop/Wiqh/s9ebIEjFQ7GbXZbW29ET+bsxwXUyH
`protect END_PROTECTED
