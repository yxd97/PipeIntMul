`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQbupKa1XcAqmDcXf75XWrTbgP0+j+aaaIo4O6y2X3/86LcrAeIl22ZmZJXbQ1A2
r7kh1DgmZbY2egbYkpmkHPLzWQzOSY8UIBxl6L7tDAh+Epny05Ppuf7xLZ6Y5Mlq
pgZvLIbF6TSkK0BjZ4vo9BmyhkuuckoUdubNRMwC7qYtYKHok/jBt7M/OLLsF5ii
WpAjSRHE5ZuDlbjmN9lPCAeU5FZm4AwB+vDi1wJlQWUu08MXHZPeAsKR2DE8qDyb
72ZxMuYaoFg5juUMnmlI2Rqq5AhOANughGWDOSCxJ3SR7sJiFRVUVKlcTwQhq7Ah
7LR0jHHjoESgwgM2riwFDQ==
`protect END_PROTECTED
