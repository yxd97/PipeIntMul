`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yS4zDyuV2jv+9MOqAYLf6XXtuO8HIxEy403iONj2fMz6FeyNQT02AMADM9wqV8d6
cS62NRi8gQR9aGycMmfpt/TiwN2ahAjDZN7LHwosVKi9nrRadBQmZtxm12+D6tfd
+jnGc6/CoDF2cue+7eOvyv2YLDF1byRIgx8MpMMys1z8PYcDhRZG8m/uDdpiNWza
B9cLDstTkzM4tebhqOZ6nOrBryCV/5StJXYjVHmv+YdlDNCwN7DTdttlKWtBGTKO
uC8TbQIxK/f80rE/fD29JYgvuJfbYW5oefORrgGPk8Enb43ORx3Vp7BrrPEUFo3n
vGTuhr0bIdFYT12++eRKLBPxX+kkYLyLrC+YqNctk8WfmoVCgenF3PEJs9HvJPng
VUbA47ptwnJRMleyKno3nLWX07DX89bhMFvF9I3oJz4yRPjy2ARIAnYUA/XubVu0
cI/KvPiDkHXlSwAX++/U3PCvLVs3AbagjVsvGnqjYSA=
`protect END_PROTECTED
