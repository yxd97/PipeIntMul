`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FO9OQIABTBIUZ9yRlUJcK1rAapQ8Nuz1BUQGPgkBJdGbpafOYcFY2+uVNeamp4IB
H4kGfH+dTiJuKhTFSaukJK1bR/BX3HN56mKb9SZv0m9V2PAPiuKtBw47C6JzIZwV
xNQaBlr0T34lKWzxI0fZIVILX5m0t8aKPfVUjM43EKnlWxTxfWStm3AEEfLLfDYZ
a41sRrrMayq4O8CFlbMTge0es9N49Apw8uHPbCXiWJzAhXDSvIk6eIplI+fpD5db
xO5YhZQj377qrzkAMtepk/N/YErjJCHqWCD0JX7vMg2Hrn6hCr5m8zMwZmp/1PPb
NCP/5/SIgywP/l8sYHbiskfSrV6tG9m5QEFN0yqD/gS91jl/8zbtmmjj228cHM62
qINb3WBQMSrICvT0Dx8DAbDctNxTGRmBc6xq7lKHo0okqk8/xMvJFsq0FIjIXXwB
PTe6Et+ov/U0pJBR5b6tL+cMJzE8vU+LVO4hssakw6cpHW8+9/eXXLTRZAbQFQ27
KjdhQlgqTshIw17u4X+2VvXbwZyByZEeJjn+3uFdNzGhNfRUN9EJ4wMYDE8q2KBx
aBof+B+fvMw5ch/Kqm1fzXHZdX9m6gPKmPdbQ7K1dvGp8/rNEm/ycK8RStpPaODE
7xdb/DiGnaG36xzUBQs1K7N6TNlXzasg0ZjsJQKlNfU=
`protect END_PROTECTED
