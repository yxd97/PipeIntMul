`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VhDYbiZNdgIy9QzM/DmcFiGK/69m7m25PpCPcJ7L8D/lkhho/yp1Po/i5DuemZWJ
l0Hs93dyN6+crb3QtVF0qXHXHXqgozmLv1kOhSLzgEL17JWN05rlhg6/AK5/aL0Z
IcewTPRXhV73NVDtGi/XY8p4731jsjfi1Ubq3AcZqdzXUYN8j8uP86BFfdsAn3dY
o0w/XQzx4ugVjIcz9V4z8PR+BiWlddw/msMSLxqzci5AUBOEAD5+enmV6MTGuNM0
pYcYsayuX3OgMtwvReIbpdD1uScdAk8afv8y86Jj40MBdpYkLeNgH0UcpF2KMQz5
`protect END_PROTECTED
