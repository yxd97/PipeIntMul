`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9e4OnyfVFcq6rUEWU/Cj48PYfTGf1gSfCTZRMv5XIxq1xqbcE+PWXwIUZxU5JVdj
xzFcjuFP1+tCysW09fn6E1BityIQxIJEkFrPofvvSI/HsRj0ENsIdNHPhkS15Nog
tJHa8re5pn2HWF0bHGo/ChlSwYI1YnLe0CU5IJ8LQfHMwpSFtPJZu5lztaxnNDwV
KkN0r1ZWwelMdNbkSNH9EQHyxXViujpeTS20zydZ0dGPA8apwtpc7I57hh4AIzBY
zwrTTt67S6yxmD5V7bvSlvj48szl5EX+GaC10rt0GmQK9Yczu57S91lhTgXCZgrL
r+Kl3oHW26mOqLwUPGL+N40n9Cs8Jl/j7UetpVKE63YsnjMNMEcuowazCKCbyNuz
S2gfqcvVnRonIjQu9flnzF4zfzzHi2PLQ8dURoBPbX1AdxG0bpjnUPxgHrh0Y9G4
AK1ZdDNxiL99f8FjozzMqQ==
`protect END_PROTECTED
