`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LGopGBVwkQ7LBY9z5hQ6NdTyHPtIq7OizFi43MbnjT+h+v0NkHrnfHPdNFzQMoTM
pMWUA/XTr156hcUKovzJkTepY7lYpRCimU+xxJGZY4f47B1q/7F1j8FhDYrFKygi
af35yj4+snheescWV87h9mo14cZWkL1f0wDJHh6f/TSkc11yqCjlYeXQGPK/dzFe
EFePkJt09gcOOC0StjvqJwiZsh/t7c8iyjPFSiUosprYq37PAiKuCj5LuirC3Psp
fZxtBihUURXMgtdJUD7TC02PgE8Xo/cg6Vm1qrdAa6eRyZ+sbjPQfCyx/AMb1uE6
43LneMRkBu/baMC/SF9L5OJLHlDUdIQN/gSCSlde0Y0=
`protect END_PROTECTED
