`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IicFlwuwMhq0lqIm4C3V/QER33n0cEHgOZ+2HBa9QYTZDRiTVeWYcR+yG7/LMRJ/
DT7t9xZ6WlNCxfPfoJijyG4d29cXQ9lGXOElNhOrKA+GJgtCffexTe1C313yPuF6
DAy7QC9TBAdBb8rGEKhVBs8+LsihnZvCBEJn1Ia+nFkGvp7QlRa0vSd0GMiSOeq9
l3P8Jfi/rJ32wVZFmWDfkvIQh0U5iKtHUuBv5s9xGqUC+LFZPC4bAR1cW3W0cmgj
/0qLSUMFuvLFcRvntnvLP/1ap092cegwvenPedNXMTfMDTMgOhqoBpV7gAgkykNi
jF/NbotInZ51iuCQLz9V1mLiZ0LUEOKmWdn4MR2gnlHaq/uGvC4yF9fJvdiIvN1R
dMLR73ly+52cDZpHSZXmqrqfctLuwXjW20LffvUoc+I=
`protect END_PROTECTED
