`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N8aeKk1IIxRoXWhjbJBrYzoQdUbDrW1POc6v29evwctIrXkLUkumEG4gY0eD2mNq
dw5kOIspATueKvIQPX8qzl8bwMS2CtKSanVfVBk8pgUAuemZBgRQO0BNKVjookvc
nJbR6P1syw5ERLyJ2ntz1koREKksvf2n0W20VMiQ+BzAnaOi21kVwWjfazYZnHZF
yLNtBOOo+K+RsBDm9wUtg+rkpMutn3doY9WgrELl/Gpamg+D4xkmSAi7jdleeoQ0
RyWlovihom1B3SqI3mDHbx5mQz6ruLxpgAywqvAJadVedDP3baF972TSpGVu/X6V
EPDfYOxfdSNZXikkyFXRjG/jEW+d2EEKd8r80fS/RO7EyPd+eDU46pLg1J0JQ2Lm
NDYYcu9DkyiSECqkeWnXcX5cS4zUXtuNuic3JIcVC7j3DzDkQLENxGSFs6mubVv3
`protect END_PROTECTED
