`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rDha28MPpkqQvGFvhBEi/ydU/1GajI8qzq927MB2JNto1LqhUFX3e//bq/AZah58
M0SVgE33XebD9A30PCI8k+l6OKsqIy4uOhgnZkoLxhutHc9zGUwhKrzL8EdGS21V
TMb7uob77IKY2X5HrXthVzhPj1JooP9fzY6sTba/fiZJLpVXU3x33cc81UdpQg2C
ofeWyRS7LAkouGTWUTtX1PS0AfwE0DTtIJCGQItXbux1jz6rtW1NG929Ddj7MnYs
ZUavvunTsMmqsVM+gA58kE+4QJ2Y5g6Flahdbht5/xjrl2GjOQW5tHGm37oZ+Jzi
DpDmZJUOTduSXN6PNWTZCo1qf3uywQSIPr1QQ6E7mQhIVxEf05XLif00cVR44x9B
qyny6rzxvC1VVFY7jW6nYvbk2YL3q8tSjVU0OwbtozmRyTs97kMhG43X1xcoxkF3
hx4MH9Bl8/2Eh64pqPMO2cKp1NxQC1f5lm3DfLIasOpt1mbfLzMZ82OtSzivQpjb
MV7Kc8O5/rw8/6eescu1qZkzSUWoPx5u2NT5uXyLqa57plCU0G36MCjgpQxWJiq3
9U8tqyQrJvcr/6peYmjp9HeeZE+ByP7JEBWG848YXsqd5qeZKLs9hGhExI0aP/0b
OjkI9eB6sfrXF9Byc+cVgEnFHBj3v6PP07W4P7On4NLuiOph96ArYp2h2M6Xook0
I9ph/vUTK0bF9Z/83n2w9dYgObPrXzbpH7RraNyancBSScR5GWkzVcDGoTFhNL1i
plOjnBWsAWkfC+4ZDvh115am5i/8wZ2pSt0/4CNpkEBqA4t6OLRR4meLXWBOCuBj
92gwpN0q+CfNfRlW4ZQJAcy1DXYqYQC6VLn8cjKqzvHHlhNKw++9LAkR8t/N9yxG
B+cQeEEx2f/HnfjguguAzIVh4cu9oK10sq9XYSGJX7IxeEhiyRp59LkbZqoVCN01
oUs3q7KRcGnJBcEoG3Eqe17BKblFIFw1LHuUrCPxitfyENrYSVfPVmRVPvLbpiOk
bzMn5hmp7f1vRTjzIbFvRdxCcEAK70Q1CiPUGiznza8gnU7CcG7gqAwcgbMyhE0G
Wv+quu4i2vg5CaPamMVrtqaWFnkcLCHRXquAAVAOC/U+QZq8956r0xsdwbDG8m6/
D7aEhvUd25lop1SkVWLT+T05xarbW0CxzCHbrRkN6p8nARHFFQvOvLK9QZrWTLJV
hl5w3PJCavhVDT+5okC+Soo/LvgXOuc0BB2GLoBvDlGRaAUvaXDzeHJDQxEMSOS3
h5TAMNAjfzLDGafkEu4PRM2lExIIvZw4LDnTg4va7RJ01eRVfz5Ar6eGa2jmK4WB
nW/e3nyBdWmwL+vJf86wqwBMBxEMtik+aBnFTf0i6eU9lhK00UrvrFQiPCt5dSXs
C+MxiYStLNu9C5fM2MB69FCggUw0uVgUGfYxtK/Eeikz4QhErTduwySyqY5lug/p
grAHc8bffH8e5njeZ04WTW+qzBL0i1xU+tC9c2eWbd5Qiv1zxEsPABNb4PZvv1Qh
`protect END_PROTECTED
