`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ish5Hg7xWPdwPcf8zEjXyKvreB5z0C4WA00gywsA8RfdwCxUhCZdTy+zCOF27XYS
bgf50dBTD6bR2px4H/VoPTKiXXMTWqy3CS0fKUm+O2M7fixG3T/VQGL/fYPbPKQ/
VB7NruRM1AITYJmjHj5IWv0Y8JkRmJsob5l/QsaDSNFr3gwPBR5vCOEoAok9i4Mt
hx2vpeMT+pWOOvSu4l8hEKcDNGTJN9HphPAvorpy5droNdRrToZSQEhaEg0iYSW0
5lttD4Aa0BUf/OTlzBjW23TVsO+w9zaUbxDN7i+G6JJM2D/AEDC2NQ+3FvLwBgCk
BeuxDB1t/1ydWTcIMQB5mSlx1H03maQ0ekaklwyCXeBdjJs2bomFNbQrdBy6iATr
EtzbmDebaT2PIQrLjCwygNFs8AK+ok86oRXPZOVrrD5ai/wKz58iswoSVf1RNVXo
WpgxL7zYruDZbS4pORxIP+7RI7T+eJzBXZa9fH3MkagQTW0UBqYOmG8TOkPRmaGp
`protect END_PROTECTED
