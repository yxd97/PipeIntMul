`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LXcfCm8wYcQp2ImbhvPZUgm82BijISUmVCfsDxo9yW2RU4TC5YeXQ64h/e8YhALY
x+kVf8qzpWgoqLtJRo/nx4C95GiBprxRckf/cXDUhMzINgcDBprmGUyPeH4rqShU
yT4x0a1D96z98ZmwXuKkXh4xoOXR3RtlkJRz8pWmVHrlXFR4Eb5JulOQdNAB1JlL
9rFYc+i8z0bcw+kB/Lb0eH8c+rwKgWAI+1R9fWQkn4SO5VWEw4z7mTkeN8WtGqiV
8pkT/XRD+5Z933Wvf/FM+w==
`protect END_PROTECTED
