`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zH/RJ5GtO87eDU0YdmDYmxm7p215+PA3dY1SjoRD0mbTMPgKejaK3VUOhNwKR4Bg
A3XvpnbdKTBoTRDNuyDmnG5+BLqgmQjVWYBY1TyRbaDJobxzsro81v1mb8OnlPZ4
0kUjhaPQSaBE+iTcMfKUWrOCiclFdwwKcyJXklfeMYyqrNQDP/D/GCzdfAlG1407
Cpsn3C9oNkkRr/mkwGh49iScKrCEy6/clGwMYVdhIYCw/zBgD26ybrnjDXfr0mcA
`protect END_PROTECTED
