`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jeSw1jJFSGHOhCoRYWxiEipIScpncXWlAGICkvUvU1GE/5ipRtVfAJXbu0v67bqC
qSlPaV8EHsb4bwPcZP8Wtp64WT+kG9zZkohFVGUfMwpEwvjjeEEH9s0roVo18ggn
OXRP9RflwGahRbEYNTMkYanvvIkz/E4X5Iiw/NXlGbnVnHQtxd024RydB+30+mFs
jBZRD/0MS9E0oOIMqf3U/POZS9wnJ1pDmPCCRBVp4ND+OjYcI9Edkku+7cg1WUeF
g+QNRMXJru2yMo6GI4OiqYbyRMb2GHKdTRMMTnmNQIALXlkUCYhdno2xynM4rLv5
Yg2BEV/0o6leZ5H2+yAzLA==
`protect END_PROTECTED
