`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JW3paciDUSW+uFPaqwhgtbCdlubb5euykPWnsr7llW1r0O7IKYLwaZRWH7Do1i/Z
m3kIZLxozcS688FmK7D2Ib5i2xvHuvlohUe7ibmkXENKVhCpJzzyxFVE+HcHmnba
qnpFTiG44zOse+dMzpO+UHZzkG4+dycCI7NmdMN/Y9buoNcP7FfHYse5M7dlL88i
LFqXYZnI5stL4/+mpG2AX9x2RKAojvkt+mjZP1kElWU6lZQ6h+gb4nLth57Sk/kr
MFjNY7E1+8E/6WWz180ELvyP+GvLvh6OdwfBj6HGYtovj0/OQCamgPt6orx1xIjm
17E83WafAaYnen1nXfhpCHYR7aEzxkIQjaDBvjaWRMgE49vleCYqKk/SBtuhV3NG
Yu+6bGFNWumhn+irw6XV5xvrzPrmuX3H/qvOwR4RVjqDT0O9PrnEYOpdVyt1rwEC
q/1eMT1C4RwcnI6V9Nu0HxP4DKcDbQP3kMB+RXGXAkTxWM//GzEUwqJ+8hM1IMMe
RzlgoW20h+hzwiprdZ+Pc/gTeQeF27BlJ2/KGemBoZe2Jwgh0+UZ40lGPRWC3Nx7
pivRXTuVrAtsRpsk6nT8k4h/P7RnBY7lB8KoXrfe/p7584yb9efXomUJrtYs9x23
540w8uW4OheAHGvJG63D8+DkI/ApZ7FPitFSx5ABDZl/G1/mxZuce1WwgHbCRq1b
3teAC4qRgO4DKIbRJo0SJiuriu0ChWB17d39sQmTDMnwdFMl7VD655uesSkDFfU6
3HSeRUfu2o2m1Ef0bkGBYoveYiaO0BrZ5uDI9jYZPrS4t6LBageu7tJX8RtqrwbG
Hm+8AAbVhNqxG3qI4QOqNfnHjH5MD5azpqLRGV4XYlRodbmTYE3xxQevo5wKKkF6
euNdxwerp21hCFKNBTdsLIhTOkyQRfl8/1hITlR3s6VPoBPSvxhoPAuY2Q7TDr6+
NoM8fSVb2pDcoQBaDii7VaoSNxP22iaooMS2bxjVU36nBXiXRBkfOcVRgO1I8uq/
FUonJkmOnUxUOj0OOAU7Z7ePzgnszpf8Cb+KOkjnwZvFMkpVY+QxWANik2l3HbPs
jBHGT+bs51wDXLQXHEIkNI8ijTkMY6F6/pEQ8oWhjLWYQeWvtwc/Z5KMCz62aMmc
v0HQWWUcr16LV5qx/NyjyFc/16/tDPZo7LLzX1k5HRUgaE6Mm9giIZKgPM/8ZQfE
52i4yQ2FkFS77AenttRW5yKD5O21rF24W7ZBuNyxzVa//Bn1z3vst6Z8etL7YniE
PeLMHfyzWaGAW4B4X9eGFneZ23tO+i2Nn8pwd/GpuDxW4boU8sw+pTN3AB3FNKZ8
JNLIXcdZri6jHD/qf40k2MTqy3/5rZvsPW9TFALtrEz+j65yTu4Drv/JtfrN5fzq
tKY9a97cPfFZbwkwytsUJKCtznjw0lwnVPvr8NYplnBYqRNJLngdt25Q+mybrgep
irQqR5CAw9m9gvL7FwIuNjHwFhZWJojzvcWXK3lmNQvXGnznmLaa+ZdVl26cYmZ9
M3KORtUD+1aca6ZMxfTgjZ5dQk7do6dCJiTda1I1qWejpsEvXG0ZVV9fiPexShik
x95Kv6eA11zJxN9iIpNtT6Dm+1pVMqwfsmfxy7GZs7J0vPo8cRHil6zLeIt3hRY4
lur8JXcXjodhFlFkwqcoQoN63V8xc7IrCPzg+YDXR5FFUZBkqPIiSm6TmHSWFDzm
dNm+I8G6DRFzId4z9GBp5zKtMqp5V0Z8ZbVXkJRu3mfWnydq//knT5G9IerZ9Pum
4Vat3HXByVcmieC+CDffYP3a6J8ttIpCfQUd1iOif7TErhXW1sbN4hMyAt6H0wd0
xzh385uqfJX3N9T9OZ1F6u/hQb1m2qdGx8bFReXKEmLz2qzLxCt93s+e+UctULRq
XT5yVS2MPXylQomSaG9+Cvbr7eTWnFQcyqIGCgHIVmADPwyQKy/Y5/YiV2nN5Kas
LQslgPnY+jLYsIDZstS+D6ciqBqtL4vJgzZ9ychaQozAyQTcJ2abjXcesgSBAOcH
r8nn6Wwh1PRIBG+PfF6dMo5eUrQbmOEdnsRMsF/x91mVqaLuaF7CToHQIe8QLs4v
W2qfAuO9PttXynkLIP8FjhAmFXB4XQl9VbjtsXVbCjyvCHUyKtWKOsG8+5FIPhUJ
WK/VmolAkIyZOaLA4Mi3ekwg5XDdIIfh/M7TnHj4LhY=
`protect END_PROTECTED
