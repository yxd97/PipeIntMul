`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0RDgzDHjXPhSgLd2FrUcUnQ/iwKkNRbV5N/UYGNuQeMYGVNMN2iBqR8q086E+Xw1
2jTZJqDHe+rqzP1fbXLA5zLOONTh1nAGnN19zMlVGB3+6Rz/FHApV56nkhNihw1n
5hGkIAVzqmdgVR6hM5s+qoiRJJBg9BrVwBjU460kc/i8c+c1FOeLofXjsj2p/GyD
lTIfYGoMKyQfQFAMfJjPRB8WDUnYCOE4RaHA1MjrPOxSYM6GwFSHrYyREQFGxbFX
7MGaPfPORr99cpD0DNezQ6bfyMmAyS6x/CytT4OsqnZukm5jjoA54dcpGdbWiwbD
`protect END_PROTECTED
