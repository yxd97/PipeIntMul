`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
loeJBWv2kAufYOG6g3bIzPNW+gg1LZbXKjFosiz9MrGsaCOUkZe89sp5pQxptW6n
ThKPZ/1ape71jEQyr9asn+4zISxNQfjedVuh/dE2sb8gdAiVU4H+gVoVZ033nQ7E
N72tdT4Yg4wnga7DO0mzw2AbZDcgXAnhM7oiEcE2ZmYgecqgD1ZXxR50jTW19B6O
sd/iD+ZgYNl5UJDHZnfuD2mTEn25gtp6RnPx1Jn8qKLO4pJod5dCIFtRfhDm+KsR
H6kHDx/0cOaE1hqlEJMuIpPSnq5T8t7+g6HqGPxUYLdd4/Mj50ZWC2ZtZAaUX8z+
NovcpElMEtEzSoyWZ5AgcT9ZLcjDlR4AX48AORQB7EpBBDjGLIIVxO5Ouya5SKXD
Vn58c2sSWIbL25FmX3oowKBdrFGRQ5d3Z4CNLe416sy1OXcP/8wpH3/XaNNbi7dY
jlYC9/vKjmHJpE973XiP2Agw09fV2yiYXP5EFFRmTva7YVxoU531HJMoHrLo4tgm
SGHqt553ax78U6Tb/V/VVnZ3E4Smq1/EoEaHX8/xuCpUOmJKCIdRiP5WCnXf6bwR
wWp1z6NKuB3GE2EaPsxrlgklPciIEIcyynoRzH4tYFfjPsogX0jYrygTDzYxLCEh
zBpaVnh6GM1+r44hvlE3rUTLHPaja+oPrVFEMa29XclXAKAELQrPtRuamG0TB0ja
gXvrFLDXdqRXl9izJ2hAVljfeNGXVh5fkbNd5BprLle4Mnm2OHLii7PhbfLngo9s
Jl7C5ZIgv4NW1pkN906skpxPoEeAQ8PLxLpmzIMXDbyrNITtB68k9eg9B0wlfZ2M
`protect END_PROTECTED
