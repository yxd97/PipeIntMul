`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Go/H/Vs0O+gNTfkUivfku2lRHmHB1QKmlU9tOSriUhaxMkoGrNEcx1Kty+INXHXT
suUIzf/1wfYFlWIvqpwaT8KERvp6IJ6FJC5Tg21LrKjykgrOlPWcvqveOdlsfu9P
i+yBdJpLTPRMT1b7xqeQ+gsd1GQ2M/8WZRDPGALkOe7Za8zs0PWRx+AjlttZ/0Y4
mg/n2LtaeVFrfGsoiHVhGd8HVD8lMdd0uHY2tOEt69rDHU19JQjiGaqj2Cwii76z
fg30Oj+dFznF8cb7JJSOwW9QspRzAB16VVZIXcynxJYfvnF2pDyKdPBqbKwx56lM
055WUdIqbyJ+e5vYqJ0u2Q0x3ebnH+HJnXn2oVhkUvaMCB3ennh7475q2T0eUI7Y
zrpS2Oy+5S/H9LegHmAUocB5nmDc1++BC/V2mY1GfDNdV4QKuASG99eCCudi0zcv
Aw/70wHmip6cuDuiTU2rBkTEAxG+67y5Of/73ihOGPdQhGETXN99ULWIBpJSbcYM
+csRdHqksnCoLYfhgH/BPPWz5xSZfvOgLs1dAaV8h9J9Ch7mBaYAaEGuH5shgNbt
X42AsJ2XEh1zQjycasdXgiE2Uk/ntuw2ksSQPVhyrlUeOAGSj7GgdoloTesSAdbU
KBpVHq+JUr7plZ4KeyOJsg5ifKLv2ylzWMI/IRWqD8dtHGPgDhxqeOCOfFg55/UV
V5elIlc/DEUkEEISOGKAOvs1s8pF1gLHsZGH6UZDu2q+eNfrt0FIGdSlRE92VlQ0
VGFfJTKt6UX+GYs/5fPwguP2WLSX82vLWEQkdJmjs+6cXEfK0XFhyOvolKjxrd9E
4tFATePfhnu5Xa54ntgIrEmeEmS7Gki8CE/XxDRfLlZATBGjEO2mYUwWspH3NJz1
Ag91iBLU+3SbOar0019FzOjyRqkrQoRG9OcJaFF6UN4Ai01HaQugQZpX40VULoyj
4bRihIPWbeD+lzqje4okAmZVeeX+13oLDsOlMuV255hINc7qureTljs8rQjlnrKx
PvoX90xb0Bm90EYgbFFgJ557FKEzEKdkrM3U83fg5DPLrJZHk9Ftp8b7is2xSb0b
zioZkDhzfMHDE08p+t2rKSmRcfeHa807loUvHtSkFqgkKzNGGbZj9totxA1GZuC5
rwI8ZuXsxNvEH0hpcvEGE7WpZPPREaEn61aFy+U5Rpf7kQ5cDerSGE98pgS3qjdw
WxYlFSo72gO2TM13Ac1Qf5s/tO6SkK20enkbEKUGWYNNZhQ7/YsUiaIZG0bhrWzu
XkbQ2mA9ugrL/3wvFfwksLaj0bUrGrUrQIcUQ8DZvngMSvo+9kLWKpWaUkOEfOhz
mCTj5NX42CYKor5EqKaYWsDRJzTrguv31W7Lq7zkIXSZ4tY9/CQy3JIJUxihch53
BaZYCW1mjE4q6Yrc1oNBmVpR6ZIiBdwVgOl1pyiEgYnFsDPUzJagNE/SMDyNGHev
9+tMNpwvCbTns+lXGWnCj7ITjaq/0lawcnzzVo57+h/IRwkKTW7eziyCjhClMDwq
N4dofPb7w4YbCT+1jEnpOHYH0l8ViujNPGwtPIVjlipWYpo4Sp5hrVRScjdVgNyh
J75RwF6KrrN5LlLVGZxuxpP3FM4xhjxvR3CNjVR8qrfnCTs5T8TCfSRW3iCLhHIW
LBCrYkZxwcskLcKeFm9o2sQvPT5eKwSsn0Dp/4QlB5Nx7HZyHXdxGBAwxgeeOWMo
X48TwzhOwMOkKuERTFInplmUS48NJqsCqCRwCtFIuOBO6sMybSKFROE0ajUh1Afu
SsudJk7JelgoHy8nsUyXH8X1/44UXM29hFIOBOwJyqOchRK+ry0BWP2gjg8dtdT4
u6kYgFTjud7gwvtO07SpB3YkXuJeCk4XATIfy6tNhBN1M/pivM0lkv3vDOHUPDW5
ASrswBneR1vDy4AZkIq3oUTplJefp5UrKLLWLeno6BxoE2AD50KXHoQx4lsBbIto
K/V6gLWehMXGoO5uMLLZ2ISr38+ByetedZCtVbxdoLN0ubTVsSQeMq8jxvowalGD
G9I4a/VX5M9EwTP0fdOLVTg9AoLTq6JqIclvnFgWWI034FFEua4lWeYs/lfIUyMo
3b3kZBg8aPFFPP7magQ8eZwBuuT1RFzx0x5TGp1DSGtTrZTeIaZkBcXFhyZuhFyR
GCqiYc2c/sPynSWRt+yRk9NG5LN7H8+JgFvUgbJQO/WEHH0a3DkNrA5mqXcKaT45
+lBr/xKy8qoWoYqjVWOS9nmeDCrXOBflbv+aWYP713+MbERU9UMJ09zMffvJ4zcD
EMtndp5j8IBoBllro+JZ6wF158Z8FeU1WpkSyhYFHgQc3ChbsD7fgKGW6tB8y5gi
SZopsqqvr6IQLRNjlcaO7kJaxtqWQHnzxJWlaXy387VGuRyPiWSjoaku1YnNabnB
DxN6BxYXkaERYuBEyvP0C/HRFQQf9H1VHpP9SI2hSpS7UocylJRkS6zsXwa6uPIh
K8y2z/CK+hWT1vHyjn3MC1rtk7YmWK31Uc2T7Kr1iI1MYyMNQL6iRVmoKRjjXcKM
qDbY5Z8Rq1Ef5sVLvWEVyVU6dL7a28ypj4lxj044RmGvReecKaX6PN5IHUBSkH5v
7bcOyujS+gUg+ozjpIRnjCVuGPHsK+SL7MqfltTBnFmCaFiSxvNj9o4eP3EUlr0I
3y45RCaP2Gg3KcAwnAjWe/+NDdIyVFo3X0jGkcUxDEN+hEnF41BfrjLRd29N2102
gu8ozCDaj0enFBykAiIRPrQEJeODLhi7fQBYYaWdE6wV/02uUXAzLSpZ0xrfCRJJ
znZvOuPH0Pg87UEsov47arvc+D+01zh2PxGvO6Umd0SfSjh23T3oSghmGzfvj4aF
5t4lEtSkfqWXQhVZpwmdyOLMe70HtrG07eJLlzo+NWlRVaLQw8VQtkca2GfHRj7P
rmKqEB5jRvcqcgu62ilrWH7u6XPxfOnqaoFZS8fFeZ+uLHXgH7/joIeuCDxlNisw
aPtx4hztfWhC/ch/vczFIvQ/WcJH8RseBuwpWz+lmwRroxJ3Uxkusn/4D2qSM0Vq
MH1UzCJAGTrv/nvh96Bl1iOHt33cWxkh6GAhjh+IaDpZcEP1miePSSPDn6+gJXBr
xUWduphpTE4Vs/L5uDy4YeBGzqW/EYcPbapmfAUaw3Z1WWW1sYshldaHZ3jAiYKI
u25z/m6WRQ1oeRH+yFWlyLEDaqADZMlc+g4nmNlj8ietzLwwR60KbAWN3+C/Cyl3
eGMqHwqJz7PVuq80xRznnBHT5dNmYKGofi35u3JiaIY5DzfBDDuC0P1+SDefXCtt
J7biHL6jq4u8OrsX0Q+mXnw9lTxrJP9jkl/E+htrTfZSEn5093tdGsO1rL9idHOM
/r2MPbYMgQvsNPJk8YYBklirD7dpuU5EBAkrOUIcp45G9NdHZxi8oJp+MrjlVUE0
IkEkaDdABsVhHTN8Sghx8jKo9jguZROL+kueq4MbsvFmGZZB8MpQ0960NvVrak+h
v8LzXebq0vsUA3JC5jarzTQ9Mfp0svNff8YlV/pk4IO/Ybq7GONvhmxZY+447qAS
zGYa75ytFUahTLFoVG+lC3Q4vcOYZUljpNBL19shoN9IJBhJ6Jl+vGeb5SE8NUh/
XPVQXNLM3ztRr4eMl1w2E6x4HBxhIyDjsIgpvjuSYKDXpcXysHkqdnG6aJa8yNuc
AMVvjkn3vF36UHwqAD1V07wD52zojabsM3gvBOyIgb0LuLfqqAUZIWTqh4IYUdDv
3XTaSACZZZyOvMz1HKLyNjQ2qhFIEfwdW8/dCOs0QS0blo8H8CraDCrCISCzLvNh
ly19mwmFQc2MZ4onkzPmre8A3JbJHF2PCnJdEjcwG3eRWn+5qD/IxjNVxZAJZyK4
Chw8EtyJlntD34mNaTvJci0HMJ4LhaavFyMxVZazbusun3Gb5wi7OcyyZ7ZO1Stv
orpG/YmDH8b2XizDxJTg3A2Jw3CoYkG+hihGDazNkbyHc/dZnAnmnRMYVvXP8mFf
jyI0SW1qLkc20oqA+t34LLFUAz3PcjRMCAMMDiDyWg3nSavmDMIbwbvU0zVbLCbj
EYpAlgM47wgf1BMwgihkZwFtw1tHTvXL4em3R6EDoml7NYBJuoNV+kpN2HTS/+d7
1mvsCrJrtiJJydQ/nXb+WzkiSqUTiFPFD1JsPpHldahTCaupzEMfYzFD9PIMXvNg
KqNrBICfppKT3r8yFm1vXaSfygkO7AEyJxSehIPEKBRCrOQSZSL5P1Se4StNdHcT
1dr2boC7sGTLkcUAw02h2o0BcTfDIcuPtazF+ftyEucTuOavbmj3aGaUrlcyFtKk
qURyl/8S3SQTVnawYpdRiJcjscL9tikyXIHlGdaq6Pb96enLzifDksA2qilVF7dy
9E1w19P3QCmD0nhE8BmgR2hWrSQKiIyWYg4SRTMD8UHSOp1MMzTG/3857pbdTjl3
OmH05PAF4TLrIVJUlLIPl7VeyYaoufHH+wS318cTW5GxUKoR52dzZTMRcT202svs
wSSPqBidvQW77Wh5aADLNISnSsS4zSGKS3Zy/eKkskz/dDHGaM/ZfNWGGTrV7544
9CcQySDx37xztphogEgSYpJ4ARP7W5ZKuQ4o4XJBWhqdOTOgI9qxxBT4u+6yPGap
MuOVH0gLl0gnD44TPt/UvKZWzSoQjFnETrVYviVLvGZt73BwfqvfIzxVEaAh/Uez
363KI+fOfYoXa5oNOZC2uCg/ApW7n4c6oY6godiD0OPbCSecVQFvNQ98/320DVZ8
bFy56rh8ygHefcpfD+FMKFumnuHb1ZSuogehtxoWVBNhQsDy3jL/clcDxZx56042
TdM+9LObhXWn+GXaSGJsrqdT8MfH1SnlJQxq8vuu3KR3bGFhMjHt2dzTUtPVcq+7
AChCwhv4QqB4xf+DkiX4R85f08ZtevvM7iXLHxD2AsxnG3DniJPCwN9C4jL2Wean
F1mA7q8o3V01BPUaOT+OEaVFNXfSOHbCPFoe4W1OJaB2vgfc5N8Mh6ajH0jFxPJS
whSbgikF6T8nnFM5TH31BcyZJK6FbSLt4HdeP6oIRHtvsqVUsSct9vqp+7ZDAh2B
2e6Qnb8C/mSw420kLxHvLKMQXJnRVFDam9K9NP56baaNFEZxV9R4tFpKam7N9jKN
pWQ19QrsOq7W6rhRI9dWl9M/W+/t/EzFmGuml4Tvoz8KY4KDp1NHTuoR72MMs6BT
KbdhceQFcq74Zfe84cD0aPu48E9Zc1dGweu6SN6bGsg9+Sd12secF3/W90ivq2eu
xNpJUCdenihhCG2i2qKzeZzinD4Ku6eWEdWmLY5GskIOHb8bqJOxW6hqLBQYSZVf
lqLjWG1S5H2teLEKbpvRCVcQN5NOI6KUUrZPOZcd3nvg3O+j0NnQWfeJhoKS0bYU
g58H5jDSOk4F38vOzsgHo4sn/oq+B9IH5i6eAEW/Lq2RXXMSoON99a5mT+uuINJk
D47jJkCapFm/ciRWp59n7qL2n5DlUqPHAuR7cmhH0cFK+3mpE/8XL64JIi4pMpiC
j8e4HQdck+je6gd4XprpP+Vp5lOdQCycb73a5OgqKYo0P5gnv1jDAxPemWEMKKW+
kSgQaxCcAA4ovYNU3Fi4+EtzQxUyxiDTld193FjilrBiUrFt2HF/RiL3TZVce2NS
xChgP7f8uhjvYN/nb/oLdL7jAtNPSFdsVLOa5QpCQEveeMzY+qjD8o2oLeLZYq61
rhrZ3l1heWCIMOGct7FkFnNhXWbiGxjgq+mXlp0u5v+6O1wkzO31OSAnVD3QbAWH
LA5BMoT1sXdeNqKLgynbCDVXqU5Xe620yMM8Ep33ZHz4zzDNT0aVh3PKTrQPiTdO
ibcmPUA7dTpS3acw7u/RVjvcTVsla1+K5esn4Kly5eqfVAo3oB4k+l52cHUTiccS
odYbzEUpZ/NLRGcw+lyjuvOJ7YiQVJzunZ/lMGXQTdWAR+AD0fN67+fpWraCEWxZ
IBipUO7RW6ol3PAc5DaA/c/iIo37VAiY9+yfNKdFu796rkc9EIJsOvn1VcXkImPY
rs625NgVMNGjWtOBWyMBek/F6epJrupLFLhkvDDEbKH5eWJYMWn4DyMOOEexZN7l
y02gZnbKfvAj70/6ahhzZHZW9xsrwUnX5AFife9aQor7x4SUgiitrS7tLvI3RTVN
g2cu5w9ZSAdE7C1ARlzYN6umi1Oc7mvVDR7ipTKShsLpyK1CkRlddkbQo7pPKDL7
nr0KUpxiqQmjTwE3wYSUKNpv/GBPiBqzqDaMc5QmNDwbQt4W1WB9p/O7idlicdoM
V+XvzY375AQ6pEIRdJa+IY/8VvDdk9id2SbzHqUQCFP0etuqVH1TtloOYInjnOSi
/xmVIkeC2XBsXvqHo6cM+xtsEl7X3k8my3lK0dT4BSRM2ZxXgi4zlfJHcsn+eG+m
fqyAQobn5UjM2e8x+QZLw8HZEPnS4lGMYqfU1FFh6xij0hbtURPhAuczYc0o2ZDT
6tE9g5fUHSSRa09HmCwKTZN7gOYNrc00foS4cu0t2Aq9M9o5/LaYSCIOyDhz4Ep6
8cBBMwmmhiIUR3fhbIMn1+/skjIgsTr0l0WkTu4GuLpcy4keO8i2a3ftVmzZdKcE
j+DNgOu/YJJ9V1NdagplaU69yOHJZSLXbEaEluznYf6RYebUTq8HQVNxB1No0U18
o4OyrNsTzcXbnhSybSdZblKyRoDnhRVSg7kv9GJXC4UDlqLEY0rb0UZsjdaocqYf
jS1oeqGlYjeRxgdaFiovieznTYSoPOu5933YihUyWlfEL2Y+Ym5/H2baRAOD1n9U
qFlcA4Ef6Gf6V+YJsjfoX7pDU+TmUCxRKDAE6UCclYnZBStacbO+UdIkDcRqogpW
DvVanaBLrYQ2MAruACXhg3pLi2tnqVtZXHo8LxtzyncokehrimyxVqzJpJ8LXv6S
QmaXOqemIr4Ruy4kYPfJgNB2c+iRZDibXIsH1oY2+OpMGMr961LQOZVqBTO6DcXu
AckghGUPI6rux4g+e+AtnOPskGqxUmVeutfDJzFf92etx/FJ4YRwKkSHHXirWx5C
ub+39zMlrbXARJ98peDW4hDGfvRCsBvfWTKIJTSSuNPXnnk3dJ/xSHrHG1yGe+Ik
MmUGvxP8XspjeVeV9J4pbH0LdRbR0PpFrluiy/LvW4hJUv86eGaW7eR9gBcAem3n
kj8wfwENd8wIX8zBTUsSF4Zk3P7jjNlQynfXA/dR3q1I7SnfSJbRpYa0clk6OM3b
dAWNluUquSICev23ujN8IlDPcAImQKPmK2xBUttH+0fhAxDxTsiq+r+Gmki1znMr
+1hCkX/kfLZ3u1kOMjQh4pf6Hs46OdgGmuQNIo7kRWH6IZdq50gTpNVmHGSCSLdZ
AF9WVbGUSflMUjEOFYNCs0dwlBN231fGMkygrObsMLmoaepTTGBCb7j8CaI57bt4
gGV+DD9Gtvf6fdEn1EhGpOa5wbKauBBwgFn213Gy5sCjA7MTOoTotNB4QQaeXrmJ
ec9MnvKRMwRytZ6evCmJLeskO6661mdoAhKfmGjuHzJuaafhjYEaX6vDfOld2A6z
yfa23N2+SDGwKewhHQFJrflvR2LVD7+Gd7J+nmimslmXI221YmYWPIZnGfjKYFYp
/2f5KJwPLgcoLvlGcpG5vmGof3fNkAV9+QypHEE0pVzWdPMHpQmYlxYRE3tFeOE8
OwAXoojuVjNJMYPLdoYbHe9RgHPZNBHzG8IjNLF98qvOtE0invtAMxc8pbzG/5Ml
7SuHiY8k4GNkG7y8762irICpmIXgv+jEuUMeWDCQKSq2wXapKXvQ0Qik9c7T6etg
k0bmRddIqay4U/S4ZlE4Lp1s9nLdiVF8M17hv24wU7e0O5AxZo2vhsQGuoTvPOKI
DmQD8mwX/0sZdzqdk4r9wuhOCOkS3xjjHBd624usjQciCFTH1NwZ2mNf4BFGmr1U
aSlgFUD9rEN4vadFl/V3hAqVWpcYEMd8eOX/pkCc/kgC2NWll6tsMmP6LQRxt2C5
PJisx4wfFybVbBFa09VJBCCZM7SxMDPrOMFQQlA94QmxtODabJjL/gE9nN92zf0T
fWVF0+V8dJs3OHNvLZuRovKrBjiF6Y/shdcajU64VQrmYGwENcuV9vMfgi5uAczQ
hRj5t17Hc97Q+IHVWT5fVCG+nwXicEU5r75Nout8IdQ1GhnRUf5D2AYW/Ze7HTN7
KMVy1ooGPxluUXkf7wNQ9UnS4woLCc3Cf9ukfOl1nA2a1w9Rkcij+0wtjBxvSpb6
fe3HoCgbycpmgZY2wegTjUZZL6t3EAjc59EavnL+gcHTQ9JUAKOOYkc4dbKwAyrJ
xIixPC3izRTKlF0lPWk4eL+4+mZ+czI7Z0BRkR1Oj7m2pS9yJdL7KSwPdNU5mgxS
FPn8JaAXUF6GmElZ23Q5/f6Z/JYROkTi/CJWqTlKbsbuHtlCX8tx/RUqYpu8y6sD
aHKzXvM5xNfDHMCp+d2aUJ5DFX6JbA+vXbBVRnwavkKztn4FO7PhLx22ybVGw6Zm
IGxUde7Fl1a73csLdli0IxavM8w5RhIkep5P1+eaja6sF9DZbglthLRH/CcxVkfV
hCaeq/4TPJCkwrqREcLAExFWg1U2t+dHWiH6YTPSMMoF2nO+N9yFCt30CAjq1HxH
h/1HXJycefkIZGZ7n2tcrBX05u/qJSaDQAIlg5oLf4ChHmi8WXC0Ki3bsGaPikW8
CyEOxWX3STmQ/zYWL+7RXQxLdFxmy0U4j5H2xeB1JCzU6H/KtZZN6r/wqtdM0Z5v
hL5nqfpjETQXd7LSGUimViubOY8aOcELw2vFjMbJuqPdknw/O7kSayJc5gdewT9s
avVNORFla4zkP/o7y0EoCyicbMwFJ+UeWhfozP4Uo8WBhGFMZrb0l6hJNSdlr0OC
jk8mjQWm74l3tPqySsNuqfZPMdaKIRgfnu3m7yxuv68tN+TqgbDZFvWdpqZNotvk
fBfFk4/Am1JG+bW+fxCOal7fha530RfeSXWjO9E2xCg+PFG2Sn5zFLKaXrCCkkV2
Sse/iDX2SWJREcGP2a2L+uB5pZyGpn0bEcCGDgyvll6v2t0gMcBGu3lm+lcFuqbJ
Mb/3y20vTfj2tIWpPjKvCxrLAjj1AxtkGBuXUOyd6u/Z2fmVoKR3ZyPAlOsq5o8L
eyxyDiYoTQpMdr43KKDCsuiRjpJqQkBEsyyxDOhL6JGNpcQ7J8qGkl3AAwbfotYo
PFPotqfjvB9Mbf+lm8uDlZvPLPIW+7LK8KZjliFVPEvUFbFVCURzePPldC9uyvax
UQNBwzGI81gycAUJ6ChwGDE68YZ6wHgPjfwC8dXzlHB39Lj9UQwTFMVlNy42mi4k
XvCaUKzpk0ZkPdf9uQ7202JQ38uxeB+RJQA5C6C0p42Xks0Nc0kkFSJkpgVSI/6n
iUV02NfFh3Yr1WVdNL+NQM8x4i3cPJ/Rv0riQgRY+/wJmO5bpbYIIwyL8HCSTG21
D//FIuzCS5USQihxFtYS2EoE82EaEzigMJvbuizE1+oJzupLlKZ0vlBvBwClflDX
gxB+FM91zB+fVk1Gc9sV8mxzf/ZJzfCSF7FYacui9bGZlILSkolcXnyO0UqwVlPk
TsUJEyAcUZeTqfjxUEqVHK93W4HsEVtYk9sfvjegFk+7t3oazZy9w2jNGtGd3/ZY
hpxKORGFDNtdxTGctX1do0rkXoa5j48Ydeuult1mmT1d45ENmVroNlMiJRTDOQ+8
eTRmGX6/QYOJ8el8cGoxSC7ux/7CbMkIyptmTr2RicSK39a1u/x17Yu7VtIT9TNa
ng7rcGuhdrd/EtDDV3N+vvZCPh61kwIeUlzDbvTQZo4wg2Qa5+e8SQQ/kGGykC8q
r1V+AUcG1SMzpVDYijBw1fvfrtQH8e2ir6bWk80wEzgyvNMdHOHo/hb4gUAP9TEb
NNr4cC6drvaDU8IkhgYlRG4juT3Pawe68avg3D8R6oa129gRgPamketPPXQzPD2w
wZ/GqHI1KETREBH1skfzMWr3wOpvVTD6SQMoUEZIWm3UNJEN5+gv3lVHHuiBb2JF
U6cScOGbiWy80oGgrcXd+vaosfDJtCJVdgsmlsF+0u299gTpnMS6XxgoFFqpBVH9
PknXGFMNJ4TT/cay5lKeGvs8XiDLhnhK9AblBpwBGV35Q4QZ2CtStUADpf58xvbk
hxTm/CX/WRVDTYdt7hGQdD/0MhCY3LeRq1okVifqzAZwUvswC6QtAF+g2AejMXNj
4G173r/KZkLmM54p3FUb0iUfBg5IjQQtw6GfHi2QXdzcUH2cm2otvEu7unwcMA+C
wjxxQRZA0mkIzTLJK2EsBiQKcZMccg3YarYpDKeuRQS/uFEjLWQo+BQdaRJY8XAp
+lHyW2ZLtsCv6SwKh2dP6VzOBdNca4/MVv1UKpv1aBnq7eEY3gdoxKhcKUlUH1dM
KEia2j7DwE69M37WucgoDNpTyYfUTDNpD29pSAn+zLHdhaayxvM+68sjV5E1Ogs8
WtqRDD/QmEvN76n63Yri+nsrotfXNI53C49JbPgsCccgYKuyeqZPYDkeLUIZBO/r
XpMmbDtgevn2vaLqy6sFdZEJrZ2nJ9GbvvsOiVwFkZ7oobvVc1TiZ7TQ6xktCUSW
O2c7YpXjEqKVfAijahxwN4IAOR3daPQzBOfv8bAeB58fmQcnUEEbw17tURqcB5FL
qO6omI+fwcZk2NgEhPVCcxoqHSfSFm4HJP4l2yXKjN5NO+MjFV/NGt0qkXNHpUe0
RJi6rCMSfptJY503TJ/gUS1vLP4lTOOqFpSIHcLvWxtmZIkwqwOBEpqBg/FtNrPK
0GMLWwLN+hZkllLiZPfiUb0hpkE4Cg1o1HTGd8zZyDVmB+wFFBUSEpziAhRNvIJ5
YtCc03HISQ1cdC66kp/d/xzNAvXw2wzhM85sjRfKlPyTXDTywCUwN/Gbt+UU2hLK
l49W95dHuAz/GljTTg5eNgjUDpOkFH2MhZJnxQiMPPZwC5d8tGRAQlVhp6fUPMFb
tSWtH/SBMB1I155cRxWPuL0+Weaj5DicITR4MwvEm1Ee+1Zrhxp9IphStbs4Yxqw
hQepShDE7J0JtymvhXp3F93nKDw/j6//q7+hzF2a6G0RwFDblSWb3mA8TXDb3APS
IvFvC17xD365/D1EimOm8zj4Rw1pMMZoesObbJBq0FNKXVKofT1sI46HTF84DKwP
6wPX7GCcv24wbxWSBBzKUltDIW98svZRifOlfskYUmhs1KrsEaWrXhrSRT4AD4K7
YXBEPQNXa1PsIdD50c6dwjjDssbB7eKp8AMG+OgFBXkhTobb4BGrPg+UxRt9HcOa
BZQryn5IaH6vVH7xyZ/0yWbO5halp3eKG7iF7eNJiPyBnWnqk5WjLhiXwtnD5aeI
xlsDr01qc43bzZjO/6yxcknN3x4H+kwVb4CjDhycBZZWdqEVCqhsA3fHA4E/7rOG
uv0eB0PtFIRqV3IqZQPOh2rQyMxX1edcUmqcSXOtTm4mxRJP4K2H7rYazQ6HKvQ8
bUyjRxQc1C2rOmhVaVeo0A4kjnIn+KEdchXVOf2Vd68gnt5qvxlgVWK76wIv0XAy
sA3X+Q6JcTUEGzXqVOGvx2mQhxI7XEd+8fi63xKTv1bONQ8f/36Y3hXillotQWoO
J+WUb+vfQEksd9b4AqagOU8zWWwBzr6PhLx1KzKzVjbvqUperOQgLs3udV6ButbW
PgyomyHNKpi3D0x/KUa75jPCkrZLm4Alc/xsF8st72zdpNxO+/IYGBjSl/dpxykA
nFcX8mnK19qUwSM+7KytiWa6K70qrQQ6YZRYAiUKccodMvngqHc09NWYYfDW3C6L
oHrsADHgXGYlYfQ/tObbYm4Pz18j/UU0M3IhT7WDEO2+jj42y8AMd51vByYKDopp
nYLDcgvF559D9dwKbTPc9r0V7/d+iXzVaPovTu6SzQUvRazrROmOVsrDwavat0F7
nteCyVKwZi9arpst5IkvDL1SN15fhuhJk2EVCHOgbpqxlDvMZA8Nri4Lh3SnyAa3
SkQVVnpKcfd6fJFk9ypZgIuF0hI2fNHLiUOCH3YoaOjMfHOdqXMk+ACM21PC90Ey
t8ffEIvOzpGI0QDo1K1iY9L96CvHdZIfu3DA3XdQoqYTR31SO9JnI0nVx5HrI8Vt
8pyGtkZXq65DmR+z4nvDHlWfBKk1m44xUHSCuIrBou4d71GpeK2GiIvfX+Xit4WT
JWNAgNCYjlr3oT9/E7RBiwLAE/Kz1gDWUwa9h1p34SEyuosARv3QbWjRQouVj1EA
f27WVeUHr/Ce0tHPx/hXdYgSDqpH+iFuL18x9iZvwJs=
`protect END_PROTECTED
