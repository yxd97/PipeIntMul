`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
43/zVp0ZmYhxbmZA8VeTRkurgmM92a1MBlE8PPKm8qhYh1RWpP04beTRpFdz1Yii
iwUuZvXxuOKK5Wm0Nx1BFFYlu0V3+aglbC1DPp1G+hagv1OGjSHuSDAPVw6VmX0y
sE0/gTSlKykHI2p5dIcjOkJxug3x5IcA/azTbifz7xwIAJrh2Y7UmpFYA+9dv/Um
jqHHPrq9b2whoYJcNd112uWEg1Len+JYs/nb4yYOuIPeVZPvThUqALohPljUSdPY
laucJYjYYsLstVC7K4eedh0aM+sFqS1n59CwUUq94ePKJUCv+oYVWqh7sp6HusDf
2h2BsvRENXmdKpQ0xa6UFHSPsBWf342DgbZ/U5X7Wz7IKrDrvGdQR8gaIrTKWAwx
uCkgwwSLvyolRElP2YIcCn8pnMBbHAFvG8DHVibDzJE=
`protect END_PROTECTED
