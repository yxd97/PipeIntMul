`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGn6CkWfNIfySlsDkWblKNecPTcywfoFoUK2mMtVgDZAFdDIaDGpypQiCN/MmHmf
E5PZZbkXWq9boE07qbu/8x8J5wYhD6bsqlAXOdOia14pCMniT8pYhbgLFBAEp0pi
qTXqkYnlOgBcov7N4PY0sp5xhPQ8Z/qyl6TI5Wt0wtNGJePXvE+CvkpFFCTMsD62
7FigYi7xu/4nQKw47JV0PjgTARumUiBd84uLi+/GgHviA2xtk1vyRSHKt629YIQa
39BUydISvmy80XVZkI3KVxIS9ZzNaH2wTkVSp5Ei3DiNt0VuVMnLkfsn64Fw5Mi5
+3ZLf06tdE46s2Y0t4iwQMm9GhlfUt7J/mRqIIp72RjKDnZjYWo0bSVi80jw0wFJ
6afl3sumhDoo1khfRb6rg/VjeGfzVoG5A4D1MlP3dAsqLk3EPjFRkTqvINxUa5SK
SQmDAWyXz8//88+g+XLvAYr4sQw94HBr3AzzY2kqOgwNcZjXZAXUTAguMHWxRIoZ
gYCzItB4xqHyoaAg1J562LfN3q+u4wPKpWqEE+gD3f0aKHa0wo4i6q0MXXhpQhjK
XTBNL23/WbJ1dF9aXFcCbQqCwZOw4Bi8txhOze6CDTFHw/4dMxvcO4yRzTH62l4b
mtsqli0mcbEERRDuPdnVSCHnawzeVqa0/Dwfd6pYqL0LvgBgszH0NH/37tHZq7gu
ogHGwwcAtZB1WL5pHm7j9PGKFPPL1VPLgmsO3uOkU5idCUklG9yxC39SDB57wiPq
doGrUhYwr8D4dMrO8MEGK8uEpg58BPptd4DDnMpK7t2SldXhqfI6oklywVxvP4nh
9alZjyTIBsID0sRL8i3beTctCZzQ+0SD55SMmvTyoaYV5AzT3aqWDK6c1syt5cNl
Xf0EiPBEvq1dpeuA9hAwLiH6jrcMYmAsGlBikaYD5SuvQLVnR+Lmdh21l/41w19v
JoNeiAy7aJtQeRmZMBc7Y9M3gRXiVlTy3YuVkqFwfiU0wz1OEezf/zx3iwXDvdeu
caxZwW/WwBfOoVnTC/2b/Uwz6s0alBvpZxjoVDTo30VlPQv0a2fpCVRcM0wHBRhf
PhocOq9fwosVkPmZxfKGriaSlcNKNhqSZ6nHo79urcY=
`protect END_PROTECTED
