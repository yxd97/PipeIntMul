`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htmZdqDhD4Cd5YAr8SNRNSw9R0wlOOXF1bjAn+miDtfp9oPBDO/tJ3tB+liDqufa
Fsq+kSm+x40zRKfab3HyV+43bEf3IXvQWA9g/Ll0n9gQ4QnDbEFH5wqTQVwImstm
uw4OQP+eQ1ekRUkzCwvsoE2YlvLtMs+H4J9PuHS54kkpbZTpSMpnoqri3UWmeVuI
pa/Cx9bdGNHDO21RG13Zogo2rs8TDGYC8yF6OtD0xgnKef4B4mr8E4NgoVNdAFHJ
fXWTFVqulLxmnu+0TZMq84jgsxxRMShX4uvYr4WryeOMfA1viFJ56/9oJXAmdKdd
31D9BXa/20eprMzekCIWLPIjL6MHIiuqmz9Jvu42kw2ZnqMgtDeEUnjMpx8XPUYZ
X8xYblRf/yscVtg10sE1DUYMJEjcaxJVhkNEInr+UdZE36FxS4S4k4HNhp5HU9NY
sVJqlOZ2CFzUzFSH1RaLoJonvPQeALIwahfMUZ964RY=
`protect END_PROTECTED
