`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W0qqg00Jwfw2sulj44ecErjYqodQn6dnF9k4UPEesbEWua43KiHVqlrnqOruAYed
y3lMBptXYrjFKEE6itLRXN94UdLM2tpaL2WyiNYkuNBfZDgTAYydbM4P75sFHcry
0CN7+RjEyxPnFInwJdACBBgvIvj7RuV4UTd59XnrOZLLGU3wi1KcL3MEq189LjdX
OD4rXu6+d6qSrVhXaGrS9kiFUtJh41+CmDV1K/twxNY7t7xF8gd0yIMwD2wu4quH
tB7dVgw1iVQKfp1JAa48CLi/WvW87LrdLFVBijn0UFgPEMO8gv74tRYOmpgRK+sZ
qYptPh22M+cDHji4HgpJdkJgz32TOM0bbklwiUhYVg0OhoritUjW+U4GgA4CCwpj
ynSYK4E1DRHCxA7WxlY2OWwqU1JZ/fEPK2vtc7hMcSilKLujECL5DAzlu7n5X6KM
MD1WYtZO45GzsAXga9tXefTyd2PSvtV9LweOWqrtZbQ=
`protect END_PROTECTED
