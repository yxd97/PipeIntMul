`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxPWIlQ40pNYojEb26kBtlSB9aeTwDtDvjKm6ist/d0Mor8HyCB/yVjeBaXYGeRz
ZHbhVsVtcDU5DBCDZKygN6NOEIUqckoTuCRnRKJVmtvbFOuiQvoPumLHmVHkgAXR
2VO9Y9w8DOK2TaHS/wlPpgTT0MYyakgqf3MBOtJ0rXQdLGqT7Ye4HWGnHKbT1V++
YPD4NOtrOhYwc/iG6vyLjErzrYgbzemnAu3vsJaV5S81Vel7psBTrxThe4MRleE3
SQkCMzafB8QcoDHiw5zWAeQCQUBN0DLW+4fnoWs+btgVUive2sv6+qyU9MpdQ1Kl
Psnq6ygjQA6xlkQh4Kxu1w==
`protect END_PROTECTED
