`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XgByQaEyhlt/Yncv19u0EVKVXxQMNJEWAo0ar62NSZR6+e7xWvmUBxnnT+F6VS8v
6m32RPtvMsvKpXkCWDBbZKA7aqUczpSeg24SGM739x54oP6GntDuVoWqf9/EQ7KR
jiMOflzP5Ovx09Kp7hfljt+1tO+OgxU1iItsBU+r4tK32EMOCdSe0zWtC+OGlhES
WLH1J/7rObtVjS1ZNXXar/hr3wUwta7QBjBB4HK+YGjISJwGqGJvxVRNGvOWJQqo
1NUnkR+0bLzyzBFlrkH6zzUam/QbhBjeDKHNQL/iV24=
`protect END_PROTECTED
