`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/UEUeZoJXF8INtsKTE1HwiZETf337QaiAcg0vdtr0aPjYSbHqiSJfzcrLS1Xl/8
eH6B3JnzgZbE2vgEntEjPciBSSC+P2UuWHV6iM2vCeOLjqqZQnRTdQ8kV/XY1SdA
KUiMZlCSjLXjSowWL1IJ8nUJJ4qc6hFBamaJbu23v/EBTcgL82A2zgniGV3KPEBt
HXXens8R4hlvW8yt0ETfkwkZ+vSTt5G5PaajeSc730TgXTOTek9Bfkw21hQJl4d5
rFCWwE1IoULhgPH+3OkUyllBFw0JwOdyrFSDqkNpibiRsJo1ZWDIbsrQzEVqrQ3e
8v0ZQtnrrf9PZyGKMVptJ4rUeqPD47qY7pSgw/xRWPTNKG1FMA4K4IsBJUlKjM81
L8Hn4b6V8uYcO7Y+oVfyc860vFebETCOkgNaJchBJKExrzwCaMMdLKIisSWTXeLi
iX9kR6gMn76syutrDM/HoFMaf3deSDWmaOH5u2v2uuO6XN4YB42X0ju4xHuxqOO4
18iCE0P/9LILEbOzK/GWBnp5iVtVmsmbACNeZUCkX77SfUeoV8J7qAY0ST33nx1w
fwY2O8DnPHfug14sXF8euraQtLuj0Q6gm4jVzNDJ1O2PNPwrXDMSGvtDg1PnYaeS
f8ABqoLg00IXyN+2z4YZ3zDixQSJb6C+GMt9mNpswI33d115ZAfOWUe3L/wSE1ac
GJ2Hijw9tNdK1cSMBGUvfuhzHdZnxnOjnx7ul396hF+czh79QNRjFQqVRgQQ64iP
NqQsTVoS82UoPWWc0wZv2SfM/B8AstADhNyc3ec2fMhp6ExsnIlTnoOOVs6kdSv2
iPMEQQXIyLy3GP/u6/Wdckv162Jcy/LpjIoTRY0Ty7+WgC4ymxZ0aKKzHjeMuQUk
QFb4eTNV1hFq3BZihEdvD4xqcQym2ByfnfmXMmEtdv5Rg5j7HOnqrJHfeUCZOJzo
ZsK7P3gL2XEZ9etdIr6doL3H7f0J822gwnTpjLZLJVrIURvxxOlr6gwxj/Ly/yN4
nLqkuf1KJCGgX4+wst5A4Flbu1qJQ7nIqZ8JTIabWH1CdFvEh7M/0UAHJRby9xNA
NzMSlYSlJRjOHdNWvjWlsgdQloToLPT7/hE/mbS3Y3bw9RMYC/G0JTRmONMudMmZ
Ioc9wrbHj9TParhWjnyaA0kMAfLEeiyxgoeT6W3AQtgNKMd+tYj5/A24sDaB9pEb
rJXFdGA0/4Wg5D7iZsJ205L2BHzM6/ngsa+3Mo9v96uR+dul3tqxsvNE5ObjCBDs
bWHlP4hB3t8bKh0HGpcvlOPIDYdOIogzceWA3ng8JVhTyZSZ+Y9BzHwJuyl5aWDR
RDBWBnodhjGPcwBla/sdBihsc5aqJWIspnX2xlj1Px41lZWBMHPF9pKVgJNUM3HK
C9eQdYBWukEoeqkKT4j3NgR96rPB0rcmC1nC7aR4P3xJb47t+bHdUyji3kAhl0mZ
2gyRGWcIHXDE6l6I0y3wzJw9GQ/SY3sfaec1UGUrG5Wpvt1Q8xNzQYiGj7btpLot
aElWlovN8LIHYlAm41pIgeqwkF6QBsLD5JsWx6j4GxFEtG+etgaQM3l2vZU28sFe
DLLAjYitEcPvjlylzTxAU/ZC+5521o7eg57SNnMiJZNpItszERLICfyeYa3BU6XN
5kOaa4kjCakLovO3nP+6VzSKYm2Jggr/rEWm+8T5rw0MdG+WwHPGPB5mtevGv2EZ
nYiio+nlS33iuWe++nw2R7MU+i2CK95Abdl55yd84CZgOYR8LMADAf7cVkPUt/yh
ZlvXWuIc9VBVNWJfp6zXlkDPjYOr2je+GIqcJok0yE4WP+MUmf5w232vFfrhhR2E
51TCj+Ab/TX5LrEtik3ywrQB0JaXN1p61SLn7WJnQhA/1hpCg5lLXXokypyRPFCp
4+tTfxSxzXprSBol1dvET0Unw+EsI6/ZRADfhLIRSYbmzzBVMObdjG+gbuwkjgrl
O2gQMYdMq5xulb8WF+JhAce1SJlf13ux8+T148styRHUPyymtjyzbJuvA/RllOQx
kSP7oPX4Sj36Dk0ZRL7WuEd9R3xWM3xHd3LZAGwdbp5gVGuOO15HzTtzWxoB4QhB
uHnW1eZznpL91VqxEixaufzUffnfN8nWGPYzueIF6DwXQNrFxJ9vZoHJWAWzJbfn
XeUnPE6C1lD5aFG2Hi2mr1+qeeRLbpOkMREEJDw/c8pAJcMBORO7VV0XmdsJdwkJ
F5fWNXWokermcdKfI7nHY4tbW7e9reQb+42lnEJlXjqPg24VcrD0Svu4gD3Ya1re
jeMenurzXi6NejdVvnslZWArPNX/45BlTgMr49GulJsByqKdO9OVJl+uD7ZozOKd
2rn3hdbU0x6nf2tUP1cRA5FBmxff6WEZWOj9pzy+RHqMyIWX9OHn/OJQOSsNurB4
JoyasgCwDyPuDdaqRxNm0M04y7tRIvD/oYdpXzwexddYKjGZHVl0DSWt0wQsb6g4
0SMiuKwLjSB1mpQiqxqXfTeolir0Oi2itpylwMJYhfNZy2v1lgTtsp2PYhY0Gx55
UvNK0BC2Z3SQvvg60uhaLm8rW8P9MKE9hLRXlC2RBtF1Fn7r0kXF320qnGm35DAz
F9VUmdna9fRCnM5xTOKXMw2cKOAv3S1v88rDySTqSl0S/PPsBCTDih9nUEV+2VDu
IAFCoTljwFSaBuAm3A4M3aNaUCNbI0vnfZs+68mJz569TXRAM+6i7AuYsoiWHwCE
mwNH5ig/yfd8EILtiyh18b9FhTZZpqLwrCU7RPsOZT7ctGoXsdDlNBZ9KAumx9gV
n3EVb00WIImqroO7P/CzU7JITIyIqf2Z1UYBzQ2DcreWh8Aoqnmm7AHi+vR38MJC
qS47VRJ+hPcXG8v2GJHIXQg5GG9H/ro9KYApp6cOn9LufJy4iEUHFJ8pP3fnT61n
KCrO3qEdxXtOldKFYTT3RCXLIHqFdQXGiX/ydaTtSYbzaHM6GEnptYUWbyB9zmeb
opM880dwP+OPJuBld9CF/zdv/jgv3kPrvb4rwHSSt/RUS2YMTvSrh/aQ/QdNQbwU
4gdPg0XEFhARr3rWE+ukVPjGZY7Hl+1yUedme47+buIIVby3DZY1gjbez/aY9LTF
mkW2soIYK9MwHMEm2fSlsP3sef/9yTJf/M8YVU/d4sldGEyIQeezL/Xc+dFq4FXF
MkKzek50TJodeXx9FMIgp5EU9arGxPMfvXgK9e5BGii8IwG71Ia3m/6CuUHylivH
CiBl3tf76Ud4x5tnEUE18FzkkESGCA5cqTEtlwGVo9MCn/PiRFfYlUH1R3eUltvO
gy32ZDlazWke+hVsL8O8V6g9tkW57hlzbfe1vQObiZrwVvhThRbBEWn9uiI429jQ
Td6k00KgffU455f/xM23Yw==
`protect END_PROTECTED
