`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXSZRsf5dwZn72/sDjU/rW9/Mz21OIwscRtEWaoGNQGK4Hz92KrI2FmE4EAbubC0
s0aaRpnxBtkKl2oQB8sSV1eUR266OJedSqMw7N9zi5l4hPTYRzGk02PFNfZIph15
O8Gn52jznHX3s3p4UPQO4wSZYNu2exzYhJfwydyP32ERrcR/ZvdFaXf/l4EjPeNH
pHRDaCMgyy3gaxkzT3O16u2x0FnuxVnF9PEzm8X+tfcOXbHeYpZicCFoDPSKDE7o
6tVXDH6twue+9qWbDuGKyXxPSk93H6Tuin2XYjPqpmjXYqFvPWXZoiJw8Wyfyuxp
9QiEu+FjO27OY2AQZPF4SrzVlCkDYzxb2Qzz1JWwX9idNSnhRKjOtIhV7EScqYtH
rjhyZQydK208g9EVaZVDUkLx3l5VcU+SWeay/93GseLFfPhxDE34bBwlPq3uqZ3Y
`protect END_PROTECTED
