`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ClrM9Ecryri3C0VzcBrKmwVOhvxVQ0fFzitS+3534hGWVvWDl8Q4CXMZjLsCr4G6
yb6ektAX65+/RixnzpdkSO5aokyzvTD10OkCeZn9JAGUw+k2OLr/4h6W+2JL8Snr
O3u8ZpGpLbg3vVhQ00LH8eRQvgp90tNP/o8TR3pJu/mMzX7AKnL4N2/rmCiuQ9LG
W/zMc5UEIwnnhi6cijU3CP7fLj9xH0V134vwlx0AITWo+lXmEJ/Di7CLGkqM8deP
7HeU7TJhAYzKPhZtKCo6Sw1VBGs5WopqfQu/4ORj2NmTjVkZetoWEfjLEGEOhkWQ
tdshTmEZp4f+Cur29k4ptCMWzHc49sY6Y7vSr+ld07tOUvhK1gBVj8jNAjjhFwFb
ei/ZVQ4pqEGwh8tubgvm1dKxk80CoOllYgdVUabRlHRcw7vUjDuupiemUEFA0s/1
zFlOLa1uO8+TnoWUZuPsqyMFVNYyB0NBKDsSXegsxBx6qc3HmSyhv+TRw8vaLrMw
y6iqTxDXteFhT7p9H5v999PcUP1jVs51VppiHShS9hnUM7sMHdCuCWine6Tdkuv6
oz8e5xV+wNRNfIZnEr+7qr7i8sfDvMojcJ12vAsvj9c=
`protect END_PROTECTED
