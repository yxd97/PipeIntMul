`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3FGObunHXjvjREZFKkyxKqu5hIjeu4WJWoDSBjUBD1r9SA50yE9l+jWW7sQOAWs9
FI7OHIkF+fm1MPg60szzWN61VxkJ6oz8WjD7FkqxLf4ma55qDoCx+uk8z3D4DE2v
r9GMKJJS7G+3hGomUjgylF+eW5eg2WZmPSrKI/kwSopCMHcEUz0LMiZ0D0z2b/DD
zM+/tFkISqSITeYpAqUDl7nv8G2Q3fPCvFCbwQXc3taq5mcgb8qn8sNOoVnXDCST
Bkb3HMkJVdURi7mKNM7oOh/m0BTMi5gdS2AIit0YmddJcZfi2Bd7sTt9bIK2nRFI
EHTxReosGy7z3UP85MGzE/7ExQBiRROwwnfWO50M/KHlpADcBm/oKy/TCdlWhyIE
P06uiXh6Du/g3H1Nhv7Hqg==
`protect END_PROTECTED
