`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nsxp4h8/jbQHbFZFdA4J0ZQqKETpJyeE11wZ60pLf7mVpOkmLJieKZB0OeH2nfc+
SrHYVbGSR8e3YbT2jWSImKc9Exc5/fw/zUKxBKZHRSFVnHR5qmrIjTUQ+2lujd2H
DmtxQSDJoYE8XKM49bgJe6B3I9F3OuOKUUkLUsiNF4rP1XTy8xFhHQbaJgsBhq3i
3xu+BLbp6paq9JMW3BPu9TKiSMpAodnbeY1s8pJQEP58pLaiK8HKU74tFE+VYQtK
rxZDSRdVI92RC4DTV8g4xDh3L156pVfDPut+DqhLDc9vW6ZBHceZKop3T2oW9/ej
EcwB4nUtKKDg+fmAuBuHpVRBl17Q2fCWYGVY10pq0Pk=
`protect END_PROTECTED
