`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6zmqF4NpqnpC/+tPE9TzxpNTUSrxOBWP00f/DHO0y1oHc6jc07OFp8j4WKIPQQp
r4P5aQmClgPKUSZHfrJWdTcgxgtuRg3Vm00DpmD9i69ad5NgKhPKfD9bB1i8/kMJ
dTFbdyay4O4kvhAUvWjL0NqaMlt4li7bar/ZIYCCrP92XvoAH7D5JbISXrV0kArn
VtwW1eALVbTucMcbjigAB1agi3t4M8Gyhos6LNadFDuY5e1y+TaQPBzYKPUc8jdR
9/UStTIaV5S3JSiXOxI0YKmrV6Dg4PdGMD2LJbENgpzYYHuuXoqra2G9uu5ANCBw
EgV+RSmxOhO4LRJi3G7NRmgtebvw6ORQ2NecqrD7YmrszBZDbeg8Nw7Neyk8scTm
SKIxvRT0OC1ud6YnLEgtLzuokxBPR+UvL/tnMJ+2EMA=
`protect END_PROTECTED
