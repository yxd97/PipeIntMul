`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mf5arB2SekBXpDl5D4bq84pFzaOih81D8hGeNEygJncvxpo9Xu1PMxz4QxQOd6wL
swvr23kQJ2h1TkedryFVBgjfLumzt1Lfrh5zOuQ+3YUTAroJYq7aW+hXZsfCUW8O
J7VPqmHXJRmGuxzue4hVvOQbMHzw2bP8XSqHebEK4/28YahlJJodFRibslehZ64q
6762P/3xgNhlqqr1p+QXIjyN9Ek5ldENwHhpOHGlAtoyVA1UiQtk6I1FS8Ve99YC
jusHNdLnFL454pDGrHWk3E8uYTeafmyPQkvv37nKKsOUvEPKUKGYBQY6QpBR9u2G
LDyepIVs/psOVwKUaigXL8KntJlVHX/lDZdaYDC9vi5N4CA/AT02rAFi8StpNmd8
6IDLvAlxS12CCAogGVkGjl43fIVV/K4tWIz7w9Kz8jTh7LDc8iXEwCsij+TJjAT+
h1cOrZJBUeZZeDwparLhCCrPnQ2BN1IlpJP5DtQFrWPvsfrHWoEPfkBFyJggzgnN
YmrpSbgupa2z3a+3Zwj6fX0aofQTDC2leR7ZDEM8AKnRDcqtD0uRr6B6C8rP/i2D
9OCdk9H0GOH6lHQqd3QvwIGWByDWPowSDJOjgxSseiBOhXH053Sr9EAMAt5rd9CN
K8RU7LvzgqmezKin0u6XlyiH/OjpYsYsRHKxg5Y5GwbmeBEszXjUNLX0e9qMjQP1
R1mVui0ZHw2PXVCCCDCLCgM6Iyc3Qu+rXEhuV+hSO3fulHHGxH3M6bLnKUGt/26j
YR15Ic+8g6SBifIrjseFx8hfOZKzT1Av6kcnKCNqU9s7I0HuPEnlGJh9q6XK/UrP
M8YD0iccVY/pJ5woxUghM4vL6xDrx9807eIRVQiOiyFiR/L7GU8mVRVsl/ZohJyC
jntZOB1aX3keL/p1lIr1Vghgh6MOeL4738kjlp7TbKhz+3oQtqVWl+EhUw4b9q22
afm+w+d9LI/9kNqj4asNxjM6cDf7f+Mk/+RMDU7Ug9Qz1ItRqjR3YqAlp2PPxiCJ
mibiywPVqQ8F2abh3k/KIzvjihLSDaZUQA5dpv2YFozwmnfbPkTFBZFQ6gxGfVzy
rKoULEYZVidVahnTWHkxvTXEnSM1AF9mkoyrxejbd8pTCcUYLhDZXz/oQ62Mlntx
JNNLrXxwis6jjxfBUu0/WHmHXmgg6H0l2a+3wXlAqlzS1vuR9Y6Uu0c+HnfZhM8L
0q6pD/mf2jO+ZLWXslBU+X4a3cFbTaxhR+KPHZyzkXjaa/hf6nvFkP4NcU6iyXVX
ERr3FgT2x1e7xtfHz80ExXTgxXheWlIy69AYEeNeEU/w2rSlRbHIl5ZLPse5ddgS
fJX4SLWbGVi43SxZQpoQLyrCFmLvHBLT4YMW3s7LcIAVvWO3zGeTMQDadsa2kjyq
Q1+rfpjZp3GgkEno0YNwfhNocrxNIDO4BLaNhUTzF/4S1aD9AbkcZ3m6jDizy1H5
8m+uiCmHtMKFrwm4+PkWja1yzkrJSetQtYgv8ORClxuWCdduhNCvzP9ydnpb+GqJ
vT56tPhNzrh6sTBdw+zkDeJTq2MhiGORqHzxUwRquw1aWb52q/hhSZrPhG57947T
Jf8ag8cSZX2U28h1Tyb494ilOCruIZA9iHyARMefQagRK1PLDReVkPA7T8lxrivd
y9ehKG0M/ZH66IrPD6nSEBlgq2ey45yI9QofTYoOG/miMempgdgBH8VkcPldY6pJ
7bG66SxjqBG7i8O78T1OSkQ+ji53bswYlqvcY0W3Ep6RxP8n6mPNGbnTanhHmdF0
paCVTJY3t4xYIn7X453q8/V1eDfh3PTrkWU7K4CxxnpVXq6/bMbHLlFxMariAf8T
V0VRXrEZYLUcgzsJ5RunmAAjZ8IRGrA37mGw8CkH0eFxoNRLShWEd0T5KKLx9KdR
a+/uKeARnJPj9ieZKLWqlxMHIAxMjDYOrHJoHRvIIZAWmoT8ZUPByCs3gatxVcjW
JQj8HWkKOdZVz05Mw1tiV6Gt3/9iWh4UBNFTB6JZjiXmUFOeqUIRdEye3O44kPpl
W9PuLs9Ebn6AmerYWKTIx6JTYu8WciLtYN5LmXTdBPxHeUe13tdrWkFrt4qa3x9O
HBy8riI7ZlkdaMZDTuETNRLt5esOool0/Nn/cO8D6I49L4hhv2DhJIRkDUngG91l
aAoQ0Gj40moaVF23HCQVje2BdL0PIxtmcUv/tbQlrOzsG84o8+Rzurqh2E6soTVU
oasPMcO8W6jSQ01vqUcGXzh7dpPALPQSS1+ci5kaFpJO7l5vQHHvpqr4joaGdLs9
/QpVjyLQth1XOkq3upqRvuFnFbRZtGAqBpUiwI5F9kquhi2HXU2+ky/1nS+Ti6rS
ytwLi8vfn0yn6FsA3TkWtpYZ4qcyaJ2etZ5FEu5ajy2bvHe0W0ttijOHIb/gliX5
Tr1BMJfmS9jYCFLlb/YregWAwhVI4pwJTh37L3UqP+u42K2RbxwFtoEWTpPHDTke
QWLkWcxLgS/bXBpEFL/88yeKuybfxAyZsBY1483eNH95p2USBwUYVLse9D93vIya
SFcseUuw3km1IbZm6z+dqHAW4dqA0nxNnYwwmsBJx/ngLnmGwnDCaFibo0yMSFYh
1u+XSMkuZ8zTW8IH08kl6fG0Wrx+zTZhKG54Fx+DL2ee5wbBiSXbeRCUfjo1MfQV
hZ7IW/MlDmAH5PBT3wVNzXebWpT5qvwEHQHXegMqduVOMTYEMRTqjOCOKN4LiG5z
7jgFn4Xglk/baPWoFbP5ZNlKnERbhgC6CqbaRKpNzmaSxnSC+9AHPrFSVxpu+3iK
etfz3B6foWGp4c8c7Z+tTvC1e8Mz7veWcFe/JUXL40Q7mHBBPFmPSDbs35ESRAIn
tT0zCC3w4mDaIN5qoZg9MeHRdSMvSJqDpEpGPlzw3T1rCr2Ch3EKEcO/pFR4TXfm
8OvrpL78yjZ5hakG6fKRN/9e07mH8LnZ3SiYku0H81rPSy59JefbtDVkpIOaoHQ9
JuypGYgzvWJFEa1FbiXAIMxhGtRW0PZR/rqLni6t2BvGoNZeT/sW7soktsL9Au7G
2faw8ICxtYEdPJ5ErgOr7tKk2qwloigf/SZOSUe2E7fc/F+hzI2800L14McBT1rL
cQMEpLwQCz/a+9y/dITGQP6WlODKqpBPr45ww1AqqRdNDODmpRVV+xzSt4i+WXz8
hnBEFg4Q5cKQHsbuL0sNYtM7BlACd2iqepGHrn/7RJaQwjMFNjnt2sXSQHSjTPQu
/OOCkYmkGF9aL2pi1gRrpdYw5Z54e98rl1dejBL0GEEVNunGWqqfzsRnxS8rFPkb
1KGOYRRiHPyPGOnJPi7VrA==
`protect END_PROTECTED
