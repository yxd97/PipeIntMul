`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TGo4uXML92tZW49Eq9MNkpdIwj93pJ7bL3WdS0vEcM1U9Nkbe4T0KmeS+ij7ip4s
7HoazZB3FzOjuB/DSnAtuv5WYuM+X/FD7kB/p2RnQ7d8z6ZlIYXT9rHfb7tac6x2
gDB1TujLmmy9dsbiQYSDw0PtKiMH5wqkHGX56JHxZGPre9eAa08/A50NfIr+b6Xc
L1laqiHPWFxqJcK9rWupZFS0ClZXQkX72/I7z9/wfcrBdOEVpubXdZC4xlUskwMc
+BVbs7VT58zPV7oe3WVyrRtDF4GNvgQNN+8/MtjrJdEmuQT1/bpmm+Ooa8S2qDZY
HjxLq3Vao0S+z0PJUfN/IDjK9mUsNkIa1mh/FYhMrzQBi6KR08pTnIbDrBjYIhRz
nWcOkKtMDmUPwrUR+9sLJzx7ECA50kIkrv7vFz2NynRIz7c1s9SUQgax/GP6NkSl
D+uViki6j/G6qQTERcvOt/XEOSrtdh4sBrOHKgCoKc8Ct1JRqG4MpDtIBmmXH52M
54tb17rp1klVCNgE4cZWoXXCfLfRU53xaGdw/+rRoG3A1g/cAeQSUXcOt8zhq1e6
QEBBpLuwKYfGeMDR4LhdkX1vI8oOcMBOX/G8cNsWXaurRhhMfA9CGY9FMwo4ZGe3
MPDh33D346lrcIBPggUb4Uy7Jqpp4it3s9cxqWkLCBagjnAzQPEqrtqB6wOTGfKB
pujCxc/l/wkGPfIrQFDm3+ZNbCb0Y5RG89vtcGNzTmUEbRi05ZHOjgyK+bnGQFlj
GoXglTYp9/UPP+uFxpQP49fS5+/twlF1R9st6C6nE/CIDIEkcOemhl/52etkGzXV
F6JW1qF+54JFetBH1ojsULuJgxU+8c9u6gJjE9Yso5M315zm4h6J+MLWrFkeKvJM
WD6+d1Dqmmyz/2nHrTjtoyYE2XZL4cwbsgTWtqeZVI3Wx+CLyxpYZ5uPB3RYUxAI
jrQmSIR1pTlnu9+SURVZRcpotOmpbPn9tI2pe/03eSyEIukY/AJkC4ETvRMfzm8N
7oqiMGMbdFhfa91cY0atsNiTa3wSwcq/V+2myxld2sPQPLfUhcWVCYIehSyQjCyR
BvKGdu0jOuENEF9t2+06IcG8mGIRj8lo29cvVtcS+CGegBt2759RyzhsEQssAfx1
p87l7eSMPP0NtcgGzEmTvG7rqeSHxIt/w+B5/5rSG0zPne1LI+eTuMDMty4YUR8M
sVF8/hyQ/YH3gfUiWFLEBUFKqiohIaQLGH/s8O3u8cFxVMVp9KTkVxvJXqajgZNW
BKweDL1Swy2UfCTIGsUPrCw3D4HI4QN7k2TmN06DcAqsWVVQak1YD5RN3mk+bG39
cGhOc/tJpZuAPH5qM5CD/zXQf8XII1JZZoI/gcFDujB/C1OauB/vRvi383mpOS06
SS59BLqbl5nhMYa25XkgK1JCFtbvcvcydj3v8vX+Mak=
`protect END_PROTECTED
