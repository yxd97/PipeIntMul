`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ujHfOUI1qCibkTvlCVwqvppSeHlig/1sljmfBc4GwhsJNel0BA0kogGW4SPbJPn
XATZbSWgwvqBnfkzj1nBticaTciL8f8slt/AaA7ui/wT1QIqIJEvj4TTDRHcf6bH
F19SDSv+M9mQCz9j515t1/oaA88MkTtxowaGtU42rzbRJuFtP3FrGpxeGcos2Ojh
Ri+nW//BBSr3MUSBNV+uvebdQ2vZV3wm3fBz/WKFH/rrVmvF1rt5FPa7YsAhj3wL
LbaandsCe9CPc4rVejMy8UNryhqXzx5+b6kfmuVcJorBLjo4tZF3fPTAJ3ntoq9h
8reXAk5Zfm05ngTfp2GX/tlXnF0UWxvTZL0H85Ex7y6KKn/Jy5kuCz7eAKEzZVkc
elg3yjQCbIuijXLyRT0l3/Hbr3SSEfi1ndq8Z7bQ24Z9BrNoJ1iMkX1hbLQ3cCGC
iUFzCDRY9KfYAsny84xA1azn+t/F7cZ/rvAfn1NGzLaceqnVR1QazJzOAszk2eFd
HaW4TYXSyCJrKHHM+rvIOsr5HjenyOGtkV4otrQPY4Aun79q73Nqtsb8+sNhmN3X
1ypRa8cCsdM9XHL4bmXl1VLorsLwTvSe+e6a+VfzWozKEpA8X4aQtIv/UtdkXtzX
G+qUKUYvsCFTnHGT2nDjjyZGh41rJ0ByXkCGnuUfXorSKCb7CxGTOxum5fQ7u88+
QlLdFE8RniruJLudnJIoBr6rFyGq5sO3Aqhlrt+nkg728+5VN05Svs2R53i0Rue+
1nOEbRW2qNSmKn2vXuCdx/D2KRjYxQfgan+K5K3V7O8cfGsSdTa/LRLIjTkWCOFM
L8HrXnmduipfyAYuPG9uBt//9pkMXCJtPvFJfX1SxcOnTeQYDyGaXV8PcC12jof4
Ww7b5RXe1AAw9emkgWQyVWbaHnCjxjq726Etmw5+sAGzgC7WwSRxErMdLr3skMW3
GrX9u07Mhh6g6LDgb2cxUrM7ldZldC8p0bwOP05xg/Db1sHBPOYgDuG/hNerNcq+
TzrM6E5nATEdhe5NqZBX0Olur7xreFlk2VytK2YAdVSKv05ZSdhSpLNYvS3fJ4bU
LTKtDqF6xs9W2Vlttz3RMp1gsImvPacxi6HZ3IAVHDHRDZahuUQ+FjAthMQpWy/c
Bb88NCjJbvK3Lcvb99qDmHmTveHBi3e3JX9HcrqNgQs0fYybXj4bKrqTLspUrjsX
85rMPpK3jzAFgy1rb/Ig9G/5PW2lxWcq3hIqeL9f/V1Eq2QCf7o/OcV6Yd69XyJ8
ccj8xF8j+EiQ8dbzjhWTzqamckwo0dcFyFFr2aHkpKAQJLPsxxGkpQlry9Q/rYX8
3YXU7O9BzCo2A04fH/cTmzrQ8amElS/iPe4F0pnJkC0w5Y4VWtjOfM4/t2PKMqRD
dkbi4dA7EkyiH7K3ZLiTaY2fR4JDpi1wLtR8xB+DobgPfLNJT46Db7QtTtU2D1j/
4sg2CSwqMCCcyb/FzelY0fhEe4V/KSFdAbKEOahjzMHUmlAEJv43CIuqwzoAFrBk
xwRX2Y96fE0McCkB5Jr3EPYvPc60C2nVzbht5I69z/0iDnRUFldi58EACq197dFM
ui/Mc50J7NYhmv6ltIbA91sLGhezgIXDaKUhucIN9L7AW1iX/7z8QqNX53JmlMOv
H/saRqKzprTp0FbyILiC+QTxE2RTgVSAIk4iPcGJXTM1z5SebMIW0ZNyeSGxX2Zz
YyKi2uW+WqNJ87Kqgm2eOkKSoEkYA9YlN1gqb1PF0YB1f03g8EgMzKHhJsx0qBg1
ezWeFuak9HAsH3whviKUfPzEn77nV1nDiwHZy2Eh8IcuN4VmxqR+6/aLMHjycxuo
/JV76GIDuVT+/QnJ9IK/OX0lkKmayaxc81FtMndO3FdXkR5RYD+EMXep0Q0EJfDz
7WwM6LMwOMnaUOMEyN+i9LgQbMGMEqthZI2jgM3ukvrKyizmm7loJz6qkIyf0zg7
bUP55/Zqv8IXrc21DLxUrrKWyImwTOhN0qWUzofG5JybXOPhP6DG4/9VpsUsKfxU
XEhGRvShehjEccWqDFexZ70RQETdMKMRBPKXlQ3As8hlKuinUgbLrhg/ziNNBpmn
cSKrEA1YGiYPmuO0Cs9ujLmfeT2sxw2JKCAwrvbrbo51jSIjdFf38rtvlI3lnak1
sIYYpxg8J+hIZ5bIfwRJgDbcNKqxFC6ckf9N9wFICKFHHIk++xmZyGhAPZMNoDN5
6Qxeil326xsAKHL3ZxpU7009sBGckpnbRTH30htW/OdU0tGevYumShcozjej9Dna
y/J10r2aqQyWo/bN2fI5kcsESEXF+fiBQ4mZ7gHr+kDdu5m3rYahdCqalv/sRmdF
n6t9t469ehEhWCXX9jlH7MvcsF3nNL63Ldwkf+IlcN6p8pzQpFtIeEeW+QlEQw92
v03OdxasxQ0RYL3fmeRKcgW/Ii3S/Jsu9otICwVvI/MjaLShN4fMX9GBJDMcT10v
9Zd8zes6nFCB7PkMDTMqoNcqac+FjvAyr0InKUKqw2L3bF2oOLITb8rVhF+833ae
wlgzqT21WnoGbMM6L192ruiL1JcivaHVhqT4y6Bz1Ydlzcbiw5ApSr12s0eOkiYi
14I994PcK/e0XEQrTQvRuJEXWTkiVGf+7yICkVRe2ep06G/+Pm/6K1X3HLH0Q3ns
SaT0mCzaw96LajStdGRJt6ERLOZAy4kFVd9lAfaBMHNIL7NKfIAcfqc8ibHll28b
J9gqjbQNDy0BNPvsWrp3m+dGuNjrTUxLWUukk/C7ciyj/cszPeP8XYzhYvJUYltR
W4ZldhLRu7mo2k5JlnnoiyngzyMx4sxuBOe8Y0vSOBlO0ZufONaRag1XO2L9Ae7f
SEwEO+2mGkeNvKF/FkQlwXGk/Y0bCfMwlLs0/UlVtSi0xrpTu4ggpiaD0M1LjzIe
qcxCBe0X2knHS+frXJD1SbV1I+gAWKMM6gwIEiloj3JK6vqiXY5b3gLdES5MQ+Hy
2/UAuN4/wai6Bhk5QrvaQ0g4fnjdDjBCpq9OpEn2Q0lO9yuIui4BRJNimuRy8JIN
QoursaS3TCwTAZrJHMS8hzoKMNuIisAf1zH+VrwWTfp9oabFtjhE60pIGKiucxOq
hidlh7q61XCrtR1aJZnyh013JeJPSBiWygMQgdKzMpfvsgQSau6FD44fj0HORKlp
KbeZs9ccpzcnXVsnY7j9EMktlS36BtrVeAcKDf46Zgqts6Lyg6QcP97kc8ZbGcDq
f2WBFz7mFs5AX3lRAW0LldHOLDL4YAgC58u4xATlMEIeITURur/lGU4AJ8VRDFAE
LHLsFRryucusERaMG7VRXJDRjwfvUZCm0De/5WQ2M2BLXnvXizuNrjjPA3w0Dhyd
eIwgOuh3jUvO86VG/CVSB5N1Hu/Q0WgJWxi5jP9npPZAJFypfr9LIGZwZTJaNk9e
h/AD0UyKFmqhvVqShmejwDKdrZL6YFYTjpqww3Wq+WzP9YFsHjwyaemIyWi3u1QE
J+HKnFAdaMYbUbhAjS+ygwRgVM+j6hzLVwz8mrlNVUxYIYdbPL0wHo1MDHh1ssHq
fQIvxoiAy2vIxQhaN3m1bXPQPfGX7lp8jGlEqunBmq16fqqNdeRzTJLPFvM1Eip4
DdwOVAZgJplRBB3EQSa1e00AoAzQOt8mw7BQVbgZs7pdWUDDJw9WMLlOh8UUXdMQ
filyRJlB4Lk5GBApUll7+sCRbangcDGi6zyAdUX6+hj54f9hLJxvBgIjV3mzKBhc
MBLUhzYpoRWeu7PCwuDtzQuYuEjC26X9r3k1azgrHxNsTMoT94DisndTP3xSnvrK
5VJDdMptGbxLNbzuOISVyeMyM4Eeugx656O2MyKxdNVAW2YbRlPMVFQM4FdG/vjw
yDddxkt7T4hMYxCB6uNH5tLGINj6PPRG35n/ROHUx2g1Wd9Qln7xedIW72YOFxe+
2Nx9xIx/NeHb11NpkMiSGa0CquSVcE6VLaT9T9/Tmsc0uHRseEYgJ5KZV3osKkL+
rj5t5nIC/DocLidHLZG9uCb+ofd86z9lOFcitbgOhPqLSpfP0u3tpvAOwUSLfQUl
e3D7kah9FEL+jHegOZpugVLPJeMdlMynIVsEMPbOUycrmkzLyQbd/sjE0KKPL59E
3avBD/6OiHj6Uxbr4jFmKVxT66I8qSB7cN1nSFB2c89qWLwJUd8wXUJRgTBPJGeC
XyaoNTqbm9qEqMFn+cfYKlHIV+vTcaXkHvtUP1eME/3JLNFi60EvgNwyGPuI/HJE
QUdeGP/BXOwWFEalZO/TxrflwzE0STpDuiZ45U3gbDKh09zoS2cCzJ9sRs59ME4h
5NW6HuASf9KYfAWB0VvDNbGd0ncfSpTbShckiLFK02ZyES/XuYzOPZOrGxSVKzLD
v4dxf0FDk+UGujUB1jZgmWjwV4EAF6KNT9KeyYO6vA7kOALDI+cOwPIqgl64IMJf
A/U7ZGxmGejGEOTdW3wka4g6Y8ttaD3XhtJwuyFvpp2RGOoQqRSvQReaErpZ4SWH
pEDqnZeRnD+9Hv1ONAwMiJX/9ZSp0jDmJO0G6z/FBuBp5WZzeRCO8xn6n4Qn+oEk
2hzqFIBlV5bE4QVzzSkojVn4b7wZYEsDGYOhYRV7GeCLakNUxTxcwjpuFRhTljv2
QbIXxczm6jbku8PBNR3PqZYqae6wAruV7ym1SQ1sBRL3tBddpf6yaOk/PLoHSbo1
sgTrHiZZtRNL2bOeRG0yPZxlGq4rXSqgwbo8UAg4atsWyN676Nppxfo6Niebxdrb
bM0ru4knbpa3mhjmb/p7C/HwyweTeDH/cQnbJEiTQ5OWcv1szimfXeC1CHVSFjhf
PqlHidEkedU6pBpMYhJBZ1pZTehod2Wh4HL80O4NER98z/mS1AxGFyMq76TKf+k2
qAX1AhX6Vofb8wIBSPCSPmTmebWqLYcj4DRsivlgj2B2QjGtsC4NxqyUJItdy8rU
3J6ELpsum1ImiPGusn3wrTUVqlnJuMh88LN8IHR3j5iAPl63lQbqt5A9PLyD+lln
petMk2iPmR7kdB7/0eD8mbhZsYgmrjhsUj/hn+slw+HtBimgYl6f0fntb2RG8YJZ
AoBzhygUu1iSFEy/L3N53eYj3bOS2owX57mdZAVUBCwM4tLdkdcwxIK/l0/Clm93
2bivTH4nVVoBT7a052u0YK1tiD3WxMBmZFJA3HbkhcilbTbq4vSNvUiaLf7gIqBc
SKziTF7wmeDftk43t5XX0wokuJdMz+y6o57zaB8t5Wx/u2gDF0jJXs2gyc23OdS4
waZIQDh5U9jSt9iBg7p7tQYahHWiQgqjtzOoiPrULVJHIUArClu5w1Vgb8oSmY15
qAwOUV4njwEcvwLcHRTv5SEE8o1aina8zmiNizImxqrv79Cb2SfoAMBm72WsWRtu
lH5tv8WV5inthduW5h4O1mI1v6Tw6/Ch3L4KqE7CQ+KqqBfD3M5oHLgG5Zj9i2A1
fESrVUDKzQyz3ObSPJpCHvLVjhXHH5YH5/pthLKtFOBwVTfCV2nCw7VAP4knBSmU
4ZAYwGGuGKvftoDhp6mUolcj0V6uKtETZZT+asEYOteFK4C5yHxikOqOIl4Za//U
yH6EFgAZxvVYw4w1dY2M3/PFQpWpvkuuqU0GbI+vbhBv4QaCzPmZo/vcLRyFO1XK
/aSn3m6KxyQN1qRdVlQRRyBqeC9iPi5/e6BZMDSoNM5ZVz28mMVK6itPXI4agsf1
4Wtw5Tpx+T0dnLpdYtF2nGAo4k6nH5I7hIde/jk8BvVTytnAXEs/Cbdp3bJHrj6/
apLznB6DGt1rCCejqK2d/jw3nMX9dq+aHiL+EtUCK/zUQ+qPe0C99TaTuN7j3VNV
EEHp/xhgakrdvGxyio8uOZUvuinjMHPpWJuvcwnQTxTYnQZnnBykDfmc/izqaxna
fjf93IEXUw9emqfbweAUefAJf/TJC3+1q7hWDQlo7cacMlnYTv1XLQbXebZMbxjq
ixqqYFNtJZX9muwOdD4bn28rFkuUYkKjWh5Kd3IbkIY0TH2rSv27mA7Ko3QJ9JMc
dAxCN9dg2x50axdKwuSqIck0Bn52SMCHAlEUcIFUq9BSB3vxdQPJCMq4K6bplF2p
aFqnEJHE8LCOHHMnb0ithDuxTNwtrd4MXiaxybh7Xw1mu0/N12lLtuefRpApsZGE
cHe5xCO2lWaP+quFBAlNgtR20Q0AMTt73A04+/qHk+sCrsx83Tv4Oe2Gf2ucltb/
+gAXzPxpPJbNahmiy0W0BOtLucJCxe037LggaubY0wjsXhMxok/kBiJHr5XwSYE2
RmkXorXjsytlZNEMveTj058F2OaU6voARl2+08icNUFzdHo80VMmt7QoSBSoQAbi
b6m7tJK1S1ml1FCBDHHnlTCW/RNqeaQz1WbWPI8EgyX3+/Po5UmVs7IXQ5IPnOw7
ZuUYisOatqxNuZm2bRAUWPxJqS9AseO6JIW5mBWa8/g4Kk9sssxVFB5lU3YfqVqw
3grVIlrFQ4FOD78ojMmS22i3RZIFiPhfqciStqvN+AcJ/BIkUnW95dUIcxMGmSK5
cBWZI7LkOFLxoJYfq0XIDF6dslM5TVitwJtf4UOCtFCnrlOo1RyXhdue/O4sYhtL
ECk8yiBLyHIfOqN7zwBp6t/ohz94Wqk1U8nWYMD4PNU58jzsV7AhQGF7rTWKnmbk
hmqi7pMDIzFzNfbRUcGL2VMgWpL+OGzHvm6tZ+Gb+KcyAGhPHuXoSChCEJxM5euw
DM5fMbX9PCm7rtvqH/5JtXZvPZuQlRKABZkNKChaWgftnTFLz3g0nKhz3NCWmI7C
PDAVvklWLX10OOL5BBeX20Zn4hB5tasXnKeMQBlk6/NYxxzUxO7vO6gqpMLz5zEo
8Q2Fx4bIo8KPfrD4yoXJGTPEySIffy9hHG+FvUwtV5KpzfJooGwYu4k5353TkH84
8f8Hzl9Xwj6dF5LTg+wwGRMZUIQsNbfu0NqJXCq4KGWq4aOawyTFx2ruD/PzN/Db
sFqJE+7qopfc5bqW8SfAAxjCzKZ7j/lkslIYpA2m2lj3GglOYiDc344Xb/bMMbYY
HdW84UdIkXf//bALwdlo1YnFS024amGiEo/mhzwpqaAmfZmuWn/S4T+zZHfOZ3UZ
fH2vf6Qa+wXaO+R1Ykxs4v4SYKWkkBa3akqUhejVTlj4PRP7S3A7XA+jpzGxDs1n
xLdiksuN2O0HRFYko7BvU1mwuIU50tdpR3Zii21vVL6qlktzRPo/2r0NXe1pG5fK
/2VG2c4PhOaP7Mv2atqRjNh9M3J/nbJ7MvNtoHF9GWmPAswuVmD5ovsJlJT8dJTJ
7ozwApdFhiYyPdK2L8EpcGlQ6Wg6l+j2r3yz2XhTwSQwxlGz+6L/xS+p99zBv0mX
eDBs1EcJvwKKE6rz8c7skmMjZvOg2slUpUgUW9EzGyb8OBl+RkOcTHGrmKqV1zQb
e+IT/V2NXdkiHbWaTG2jXhnYGz8HVQgj1oJ/jWyC76XCfTNfVr7Zo0EtujD5j5h/
ROjTEAQz2PwHIbm4khCGjWqSt5X03ZXb0RdcR9qv3+oGjk6/vfQqP36rimcHuuu5
iY5LJw7w088g1yMoV4V2K/MRz/p97FsdY/uaMbEyLMdRK7k2xGYbtuGtBS4R0Q4j
LtR6ry5W5YV61+fWmY6E7SrdBonnTo14kyi3MZqMRJ1avTRwJpV+6sTBoHEAQgX3
G41NCSaXNbBkLcrqQe1SrIoma3DBzPNts2kSFXj+0UGRlbiBLYLYLR7OkjsW7BWL
/ALb7oMjooFUU7dNLIK3xGzn5XjF0IzEQyXfYZZS5HCsc3mnJzReNO1Tg+xYD2ey
KuVPq1SVHkM7QzMIH0jXTAPCXD7SzVmEPpe3oDZQKfG1IO8JXUlI4Gt6ktN+QRXO
QCeFOhpvwKzL1XhUr0BQz7LBSWXPOo+yX4YFjPLjsj+WjU1BLwf7IFI+y90fyfJB
V+TV3/icMrBOGYYq13WIeK0P+DBCCRmL36tSfCvOP7dM3lb9y3SyCIPAVOrujXlw
/qaayKFYS7knUh4KF1B4fYRG8Mfd3oibR6NUF77RW3ni2yKCBvd52z85IrAgWznb
hvDpPcMsfqBgXD7fQ7F47Opmxgc1e45WQ+Eukv+SS0ncbsmGbAcJf5LZznLiEmEd
Pa2M1ewQ/rhQZgTfxVupPzR0i9X2VelX7xgrTdspGHhL/XNgp0xXGkK1ylPWu79b
4iGeYSKq2a9FZYNe11uL5eCi4WneyqzSdAUg6h6Yozz9KyOzbZVE9a/vPpCUg2r2
OPuIUahpJKIiHfHAq4jNCxp6bs2sY+bXKvOvzlFQveITpY84dxz+huC120KpXaDz
0IlH9/YTWPGo5Mk7J1RNuJLb8nekHJSrERaP54jp//LcpAj/tiEy+YDZoNNZ/jau
TsCPXZEi6DJx2nh3WNhVrzJm4+KSQbPN2jXjXD7/rbPzBpYiX/nl2rGq8wSqgbn4
FlRa9qEts9+V/mpZ6JwfQwTKc89TcmOv2SeIlTNfihWm9Fbo1oFgRiQfe3CmLjyX
ZIGHatF0H3IEYiSgVhqQBgh0XEl7SeCJm4543gFWOCP/Pj6eVWck3jNhUkas04c2
RJyMdO2Cj7+AuU6J1ABCeRaQi+iox1eZE6s/NFE/4MKepFamDhe2o03PBodpjnW0
xMWXRSw8r39KixPws46Zyajjzc1nNypBYnzm/p2YDXSMp/pmcaJGvMY3TYFncWfM
+A78Z98ixC2RkfnVO4CqVLDPsPs1MVuWg4sXha6n1T9t+c0B+ZD3QjfZTbVOxIFc
kHxjEBRCIdh+BQLuSj/9LyCDAiPuVkYoHH28rusY/3ohSAWd5iFQkywDgpBx9UT1
uku7CCMCr3adJfpXKLvVPrzbpepseR9xD6G/9QrWW/l1ifLrYAocGds4QdVOudDX
0HmtB9fArw5dzMZ9EVxz5iT+TS06c7YFadNhzQTIRHMgVWX9l+Jo3sz6iYs3tAqL
fnsKP4KNYMw09UyFCsjIq8aPRCLCgtEXxumAO9R0YKqPZFmpIoKuuYBBBeTwYVvf
BjADl6aXdtKjwwy6ox+h+q9d/Z2hQwPEXzX0RvzYedZp0ZDR/Xw+rXEjgIvbwWWQ
5pBrLCPbMQm0DWtD92Sc85eCqsN5rFcLquYf/72wit+KDbsrDgknEtZkpeJxVs2n
GewTDv07NmA6DMx/XzFx+L3aHHNJxLx+Qes0y+bo6J7wnRNvBtLnNprdscH++5G7
TKM3+0jClxY29SLciVKw00cZSOcGyjTElQ1wwtqMVddLXhg/I97sqwOFbH55O1SW
ByLC9jZ9wzOZAi3Hoff5IwJgoNPre1S277uu2nUbps/UFUV9MZpuRE+ZkGJJs/up
l2znCkM37MBc7g+rT7e61JdP+qtekqZCXqY9IlPLPUUFLHR1li0/Cyx+n9dHP5Kj
SSdbk07oqIKGUazYk21T/QNtLXI9NTkUqBk5XX472E3C84XZflvKhCiSeXSVwdUX
IHGYF8iZAuNQxDjAvkh3dmD4wIftuGW+1912SCsyX55Mo++Ftl+OPU1eMY7CWNZc
b9BtkEIP8hWNLdaHBa1j1zw3jTbfYE+l9mNC2WOP+cccZs2U9Op+uQH04K8kaoM3
IPmRkO+qN+hfn+NLYSeuoR6O+dFYjP+KIVLWNwtFSp36/ZLfEH6lFJ+97jW7yTzm
JXOM92oGkOflrpvfQOxr+Fljm1OVmnGMb4YzR0eNOpBOWSUxfytQgB27DLb3Wzue
ChowG8O32uBZCkV5GczZtjTGQ9iGJ6xmgUDx4W9YuEeFypivlndPSODQOfA302rC
lU1NlnQPeGSuohBWzhTDIu/xMi9d3aMZwcXWM+r5BxfNhc0CKYjJhrd9cmsbverJ
nLh68rNzTMeETHBCw3VGkmtMWd3SMbqI0TzPpJ8Cjp2izzvFWSERE1zTdsL2mqvF
p6V8RV9eZYl60EFqNHMhRdjjKHazwQbL795Tui6Mul90eMBnB0QFW7fTSBW9FUJw
UQpwNUP1AOg+4tDsfDWs33+Shjywzj53T3A0spjRO5exvhwn2eSWY1VyjBfKe59B
mtgn+sXPlBS8JCc/PnhDPy/BRUJSh6ki7QJ0oKEhrVVZIU5MulG4hajYypDk24EA
EpmM/WjHWOSGb7vUB4WPBKAVDoxLh+lEm9WuKwS+oLCbMRnWKCSclwOdpJiT5Nlf
JQU11CWXGp5cMOTdhZntXi1XldWZqxR5Kg7jtO4W4Td9VvLnPvY4STDt6wGvEBCh
1O7HjANTh8DIYX1ycH2R+4xjxDgBlS4RhmP895FwOi5NIPBoQrZwoeNHHL5OpMd1
f5k/QI/DK78Kuclvxway8rPPgVFhmuz/fRhBKqR2o9JQVt3UcGyimjfAmBQTOLbl
dy2cmew5g8Tz5sVSUpXfhkWc2MGiX3qljVoQA5yZfZwbODCvFPN8muCHM0Gnymz/
EXaTh8wt9HVeYL9JyCYS7eibX+O/q1hDSdqfpLzV7AggUA98o19rl1+BLOQct4c/
Wn6+8eY+D9BASSYn3N56iUDqjaUvk8g2whc2IoGv2j0CXrrA6ZkGswyffUahJX02
gfkwkD7CO5rSgGvAK3Va4uCnZgnGfybTwu2L4mqBTrrrupmeGsiddP2oMnGS65zM
LzUtJ5vAUtaneDY2LFoqNy7hy2Wnhevef/heq2JvGuj2+olsUcHngGtijPomJ3KC
x9e3XYI0q9oAYvvqGvEXtyXk19Fldx+WanYH/MZpvXEuofuirG1aGHSby+Ci/Hll
lM9IUtLRpGI6XY1Iy5ercK/OdaWglOsxatCC4OYrh8wG2XBZ88ccwi5CWi5guzJv
HOrctYwIj0WRURd1KdhLwhsAWEOiYbTwaQMuxLfCkAPD7ruy5mVIQamSKFsQKw+k
Ex8scxx4mab1sj6mSlCZ/nAyWDR7DBF9+mpavr6GXGKJuPFn3uLpWd533Os/CqVG
MpnxvJ/lk44BkM00pVNENDQA1lwpF8+d1XFt/bS+wZtS4xX0lYCU2XGaekZD6+vM
L3YK4hvziI0JK5z0yezmTJPfQhMA5ovuCpCqJddtUGS6QHFyMdFBubTHcY/3vLxC
oXb90PPVeaz3bnElhPuTicNpargonoOOS6ypr7SHEdogjksZsUmHQMrWoUie/ufZ
5lgiz75zGnAyWf7AK+e1aSmrlhS581hwH4UOwM0kQb9S6FvsMk4GtkChNZGNaNwO
e3D0O4VdDwYbSBNsUByGA09hx8J3rB0RBzVibO1wAUXeJ93epoVuO8nqHqrDxSWB
hgtgGMzp6kZjvdYRMzLTcf5UT5zubLDE+YS7DyA2xPrr6LNeqEcaW2CV32Su+4tG
CaOouUKo20VkEzkkBcrQBDrlWDqQao5ZDjnsVJtknOhVZFJ36lcMOSaMBjZyNvEt
P/Dc02yw1qg4j19qly8LcN1dvz89Eoes3lMzgi/nKVSeOizsLPm1Ov77bU/wPp9U
dTgPyBYJnHTozJ33IqZQtmqZ5IZn2DJYadTb0QYmjtz11CvrZf991D2WTra+ylEr
LENrY+jx/Ymy8s34ez6UQgB6gkmO0Bkplh0nRcQ+cP3EzA8pOxdcy9kPc8TL/G6J
MK5rmusWg3J5mCkGdyhG9/8soSDubnBP89uzZY+gapA1YdSajjxJwg0B+podt8kf
gyWSscbPvDBQ/4szWLYwBLFcjTWs4/gX+XSX0piHB6l4E2//RXznxmPq/CGWGj6j
eUxBBgexP4B4B0t7nWp8C2rDvYinvIu7v63VqrnYKfCkaAOdaT3+TlOqar/Untyq
z1BcmgZr+WaaltYIAgRanFFSILvBqe29jua1amSpMUVyksp16488NxtyWOA8vMEG
3V4n0YQV733pH2TlSBODdW4ev/lFjBAPBoSDivQJwKOre8mxxZ9jv+pIVxQ++wo3
kPhHkv9LoQTVIMte6iDNY4lCEaJ0Nx6wNGznfwgOdab92XTPxVzlAxx0JYBRonWj
J/cNSAco4pknnFn4WLZoZbqNZnOJ90nmwTCejygv25DsFC1UGdLfjPfIylLBatW3
5cvIZtwCN5PZdbkPU+6T5TEJRYkYoUUMkP/1ChNaW33Wlc2L7iSbR7XceDPQLZk2
WdK1pZtnqX5L6Gwt4QJ+tKpW4PrRKlUVM69Vpt2kOhP0xOCoxbXbmL5eEwsHww3Q
8pZISW1T0C7UItf7yy/lpFsxMuCFOkuSBxW/J70asXZDAu2XKp08CTYS5LpgpRpW
1XmRsvyYx7oOwRuWWSFJ5rEygn+D3aB6U1Fk1QosbIBQV/BSnPQfRbXf6Nex0E+2
1hED48M2D4miHc6gl78bv1inbQPoRZ+LDo1Xtm7wrL2Sjpxy7n9TSlDD/IjHQ+FL
DrTx6L2mcikHk47zA8SFGrRJpIuO+gHKYHPx/D5s6QLEQANyW0Y+pxckbMEz6QvL
Gf/9wBhA8iUPnHBzIStw8ecqpF9/yiAuBArkSD7Iunar2p1/epVSJF9wN5In+hk6
gtxsnKvC6ryWl0MKSnSWsZNq+4xeAeoU5WEkQGui6aoLiYFm7kWi/Sd776q4spgD
OwBoTtibhldvn/XGTcekAZyeGAVwhvIHR6ZEB05I9UDe216ibJExDLLJSGTfL7HB
hiVu268DC2qeO0ikIMfNoc1q8nefZH7OUMUuSfFPxg2K0y1w0gWCFGXPVUJZXNOk
RnlJiMSakjW3MvIvyCJgtlXDx3Nzvey6p0MTfwWlBoGhc/lmWbV64cJIjPNKHsw4
I9FwpDsYdJHq5yv/OC8tLIXjjusVGargtTaFOxasWK50A5W848P/CLdqrk0Quw3Q
358yIOxyY8iBUc+MWVTFQqaIS3uXSvwoMkTCeRyOpfu4++/fn8z4ZBZPTVm9AjZ+
0olYSX1iBO7kX9SH+WFaffYAN46UCrygTaTrWCr5gv98gnQUv+PXohKfYP/XX+eb
nuXASUSKWNyO9SyL+/pWgMd4tn8j3TgZGpTdmhI013PGCdzr3vWejj2+2y7gujqU
/1HnUE/H5quvzf9MJEl3l0L6/AzQixRRHfaDsMHNP24oa1J/RLTR+PDoktCEHoHL
ZHMMDKyUGGWScpdXrV86t/WWrzPfm5VpqP5lgNwSAyWTcEmJBmnF7YqQ3uOQZu2/
d/+4IL2g2ISz54gjMUwJ/2tm9xGBazQGi24lY6Upni7g0LkgCZU3PuFHJQsP8RQH
UKv9jX+oOTayTrK1fRUWyUA0JOi0t+14OYU2C7RUtFS9r+pWCRJ1BA8E9MF2TOdQ
gyU666uQoIzXviwdRyKoWH6qOk4GzCswwYV+9qqDPQ0QFJ99f4hoI/U7dYnppvWC
Hbtn6HvMOCmksHwoz+phQIC+1DfRVAezMVs3eYLlinIRbTuWdVvbStbjgQvydygD
+ro6YrLUjALbPDX8tWg0rTXHYvVLXemmo2sfXsxfOqRKaYYLC2rTVshbw7uHjTCL
lHZmiNSrXdodsCiOKezECgQBjrGyGiZb/PmriVuZQH4ZlGYagCh13BnIb/8M4b0P
54QPOLOElboDpwCc1O4FTyADsHVR9CLQJA5v1uKyTXbBD2QftagTwcai0tbVYkHe
6w/ZeCmLpqTAxWWcyfXk6vK/SWtPtLYrXbwZ4KdQ1NnerDoFtSqeCfsoLZCRGDH4
aPMWE04G/E8Js0d6olfoOxSJyYNAjpHIaBbzpbS7/pi2LVnW4deJ0s0oa9pkGeeq
c6Cq31EZsEOkv3Q1Kx3vYWXL8BlCBKvLZdKCAuGmQHnRauyjT6mOovcPLY6yIydG
6U86hy3CRNUZTjnvJWfT9f0RG4MjJ3FuRZMnTefE1vB/3zlXJWpikpsHAO2VLLx4
fC5MgD+pSaBDiIZ2qJ66aA73OZCVYsZApzpJCzxfOn1z8QWRHct48CkZ+VBAmx3l
ugAr9H8Bc5RNDyep36cuVQFVjxPJUiinU4QOU/pEGvD/Z5PQDxFZNzaMNmqcWWwn
P1XObRra+L1y6IhaqimfhxgpR51/NE97bJN5PS5WzudpGQGxwQjf1LfzgH8UX7LA
kvf5JAjzT97hStcaoLObtzVM0ebf4Y/Hi5SYVPc/SQmd/FyalQZ6GI7qlntFiPs2
6ob2yMjn6w/1N5Pa4MS5lQN9oARGOkpn9bac0tcK1ylA4tAfgOSQdFpMX3G+3ArH
PsO/Y8e+EQZDLnGrmYPkKAZqO3wH1LLx9Pb9l1PgS7wa6SSowgCwcyB7lqQaQ6xO
zQ0hb5dHPVaxdFSmio9+tf2GmdAvrbyDNb+J6JSD8xFtE+1EcJdc4Ap53lK7W7mq
TwiDnPBfhh5xNE0iqdsQI1/JeqIDMCMyvmnwWQmnx2q5Svn85sZYrq7qeto1b+Qs
ZVJ8ZiuD4tBftlsgk+oPi9gWHc5C1mlhmRTzQBlCYhHbE4qDNrowhulclkdKMQl5
0ACocibbGQmto+it4fyqUG6PBLf7Ho5RBdlr6OrPM9uvHkkdCUSRE9ykPYnTmsh7
7Oz2czJn686XmF82SCf+yaPyXU+eN2ZELl7wUcT24z5z2X3FvX8aGRO6JLiG7N92
EM6TAbMN+2cVWUj/ZgmYci1JQfBu9ML18G/97z4H1fYePxk031fzUOvgvdHsSDmb
4c0PJfyShlp/ZqKmnlad1dSggQJGpa1u1dAPaVz4yO+Ne4iXWFlzTdz6Ce9u8rm7
CtWogxcPKGLfb1cX7prgXS1WUCDxp5eg8AsdRtTB69J2WfnX5cM2FsWPBZQ7PQ2J
FyL7E7abWBtztXXGQDY7qBe4oAavqV4/90wW/9/MiJ94zTPan4GLnUXR5mPOn+kB
SKCk2OpmkW9kJUB2eHTkL1jBIZqEeJkVGHWSiPahuD5S5ZrUL4Ov2BGW3CqTeZ5X
l4HKpHJuQWovoBP2PO2ky9xKDalg1udI0cxl1ntxVtyaNjeP4j2aUIywYPfMupD9
UQY/G57kl6z/EP+pj5xUWolvXHJsRkYuq6y1PvC1W1HMrkByk0MRiKMvIhkvGXjr
rHJ5wwr7jGRm6CKy6EsEQhrUurqgnyaq7q8hPq51fSw8D8JVMuP5TMDczZerhTH+
ZvZ6lR+Wn149tBNYsQGmtUjg4zEZViSgqV/Kv8Tuml2oqDl4qsV2ETcDWPzWnZp7
VBROQLumoTQmCPhXl1QbZ8t7owV3IMW7fadsB8bpQZ6qlrYUh4MgYrqC4MybarCa
DGdf/efoPsbeaSZJ94HlkINUBafbY7dV8bLRvCougAmSt7wVmkqmEYy/8Mcgfti8
lzV03UYjWBJXm4p+DblglRCYZ3MQNrL0YlHib6yVnVxWmjyC4ePhdHDxBbTWGHIe
bW0Z4XWhay+N6O3PgGVwEnIenLIylr92fgRfiiJbiU4/Lei5Pcyf1uSRY3HJh534
r99sgKijQdqT9O7VMj+K2MasRITCD+AkIBkQDWKqVpMvkdXbBrtduiA4Dtqd9a+C
EDK5u+BN7euoLaBkQVoyhEvVkfLuukdLlz6FZbLaEkNC0NbAzG3G5Vi/ikZRZ3HQ
kHROSgqx/Effu7pbGldSSRqgjHbEc+GAXysXkGUCbxdpIReRELTmMS7kp7z9DULs
2FnFuKt4bw0jf2wHriBK5UZZb125hJ7HWr4KTpCvV/PHEMmDF8md4vT8GCIaXbIP
PQ8s/yr6ptX4J5jeWt4mpMT3YmP6ntuzTIezM2eEvsLrKLtbGUh3F/FoU6iG5DEH
RPKEHqQM440OqBAKryNNs0hHKQdA/shqRm57DxJE8vca+NlRv9GrVC/MAGTbg/KS
h6Lr2bKH21O/dNfcPb/bGKHttbtD65tY6JZdQ6edqE7TvYAVgifcbTeTHsP4dPoX
acUyNvoxrh67Ic8MChaMjedkb2LckXJbhNDHvmwSnaqm5/dGAQwoT22/5HQ1LkVD
lUMZ52SzWTRO7ulj9jczAX8NvuuQiDpHLwjpl2bJC1M4qRE/F0QmHl/buXVb368Q
tRFRDgeqwZN7vcugcaUS/81AERemsLrrgSPRNQ/4R1PFnY2MbxobLA4N9dFZApK6
6lLAMMEXW8VswGh4NBd9EnNspYcjSns62eFDsiOOqLTQfwEnuwg1Dxuud6WzcYOi
RPl3qNhIPjg8us0PQw10WNCrEExJIra0vuuA66j1fIYfq5l2/v1WHWqq0LnlmIeV
b15oNezsqQGhEHY+gbNA14lMR4LGfO5MTsud5r6x3MdloMMs1f6lR2m/3eYgVr9n
+cnu2Gecr+7Z0iCuVJN+8d1rNI1rlv/tPd69xhXjOroDtnYr7vYC1i7EC3akLQ5i
j/99Y+cqmayznKZX3l15hmoEZjFtTsERvjQC8AYyEtr3WuO2suqHSp1MsSA6FSAF
hxZJdSQRT0O8Z6k7lARUPgR1qYMu9Jk4sMRIf0YDlR/5rQ4IUJFoXQaCCVbwySqh
JYyM+Nklf5EMAueuQkFMvMJUdGfCAnW6Uc9L5OgGEjjvIuZUxXHSQl7zIUAETfRI
TjKDMpDjioGkEc1uRT4nLKhZYzzH1X189WyoSNwOqys3t+dq0ovGupEy149iwrKQ
2woXr2ZirnxAAVKg95fIwz6hl2qQLOsScelFN881MGmwCU6ZlnZDZmFOXafJiU+y
6BJfNc0JBrxAN9GSaiIKEicHfVlYhIgyitdQrGncY9itfm0tRBKzFW2tmHbJ7b8J
pUYkZWi0k/Q12W2Rhqvxdr2M6MgGVdqzuf31prBolfkvkxMffajj6WYt5DL0nJQG
Qq8lnrfa13Fm8Uaoy1NH8qVA46eHwwZZW1PkuIvsXe0Qz1Ho1s99/rUfsW0T9giB
/GYEh/UlGXNEmRGhS9d/eVzqjUdRiyFZfvdw5UQZq96m7nZnkWN1VVrw4fs7ielt
jeTmAsor1zuw9u07PMGWayLxsRM0vYlf7mQYGPm/UVPxp9vhgXWFDp8XL0fXW+2z
VF1GhfMKEqkRpKB9JcmBhF7M4dMw6uV9jQOoJeck6MI=
`protect END_PROTECTED
