`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SsUKpb2k1mcLPcDyAVL65lb3EhwqCCifgQ4wF59Osq8LOpAiV+VSP4iKTOZrR0Cs
dfZd8c0jHbuD9VDQmwOT3JBI7bbCi2RP4QyDu+8fGKJRqfP4T7z6faHUJ2c/8Onz
CB8cqYZBygE7aVu57yJH4iz6QAN7yx7wQEQIw4G0BiMjBtKgqnNhjC3wlhl6K6bx
6FqWIo5RsHVimCeuSZnbo/Kb+42OKIEt8GHq18OKpTjcQV8BHnByQNQ6zHvAvnNP
35RWKPRRq6xLwR8F0nwoXDxj86pjU02+Y7pjF4Kr8SfaWlyXVBIkjcL2LHSyYzJs
GV6+vcypnjrqfHWUjmGuox9cIJFSkzkViCYg22T/L/zhO2GVo68tdzpYWyuokGrj
`protect END_PROTECTED
