`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xFFjV6ZlOPkQibXkA3sLz3apNN3mTrZu7QxpsgnHDx/mEZY0+tmVbEEvU3d54LeA
YfCDmiTA41/yU1fFyb67xEG+esFFKL5W9uPr8FzJ8si1G3232KgjDkC/a3jjpDWI
WRfn4lQA33i7zp6e2ijKJBj1frbCy/7EbRzhQ1/phwYh3jXJy3nN3lOKfU0/z5/l
WCtMw6rW0uYaPkUm5cF3LopGVJO/qGHLB+B1YTAqTcRPKeLP9jzQJtsC4JmEsuL8
x1Y+R7JSuYjfWWCHiO9gByygiqNH068vqzq1oqlVg+CbaIpK2SBcCPl755p9puoN
7MuzaLghaHVGLBSLx9e1Eh5dOBih7/IHTRlhl+Rz1tENsY+VjxOGnFARyOlzJO13
WKv5EyBSHfYBD8mcrZ0+WjUfVAjFNlNXcvhoWgPr7De22tpztn0ENLdo2VyuIMEm
aRgYrT/UXjkS9CB+k38jX7x7bsClfm81VGJBKXwrwC4+DzsIwA/xhg2EHNrp+0u0
`protect END_PROTECTED
