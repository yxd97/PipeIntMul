`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
du6gX6fudU8u7tfiV4QDMwAuokPcuGDIArgAb0eKgHTib/AhrTVl35xAO+WKiCi8
SzQ1zHxMf0/cLDSyeMyfiqrAztwETf9plFKpBj+lRCK2FC5RrhGaf9C51lE6I08T
qQ7DvS8krbpIBpSuY0X+AOtg4ke//LNLyVDxjt3tsz6vatyNTWXD1DrPGioXHYKU
YV8OB4KzH4/jmAeUdX5JqMQamZCo4zhjMZSNS5OLLrffl5C4WG8qDjQeFfcAupCJ
9a8a1NX6Ye8tZnRY7686cP2ApKVsh47Jb8wkdQZgAuAtWvBTBcvDHFGNPT+1GhMB
/5g0Zys9KyVKyyTKjBUgB9o710MnYW9KasBLxJgSyoEQfMwOYo7v44xXIavTQUoH
`protect END_PROTECTED
