`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCBOq8HQP0JKfkpXnPXD7oGCXYgb0h/ItcKV+SihkP0MUVW/3xX9CLj1gm4pGgx1
zKdftSLzrNmNrvB2qHttyVh84efqXaTGY+68DpMAlg1R2d41qSQGtsAEAGICIQ1F
+cdbmpFcm+OeNw/Aeh88CUElD+TNAC9reOgXR/lkH2+Ew50ucjoghJrOl6tz7NbH
SinBveP81zF9jB4hk8NkUH6SsZ6+BHmDL4Z3mAe0upVgacUwyAo2SRZTSZ3Ba9mn
eEJujoPuxSQsUaHGGeFeIw6+ZpWy52txfwbViRvihVxis34t8e8XmYDfq5GbsHaG
rfSPGJaNnJd7Y26DSNiCgD5ChfpTMd6s6TorS4cbV+4B44AXU3xZlJ9++txmbeMr
IVz86tmUAcvfcb2t5131vy7PsXjsSCBsmgSem6riXKPFvlZvS8RB9LpdTqJW/I+t
NV1jorHoIPD5/qwKqjeaZfEF6IBhS9Te4hvU7KFR11dGPl8tyZgHjJQMm4L4LyIQ
RMBpovq98rEPdSqF+nVjcN9NuifzuuhejyjyotinkNlR1FO1r2+DfKA/fCte0Hem
T6HA++Ko9J3f2UJEa4KXUK8D+rZ+MMEf0Ktzqaecfn6/RXkv05dJraaRu+eW7hlM
KPdJbKRjS2+dw5wIuJC7tV6p7h7+D5QINslhAzUQRRFO0/PW2Vhi4AC9XKIeDGtA
bF/Gqt1YWyJKAYFr/BCg8qET9x4yPbhlU4ZnwbjIW1gFdV1Q1aK8DO2lxAgKHYSw
wJnoSYIcqof/jMVHawsbO/GRDtCM4gkAqZsm+cd7NQVQ1vQiIfUnvTlPZcQsjtaH
G9PoZ7OS0IlojlI3haUJyRpJ6PnyDCiIK6u5Xx6k+RSm9MyHOBfHO+r6sY8yF4+e
H4df/SS5WApeVGQuzWd6VQu0BKAEKYa8lS/CSjP0DpWHBnreFGNjgpdOXbsKhYhO
019G6ZcEIlYs6lVcI4ItYAxB6uppDVw8raShbAa8MVVB9ShrMlqvd1BRCw1fr9Z9
EInIhUesP7eJIXDZbkav97XWbB/fo56/8VemUIS2vuhLouf0/EbsA4iZxBkymeV6
h/Co5zgqcnCX/NonsfnY2PJtd99K/iK5vE9hXDwyiOfM0TxNJ2j+dOX+h1sDQGqG
DOrPaUr/XifZd30I/sdZUqxy0YAMZNpKzY5ri/NL5DvPmXR0UUuFphM0ul/9qbaF
YULnKhusr/27uLgl5IpzJOlX+2R5bxzSLDSS8tUHaADQ5gsf/pMErpk7JiTlIky0
FsqUwNizSbp9ftZdzLUgqNv7KA0Ddm/lhKVzYdQadi2wmr9kWAgN/ligIPRD44hT
mn3II16kN8KSvamTNEePYkKCjzZTqRyPyHadG4TId22Ka3KwJ754l5Vjqmaz0ooq
6qAyLGvMt0qi7SPPrPWPYRE1Gg1s1GcFItWlQeHpRzWsRW8liWSKiPlXMrgcRUYO
QHe6lHRmPP0nkyYglwXsBTjAAche1ZbqPkHbmFQpIdG/LRpHMQlDsBtCBXx/Pwl2
5NUOYxa+0I1B12fug+njYr7/THd12kUoCf3m1L7kMSnsBvBkXLG423TGInSYCnHz
+iFR7tlGP62v95b+CwqsGFx1pp149DJxdtXN0ItsY2yANes2dXxCHiItzABIRL8m
s3lwxhDqA+2FhVOhaXWVVX1oUxsJdYUqvMT3m/sIG+1FWoPipvqpgGyIBf1hii8+
ykQqZLv65Wv8+bK2mormseKKAl906MDxWYtaQnXQ8t7hyz+Lh8WtiUBFDepDs8Zm
QRXZkMDsCRJFr62gT40fwhUQDrYd5e3wolzW7zg1enLI3m0nRed2rLB1SkGmdRSw
hoKqi6j+EkbzwVMEY+8NQHAHHl1156NVRY4F7LIkzFqjs6I8w9CWPgqyWH2wsUdu
EpMCq/lwDFcy+N3NuhhLp1VHhpo2bFmAY0SDOfROthF5D9hQew6UDWkPV44v0LPM
RruIruESwU8UVkcCT+JCLrBJ48aK6axDct0tIEx3/TsHh0cqJBotjcS2RrIfkzZQ
lO/z1RIL1OMR4JaLj32EtgRBKr6M5aZTMYZ0AmzgJ+wQ88qTbrtOZsrPGeLGGFDy
hJSPaFrYWyrb2YBgLHMvYeiP2pDACuGd5vveAY9WOG1OsgRBEce5WIwPJWqvxyIs
TM23eC7bw0uGZfDiCXMq/ASXu97Jwk7dbAtZpfsOFG/mwmuucBv+VAfi6AyUCi53
YM8Z7dhe4HrtSAXxFUSHX+Cv+0s1sYZtiWj7S41/xnuPYeR37GvczoDZen7ZRKjc
oM5FtUl55tpUUx70vDy8Jj1J8XmzEPTghafULUCoZoRrHiZo319TLBboY9QR6RDl
irKlmadgPTf/wCWYLeWDA3fdDy/SNu0IixaF3yNT5HeLN8KcvgmgkKLncoBhwht/
Pq3seG9Y/gabNlmSVfYxagypR17vcklNmrjhLMTIbdT7YQWFvs1uv4wGopq9XpMJ
3iZocv4AHCp5azRWVtgbgA==
`protect END_PROTECTED
