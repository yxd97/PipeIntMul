`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IM/MiSuKEOnyH+dY05NRT747yV8nBS+vdNKEy2GXxUvxkMNnB88VZ+ztYjKfd2zu
qXnIEdmJ9xFAlOTHDkrOSuyMGOAHOo3Ze+uEQ/XCQV0K1dIbiztJLmvwKyb5Hf26
FftPSd7purHuAwbLZQ5bD8kBdBSYn/j0iOOBYjpIJxdO4CihfHzQzR0G+DWEgBmQ
LUhI8lgRUp+RDQ0WTa0QpopVoEXMkmyjfWN4eoVcaUmyiceI21Cjnbp3UUH8wexM
dCOALEm440fNxvGNBhZ4jhvRmzMQToo9hpSM+f/3Ima3bBuISICi4ZGvdSjkh9EQ
zLB4lfzN69meqzEXNtxUaR9F3sZ9fLTvQsk+L9JcoukT0a1u87vNQA7Ecd7Sd7wp
EleebjbAL1YnF4TS5DxjuF0jnyGCnHENmIbLIa+EpgfqZDCEHXfu9B8NZ3Bpu7Nr
jpdaAedpiYHQGMNzGku34sPJjwhEdcSs9UGLyNSy6vbjIy2XZzPl4IBv3pxmikrA
YxCQq/EOVjk53DAdkuhJIDDIuBvKw8tiHYSNO1I9Zj6rN8pwYadzxRxOa/i4nfZE
9kDWJAKaxUzhNrqlrxOu1W87f+q/rDKbVdYU9eXNPgY=
`protect END_PROTECTED
