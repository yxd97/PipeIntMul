`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+sX7qVfHjzxLiVzfOwwPSRUyslz5zYa4gYO2Ufhnh6gVymsqaTOb+NrRUDMlxa3u
EjNAbiUXhdRU5FB75uHfekovlpLnoo+euUAlhjDeW+18jXWdRWthBUYH2dddzJHR
KuIyBUh+Z1BmUlei+Twm3X+Q97ijozK3JG5tOsuN7nEWGMMsDfZHdKi1H5CvrOXG
1yNvn8ZDIg2hOPkzxJPK/bkKk0UHvAg+xmi3Y5y/urxIkcRKSjnq7odFCabOge6f
uL0p8dNPlhIraEuXPNFFdUPVoqHe5AdCab+b43fVLUEDOl8JtWWh86AJnC8GpXsi
QlkHK2AA6PX7Msof3CiaO1hxVkVxmZ4g4PNfK8N0cdRbl8JRfTy7gc5FbqUO+GBz
ATWi3JxUT/vsGXS+9gBfuOFizC9f9gUNFS/9yo+b38vvA8oQvfBHlV85HpUwwlrH
eTs2ftcJ2DCXFOS7m9xd1B6oMZ+O5V766MN9mAuVpi3kjLq93VjpVKkGymV/Lar3
pjo7Mi92R4f1HZ3FXZm4tjlJ3dChj78ndIJ4Q0HIsx6buST4ihFGH8+nlHMi50+5
ybFNCHh6lJbDQv0fTfJkCBE+A5ld3YH8QXssTGTHJjvNPRuoT9JR1UbgNv1sPuX2
/kLehobAubgzfP+WzwoqcuBNSj4+i9+Drz9ZqxIhCFTWIKQZX4/ZuTrzoqIKMiwW
KfKNMVAs2kS/6uzkyh4ktcgDvmHrfvr/gRKa6r9RRaKxGuWmffNKzJO8OKKqFGiC
OCVGqG50XyZHnLF5LIk7MkerCn7IUWPHIND/8WXosp70jid3saLqtID9830+VZw4
+l+Xrn2vjLaQH1SI0aGgPwDEOn0kJCaRAO7D14kX6buHXAaHZLrXZzhYahFCfwHG
8RwzkcVi10nD2tsHkcPuF4x0a2876dsJANqqF7UYA+am9soPf41BelZfJH/CJ/Lt
QEgz3rhzjii1TD48UzP88bTnqm/CkRMK/ondqNb+LpjXROj1hE9BgfVstOSknDK9
yBoT7U2MytC145GDv97TeDDSB8IpADzDsyX4AK0qOf5TUuf1cpUnOLxqnGgPXnj6
gsZeSfJ+/siHnXZHG/kV+Wip5OzvpZMZ78glill3w/JTVMFM/88FNVn87FpPoVj5
PFhE3Sa8EAPwWisBEWpC9YVft1C/g2xVDxvrwAhQ7tQDn1hECB3aCyK1Zqw6RU8U
BWiYLRsAF1RTofQhrHFYptXgDrOuUjUQy6p/KgviP+ltTXZBc0U9rjNwV/u0QH2p
pCsxyOCJdeSKuSS5PiUlSLnLt/MmbuQ0XSNsWiqeIOqgISfoyIFq5sx1Yd3TY84b
A/IX1n19jYg5nw2rPGCedKvC8khBj/oIptM1FtXVetMkJvaTPtjzOB+sB8javjsz
Qxa0HMd+PYd372Siqlwo0S2+pEDoQzTk6C0t/FlYsZ9qhqwPMO+DUDuaP04BfCor
Vo2vwWmFXUYMKPcTab7fYr76xuaAkv1LfgYrRRszn0GqQEsKGMb6Jf7HiSpFvY3c
MP75AMkPt8zIlbKHhvNoEXi6jTQSHlTwCTz/2CMvpw26QyBgteUDEdzLseTZXdTn
Qwb62C6e7gHztR2WHtD5R4y2p1k9Hb20CpHn+iCHZFPYa8otvnvvuKuPuphaKbDb
53YugaOwEIT9OvHB/FXBVLlVMJfAzu33EkcNo88sixlwLUHZO5VJHSSmi0utot13
3AFXPyULDSV1Z9Givx+f2qkCW3HyQCK/zRju5jXq0CV5/oadSnnAu21Ne21ljP+R
bgtSxEcieBTsw7CiqcTT/Q==
`protect END_PROTECTED
