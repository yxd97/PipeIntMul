`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QlcbxW5ih+QDuDZI6zwCsA/8Oo0iN8xRbEL+fkRvVJoeoFonO3Fav50hv7K8o+4r
ni1VyDTB0uNfiL/LNU/mxtUFCz5bCajYNZb4cY3SpVn9d9iufHvSEhAOJuyMtJIU
CJgl/vidDQWf7DESXo39wDFBjihrY9PBEefDlVExiAzFPpnMiKv1LbShLjS9lLtv
BZtRQ7ulf0s48NIeosabcwAosDgcmkYvT9R6PVS7aU5agS+SSMZt/N5PH2n8ofTP
OIWd2CXWTYecmKSCZwOfKcbvRwvjzVAkrHbMBmNbVPq/+SxdV19zmsjHeldH1EGW
RKgx08NgP/XSKHNOhUbGEL9DXneA9CJXXj0tQKmpL83w1nnNmyrOMcP4qWZcnGzv
fM2ZTbeSyeJu5nQoqpNbBm/vjD+kEizQfW2c0vtyK1a2nbAOQhdDh/+LsXTWBgdg
EbHZrNf4LQ5xHENFvGj9/HreFk5qJjkgdwwFyuSQ9gPUUxbzcIAbOrwwNRrE7ctl
5aYU2ynBU9BV6uK4Mx1vnZ6OYaRrwfiBcH1VxcsF3d8Jbxa+Xwfr3YXtOTd8sqNd
4BtGYHvg2yFXOvyqBdF7x/TJNLVIGa3BKEq1mOEOBPpNvxvamL176uLGrBODfS3r
RJPSozHFsNC/jYVX+IM2g0YnFr5zEAltNsp9y/QqpJ0yP3nGPvHGLY3mzaVMyHiK
HgGqABOq6nQVEophVPifk3Cn7+nFdovft998YTG03picJ5ud3c2/nY42fMp8+YBB
vtl/fqU6SdpyGHGppv0ssc7+nin30Cp52JBZm5CeWW0Dq1IN5prvy2ttQCT/V2WG
ICT6R2H5LjTkKWuIQVsXng==
`protect END_PROTECTED
