`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cnfZ2POPQ2Tq3SXRzjpJE9HkyipBqLtGYfXbi/WNpm4CVn4b1wGBSFtdM/ga7c7
nn7rWizLLHPj2kXSuZgwTlEuUg+8Cmp/AAXo9PIuVoJFcYolsFVdWpygYqKfeRlf
weD59iKb4zE8ohN4v2OMBPzVzg8Is4xF8MmAgr2r8aQ/ebN6qhUQ0P7AyRn0oAA4
NesMHbQQrVWZadxfeHJE7bTE+TVyfcLvhoNIGqxFeaOhzfaJPtmLO677COM/aXRL
GqyTuXE/OJQ+sPCa2iL4B96PDxcKdb/D2RWk61Z0LK/7NjKvZ+g7e4gY8sk18odB
COocqr7XJZnNk0fy8JjH8m9E7Cn50RjpeWejyM6W7rbvpZmF8NqkqoLWZ4ryMu3u
04ETdD+wozbeEI1tLJ8KG1OY+gNWHfRGrh7PUgUzAQ7R4v8SdeGWqDJEM5A4acCS
CPGceTk5EqILn6lx6amf3jEKLnDlNpPIkUGr+VUa5H9wXI3b6tiiJQLzhysSnSH6
SW2LgFMaWFZo+9+6NdKEyvISSa1VmLLGz9oQwabhP20=
`protect END_PROTECTED
