`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHMRNNpVKOx5PUYbNxu0jHFNz2Z5U25vw5RGcysSThWpo9J3uIXv0c/jIx8LDynD
MoE+6zXTaTvcdheg+pm8R3Un1lKXKj8TxoYTBoVS1tNypwdXbS+qCrtD7Cy6s7pv
xPGsAoehcVVPhQhsdyZ+64xuQZUTKnuHyshDM7UekOSvYJhKNYWuXhZh7QnjL70N
eW4g1UffJFp4y0S4+MoMkIfYVFvQWN06ufOcVWJX3d0LODHn2+fZA0G8qjVdG462
S1e67KtGIttBlOKAPCgD4TS7IE1CGVq4SKzQsOdW6D5TdBP0cvP5LpqyDseWtuiz
kPbaQQiKVOrgGvzgbLnjgdyrZDja4A4UVx3AJoh1WvKpaxEQlWqiOQ9QEgKgDtdi
70HEsqGOdZNn0ei/PECpZ65K/9N76XEhV/rRJgwDpxbkMz++mIg3vssajQP66CaU
Q7EASBcch6nj1zlzRtxb4L1sBjxF+B7jVKm78cw5+4ZmW3MukMD/SSB4xeb53zCh
ussNYK9xhVOdj97A4+9p7Ai+VGCCtKtynJ+F1q9XDcadb311f5UAlMoKQRiJPVAN
MXlrgEcyrRtVwPE+XFgRj9mZQdvU4uW+fnmSQFqIv8o=
`protect END_PROTECTED
