`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xF0wzYpuXbMugSx8KUyUaO7WRTeyEgV7kkMGFQ4ZZ1Gy2dX1M7TgKdVYi2vdWXpy
4RI83pFvJ8z9gZgSTDipInr+hfwypEDhkvVbNaTnwALCsPtdLMSGawMK9IygN2DP
3N++/nsc2FCUFksU1LR0g+UjukPaAhaTUi3Y9IhlUzb92SPc8p1ftVFxQX7nGR/4
+Hzo/xVd6OVzExQty2Qn/lKnZceMx2fVq51+W4Y/Hb7AltlDPFYdjmQlc1cimtD6
wEPopDGcz2JfzvGxACtEld1b+bCZjepV/y8EQN0UnPHb7oriQwq8ifi/qvWfAI8T
lwuku49+UlkTe0Mgj0jmUkPsH/vRXH1NVmOqEDtgg3EOjfRp8Op0AUC7JDX751DK
F9eRddOBz7ADmS6knMvb2QncluCaldEH56qISiliTW088eZnOJkj/w89zkE7jZnf
tjm0kAIunu7rA0sXw/j0B6/idpHNS7cujK2n7hV9pcgGzVfTp95n3C9x2TBnCFBH
ygO8/tDxTQGymTKSMq1DNlqiQ9jQnz6INoYerFd01gR2KB+o0S40r06QN41zIASe
9gzoFsuKDwarrxFHYaS94wGdbSYUg+QtxQ94DMwIvQDou/+4X0SBu1MBbfO2FCfL
vMdU8fxJdnM4kBLYMy6E7ZEkZaNMllBrwGOGzSFphBVZEP94GStOU3ENZ4jAf9ir
vx+2zyHyGxY38vsZEpVvwzqQJ/Klmxsx41fAT7I6KlonvJuqwCbML4EIgLZcFkaH
aq/UHFkVcOG7n642Zh+jznOx1QosylzxCGm/7MbhVL8nysH4F0QwTGknGD75fPao
lT5/jaqeyVT5hzBCg6jEOCtXbRmh6KaJZd5bFg9hKWqSb9LwPnmc2Y0GzmV0KaIV
AmzMeDqYG7A95UrIONbVGJcowPMKlP9czgPJDwW7K76fpTToCBZyqJ5YqoRmZDe+
ZZhJjl+TAg++7mthnslgWgeIOA3u2T6MOdQ2/2rPQoRkFH6qQlOBjh36NxtdNqUG
Wp7hGZeMf+84j2+nOEgWHaDTJJWcF71l2IKwkrjQrxSwsjQgeLPYlJ/YcwKl/WXR
LfwDF5UN1Su90tMKTIqR6/l6EgX7mKWQZOIjvne4f+eqzaD9BrlDvel8uz5qlESM
1vzPgjflsak+MtrZELbvjR6QPeYdOVMbqAA0QMb1OJCzUqp6QfSHWqrfNOtsAgx3
QlVkeQc6z2HUcP14u3tNrT3CYp4oRnx+A/Ls6SwOVQlynt24eMBEeeBF2oMqeL/B
xSDbfBa3b5JWvlhP6u9NWT+n71/PrV5geINwGFPeC4lM3j2QRuInWYkggajIJjoP
6QGbA3Ln4kfoH5lQB1ipRq8htfXZ0v4IFQDtkOLfYqpNqrOGnFuIEPdijpIkHR9O
8+jInO1zBxPBQqfQPXu1vxuzwszeh5IjbAEDlNy2fnn0YOXrE9qzHUm9dP+g0NYc
2kiYgMRYQueVEvsQhCXeX0sQibqZTYnNV2HZqDw2aW5lUz9ESEc6GQFnBxzOLkOj
ITOjyJCGyVpjPielbBGE7zTA3qb3BCr/mYmfZcO5MgCSLMZd8/ih59riTAxXRM89
CBGqGVl9EL0gRnZ5kiHDlV+8t0UzQBdKUo6lDiljHXyKcV3/ZG5i8h2AJnDQwr00
spdtwOk5VARsogya+aUnGQxdrACnGjxT22pjNSiwQXaaOLi+Tv2QA411YvgbMFhK
9aoXw4th9TbQlnfJNWaX2HT0Nl91XhSovnbM87x9iywlm/xLJ6R2VbiLLrvhgeRi
ih7sXAdEtAoNxKQvxsHrBvFvaavj8VW7qwYhBAG7gfPN04LuI0jC7VqUcz5my63b
UocKx0kjjy2is27JUIvGS1+lodN1OKgq6FCzQNfyeoS7KxH5bR+I2qLQqfqyEzCa
PeHQM8Ogu58QYuGCO8K5/w2XKhH9G6fGykU/gZoiG+qLk3LCmE/WyEGsjBuSWuBp
`protect END_PROTECTED
