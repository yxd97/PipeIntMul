`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n8bAvAGeHyAIyyHvfR8igVBNUNojmnDXB7gouuwG3KAMVjtBHIUPrWaC1XcqBVga
hdiPDml+j8hCdKLVcvtCxtkGEYCg2gEH0bnWJOKY83o28OoXAJVahz462pdVZfvZ
Sj6V/3k9kjrPLlSBcLAissI/BkqJswnzbMW0i53zUBidm+Zul/XFN6mKY7dMcxCm
Vuuxf9DaFazDaBZYUsZJv9uNDvDh6ZqVuL9q52H1KhY/neLSJSbERSoDHFF9vQnC
J1fEQ35xIHZKOKVzpsnQGLBgt5AH7p3bi3cRsTNiYL088eFhmtFpCSJfbbZ3PK06
CBsrPabHYhPpLGwx5x7i+uQ0yJ48WZh7GPgHy8IzXNDQJ0YtAGF76AwFpNwKtSjT
57ZrXyntE/EgkPWXFAv1xg==
`protect END_PROTECTED
