`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fyMTjQcQI6JoT3rtKc3KGTCGxM1SY82MXecd/vwep08dOivmk1x2UBSgXPXChBLd
w/RboprAl/bwh0KoGEHRI06dacGcxEN31kq60k8zihNAUA/O2JlAWu7WsWNL6XhJ
UT2lX7tcNGUQRY2QQaPJQmxR5p+YmQCEnHKbzGY1jPQ0RqMapmGeY9W/cHEgPv10
AxnPgTCZMxENUGAyvpJs+lUQfMS6z2bKZh7uaUkhS/ydJMFEvvmd3QU9VjEIdCc7
HVeDqnDdYWPo3YE4MYulSxH79+l/wBldAJYVL+Raahp6UY+x+bRxyp0tV7JU8Gu5
7xaOTcpmA1MT+Iqjf9k8f0o2+T4xw0Uq4y4fRROcmMy46q3TQRSDoHpn+jdNDfE7
`protect END_PROTECTED
