`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bEDTD5uXB9dghPfwwK+HpBeDNWB93x+6L8PLctrFVjMorPpOO4PguJwXaU3/RJP
S9paaEaf3sPCm9/I2r7pZUG8U8IFyoSqEUVr+qlWAtexQDfQ/3jBrtAHBNj9Xbtv
DlgXf1bSIcF71fI29SoPsuLH4UEA6nfARFy/AIgD+A8dBB3YFAxdOM/UAIhYS9Lm
/CwKtZ0NsDov3gDo+hTqYKfQjPEC323f3avt1fH7IdpfGoHKESOmTKP7BU6yQAeR
9oXygUGWkX4VNZWFE/PkKmVzJU3bUX0Rlm0Bj5PKYx99xFen/pZNWuD68wS2Tyta
7qKweeWbN+zheQm8Z0pcUQkdw0xRcNP1dc6yfadKYPmH5oPcW3sCnwxiwAo//Ofw
SXwPFsmi/oA/YwvDmbbRE9bIodQH7SzzuR1WzR14rr4yKhTTW5Zj4JXWuJEsXBbC
ryTByevavHrxz4naRt3kHWw5DRT0CyYC+8Wq9aTnyBRcz3djA3iFywS3RHSC2cIJ
0mkJBokalQAJDb3NZqqHCrw14TcFqK9EB07kzEB+8i6OTom3z6hQxL98tDCqxoCz
eGtAugy+WYQxs9P8uF3K1pP2A/yILNVgv/19GPPBi5dSmYDVe7zpDn3fGVY8kj2K
`protect END_PROTECTED
