`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZ7A+wbpY7NpPyIhqMcgThLHObB28Fl2gmA19aRjj9tXhzM6+sNRao3UeKdClxRa
Sp0cHFSvNB/OW0egFP9+4cheq5eKWv2teeTcaN+1j1cweicDLsKlr+VMKqvCYuaQ
ZgOIyuiT/17Ls016GEWBQySZHhdHTr7IDlHbJ6NrNNBZV6vL70XE8NDeN1nvzTPF
x7YBvg34Z10FbA017kcBWGQ6Mr6Cfge9JKol90jcu8xUdcXFhPwck/vKiegYzjMb
R2b1nu5qgWQ2W7yFVMgFuhzG/cG5cj55UFWY3QylXpCblUubZ5dTWGbtAFjVOPac
msxhQTUSkMWdZlaLWF3WB3rOK3vCuj7tVMSebd/E8LTudiKtUmXVOVnzYh1+CwuN
jEFAZbyb7U/hMlxdE4SVfuyYy5eVlhw3lOcF1QjLeZn/WVkQF8Yg3Spox9Kba9ns
k4w+ybo6RqegO9141iGkBXr2TPTxa0QDS5vt8mkID4HTxfQbsEc3pmQF9dq/ZrBC
o8qwBQU6JX0wgcrYDASEWA==
`protect END_PROTECTED
