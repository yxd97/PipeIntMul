`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KUQj+9k6i1kygs+yVKF20PajBGEBrNgnSj0Q+Nq0OQQY+7Klvhu3rOCitnHgvGcZ
pMs9N+jltzBSUA7JK5+UVg6GlNWJmqWGKCYtMGutNX4u2Q41UinCS/DijyEFKSOc
AY89Htx2ACyl54BIw2sI05UO+Q9vjmbNOXLNCVr5f1yxyv+iDgmcbJuiLOjZBFyA
5DTRsyV234xUH08wcNA8iYk+9mztTimW4dU9Srvl4/ZOH551TwOs9KesbHWcp80V
q/1Z5tJrnU/iGi4qNYS9hmGwx8h/S/WQXl3k/0MGrkNik4G6itYOVEeLpm/K0iiD
b2IA2WJP2bc9TWRWKNMRcON0bVvTsIqYX/GQw/wu6Js2YXSReWLXkFVn5s8EYFld
U+SJGNhEk6QbeHeWeI/lZ0uMcJCnFHjMGcmrsgX4J188pjs1vkA8buvFrtEKQmsb
WmyfIC70gyVwR2eZJdhmzeS0QJgFv/PuaaIbB2giya71o/FQv+Lo1vlThMDlDqSy
5abxM4oDnoMBjYx5FFkHWZ4cBO8cli7rf/UVt6E2wX6R47ggInfKZGSVBRcHsZMU
vgka52AUitaCfqXKUgPu3RQm+QA+xWDjdC058pof8Baj1kAFKrgW/A7mfTDfXDrv
ywi2OY1TwkPxgNR7I5TZtQqi+SPwpypQnOQPB++jYglSdB2o50UZ7uNcwSiav6c7
kEMNEtEdEMjiebpM/PIfNniuAJQLbEc4fX7165xw1ABvwLOmaG68P7UnF3RBTbxj
t9bLnJEN9GzkNWR7vnJemrzQvJiIJM2d96l7iRLXFQph7JngS+wSkXsWyHSYTX4B
zq1R/o3knr0Y1sTvwsXtQ2xun8CHtzwqP56vDhsxn5MWSB9EJ9/6QDqdgtQZdZJd
JZzhUzPQVmUbgJuWh1zr5R5QCDCnqtrPkiqyzHrjNzfKEm+F8JOG7SW/nRzN7pvh
G5+Wif4Ho1cu27gq9sML7SRrQowlpNgqY08HJUj9tycO1cRAoDqtK9eMqtEmcfua
9S/WTwWqizC9cFK2hW90Pqhd/jSuvdFX7ZGtJGYxjYY+kuKDaevvxeKwmYwtyJCH
ozptVkHf2DI2wphl4bn1H2NlFRzTT5ZW+ksp+xFp86jb4MiQJI1vBERVTragN0/H
9p3EMqA1t2yP+Co3xNWYsxp/3ti8DCK7E2IY9DzzBaFaCj6UeuYNXkjMpBXM5N91
3qFA7L7GE4idKU35sy8aFR33ipraUcTBQV7jczuSmqDvfEkWxyhnr8VEFNpRy71+
Ymu1L7FSYiDt6b6+UVkMNytprlra4phKxPNUUKLzcml0FKMMpFi4s4HOsWKrwfQ6
60xaSyZ0n4ANwnJ+2r35jWz3NAu3NwddWdLJ7EOcEhw=
`protect END_PROTECTED
