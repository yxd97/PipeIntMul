`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QnDtdp95NL3EJmzJaamIIuvowFWyAcPUzYdu+zeOk9H+06K0OtKAiIfvRiv8wra/
rjoSUqdl1xU5VsSEzERv1+AR/3Sb5JX9RpE1qbp1vomQb7IwiWzMKmF7iE77OFDJ
IjqvYz1p7EtAqB41fonbiuasHgktOYnbphr9b91xT/N2KnK/kEupCy+FIgzgCtYp
G0iIX5ewuZvw2JsR9ifIlgGBsXrdokWGLNpd7RtTbQFAQOSubtxwJuDefSRGPGuq
PvuFgMJYrNbXMwgg+Ku9jUrTppoaYHQ2ayhyzZtGWAATDP8Mdi/eSt7IKywhpdef
jcPqIeG9yX/WpmyRPDA1W6vQLaVhCC8tsjX3ADJtXZfmG9Wru8uj4u7dbTTWT5/5
D8u4iDq18ustI9wSIzO8WV2oMmQ3gWP07RKqbKv0cTdiiQjK/GO5w8trwI/1elXZ
l7SskYffRtPcnVtxYYp/Mi4kfPccQwYKkZ0fw3N3kDdWk++ZTqaXwY/pKaxde58E
K43frPujjx0WvfDVpLShYAEH7bQyn3k+PqAWX6nvP4w4kZ8XurCl5UvGoZKtV9QE
LBzSSU33QvgIyISq4Q0k78uloyFswMYvgnnb4A3Zd6OCpBQ0YHEE/5MWMQGyQxBw
w3b+SzcTESPrAiJZ3Z8RMqxWopUc8dEDxttN/x9B44nR5Yfbt7Mfz55PVYQjejhg
6PPD42OO3mBJaI3gk5jd3gA54wHczZr33voInJl0HJEo2b/bEfZ7UsSZHMBmOyb4
J89Pwh8FK/1XTR/E5FEVNrafzwBU7rRWSZCu7ADxH0I=
`protect END_PROTECTED
