`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7oiiqF2E/AFTMx8A8Y12GeAu0eHGqEinI5ZZmfvvnBYxaOEklQN/44D9PPxfckmw
mrbISWOZg/dgu4GqEiA/5h0mOS12qMZCwvABzDflRoIgbMBdv6h9OXt4Pe7hdGPZ
muZ5C1R3ZuwjJDvvuZu0/8RIvhS5vpQ3i69OGQdKmyVHiLIZe+Jjpm9J5r9+pVB6
jh4DRtxHXgjCFb8zKKfSTpFGqxad5XhSU29SUxCzL8PNB42VcUlH0iaisxh4VVvO
QaQmX47sZcqltcMcM6tSPtpxguBWNjCR2TObucTAu75Enf5jLCLrbBk3AK4ymfa3
gmUgzjBx1YTC3XRPSxgqrs9UyzPD3CMdNGdSJRmwdZ2oI2Q5BGWzl/1vP0QKYGII
g/43nhk1MokwYbGD+daRRAScqa65+xGW8HPJnQTF1InOMi/gPRjgDTk3Lm70DxW2
dU9QRWfT9z7K2IsJXx2xWHCXOJVgIszsmeHsuqP9n4ReOLLhvWBXZL48WHxm6rK7
YrEK90yQkFDF2AIBqQiPpvaTVw1OuiKiKzka6Fe3WhR3LkyZTWmNKIU/xSRXTf3w
YNoYprkrI0OHqcdPFcmcP3Tl5iaPUDLpqlMyEXTNtBnlv55cAHQemYaLYPQI6/2u
79ZGpKXcVRQuEAKUSVDl8dvT1wHgVZqQW7RiHIR8PCiT5CuEURnOkqYsP+PUU5rC
jp+ZmYp0f04tdsZsI/EU4C4QrJiv7GbnzDoWvs3/rGoR1zKGucQEd0KK6RXb5bxd
UaGA0hoEIB2DfTaczaUxo/et6Gqrh2wgHENtS9BVbWUn5QquLy4qZvJK2G5BNlDc
FrWFKp+27VA62bLvXQeLbfLTG9untir05xm/jgGMA+YCt0s+m/sdB9bvbl+ejrgX
zPGD0LPJRzrlU5cpK5o4bzWRSrGBChGGQLfcvgKN1O5FaGOpjm+YPeDM04bvjQch
zPHcwDteWquWcvmKapNgcvqlx0m7Xu9ljbxr+1rRMfA=
`protect END_PROTECTED
