`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GA1p+slXE9uQ8+Uq7mFDGnsYnxO4EAV3PNNnrius4kGri7VejdJXUCMOBcaIbr22
6POC9grbtvWstgppe/9j/IhiKLqnsTR3YMSBR0MhjlHze9H6l+vYSxKYrcqUi5da
tWHs1MhV75PDsQrp6HRJUyg8kIOMkdJyhHAP93XiQcTJiS6x54ayNJesBGnOOFVy
7TapKzG4HPwbBdHcUNyA1cmikB5CDVDnLhSNSIUW8H3Lh0LVzV419whzc4Pt0DbB
VDH88zQb31FTEzxd4N6dOXpgS4fa323QrjMyMqE8XJnhbyld7CZpf6eGlEDBThgk
gliYAMCCe62HLIUtoDSHShE4gKKvBhDnkUDOGtjcAXrcwLaLGMYxEo0iBuCdr9Fj
zLM8X8s0Af2tZSf9cbey5SuNhnmue+m7KzbNF6cF8lpTHo9PDc0hkcvAhnLr3wac
hxRpTbsktL56Fs4UZ8g26g==
`protect END_PROTECTED
