`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l9lmbm+6hyks6eDaGuQ/X8vfLK2VmSlSFFw4yolGDKEetU9a9aEiQOIQ34q27EDV
MjrPO1VZPOVHnVpc9mazSBXnBd5qc3IPklDILihMLcwllNtqnlcXt//LSaj48PDd
zGxy4eNTnrJuk1ogu5sfNjqyaiI1uWYC893y3IRrT3Pab0rwbBdsuLkE5BOFuPlv
dfOLgWVqB352cAPCTC2X1V0NbzRF9UC4/2MDZ8t3bA6JSJ0py+XNUwzGwGTS1uw1
rw6J3L3hT5aaFHhNWa7E0IYD2c3jlTErVgYUddpVFfRUyU/LsOicnYw21rhT0lRv
h8i+9/QJtlKY8s8HTcXJAUPGr8lHzjZyE8Qzy5wKpAu/N4YFJQQQEHKgIJLE+R/W
kk5Cf5jOq4lhx0pZVMni6M0OwiD5GN+7Nv1lUy4dP5/YofaCqTlKJXE3J2AU83U5
rXdFxDYcbf6vJc6DFbBXALUT144jITukJlXk9wK6AiaNlETXHdQwonaJ0h+qivxK
hPmGAd0TbnfXnG+UMDCCG1ydyfqnrbq7oFif8EreOVnK8R7amORnEpsza8vQ4VhZ
shH7pZrL3QXUNuPHKMlca3FJjQhtzUSNqbkeZWpvrZjyEzXIjLeT1AF3wnk615hp
GY4V7nHab4mmVJ+LT7IwisXgu/96ePO7sVBZ31dIXk4G8j1Le+5WQksXYI/TF0lD
ICJDuT/EN/t1UwWuw++IPV9OfCONHE6qQE0gTPTDL71s2LDBmFR4WnExB0a3NX1k
7RzaAtodry6juaopBmhiLxlBfCHsJYdxSl5N6WoId4cmraYaAGu4DbnyozoqWAda
LMR9uHBhMxAmA38aN4phY7Xj1ww7PgMdo+mwdMAAaGcpH5VHm/ShMxM7Fao6PFKs
VItBq4z6jrtXwVb+mCyzX+eefKq86R4GadZFEsSpH9XGE6f3QDzWAWq19QLyuzSk
8SYefvJFyuQcDmoAqU088m6J69Rn9P6skMl6xJZeYEMD+3ssxnw0rKzoG+rdaKfi
dDg1SZgFpz+0Rx+oXV4EI8T/wwaeRWPtGTvulFUjVIzV9YrOWxJxI8M6Qijn8aYa
UaSgso6MheiiMXgBvKDiVZnQ9fSPEO0MGT0cycAOlZnu93Omc3lWB5nVmrzcyvc3
Eu3od8FXFJoTqGTbuGpwfHBMCTTNhmGaMOxit14ZxsbBRh6oeu/SxQWjh9OxW6fT
VoQxNK85jsbfsIlrkuvazLW3T5l7uxHjHtz+NkqIy6l+aAgK9R31jzSG8LlN9J2f
NBt4VFxhfn+IAwNg7j0NbDMvpWl4mSXo9ZvWIL3Br79G+7/+cjSYWJpYphc9F2UM
3zYoJ7gt2YWzumm+Vsw8jw8P1WMlSFvs1FI/2xMoERwGvaftDXT/9A68oG9YoBlP
1RYkwgF+IsxlS9w9m4YdhdadVoVPyt1rwcZT+Ae+bauJ7JsIeFjC758x8l+0kIro
eNdS55AdJt8rdq+fHAOG/V3pxKjDyGSRpBuYrEk91h07N0nWwhg/XWio0tBiYj88
xG3bTZWeD0PPv42b/prQspwru2Ylzrh02/mCL4G8XN2D9HtE6t8+IGY8FaVfiqk+
oLnfduJPlu77ujBVu5alVzxXHrss0hdvVOP/rIU5iqcc2LUA2sZo2hYxG5lLPoQe
Fhz2A3JWee5+HOJAqPTcoK89ddnPLI464org1gEJ+g4mygQ/ecq7XVQ8rXk7ADZg
jfaTPUt9PKcfFhiEIffiStcVJsgPRh1QZuWbCY0QaPNUk4DOlEfyXjTVjLRukgWi
hPtlIgB/WafkIAjQriniryJjLHt/0+IDSF4Y2WGwwSl8pg4vZRO1znLYZk6lOHkT
YHNpZgliTzX4Y5yXpALEdnRWw+U+jtwKvfP+1MZFA3rpMAxt8SxA3RCcNmKb8bpB
Oh/ihpE5Jre4hHdu5c1lZO/I43j5ut+YyX3flhqmej+hPsWKbSOGjnMiUSHtmg3q
5ZYyCEgCmHbUWxo8k+zAp+YTiqJL6y6QeXbpfkD3tmTqPt2o6I1ecbtm/9hMOduc
pjVQwQDuu4/4audI5ET0Gdvsn7w6kh7+y+2GiFC8LB0JONovNe/qpWysTdrjAW2R
vwoPQavUrqSRMvBH1zwFkD2sz/YTJ6fdGmIsOL08ZMMB5RfuQ+UmHxGbu1tBlR5n
Us0NWaohvptA+EIPwZEDqVOgcXp5nngNpz3iJNIR9XEn3Lcddin6PtGwLWAyVk2C
k1bAtt2Tu0YD8j98MrnhQczeNJXXpJFugXNf1slOrxcxUuVnN3P5P8sNeivHfrY6
+Zt+0jmIICnnWdmCQ5pKF5b38F+A6QxhSIsyxjEQm8OOKmMIB8Hhz11NeR6YZ0ng
A9h9kvk/vZXGHTgYTFYhLDwK/DKk1P2dhex2wLxlgLMHQ2Vlr/3b0eiNh4w6j54A
`protect END_PROTECTED
