`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exP/CAbOIDXo6/tUOaqPxctUiZRJWMj69yCiV+elGTRg0P935yyS4XuSCjgfQ5JC
l8YdVpYkFruiGmnLiQIv570E9pnuHtuY8XFr0/O6HN8TCNTOdbk5yxtwGljFXeYq
ehU8tBdvKGSwy/eRD+Py83ncL+R98mIGOoajKYPd20gAwGD+ZMNisXirDTIdgBJx
fgM/3DC28mQJjTe5vfAq6PJ5vyY/jTF9xgu6/QSnFqvK63BP367HaEVTQ3Ga8Iby
iOWvuI2lwF/1/3WWiamrgrp3mEAc1QUC+RZC01LDSbgyplhdLyWWg2Zn/J2w0mMj
leGRFoHm6eXJRoqq1/KiDHWjLdv8acagy0jvspzMfSQl2vqNtyI7Tsgp3L976T5c
gCrEX4LU7dYcxn97gouVbH4EQbKPr0fW9Q5e8fO7v7610jNmsmBOAfEOynsucoOn
7nZIbmEZCUwKbGMXydrjU3nyjtCdNWH8t6Hy1aSfCld8omDKQoeVzCGVhK41ZcNt
`protect END_PROTECTED
