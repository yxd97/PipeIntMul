`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kDIPPXjIHvrD3utxDTqsdbcr6zHShXqxfBA6mr1L6XLW63amW09u8OLUw3zYnGd
gRKfoCoDmU7Kpo2wm04IkFhRdThmHkGM0Wnca8ScSpF6VVDFK9YNmLiVzTEKIzLd
sHGZFqmMrxUOKWCxS/H96L2pKeH2odRwC6ruVRx9MHmKMtSOV+bMevTiPQm6EdjR
N6oiWvW7xDzsH3EAkDbNCq/qnFVY0vxbzuQVgqzZHYyP2IuWwux+AqgsDuhR+2Am
tFXovttI1fafwi/k8PkJh4W9WIte2pMWIu0EyyaTpIiSxjJeay2YsMLAGXMf/RyS
0bcGmdBlfip0joyi1mjlEu9hiHLhHm+7MXfwYdehcFK+UuIcR6EqWpZxvcFogC7H
fTrJe+PzejHfIjQYaCZbRabZEdOAOduqHtwlehrbEBUv8edwUvIDZj6m0Q6u4MO4
qqMzXBwaGn6oKcCfXnM/mAQPyvXqrTl9CPrtG1hsEzt3wX2mMBHaN1XvvnItIYvQ
1rOWsKAYNKUWeVwiey6wRrq/VxbKcdf/JRL1yylltI7UeGZkYID79T5G2qK/PqM5
`protect END_PROTECTED
