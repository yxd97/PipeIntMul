`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cke4KMgUESN93zcQCHRZsYwwzW9qd0PtTlDUl2koNd2vnHFaX5m9VfQbSySoJGbw
o/pNCz7sdrPCLQYr0BPoe6zJ7NxR3QxL2KYtgdNZQk64Ota7f73AgIOGbhUjSF4c
m60t3MS25qL7qxfuTX5L86qklXgUVJVfpxs5Wc1Q1YMYzu40Mh8FvH5XRFDspdW5
UYYzCmE94fnaRX+TpHbWXy1KfQzTIK01QWOBqym0N4PvORW0EhMdX2x5tgXhT0PF
BvVZfDqM8Y0d/RIeVVt+zOXj/gUfe2Cr7BGJAoQy7Jsey/SX/YE8uIFEfO25uPVI
r0CM7Y8YouXz0KwT9aHm4By5Xy7nnEwRFaZq2l5aCs/wWSJMQWHmqJnu8da8ZZMT
CH0BUyB0pHK0Fa5QWzpetIfbi4q7UyV5gdCIIAW4GNleb3WL50sazw/SaC7Uu7+z
j4jdzxqU4GAoePoJhrWSLzQ0jwwzPHF9FE9niWGklW0tr0DlUe75y+njoUYYMLlW
4b7eB5DZB6rP9lQoY7rAvBVfEHL6kjgXB4GqrbQWWxDhObURKMaXl6fhlttS+OHh
5x07mXj1KeRIGQptFl892wgL6fCcRYxiqFp+9vyFsN4=
`protect END_PROTECTED
