`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m8o5nDlg3YIn9BRVh4r+NSrN3bFZjAGqGQCA6pU3KXV8pzos76d20+eZjfG0D4sO
V1eejiFKuZJRPAgT1o7G3TxhjojO0D/8DwMZkMvT9N3UckBQShvoEpU01XzQZY+I
ZU0sbdeBWbTc3MtuAEtiMDiYTCQLlRs277Fr1sEV8BCSVqvVLeRKUrHqtkC8kevY
CmAoMu90x7ZC1GbdBj9sgCihbf8c6u8f2wTr9WAGHtpanLg0zjkLlFjMwHaGpMSj
8Qp3m1PhZOcStyH/36dWx+QZKdrmaVu8bEdpdnQ+dAj0y3KfgHO0REPySHWb4yHG
Pl+jFw5Y4l31aKz8GF9RUnOu4aeMEvJAU49eUFXtQbwlK4NPuaYquN5jw2kHUWwX
zk/VCsp66UOOKss/FXXvvcuaHLMCCBkFvFrHCuyG/HsiBUk+nDP4SUhXljkotqQ1
jfGFk3gc76HElySiBtXxjtKmT7H2FGsijldttakuUDPwgpYqL920PhFybMd45QMm
zyrYho4m3m1V4X0qQ7Oz4uhBgdXreK+aFbR70af1MlZOaVW5fT27F0OQ1HymlaSQ
RFrGKauR4OvyLGAuJM7Um5yg5b18FOxFhwVsEZhJg3SM7oK/OaEThNi7OpBSQO0g
Zg5qlCRn48KBprl5Q+Uo4C3dS8U70idT8OcKRGGbTvKYua94OtR5+LGEysGAmPpn
OrkuELulk8lzlh8kSQN3Y9II+cSDkwl1E6erI3X3ZEOcByorBWSSH+oAndPqet57
dOjvwuyCMPJvYKXPxd8Z1A==
`protect END_PROTECTED
