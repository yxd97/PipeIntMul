`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfJElMqATsGTRHAuAvarjhujbrwEF9jtbdi8n5zdT0m8Ngu77Dtv4i4H4rT81unJ
3uzxJxV9A/sR81nlWiC4gz8E3bSn4dImF8fiw6/6DS4gorGq2xP3mI8ySzPSg/Np
lz4qPpv2rTmG2ub/P2sOZ/iCR5A0vacsG7ZB/LE2OXJVTA+R/JNagyJCcm5t/aiX
8WuZsJnJbKq+2gtA77v0UU8kQHsKEbbpB6yxBhzUQ0w1FEu3v8yEyED7YMR3TRJY
6sAh7bGE8cmJkaUG5yfVdbm3bjhlldIbJRUQkwhsRaDHezzW+PNcyxA0dLpufWei
g1kkpJGjFs0TNigNIurtaudprJTp1BeCcFgbLgHvEuw3s21Yds9I69qjjN0mhFbL
5520g08DZZuSQMZlR1ClElDXcYSIbFkgTUonZR3Zlav/fZra347ugpdkJdLV7hQF
l12jMeIARuWt0hA5PqBPvwtPVeEjhj/p9+YYssUyjyE6qDan1kJSw7oZccuLCjmL
MD+IwiPk4jnLINOb/zyhftNBv6n6yqpwvyIkbsjTd5l9kmN3zlVaeQemA63Q80ts
kU/i/9FLuBoQ0LHfsU1t1+sNJs7deSUueBNma0Li3nU=
`protect END_PROTECTED
