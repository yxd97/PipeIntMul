`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rTkoGtKK9/ID/GrE8SKmrweHMPJS9sJZ5TZTT67b2fKjhPGAgpVHfRjE4sKBWRj0
0XqDL68gm/gWuo+nldGumT1Cv9y9PBvA4oF59YYEhOQbTwrSSH1HrCSAtba19PxB
Jq4UzqPAFa2wIActce8KVVGxeWY52kBJlQ7MWefHpsVWNnTO5/tSnwSC5Eri41mf
i2A4qz30nrcrMR8GjvhIONBRhNUucRPegh0tPbULORCIKvD3HkyQMEjq75rExAkI
XuhU4MvkLfFSC2UkYCi1F40wvu8dnAEahUbBcNIvpNrcqhNe9coK7rKIdTgdln+p
kVroyhr/HMe6Lzf9ITNDRVyuLZuDUozLjw3YXAWr1Mgg7q7OB9ocv56DvDA6n0ES
fDhvhX58K6JpfRblzcu/VO/re/Y/5m+byjZOYTcuxC/SWHqSGFhjcxFIrdYq27F4
uWm9dVERe7AHfiWSJGaRTpZS9DEDomzMWpqn7W6N7Ud9bZEpxAb0p6O4x86x33tV
gjaBhtIUK7q+TGTi9KeL1HsPMPN4zcutBRJXVkzV3vuhMZevZSDBrtOLSxqP+i3V
Y9T8DsrL1ldOtbTlZj4hMTAN8RzuRuWlgXOVXxakuRHrIZSaIT6yG/EgRx39/yn0
wjBrvzs69EiUGhfKZhuvcOngyYuLUkIQ2tnWAm/5I794krdwK9wSuIUNGPbBHKKB
FPx9D3dp7v6yR6TnO1hX0ZBcnow4EA7U96EwKDMkQiTq7J+MbMulhzxcgVG7nDCQ
+o1zXR5zmw2sCPURfASCZA==
`protect END_PROTECTED
