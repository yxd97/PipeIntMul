`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q7J8g/wlFKhi5sXDICtrWiTGrGR5J5sVmCBFYJ0+sb69svsDa1n8v9zyW4rft1NT
Aon7XiCJtrgSJxQVwoE8H/X9t87JkSwQYoDMS+enYHxlQCkB4VR+9lCfIaKvNT1a
g2bmC+JEnnsX5gttmwC4PK0Qr10OL4eRcfnBcHeScF0w42eMuBpvgIUHIu1CilyT
b5u0EXWd4cPfK00+Rgs8jtmswfa8ZCQTbhcRVqo2QcRVBVNHQteEBIF5+U9C5k37
eCiC4LzVqgo/0NNrEtFl6aBd7Yijf6EQt/UMucXxc8MHePAhRqqhJebNDE3PBuDU
L15K6cvU/wcIixNXfSjYTzot1CK1EKt/5Z+V8DY2lteuJjt34CTxbAZ4UNugcdh+
JsKpOunWwAML2KbE0OBa1QG/Uvi8VMcihnTSDdn0QXJuLTO6D84cbjt1rgaZCr9v
Y5Vt7iGwJ6iW0vBWoUf0CCycrMOn4/ldFHdUd9Umn9q5Z2h7MGdTgnxSs9WgHa9L
ne4redukd0n9p6WdYmvTGGzBdfZ+6/I4yN6GhzqoGi65/jxp+OGAurpy9fspUf9b
GHbAgV38L21mQ8pfKKITLkbwL1f9W2zpsdpfSxT6yeio1t2Cc+BhdJqFMSZ6qHCL
Jv5SmikExx9AhOr9aQi96zVG4AjcsaWV/uWgfsf2wZbwmvwxVNt8CIp3R9W0z/QI
qaJriChrYtwTHkM/+F1Yu6Jv5EvgudxFscFzT29V3iYjzmkP0YCZXObkTlwMmN/w
hy5eN1KdRk09nMcIImxiuzj84b1SKSuigRoLP2BcIOQPxBIQeHNI953U1k/xHKB+
vvDwyw9yCcme1jEa7MfY4GirtNFpb8SpNCUIEMbhvVX7QRa/nYROY8EcwiFkEPD3
rY0CV5IgrwUacBBprtZZXA==
`protect END_PROTECTED
