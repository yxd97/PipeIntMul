`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SsKaJ1z6o+ocobGXHCQKfr92sVyFdxwTVPQhT+p2Bna7KnOc8ID2rt7t1KT07sZ2
AZWjZMksFXtpZdVo0E33jYGhr93JZ0/3wM+e39G609bY3p+4Iwib9OvGqI4MDf3P
DEzxAA5XKpcXcFMmEZLb4lqLw2cu2tpy2Svzkd6NlmZPjR7AqcoiLBID5IG1GmIW
NMRN2xFOSZtGsZRrUFbSP3dAlhsW+MrbnovXS8Vvuyi7lIkVI4d3jr+gCFy9pKF1
YUDzbvte8IB6rllcHsF3WskaeRmPIRmEM0FOBnlqEzrEn0NQg/QeOuSznJxxwXeS
9OA1UMVXxTCYr1reQLBFQAB+PbYCUukk1iY4BjhbBzGHD5Xay9qHkg5q8jp7+d7y
N8TRnUbnS52gvvVv2HI6Dw7fZEsKa1lkshARMuX95XWOOtn4Ma5r+tvSu2acabKU
XtW2E3cQBA/FJH8TjW2g2SgLggR+ZKhA02NwC657YzdXOJ+7zFAWmRCvGy8vUSXp
A//VWgo+jiqn16UMeJI7ROKDlb9Yc3Hx36EtWJMEThfkunvSX6WVsdkUHcMRLQY6
D9Hqsz21jgZ23u4TSZ2w2xRU63GD4AtCkBUFr0kI++ESYCInhgPueLtIpzAhC6Io
eM3Ij1a5jyA2XUvvNgltlFbCkxpXQwMNPA54S3COpfvoqfjI7xTj+MFES85e06hn
y7wFrXNhen/ShBu7iPOxhNa7wTMrgeFkKB1ZKbIvm4Mlj7Wk8oFMinJSq/cDaW4t
87xr78uriUDB4A8WkRlzAAAnbzp6PieTalUH4jvWJ6ugfPCv3okrkraLnKgkYCcH
cJwzOAoSvHu4S7HsqrgkNvQvONUtAsl1N3b0XZllqlcOT+SsS2YwchqFsXAc1UUr
aOwH1QE738FZIELS42oZWohXECJWJK9dIX2jQ1aUWxwMjqM1bBVVt90d9HUjJFJm
A3q9xRIn2H2lbwUr26DKLFoNw/w7/7Cbw6zKZFZN9tSrniwi5PKcaiiqOB2VU10U
/dk2E7EQdAOPUePF5/JENLl6aC7s28RjyCX4RrURT05x0m7nBXzqTRC2/mhzuyrb
I90K66EzUnMS26m9dwz8Jf5Dy6KPdKU+0l2EVd2++aRUHf/Md+C3W42RAHgckyBx
gQTX7SDQoNSsy/M1CGkMonT5V8zqJEwxzZEzT6PIbtSqjI9ysSMKroFZ7boIhXiF
ACyJSAqjmQpGL7mTytCxZYlHTV40/AS6TxnivqbzbRoCJzf+Y1m8gtKoMWksCzZj
NLJmUNkoympFT6R1WFXb9dFH4TXDT3QSrOl187ExjcATLl5P6o0/iRiSTgeC73HR
rBFiKXZyK8LBVppdUxcV6r2ERb9mgepcUIDimXxJh0F2GTNZXJyB/0FQwmXUkzcY
Qdlme0uAetKlqow9wnxsnsNK3dexNZp1pzKIV5vgOku7HCDoeMg4ykb3ysSUbggN
Kmh1PEZG6XEefYLCbAN6GPeJLXwa3CF/SGMiiQ9JHYfPii2BnbyHjKl2s/87LAOH
xgQPFFoVKYsUON7+8HYlNMwmwA1XFquoZlYSPHL4iKjgIkNa/aSbT+6z+hs59HSf
+IR+3Zr8foP/Xl2zHuI1G5/UusBLa46bv7GdXXl9q0e3FdstMQQt4jCrlIQNXiE9
4hBossiqhn6I3s80mndtxw6DRjkjG8qifojMCvwOplRrF+IRpbF/rKZUHXYeTrlj
hhU2gfRqEp5OLRCK6SghfzmxAm7o0fWKbtdz7kCLue+fcBGxQXm+s3hDKXrH16ob
9FvWo7VVox7ViJtCYB5ojQWB9rKrFwhNl+88DWyjVRlUDJg6/+LSBe28EQA2oZoM
`protect END_PROTECTED
