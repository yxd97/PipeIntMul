`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvvJx1xxxfPn1AQcB+cWda5U6cAiah17Hk6NOKRTWyU5Y4xjCzTw300TAFeACql1
O8i+gOWEB5FPlR6E26SW1KaSh6PGmtIpN3FcudUaNHAYcxwx0VBXf51WNweqe1Rw
ASQQ3/i3qv/07U31B7E+6MSYbcudBK88+Odr55UFtRo6PHK1PWmR023eDQkWQiF/
P1AEK9MSThO0ZPdVnY6/+sWWxqzPp8+eD7ikYK8rCRBbNaeRgcZerdEQI0/7Z3gl
Oh9zYV9vfdQwxPNFo6tWWkdXGIIaSxx+JvEM1MHQOP4xmebnSEp+Zm5bHh465Szs
BtkPzS836qCg1UESvfuXraA+MCLOJq/8hP6gdvZggLoqn4/Sokkt3nj5C4D0Byaz
`protect END_PROTECTED
