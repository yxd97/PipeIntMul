`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KHsgXAgLhjmo+7XyHovbuxKTsidwXYdEJlAxQb6pe5pp0I/Vem99kI+OBHnN1+t+
Nmu+IIBEdcukD92YxySgHDvnXFm+GbZ1PSD4B1hN8NTY8ng3IKNMuTt0FzlnHtNv
zZSwomkIxfORjLLlO8mlWdXlKlxzwbbDAVPojv2TkwkBOjkSQojaioVkoyOFfv5W
Xi5wGoVlXdTKuqCOaH5Ay6vyvQPpLkQ8HeN3/pfd3OBvmb8iyrKaQg6pR4z8bl4h
b5e16j7a886B0SFQxylMH/fq4H/CD7+mUvx1N3y0OQukzV2ql3DVuBXEtqNtCHn2
fWD233CISbnLfxAqRrFjL1b7UaICrtyv1LOXojk/xt9xFQsLwmsRMMuJQXf1C9Pr
brno/YFc4WJ0kyDuDj1kBtapkokCCMeTKphIqJAa/OHjNUoOnmtU7Aig9MLXxvNE
/3UFeTXaG6t1NzvqIy29Wk/swvY7rNYJ8BZ/0jXpOfcc2x3tm/iIS4nxVa/Pu08J
hiw5wvbCpVgxQ4pw68mGNKPSiyrzPTYeUDY6TLwqJK5YWMj2XY9gHthJTL/X5p4q
3oenW96c6FFbkUpYHYTuod8dPRU7v9kSjaPqqbAH3/sJD7gr5OGLSxB4nSG3KcZG
jhUEWit0CZdd2PIWHvIZfO2HFYefew3ElIM+HyP/GiyPMj/kDs9tvz4QJYA/yKlF
ihtdtoT5Tq7SpzUcAF3KTZdB9WBwwJMluZJsaO1Ayi8ycynjH91+KwlldI2n5TP0
cls7zGVgr2eSGZIaHkLkt5O40xuZx/xzzPPCNpENIH8dQGgFO3y2+4IjcrT1SINm
LcbQztaMKCMuEO+pn7ih10+mo23XGxVqHUGUQUkzRzpAUKoD3I6Rf3RNAqdf+xY3
wn3jyC6mIcBJUwJgPWTlA7qCoWmhyOvMQ+s68Ys7S0dzoqmoKnXjBbFlb8qYrpfm
32S+PQs7GWovC0nLWguuaZCVMvwT78MYOdwftih15dgnqxE6XdANUAdb547lRbWS
p5URki+A255uHT0IdcqAZ14m0WIeqjf2oh3cSKWqNeYybsFewVBQLVozojq4zuae
rtxb7ORSjE8dHyWLaGB6/3ieY3zp5WCwxsEnujrMJpgNp1EfKuTkLRDhwfnZiJ05
hn56is2m44dmg7aEva7/9LquzXLtOp3DmKA95S00zXzeZd6gUdQqrmEvh1IqMwJU
9baAOC6dZUaGtkevaKgKtXOC6xIMQMlABJkK4D8owDgwkzVr24y0gQT84PgrRqTc
1/IG+tDFojLtUN0X/lEHLULP1Ie7K3g9yQShDN5etyM53nmW+7+Ze4UVP19mLXmv
kKt42UnhsXv8NgCZz/NXhaJnMR8t5A+AZgxloGqIhot7AYYf39J+NZh84QgnLrGT
aqlVEaXQD9/yUC7ohqt+dfUsLzpY4R7J7wJfI5p9Z5ePsFFHMXPWDDM7LlRn6PIC
T4KoIykFlXMtFFUtN9/a4P1nz5QaZlfHlw0yCc5gpbrr+qHRzBGh7vt2EppWdhK7
RWeERtPfLyfLkYnmdUC+EOMQ8g5ojGwaTnGl4SB9MpPcrt/OmCnn/NbsDGaABGRW
nmbAnYLdL1s9E3axT02fL5yRbtAgqONNUn4yTw89c8rYJ5M/KQDwlv6O/GMt0ch3
FS31wRviefFK9FlLDVD3+UG+/7u7wB/I7BhlUzqp9z4GDYSMUHq6LZkoXURxSJWg
6Rig/Mnub6+JWcK9+JrgZySSvnUFUBeIgEADmZr5Jwh4kHTr7sRPoKh+CtQ8efSZ
O1a4amnXiozqPz/6y9Izi3pIYwtekjIKd/lXLIgKtJBaBwEXeUDuIJUj0OL8N6pU
+cwOi5qmJXpd8mwhsyDIxEXKJNxtMkA/wk8CPjTMER6DIYkIP3KtxW90IkjbP7QE
wyRRfb/CB+WGBlUUstD7MMDpavIGxppOXwsBa/+xSzvUTf6Yihztf7+AvzTQ0CR2
LRpxShlyVMkPFfBY4Rp4LazOG86pDk8hwvav5CFssBUj1n5FCCn2G5ZGJQ57TE81
7sdF5MtM7Yc1W59EVhk9BnXs704I1LTnIzCoYr34AKkWUGewfmdEuhGgP4fVqLVV
oQNz9gLc6Tcv/G0O4LmZ0f1deDmJlKDtu/Jl9zLtZJHqo8+Uudarqjm6kWtzAIXs
RqYKZBjEodClAZWTiKAatZSZCFzCPkhrUy3KR/rqmrPMYTDmCJb/6skz7UN0HCH7
2gZWFBHAO3YpmVQ4KO0Qrw9XOXnEHdvaBhY2q8PYLTH49pyAF7Rj6vv/uFHKiKGi
X+RnnMaX3hpqPoDzDATeZoHih9eW3XJZtzdHS2tNG42HUMOs0IVVLIS4CyCYZ1T6
Qh28F/YyKc/389YMwdaH5ybp0Wih/azq7fBdD4vZqEyDQIOAA/8/aYXpppjyPIh3
M7ohO/6QFtJuzmatrRV0DttDYGfxaug03N8QOg3mZThXmo8k6pqiRd0TOut9DTQb
xqDsTfYD36f4Kl35P97LxxGYYIxQ9x2vWhUSQn2Ts7fAdvk4iaRfi6qPd7PsjrZb
AsIYQ5Ra97GypMjefrLFENWevKlx1N8B2S59v6tseSTSDQ9Yq1dfrsSn1bg39suv
Lt3e+Xsmwxw+7hXKsJqvMW9fuXNvk33Iobgt/qDBXvgl+PowUDs7fOs2RrLJsQaS
yUqOJ7+1GWTsXS7EHNsKbArVt9+FtZHXqRryKScrEsXwOdxNI+4X0IxSWp/sPP4/
pr6ldyiZh7cF9DxMW5ERDjVQSrAlRmU6m/HquK3HLhO1o8SOKNuqGitt1V19Y8aP
icfi+wXuCsQz8OG6dk5RKsrVrLlztnqeLtApUx2PcAhEf9GtC3JIO+5Vo+WSs4KZ
HOR3OWx/bT6cGvNkO9D8ByhjgCZWrzfK2at55Jg10QnxwZZuvdmPKxenujiHxGms
/r10qk9LaUjh3KmqS2mM713coaro5QAbqreOVEkyrdgh0qa7UsZUbpw/WB8VIBlS
a6waFt+ro7fJyzdJH+FPnhnTukBg+hyeZ9zBOINkchMb1ngDfAVo5IwPee8lVie7
y4LLyjoykHdfumP31W1a22H+OOtmjiP7oO1tMH9GV0AoXXcm6O4AzSctGDgiyehw
J2c/l2OaxA5JqBWAMdM8+xQMtRbOqr9Qpg6wP1V3KJUCL4f26YmMOe/XpPkpjySb
GegaDjH5E1oOhdsYzkZmMvmozbNjEhH+w/sVVzOgcAXDZQGutO4kSK7kFFMup2Vh
/dAj3Ys/JqM4gfQmBs3td52jB64uHVsKAy+xfbS1GeNpkYT94gGWz5DATdxSYD4q
xV0jPMFG2zqVsUMQ5wiPUL1F4H1xzv4GH2gB0dZghFzaKsIuPrTRFlhhdVkMYNYz
IXLMhLr4dBA12xJlRSFBB/Ac0hFjcQcFqzVJf7ECzX4AvZ6r6FB/i+LCVXYFzx4F
VMVKP3D4xqo9b+qkyxNUUei+9OyQzMPxHp0dXtttMjunOcckasQDe0DYfLXiJr2M
4hoHi8+Yd/wNYHYiUhuABTpkuPzIqlG8z0B48mSgArd5haXtPl4Pp9MDkN3FgIO6
k+M0TAprDf3JWBRsICdjz+hYEh25dgvaoozR3QA+VvaXg0E9alUK/A8PYO3TU/nW
HWE8SjySBQV9uxGtvkwPMg==
`protect END_PROTECTED
