`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpiwG6YI0YnnNFgpxRzpzaUZH0Un43Ww0JE6V06UCx4vNf3gQjQjaMTRneJkwduq
VDsRrgowO786v75/REA3pw6MWS9vGhtzDniwb5w4ILWY1okxAjFUfSXjj+5bQsis
TPuG6ktWn0w4KWBmZh1ErwQvBUtzCYgDgCv1zae/NF6jtDrnjW1dxMx1vG+fXXhO
wnXMilSUN1gCy8utywLqPiytc0POBGK+vNxVsip1wJCaI3ZgHSriwA3OJuVDj3XC
ugVIVboOQQ5hHidXpgUSMic9Lg5q0uG8tT74CsdhxibJYkkY0+gdB+SpLDCJ9cDy
v1vWF/H2LXeR2MxZZXU69KoPoIKlnT4kK2R4nFfsJ2aawr/xeB7C4rTlR6YBUNsp
PQ1UPwzMxQj8CifVs4VuQnmR7LUIc0JejQntYmCArHzVti3k6aQTvtNHufZzh7SH
jFVA5qSZ2c5s870Eh2d1FXmmKZCxAtyADeAHhZb0kYtc3y1e4BHH4ffEvNxyLE6f
PwKrVyNHdk8RHG72txBsceMVaZFjhq/8WRQ3fpAW+hFDj8rx4CX9XEtLOwIApX6X
Xb9ykgL60+aLzw45yUpUcU5f9Tx7bdlZ17UcE9MEjeu8mGzoQOLU+hn986kDOCkl
X4GMvF4DuYWKkd7jxtTydw==
`protect END_PROTECTED
