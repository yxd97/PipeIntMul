`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXKN+LnBdJwPhHl65azWzXHHQxfIIaTHhv4tEyToYPZBPqIMB0DBmaVU7nDIDzwj
vVHlwRW9GBKcc1qbxcD39hzl31QmxW60N9exbkuWgdv2EDRApXvOjFsSVcyJLgom
xxYqN/5BWPIJpdMIMK5wZkzL5Csw360+Hd/qdrngkjbjyyoo8D1dsabZVxEHW8Hy
vFnOnBAZR7u6jjzMX1F3ru/c8FOZnvjSfm2K2053Y7YQNt/LjHm/+rWqrXaKBv/J
vy6AsCaFQS8Ub1wCihp7ISlC3LGpqE3WhbvXA+C/V5vVs2/0WNNGGU6jjsseZBY1
gAJPklNMjS8r/sUgPQXzm66oP0X/cZyqGP+3OW4vxD49JdRcwSVI8FpPQiWb1Rdn
KEtL9qtgR1+amxfF3m68vl7eLkTo5nUDH43F2sT6jbAANHPyaiJuASFqfZfSarBp
`protect END_PROTECTED
