`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fL6Km6rqdzr8adUL6Tt/5/HzpcgBAppbWvfxEH27RbGGPh60rQxy9rpe6X15/MKA
BtIZT3301hl+8j2x5W56TwMFLZz8VU7up4RKYhoOLLCwWKwNfIX5oapzxlT9STCr
KlrgFKSusb/A22l0xpJJOVgPZTyayElVTWnZ6Cs25L8pCHLP6nPSlAVERZRNfuhA
tMXkbyIXrLLYz1BWgII254afNIwBy4DtVFTM2bZpPjEHm6d9tWrr/iECn5Hx7jdL
MofkmdrhNyBe8INVgSzORDHgtNg5c+gBwry7kIbR4z8sNri8Wk6mkO+/X7tErKUg
57Xxph34Uu1GFPLeaRYOlOof8yN8YSw2bBb1dMd0qRo=
`protect END_PROTECTED
