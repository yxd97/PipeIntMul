`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQ3/snPGTI46Ct8p7k3gMnyAzJ2u9TXx0x/PFdel7W6gE6fGzBnZxRFDWkmzyRw5
X15wYYxWgSn72HaRrDfykdsorl5wq7Q/u3z+tHo8/b8z60sEMIIdNYKLZkTh92/K
huJ7d/Um48YOh/wvZWqkfpHQ5jRucG+yCRL3jjvGVFRznAXtJeWBMo5OyTZygDgN
ozPfTh1kShBfJ211LzNQdIvaCYQA7TaE/PpfKlIC+hp9Jh4CkELT30mGi89wl0y2
SEGF10gcapTltNPL2R5LJX7hj/aHVXxI6DOcGzI26fC+9K2XlM/+NjeWtWEQtMEN
RxBcAO8Np/W/cEm0GdoasI05iDE0bH+ufiy/ZfRrWKO4sxeAQjl3J/Obx+lyxVmA
WNgp+U2UW2GTJjTABNTCL9mvgSr6APuRuvnhx7WGB/j9PTUJkyrfRjck+uRShD5Y
mIW1BYwHAyPvYsZukLU6P9Fo0mx1fULjOM53F4eYYI/Dk2LwzpboVoxmUIROUUXV
0gzy4xnFDawQ5q0Q6DlfcW+dFDUhk73DkczWR4ov/vUBMsUfuqFAH6qxV11KZmRk
njs2PnPmmGpm8BzsFr3D8Ei+zcbeoltL4cB/Np5zwDocRu5c27SdFnihM9W3WPfs
gVzErjpYo2yrlN9JG/hTe2r8fpUStgI3C2WQ2UgbpHa+UsP3cOP/2kzf3TLCS6ag
NwuocUfBNplzAgYAkv9wH6B39SpFDYZ8xhVW4Oo5BOC1BTMZpTgsGiHzSI2VZOHO
Tb8n0HBxOP6vrG3yG3XU21znaSnrqI9Cbf3nvPyiUPUxv3q03rRsddlmXzhMdCcH
ZLR+07LfrqJz6qj2/N+G4ZbhUltQyMaVbg+pgqSirSxLwZOA8aDuHxTgDMsGxQB1
+DxDOVLJNPCFQgm/p2UYyA1wKDfbPx/gQcPix3D0wSZNITDiBEWq/aiZZ8pmKSqW
a+yJWtjoFUKqXL5lQIo5bEX47HK6OCOvsd+qmCtBw0U4Ww8wwDs5XWkTg9UT6MQn
Xr3GM1qiYXrX1jSDnuxzwdUHqF7+7lj22/Q+dUYUNfR5OKG5nAdecwFBrDpvgwUp
EAxONCtSxPG/PmmLI86XezdBe8Tu+smoNylAvFwbWhKi2RJz7ghzYcCEVhz6Da/c
nePdHqAya+d4kx0A/IvyNg==
`protect END_PROTECTED
