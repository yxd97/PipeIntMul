`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umZ2i+AUqXrsHQNhsrtJaVA+7VepbWD/WCD1O8bJ8iqOYRtXv1eRLF+kliZrU0Ww
goQ3ZKtn5UuIP81Ftg0WRnyKG9ERBAj6DJ0ypd+4i7dgWI8Z9QOLM6jPLjUWJfIP
ccab0eLKz93S7kmN9x4ojkyo7MOdgDNtesXipC8jUnjEWTg1raMZuv8858XA+C4Z
DoCOwK8DFz0q5VSAzeFsvcM64yUZlYqrn0+4XPkqHVRbdvBPc4Gij84y/vO3A3pH
Syg+JVfX99S6JYJkJVFSMF8hZJTJ2maFKaPMDHUuVknLZ+49QDyXxBCbRhGRNMSq
QWrl5n+IX4/BKoD8PmCu0BZ/c5yOXBHwSFPmjZKK1cZb6JFprsaVo7qNPCFtauoy
3rLYGYcykbTP39xWEXdQ3bIhZIDkD5Chln2L+sBf4CikPQb5Pya/pyMuxMsYE0Oj
07Sqz66o5HabzawVB04PaNbgDaKGeeLpY7C54aS/x5HHlsdXPDhhUFnPwzfSbmhi
WWLml6M8cIjusSAL4RMn3g==
`protect END_PROTECTED
