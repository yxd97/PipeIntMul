`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6bxVcN7vYCdX4d6V0X6vUc8ggeZvxeexZajE07RPNF987Zt25LVaOn4Y64DVBVU
m1318EQAxWDsCuuI9MWl47ElEoMxOARPMXiDDGAQ5lujhtOBLeVvRyZJT8VXPwZD
ViLCrjABndS1YxHy0yzkjAlYwrgMMi88uRR5WzPEd51Ft3NwmCLKW4xNR6nZTQCh
7QtFidaoK0NDlBffG/G3+UoBD0zBFsmcb7fIN7FlYOoN2Kpurz37/IbfYpdgwlBC
T+XRS2N8rAT09iLJB0bVtg1MiEG+RZ2iew+YmXkiE2OOvxGfAaoHjrOB4SwdbBSk
bmgK99RNBFktZboyH5FE4WT+RXlp7gsr64Mz3J0zV7Ay35VvjG3pazgh+lu+2cSJ
SkDBk09zB1uwHlm4xnr2xXymoPSfezzJdUvim8E0F+Ed620MpSJ42uWSy5oSDuk4
59Ix9PxOtZifF4h2/2sSyI863jXhczwfEx0UEI8zC7Mxpe3FMpHMCJZFhhSKxxwM
EbusO4pTYCEZ1/1tEQu3AJrYI5JSXQP9gYEoI7OKahiJiKg7S03GnoIMeXDJd4N9
gvIVmBxXndV8a1gz/Mchcimt77F08l4VYotrrsqFPudgxGyrT7KNKN4Af+/mTc0F
`protect END_PROTECTED
