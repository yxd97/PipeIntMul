`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VyMHtcvefWgRwys7DAkMjfVk4Im3pomwoNIYKw0gnHoVD+9DWnl1NdpDmtQJ9dbn
M1L8VAult/z79x5LK7c1Hv/iq4PTXTXcPcyoML+prAU2DquEao4k/ZqcQQ8gezTq
mwD08wE8J0elNnKXPNFDxYrMFtJrG0jbztaii2hDcWfZqrmTPD7kV2Gubqclocwp
Le7vHtLseO/yjBGul/eQQjBj+FHcCQdmFhLH/TRxQ15XeovSMYH+DtCXBCp8DNGe
/jqV++hGFylToklTdPbwQuR5dTi0+Jn5Pb7pMMAoCh636HS3383Cnu0vRdZMvbmf
UuCPO1nw0s0TJRJVZNwFOIejyf1FCwNnDqWK7EDuOMaYNVQeQBvHrbV16TWAk52a
qjej+RFrV/GNSHtuqEQkhkLaTvEs/3LSaqj339Y/9HY=
`protect END_PROTECTED
