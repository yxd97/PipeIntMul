`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kselC3PL/P6MX2TRQUSmwFPPgz7GXh7znFWzudZyE85VA+iEd8ZKXP+KKDQR/XBP
S29c8mjqJwk4pYKXg5HTJbV3cKaz6n3XbZ9pPvw9Tw9jHS4tQdbJ0t2VbGv19uGz
9pqJymN6P6Y+EZ2MBtwjdl55nR6ZvS44S0lcq5avIs95OAAxzpUS4zU4N2bopxRc
L9ivKV0otnudPvwA+SUlYyNDpQMmizGcG1tj75cuVVDMiy5tDU3+a3gIDg+OMMHd
svpe/OoNC4JQA8tgdRD491+1DUZAFV+w8XyPE7ktp/UHw+VbVYffmM0FVWxbqsZe
ayVl0uzhc1Qyd+l0Qav7U+rvKf+x6qmDeAFp1NZG8f8SAftDkEdBO+U2kkyJ7HLr
hkCFzCmc2Zm87EK84moMIRziMICDc/LskrYoKusLY40WxnNT0bK8RxfppgNZPZYq
fMPzikpvyexfjF32AUVPeuFSJo6t7B24y+/e63eB7WFV0q0MDskAiCLDKG3jviq5
hJFr5kQNrj53+jC7qdL/2Yhg/ubBzvN4HkqiyKho3e3Rc/piYG5OZyDtXbRXyV11
S0m7JM1kTHuSlbQ5nS73yl3qxOX7cHk4wfbZJg6DV3ZLGkk1p7xnFoI5iLisD/Ng
qwS/KxmGu141Wk3f2rqXTA==
`protect END_PROTECTED
