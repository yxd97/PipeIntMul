`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qu1fMt/Aom2FKvnAqoF16ugK7zQCARn+F1iZcABv3zHhfj65HvLFEibASTCPb5y2
EBubSlJmxu6I0pptJpv1wttc9WPzkz4mWmoyymScjlxB8qjOdUyHUdMr+uVEvgWj
gf4qs3Vf94ca+NMi7Xvj5ox9tQ+EyMnCE3HBnxvkQyQSevwMCdg/5T085OtSVb8B
GEtotDH3JuYMeplB+1sHQJP5VKjdIwTIdHWi7ztcIx7i+Jm34rG6GeAbwh9cAV/7
B0+Dbnoc3upgQZjFT+Y5MVUQts3yWWLVOJqV0zIxxm1+FYWWB5QBrKtnCpK9sg0X
LTVYXWIIZqePpfnRtlqdSSEVbi0ETRIZyV8XoiP7BztU/xn6//n37Ujr4tCB5SRW
3iiTte58n3UyZzJqeGA2insUvrPOzV0bA+2JXUo/T2jSXi+ci/DiKfmuDGx7zKyG
e/CaWEXVhPMrXBuznUBNMR/t09U+7b73Y2M915aINtWJN5ltfP8PzFsDeyNPr0lm
fJJVfV8Kq5jp94uSj5LTi/G3tL0PpGnU/oX2zX0/vOD7rJpHo5eRW0Uqmk34m/ay
pb/eAbInAt2LO0RmqtHyzQaCWqfYUdvkgBrWG0/BWFgXw3O0Zm6lkihxfcZpRL9m
81hic/nVCYGmsEwSq/wy2F5mhcaLU5br4z0kGKA53JyaymVwJUXalYvZ+HbNy1/0
DKQNyHEAZI9958Wy3J2m1qI1gZGD+yA3Ycpf7yphSCT187sHusTVy1cHpFNpuifH
SLQ3jV4IVQdGNvoX5Kw6cO9KlxO+Sa5UobOXqWWu+lZkp2z5MRJS9tvhmmtpm1Re
a2LuscYwyPEU7PHtXMXFeTktSD9EdhRQHRxjr0yhS+NHht7mQ6zSmZMUjzWg1Cno
6v4M9ifsC8gtVnCDD0/0DPpRHcKea/TQWwxo7Sk/uLyVA+E3kL+e7/lHpwfQBSMm
HjrcSj677gX1Zo1KdVNLfzJvxIutfLd8PxgbME7hwGdNJzZq6bPzA4F+ci+Xb688
5hCW/J1abl7erAFAJYJxwfwn1Bap/xLpJrdJ/U7d82rnVwQZ9UHO3rVQ3kEQ1Yal
4vWKSleBjYPEQFL8d8mCLNzoqJpdBX+y5FZBQ4BN3u2/Vd6VjbwumOz7MMOB+pRH
MicCcTc8Gwn/e3JTSTkTg+MmFH6f2Fd3dkjUawALUbg/FfEi8D+MeClRX6RSE6I5
W49ah0IEpuuypsH50LXuxj3lBHwhisnkamyLoi4thvT+ddN9VJGFRmFBjCCKRLgc
+yF/5ZFKztHX+4d8LIYFPl5UlO/unsUDg+mk8fxysQrsKM/rdncSeSRvV5K9V8MW
HD+Iaq8FYNTxMJLNcH1+zHf+OcqgIjnneKWzKD3nshhNdcyNKTqmHDpXxI+bdvqW
5Q3PDGsm2cd/ZSTdIzjqbky6qhrHyeNGWzKiicG+5XPXjjRStqrWD9bjzR6pLOFD
Obg0mx554cOBmiQDhzVsDyGtrqeT0jXfK3JfOWvNwe+q7z8HvIatztmKI2Iakz8x
9ooPcx4r7w1UV1sk6kYGL1tdy/m58jp1GAL8SJMP1sIQHci8al3F50aJlZp6XzW/
5kmFp8lyuUbkOewc7XRk7sD4hswZaHGX5QnZvYf066BlZzaYebYJ8a7OckzF/w0c
Z1kcXz29aFtEq1NWK27MRVGIWTi7ORxfw0l4dJA96PYtGBySnl+V4GwHct+MLQnc
9xCDs0NGzfRSr224Cgz5BND5PjQbGKtib0fYmUFx5jGxexLi1X2twYMYYvfe1L11
vaDsBpWJBQTC/pHSkK+EG/HiF9PiqcFujRdubXzQsbbzrXm00hV8AINte9fmFRt0
AmUfpk/Nu2sJvOCX7R7hazRRMUidebeOEj7jPVoe6RNQBwKJQ9xq525DgG/PEqVQ
Qrz9D3L66UrHMLgGJ8gT9zog3Bfu17Z25gUpJwxIRTCssIrZUAKP8P0+Kt+1Jcua
472wLicudyvBfY+7/6FScgC/unhzP+behYPskGqrK8w0qNPsOTb/FsC3VSQ+p+tl
6jJK4lLkiIYxdXk9MNAV3Di3anbxqBSKPJAX0ckoQ/4Q82ckEESaoJu5whFF6fHN
mIF+XmrXX0BEZBUjEIfqsZuFGh7FIPOcIUJJGkboPKimOKFMpgrNxelxCw5pBDdu
Mjr8FaTxubrMQld+ZQKgmcSh9gunBBkw6AYRUpMaP4juQgwZ1AXxMB9qKB3iJoGz
GA75EKiR6fW/rI87IkWYbsAdm2sn6L7IreABMy6Jqe+4w3Tt3bduYBUhhL+LQxRW
bVtCvY1p1fWsAS4jgYA4Sq0/H7GWfCoM4fPIm+8E+5ZWTRy6i7wvbOsBc20k4e4J
QFm7ixPV400iF/onFx8Irku00rEVwS1wwlJ6P/uRi/S0b1pQVkdzasy6f+1uQvrt
QOIbn2SMmCyLG4dvdkmaR7OURU24GbsS2geX5+H/UB4doiUCMIYCEpAIiQPtlJHS
rCIEWc4wyIsV0hxSwS4KDH8RRyOZXJ30uYVg+NMDpEnU44oUSFSYYnOAodkyTZcF
AR4UBxLTpJL4sL1e2QvZsf3ET1ADZnJOps+SyfF9NhuY4AM7wBjM7Uz7Jp8mdleg
EcMoGFypen2C1uYB6VhGgjlAwrL024wd1D0L2TxSf2QPJfe8DW1hDBAuAvvCQtG8
ExfugoIQJYXxR56aQeEuWPsMDG5RvNb5nX4l1XGbFQjgEc+swVgwl0Az2F6u04+V
Sqpjw1EdFyrP0CwaXdEeGEAA1WIxaG37SOijMrbIayJqoxbiyapt+6vX1sw8un1f
aYYZqENdV7oXPaCG9dgUjFw/bMVgJ5WveawRBBkp14ZIod3SA9O4mQGpWNj98XZ4
jXt5qJsuXe7bpNy+Daz5JRjPriQXV5OUAVofecXjADLwYkxxgYoTWOH9crJ3cCAA
a64gpS8rJNYGHxTHotZzlQ44mviKcJN0iMunWmyncHBMp9x9NVq6WpwQTVFK4csc
ri0J8KE2s5Aobh8TA+FHG0jSs7g8ZRkOmYkmNxkis3qjgYKh1Z8/a65GINRb8mmj
f3yVq1ZUzE61ArAk3ZrECtboQjdDb43ozaS5IOXOX8Q9A2tPOt7Bo8CWqPy7H2dk
+vbePWnpB0OtZITLQLxErvwCWuEdUrb5vVtNhfYjCPeeyoPUrGTSrABUvLQcVFw1
dxItF0MRKbGhXmVkXjvnmwM3E3CdJpyJ0Fk1ILZmUea8n5g3bxriVt1tQ3rVMuu+
dsO+dYOLi/iTVZNpgbF38l3xO0No3cL/iW0JJKnmhwBdoelVW1B09iEsB+ZwHAaT
Ggq6pvW+gLZ9E3gNi2sNPhq55tixigIvelKduQlyjklT63uEhfKF3Ohy3aHxoc1M
M+fXKRI4/FBhoO4WHHBwssZFKI5M3XVbaX0LaGEmpTlYpOKal65lb7eIHGh/yBwn
Xk7CDTjcztXRb5EU4ZlzKFQJqGVN0y6mo2AiAH+7ZKK1fGBhWEdzhXdPrr5YIhf0
1EhSdOQM3kGloCB8Vm1cvg==
`protect END_PROTECTED
