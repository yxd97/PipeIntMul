`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZbBgN1l/GqqMRxiEjUZjn/3Tkj8ZmIMyxAfgv++b/uqyzqxeX5st7qVsThdaCjS
U3xLWF20yCmUGuu0PgjGNSt+awYWZ2qC+Sr9FLqzKFB4qs6431/+0iX07O51VI1+
zrSYs5bVGl9HownhzQP4Wqmdz2QxJVdyLtfPHVRvo4BcUeLugMcVNVO4VmQWfJ7F
bXelkwmKRoJLzHISp7j5g5H6mlye4kwUTwE2ysEvncn12hEi3F9ahATYVvwy/C6j
hfA3jp7cZwc/STnMrQjVWP6cqZCVZAzbKu51R36RgR/Yj0k3OXY3KpYV3p2gP7bw
1ItRfYq96qco7jFf7Ba8+HbMSkdoW+pYO6P7e89Y9tyuOAuJ69UtS9j6KzzMURxC
/DzZcrO3e1FG0nIcdqb9i8xADxwAzmtCqnlOLsvcQs0BFXfCL0JQ+pdALWMzvoxz
k9WhTnr3eWV6k30GeTOli5eMZ1BNuS5Jx4gotAKxudqloSCUWnv+XO2AZvfyUNzG
+lPrQaYzL1+UecWxwafLTxE/GKlzT879J0qyYX36jccjTl6ifieLQHZNNdj0bDQZ
OQE3EVsllmq2OSMS+9X83w==
`protect END_PROTECTED
