`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdwLy/4hlWOsyrCja/cE45tuafbzJdoAx5jlMiAhrKNS7cKD0PpOpMtK8Mlcz0aR
C5iuqfFDIiNkQmsHqxrWHkXcGS04DX4Hx7+FLOH/y8eDvAF9OwhM9IcTWxGvcebV
4H70l3Hd8gvSNC+LUFEKqRbM5tYYeTcypp+T8t/xIXvmnWUR0+Vi6zmX+R2TP32U
7TKrr/FYKvPACQ2di9lV3mZY1Cl6B/QbCObZsR5PZcfG+TaQVDisrjNQHtUPZ9d1
QrKqY2pZ7mUHrc5Nvzc/h6+TSnWYHid9ZvHVm8tKQ+44b/A7DY9+TBl2QXfotHHO
Swv6mBA7EkbZdT+x3Lv5GvM18JDrR1yphMFN2onz2N/WV5JAWl6Uzr2CE6IbzMoK
TnVj2pDNNh7Zk9Judw48XZ0yy8TDXK8dRPbwFnnC/Rg1PF3zgY5IH9Y7tYJGKuyq
zUV3En0j0FlZNU7OzlYaG/hdN9Mk/bPW+jMFpTgUPbTO0yX0gekNCGb3U09FS+YL
JL2Ha1pEAY8X3blG86AXcaXU9OqsJDKkqV09oLN+tvVHwxlUG9VroN9qiggN17uv
XkZ0MswP6o1knR5k/nNcFDiBKOcAmDazrccYAM1db3RkqGQY8tPxwYrxNLjG5A/4
97jFcFcM8b1L4fZk4p/Hv8cL/4LEFCyTV32+qw8XEnMgXacxK8yFvsI6je+EP1Qn
4DzNNACALpi2+uHfKGvT2SsIxoDRggpoXdrd4/EF22VsB+dlKzBhTsvfa0Ow14fN
KGOyrYlbgaoGueiBw355jpveuRq/Rs4c4Wlf+kTD8FOPkrL1bQj+D9nqH8eKf4Do
JDNR6XiXcmaHS8vpsgkikujSeotLPL+UmZefehViRf5T8g5l4tyzQ6Opehnz5g5v
G0mXuhCLYNgIynigN/XV2vLEQsKmCRX7T/aoQxmvZpOrilbL16ec6YjIHypZ0aBg
/0mzZJJMLFcPyMOGjeKTEdXWgiGFSJdTaSg02Pu6TldCzFV+XE9uqqvOW0BDE2Tj
7Gmhwr//njRl59x6N2xE5kKC71VI2YMOcOJVfi8RV+kpnb41UsP80Lbe3wWgMkm0
SQA4+9l+74txVeHw6ZfLfSg4VDsvEGPeZLOrKFv2oLJ+zkXK3p9220IOs6hVCUcf
KDYw15yu6Lwb1t9ebdwqju334ihD1aIg1DUTR7vOKvY7x9yr1iFIn0e1/goeu9/0
cFFdGhAizMmhlZ2KKYBoLKCkEXTVqGbnWic9upysWt/izwHWk1JSySVAqg0sDhel
G8LxMKANJGmMTZgbVK4Dbh5f7S7SqU7flDdfZ0sgI9TCyVEsivIa04hKsB9XitZs
hR+84sIl7abqQKRgIMTEpMSCIvHVtCv4pOJBTQtJq/wp+xz8+W9WL6Joz6BiJtbW
Tcj0p9jrP8ToSja4kwbKP0PW7XrvNAyiYF9N/rfysGk1rltT2HEUkKLQOKf3p6DI
nhO0kG+AWA19gHhQQ4lPTSAVHAxUwrCClequSthSOCg=
`protect END_PROTECTED
