`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9RBBsPLJq0iQ6MOwtt2wPs1VftbnmZzJqUK9tujMcBZfcXvgr3awsZDdwPdqZv+
F87auNXHbH4BGERVU2eHyyAYTsw5QqcV/lYtkpYBmBfnyw+MHuOZCR+6xTH1AjJq
Y/IBFnvDpm4ZJH6QJ6XaNlH9qehUh6NRIfQmz+9xdz+MSJprVSC6lCZlOA6jcP4k
E8x5kIzqICo0kmGz+30L+3z+dZ+w7GvmRQ5KzHsI0i89/k9VYGNmutC4PoUjvO51
5o7e54oIQHB3XNobahircEdqT6kj2/Dxdt2RfLtpItWsFsVUc8WIKtHiz8QhEx7a
UtferMfStPqktQFFEgJf2Q==
`protect END_PROTECTED
