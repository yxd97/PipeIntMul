`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PlERyhsCc9MvGDbhW32c4GTunj3FNXoyFtKgvH+229LtNaqlMzIXbdHkWBT0Y2K2
FDsmDANpVmD5MsuBRnS4kg8JG6c0h+QZtoG0PQGsVyFtJi+y5GXokVDOLOsFlA9D
astdDiVBgXETmgh6qr3fU8sxOd9qbPoK9qgS0exKpn06zx3qVl+0kiLpKpxn8SJi
hFXanuV2N8yZ52tT+GpC/toPtCVBSvtCyxcPEMx/Ngt5lnKm+NLAlv1vEKuXQPPu
f1kpDSnanKZ83aGVy8uI5s2d8gF+ixKYAYbOYd2KlwKcD7OwsBlabyC3QDoXmxXO
if7hnbs7aj2u4RT7sXT0ISq50mv6r3C5b9pYVSKgevCMV33En4SdZqe3FEo8aT3v
uEiao2dMP5/+elvVmKS7/RWpo5pCA7iy6dzv1wUAh9RPWDVBDRwONE8BQwueOJsY
HjgeUZmCNf5Bf7w3rZE6Hw==
`protect END_PROTECTED
