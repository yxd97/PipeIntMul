`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qWg25ubt8eG3l4PuHsmvx4zdg3Dxb96mNSGthkvCzRfahUMX5QyeIJOIPcKMfgAI
sRo2Me0xf9UvX1XiabI0eJ7+sFN+jHhAHbRbCFXRLlcCGocrED3T+OgraOtVUFmo
rxFs/snF/rHu0L3bpZOqA1KUFk7PyhLMwvb94hMzJ1ef2wJFbvl9k2flBrt5D2T/
kBGY87OCvfrCvLERgMRemMzTVfHezDHu8Jq+MIWFgH9gyzBL6afAxrlkfxGj2YF8
MWxh2XiDmhbbnmfOJhAZ5oZ/0rPH4OJQ0bdUlt/Ixu0rTnuuaOEWD0rJKssnS2bk
ZXX3DrSxTFEr8+/cUX7m61QxNcWiqemJKUYPSFzPujAXlGSmpqbGcHY8MwHdbals
UZB5mos1E5DlZlp/VcVoz+J0DaT/v6a2qjO1f+McHrBlfDbNKL1PJ36GsYkt6Fom
Zm4yMk9H2BJxiigeHG4tpJZ5loZPLLUspCtmWHBJy1q/JMJ5Fmz/FE+BqbsQLZ5a
JizlI6s4a014LixIsV6DITOsBCl7wqd65GVkf8dJwUb+BnQ71g32Y5jWMLmU8tL6
7tEIzBFkgr+RlPlUs2gjCJBmsF7Uqvvbup7GY8RI3bJCjjN94wPyyVbr9q4YJpDp
vaQwbIMCKGpJmKAsdIcIyWI0MTUBUrQn1J3TCaE4sbHdmRlx8h0y4wm/krzd0MBB
kiqKPl1UD+cznVJNnJFA3W8rA9oxZLzPHPL5v8TrNu9QE8otOIpR+sOp0EFQ+Y7e
MFq0OABN7OqS6lSlQgPKYZxqm4qlnD8w8LmdulYqAGyMMhbPpV9r5fKoXQwCCOUH
iDSOpozoXGsw61Vs8CbdfQ==
`protect END_PROTECTED
