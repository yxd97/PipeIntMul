`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VM/2cEqdgFzhuQ7YRy619gfkHM60vK3lzH3JV1uyidIrHscqY+JZpGwZTR1AOp/D
1mV2uGNzwSkpLLme9IANC1MMzjEty/he6LVkJkkkg0xUvjprDJqbJ18HL5ak+Wy5
2DVnzL8JFZ+SgU9tyEoXz9nGuH0/IS5UoZqVLcpxaFLs2LZa4ih/0QAqI1QeWeMH
P3mwZsLrnY1HTcXeSpT7w7F5b/bDwClNQIjPtbbRYQW4ZC/SIMkmvnAF+ktFFv8m
AltCsHzfRypfTi5Mrxz8LtbGpEx+xWiByPGGNnwaxH3u1H2+oE60CVY/zfZbiBAv
9k1OhGgZp4HWI80wvS6cjF3wjg5/W4Xt81LAenRrZ2LbvwMImGpdKQBVHEv06mwT
fxeAdOTCA+a7h3VHz2SFV1lnljK/R1wpgq609Qj34pEEaM3FxUP9tWlbvesA4nJ1
v1XoKyjZeZ0SqG4gg3IUxVMwfaWFT7e0oEjCWPcbT1FR9TmmMecGXkwm6oLzFZgQ
/wNvQ2fCZbLSzGQChmOgUMT3MdlJxBLS+U9fku2udhkgaMeuQHdw2eVAwLfXAbyt
1G8fMdJOB8uxr2lUC/QdxPnYM6lyJ+67DOg5hOVTVxj5X8ZGvrVMcd/mkUCcHY7m
X/gB7NPE3tPWxz+hMWj9lPVLC/3Pyvo9JBQx9VNm3S5vZIoyVbt31NzIg0pHcyVC
3IZzn7Y1Q/GMPYAXJ0FYqhGg+sNOU8p7+msG7ea/ANTJ6G0Yr+Pt7p7+ech3m92X
iZsHAaoYaKtnhEc9KBPqxw+yvzN8mhTvlqNZQnslEhARvWiSd/6bznvTi8GCbM9e
iWpv58Lh1YZUCb+91K0EAt+z6PmGDpn38yA/y+M5kCDCPdtrjdooKU+CxbkKz3q7
LN//IPFKwEDutsJU0QOySsArmFBNd/NKLAOLrMUR2a8KtCNO1sqvgTdje+8xFiu0
HbHAsb+jOEazxYJ8Isg8Owa3mBdk7sOfo6UPVDfS+KZxj9h/fP/sAH6SLRw0q59I
Hdlnsbl/U5u416AR+JzJw52H1AGEdq9Etq3jwpNTmhV4On6MIm/qLmiJvRzwDobP
1B7cwCdu6M2QfmctbkeE3HSC90TtyVHJHJZCaocpbvWMfLU/AnqEOoTZNz7aqSWj
DFPeVRmzhGzO2xxtdsllQl3ZOenIL+c9J6BDubqQAIi4pY3KXVhFUyalLi2CIdkT
BgI06EI/rlXgC3XGdWhkwApCvg7D1prJ+CA7av4MPLnp+XCeOb6QReAehSpijSLB
Rkfh9ROUkIl6wPG9K56m7lA6mkFLDJo3fPAr0sdzD6X2D5rmog4BsTgG132p8hjt
rbLYGT+2z/d0cCHIU9dja6e0K+IQlJgO0zgrEl8gMUk7ADqet0TiJJGUEctYRjl9
pz96xoGZ8lQbQUn5fNphBRh/DiaHLHY2b/qC/x9iw4PWO6ExkSiL1rZJX/yfSIwt
`protect END_PROTECTED
