`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ykdxww5b6oaUVgr6XZa+T5xwmAQhNGPWFkowlgvTyb1jjLOM/Sp0xeo1ctnGdAyW
5CjAN/octp3SquOXjcIex2dv8DzA4JpCsRB+ywRk8KPMRujl5hs6w6VyGRFNHN3u
fm1aUt/XMu5PFtNTUpjNOqJzHhI2yp6+H3uWDmP8GZNINgIoHnE8/N9YeRtCBL8+
O3XW4/OEB00yRYQvd34uX3Q2i6cA1j7GAimBNK94xEkL6owIupOVtvRTCXSNAyma
jSUl6tW+JfYiBaBGMe1Ok5ga7VwoaY0L+6Yny8tImmjRRCMrNtFQoVzI4AQAiZyx
TpPa4pccMGO5Z3aqcu+jfx/He2gZcjd5Obccli5IUfQuV1CTV9y63402BtS7xVm1
7+qa5gK/ZGOdPWoqg4a0pg==
`protect END_PROTECTED
