`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFSuXziYbg1A1exrE1iEyVOCWyzxU6dWuEXPghLNldKae6ZALgloWvFQsYVbBO/S
w419MxmTuIIIj0vi1hgUpHbtREnI5DuMOZHz9oVeDnNMab/KxHypvGLlOchl9cQu
VLLnj300PZCGD1/ZU0JDWzBeOLAmPnz1AqasbWcFuDdj1/Ms0utbg4OyRjpACU95
tbBVAVqMLj6fAJAGEoKkBfGCXZLCMe1gRJ2RWomq4WtgkC7+IDIPJmKBAlOZb9I9
jr5kgCjKRagPscDWcIxRLw==
`protect END_PROTECTED
