`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ySShHGpOqb1gIVXrHRpGBK2FRdPqJ4RCoEoQEPOGyWXnBnOlE7CeWpI12TWediV2
6Surv4MjOPlFodHzbxqWgMVGo7NEgxoRwsdU7n3hch2yUIlkZJG5UnrN+KNeO5om
qw6AWb7+aB1q1TlSztrSi+qjXY9M905YLYcdKU70C7qvetj7YH2AiN5UIa9PD3bH
vKrFZHUAZGOLyikLeHTYnCBHF5pvsKrMgFhQksZRUEHQLnWrRKYLtRHWXr5VvOHz
Rqvkp1a6EGn/8GtH+dzeZIcGQlEYfDJjsLMIsa+j5ds6xMavhmh/wYlqxT2cIGJ3
`protect END_PROTECTED
