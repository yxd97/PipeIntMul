`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MGZrKsBz8NDRgEOzXh7V2NwgpZpConTwxKDdu5ZkXDs97qs0rIB7rgiNQ8Q2Ljw8
S4SJ4aONa8zzwT2OVL498nvEUpuc+lOs4IOitXHMiv8dAa0q8fuWs0xiNv7+BjWw
jFaKaXlWFHYzijczj5SjoV5kbWHfHJo9Y8daPmbAecDJjnPlMm4+QjXADm11ZddI
sxqypapLI8KczUOwXvnKOUY9wJN96BS++yjizSKiUSGWHSZ3OGKZRQZYfffQRKrI
Zd1YYJUktOR7grZfqMfLLK03AXEeYxVHsxlnEqO04j5RFlyliH2SLEyhj4ucEWVb
L7wlYpCHSIEwrZmMHp95KeOImGADkO5B1b4ET6Ywt/peFc0ozPmpkie7uMKW5XDB
3PLshZQWb5R61lMFQAEUhw==
`protect END_PROTECTED
