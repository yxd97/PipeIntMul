`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aezSkvfAGjx/D0NrowsQkkxhe7k8ilE993pTV8J74qWyWV/4sCruRT+Eg4+NlIS7
42wMZ6DFfOIuZ+U7IiS6NIxLJCG+ZkW7SfUQtERP0V75O2iMtUqosMUGt3CIbN0a
p64EGPFIWYWdEiuITQ9XUTfRt2/0Ea4ikv1NPuD2e0muSoPyZ4LcDyr9a3yRGARt
3Qv32o07hOaWi5pewgc7aq8hPBN680H3n18kQKDo93b/KgWsZZMYu+YhcaRG4+Se
AhpRLAR82d9kETi7q1o37GCSGZp7agihAOoRrsY9D/apnZ2YdEsoFK89MsDQRYMR
vFZ2Wvy9taWO4AFIHHvFqRe2wvpZHZHKzZASVqzpZpeq28Q5m2Q3j6NVAuWc30Ke
h7Ugf2eBpwb/reUSn9P1HwV+s812ueFSneg723tO5RNgoTrRAL5m/FaRBQTS+pQM
OiSf9HjpmH1v1Y91WHLiASiu9HXZmWJp5gf72+LMKD2N548eUrnpKZ5TObgJILmx
c3wiJjda6RTz6Lz78zjn/0O/ROXx0J1RcOihyTVA00Di+0vuKWyxjITcwlZPRSTo
VguMmqdkuRwuuFvLsdnvc4NcQ55jdv23X5SPB5M5ZsQ2NNYPVoLuLRxfmy8YpHQu
TrPaFNNbA6ZErNkEyQgMWL8vgyS9FmI+a/tfjHB9yZITFkz38kpnjM5PX/rrTSZJ
wfxlesemeGDHcJFhrLe+H8jdBMWMSmpJdNEVw+e9JTW7+ue7a0P7wSD9911bJbjt
9ajNmIwdXnqg56OdUQSKIRCUN1aRj0SWoFDaC8c/Oej/CP6uUTc5SZBHP0x2CyFb
HmsgfzA1YDiygfwDI/upDdfiPNhsazzISr7VuL7zsDfF4wtZfjwWxuCsKL1NyCSX
/qW0f+Li1kw0OiclR1I4FZP1pXmPFDzXPNFFcFawCQXQRNRs51cAgGQQl/hU61O0
eoa4Oj92ZAsJi2iXJe9mqhOtf/jJitsSnw6ntJx+zQyASVbc/eNt1tTnPPR65Qqj
R0vDhI/mhV+VB7wDKuZeDcFz8gauDhWfiqQA5ZzSfbAzErexob8HlSdhLMnqxOIE
BojwffrjFv08Bz3KUGt3Eo0//nSZTghjIIjrqCOHPXeeX8ztkJQB1S9c1L6VW9J9
Cf22z/j2LoM1L26PCimAka+7kYGtOwj2gZlk2LIjYC9tfET+Ed7ZREwAt/PAyZHK
felnl4lbm0+bABOhWAEvycPxM7RwtMEU0PRCvDEXcU95Xj0Le3czZ/ClcnpTwzm3
76wn9KI7RCxLfULXc3X+fWtJDRnPJz6lgjSrh9qU3XL0pu82ax/G/licIVu+yo1O
zePLk5SHWMDAKC+6M7GpIhSyDJrjovx9aR7k63yKkFNZ13l/QIwVN8yKb5lXTdjN
M/w29+/ACZJCl1RxcYlKzVqv2sXCKeTi7urtHapET1jhrTOhOVSLMKIbc/AAxeFq
UhFQgplvh7QeUgWWoTedDgXAFsGRwGeiyj5E74gLiuaopB1vtJON2VG0eGYRX6Nz
EcqVNns86xXeDIAgOlkfqRbf7r+xwmWEROos2sWMabfMQDBb7Gk4dE4cwrMo4HHB
mlqhwNQoCZrwVQHzzNF9D5Yyj43dcdbn63EV/TxUeq/j/QRo3h/aCWO2yX/leYC9
HTdMPan8RfRkioN1f61NkK3QOToA+glyXnBIA3i2ym/zrOFVG6phv4VErihDcWb8
6kqSd+Zz7j/gv06P4xO1SpLj6A0C4mqxTV8+8Z92lrHda1uPxEmrlmOsifsbtIRu
ErLjLozaSvLzvPTynQUu0eV5UxJoXxm1rRv+wbA1XnjN0lsVCVAbm3HC+AQnDwPK
UIL7hY9dgjL6hkQ6mScHtcmG3wRV72wFk1R0VrHsC6c31Yxa0hF8bKdVcpOAYs8a
hr+hEcMDt0suZcMZv6/KkQmccXKhRrwHLDRwtfqfylPg1vvQq1EGH9rxBb1so59S
SroDHonU6v+erTSMDZgHoVTbdsdgZrB1obw2OC7U0R3EqGNyN7s0flc/YitsjXel
bLvJi+TPP4i7veZBN2wUU980cmJJdpJwW7Gedqb+doATN8pqSUUsxAlmJY3Nsj9c
tlCZHj+0ehnD8xt+LB78OjD4AqkYNodMAWDAyKGpL7YIRGmkhixs+yvr6ZGGaxR3
66Svr3dcgoebjUhPT1zr0rcwJKS24g+pce/G6jryrqSP03P272eHbjFa6STQM2CQ
9VrENkCzI3JICTYCD4EiTOcHPW3PttzTWmdM/i+QpW49DTb7syzIKZsWXKjSUwyc
jsGYB9TJlpvR9a18Ep4S2LOHfGsNh3vYc8o2Jd4aK82xkDr+Q9Z9k3QH7nUTyL6U
NvROD/0Wt71Y32Vo8FZNkdcFM3G4Tbdq1fEFWaDpCYP+epalLbWa9JFbeM74HMZc
/daQDzHtwjLvpNfHJ8iMApqyU95Nch2pzGxUhaSY6FpOu6Dn5Loq9aaOcdqPs3ej
PnFC/yTK1rVCJ/eNbURtqvuJPV1i8/2DMRhqmFnlAAsw6+tC7A80uVgJxJ1xxBYg
371sdfvdGCehRIVWDpmA6gZ5Fy60WySPPe0ItbIA8Us7eG2RjIDCli4EVh+tmFA5
NBwmx7It3BTuMaPbTqix6x/mr4vkSoRYxJ7Zz/QNclWUbhV8vQ0+rLCrfdWE64bD
gFTVWLRUULmcELSdmgtxB4aRpBJq4Pogq3tKok8CyWYyEQ7aPU3Bi9h2W4lUfMiB
Sq+cO03KUnxATQP4pGIP7tRMZw88QbXEahDLqxTjVaJgFtSpM8Sc3f4xUv9a/mlF
XXkt0uzvceblzeCnTiKvJBggGwa5iXJimH9Let09hz38HQEPJAxQhUsjfixhB4Io
6SJ8rvm6A1Mgo+EISYdT85gnVH6e7gt6cIIZbHnIDit5S8oZY/sC8NQipLtqoJmC
uWqjEtO79Gad4ZInoK4YNpXVdKpbmK/KX6KPmVUjiy8hc84RfIL60DJhVenbu4Lx
UiCsl9PzbuEbOdblLDlONfpvRep4xPdGGkU+TiATJvG3yhgGTEV7ImIELtCUkAyl
RU+kFOG2HJ0RBFqz1F1e+RWhmVbyoPloLZXUbEI2FM8bY6OCfnp6XJ26a+0LTJ0p
+uKCV99UNru3eaL+XiRvsICka04fsB7BQYhB9KM2A9gcTM6cRDf3ubLGWrwmGODF
oDjl2tgPywqNRjE1RtFGfNCYkwT03clQ3RLd+LAcoHon4nG5aKSfmOvAyKVAH16u
Thr2HBAaNYuUtrlWmTFb13cfaDaXEdBQSEgXPeByXo6hqid/TV6JBlXEBo4NTLj3
RgJkxGdhYCf5aZzlNtXeA1eG7Ijf6Fh3Q/S9BIrZIH4tGdDdFIAtA56sv5ThMYh3
hbqAmSD2fxlHn8Y1dXL8clwRI1jmyThdFGpSoxZb3D/CJi2M4EeV9Ojj0oldbP30
lRmimT4GEReMIcuyvSt6kPmN/ruG0LOrPwrpTkWE+OHUTYiLapWGj7EwCGqtrtcr
rzSf375kwDTwREZXqKYJt7OBJ/jQGYcRA3d9o4K7cp8pUe/ji9a3lRPMxpM1zpk9
F8IIZdH/tK8iZetk645E1fAZd5TpQFyct0iud+IgPJVXKYXc0U/SEor1+EekxK3s
KDqu+mtiOXxZyen0ywnD0wwS93RhHrQmkudRCnBAFVGLvqVIyHdTXegS2yKorRQ1
0qNi4jjTKbnAdZZKqrhkFLg045GIAXkOPXWPcv7pVSKQSsH2m352SwkNoAg7NuYU
`protect END_PROTECTED
