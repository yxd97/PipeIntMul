`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BhZ46HlcEiVcnQcj9sCjlN40BxAZHvlIXdXpmAhj5Z7x1n3YFS7VeUT4j+3ecGBb
J4UX/z5Sh8FxVOOloY+6RKFUMado2RNxbgHfuzsqh/MG3b9yPhiDBMpKe81CWQI4
pvxnNewAZjlk5wIbKB0eliaDuhCXIvRmFZUZog3qIAPTiTWYZmdiAokjk5lFD2nN
0qmZYY0rbIMjd2AKAgMaz8QxWoU+qsmdz95sLdlohmtA6KXJf2mRxfdD81UBAAzC
Z6nU7CwbpZoj3bBs75sjPM6MQbdoOM0GdPt3Bn2sVhNTZRYmOJUgYhaYrouEUo4Q
`protect END_PROTECTED
