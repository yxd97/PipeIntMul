`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iu3KCuJsGV10XZhdl3YKea2IzSgKBR/owcEmaSHYT/G6orgB4aXyrpzX72E7dzes
QqasgDYYQp+L4dT5zWlcFcaAEQME76ImBIgVMHRqouHJEofS4TEIsN3pEjL5V2tS
R62tZP+dQqNtjcl9T7KRtujKvLUU0v6u0cU5b4WnxXLilqMgJXSsEwpSSBbP3muK
BCEts6gIoOHGGQFQQsYJHV3eqdTOO/+m06lLTaV7FexcIGnWawAyYe2LngKr2PxH
bJ6GsM9YvNVQzEE/JZEH6zj3L0gIgvORohvxKZ+BmpGHA0EYyjBEKF/0OR6OmeAX
uh9X7jyaUQC2uLt7jkxw3ezHbRV4cP0Nv8zv4dUTcep5iBq8FdPNVQeKq1j4v48b
RvvDxvrRSknx/msMmaJ7/Q==
`protect END_PROTECTED
