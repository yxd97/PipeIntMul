`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ug1SCjAZuF9kp+Bq50pdK4CFBNI6I2+/L2AXN6d4+JIl07wO89MkACCMzIeygkzC
MbI6SO5VTHXLKSzTZXhzFfk44RLj6QQJYYJFBE6615UYyxZ+OSL7IL1e6voz2ifk
puFR2MTSkweU7l4KWv/d/FgctMClBsc9HuB2Ugyvcnnpd8C8XkDXda6EG08EmQSs
46JJLVbsCtjV0W/o5iexD0KxODcR8/0QV6HRZcDtw17Jb1th9nOGVfgRimaqKjFU
0tTP26Y+l0USuwBHZp24YsxFZPOkM0Q/ARvl8k2e8/4=
`protect END_PROTECTED
