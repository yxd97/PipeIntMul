`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4V24zXfx1N+7gTuPdC8OS9uhFL8R7NObwpuHRqH3NTgq3h9NSZGcFonUgzLVK9Fb
XIrE07g2WI1ySWGD7c7LmkUxNZkaJNaHMrkQI0MUs2cezxF0o9j9IrKqrL3t++TX
YNcsrhNEq969mWCmPVUwFjhu3ayCgyKVgnZ+NymalbjfR1tJKFmMxdTlmJP4m3DE
NJJM6oX5EbpF/bQdyBJZFlEZRYUUm8wzgnDv2hQ/twictfgoMoJ/paFcBBl/CH3s
jhV4xSHrttfFliVzKHjLAIXjTPj9F+gCqjEeKaeIWD2EPgqRfehjIKTaK7aIZOL5
RJHqieqGApEivgr1zj597N2Zwp3lM/hlZNuxrt+03VboSSytplHmqsCvlWh7Dx0X
ce0WG5FskOBqjh60uDAiZSHaWR0X7kFiq9WZQkOhlfLr6POGOVWNTu1jIYUs0rgw
1fIGtubD5TP3WEVnDeqVlc3KpdPKKBArA3aF1CyYdYRv0tK+t6TL8kTwVKg7FscG
UCVT7L9KpnOSqB4DA5rKIyTfIzP/BqMh4u6b5kqX/ENrTL/Ys09UKY2ban5X7vLP
8VlLKe4CeWIRrmJfx9VUvmaqz0mQN6WwubQ5H50CGp+7o9Y4jsCf7u662D+IR1Ts
UZrGGrSVicagwby0fk8Gzw==
`protect END_PROTECTED
