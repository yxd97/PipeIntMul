`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pgXS+jlBL/vrlk5XBSYY4M4jRSveGgzRLWqrOGowIfHjjbsW0kt+r3FQ93X9Pl3W
0us1BI0F0PdFkrI8izKbXMw4vBKrKnw6QGVBcUnXjlHXHnrFWRaHJibstT/O8CFo
NbxIg4nmt5iyd4LgxAWvPSZUKJPMP31e2p6N9bZwqLpFVf3UjnbtavQ35FlH0tfM
doHCpjsCqm98tzw1Ivebvh8PVxA0nQftdGpvijuycFsAs6eFlzcS/yG8waWkfEF8
2oy5jERiCnrDxPCEEEJmY85sRcyWcopCWO17wMvMagCE2imIw8QNKqgDB6DzhxJR
sXG+0cIoEK3LPJD557ihEwVdRqrADR3uhiUak6lsmeSmws5S4DJr2zp/i1eiw1fA
hQH0ZwVuA00ubZ6ECvOZrRukhZiKQpbAQADqJXqDthBGmgiCrFnPC9AKekjg3gy+
`protect END_PROTECTED
