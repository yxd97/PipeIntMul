`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLHM6nuy5MeHo4+nviWPtS++IEan03F7FSyX6PIMWEDBPbup9NVecpususlXUpx8
PxXCJj3tqZtXgBtJbxobbWxnijVNf6cZsZYIyjUBH5NN834tAr7eqlwYoPet3uR2
Z/XSWYLdaPI0f+shSkfhy+f2G/wcB2exHiBiGoYjpqPixgZ9cukkrEZ4kCBnwQWf
2WjJdlEXU24vf7YVPamXWMtR69GOyqaiSVu2AYP/kJF58Y16D9P2lBTbFyij01RX
YiekC7vEQHEH2UCq3uJwNjRke05s9F6GuS6cgJnQIOsCGWuTVCx40xB0s8HPK7EK
VB2iuxXUbbV6FKR5ei0fUDLKyGM1chf++DV+5aDCnseFbeLIt+4VWbgQ7NqHOOkO
v4WSSkLp1TmKs9SlckRiqfKKrjWU7pPKTW8veVQK3gc=
`protect END_PROTECTED
