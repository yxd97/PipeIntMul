`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HObSBXRnOKU9zYeHW55V4WJbFH3tJpSrg0vof6l2LcJ5d+SDkiiWD0BiTWZeXJd2
qU9Fo5wZtZqCy8PHzLlIKW51VWF18AezjHN23V1JJ85JkZvIttRfzfYvokHbTFZN
45vSDDNeuo8+0uNFoRoJdl96rRB4r0273zcEvJCxVlMXKp1eG07I0k/C9qHqELRi
SrtMqTRFazf2gszcqigluiirG2stgWfZMKUtEwpIuDiznsjsmc0D6pOs6Mrc9BqK
O/X2Kk8Hf0QQebAP+41rWiF4iOjOHJ2nqKoI1XeVY2/mO87e8u+Ms5y4gMeMjcbM
UsddcZAdQXSMkPIYOvKOuYiNwyufWlav7Rs1AMk6cdiDl5RHQmhbfcHgGZVXTdQ/
P9uPZ5BaUVaTDUC+nHCMDMtdAFt50IPYzUykYPEw0WbW3XBBxGL4kROdlmIjQXpi
dyo6E0+mZlGLvnL62lg9o2oEhyajP0pHPOhR4jsr6AMJdOSzF7ljljOsSyjTWE33
FjrM6cEoVHNkjqO0qE6HgkDZP3Kwm47jAJPLS1rOoX5J3Ah597hEgYLztxkkFROo
Cjela7iVPumqQxtoYTk0Dp1zs9phppymxC1PAgo3uVwOpNPuemnASzo2d8TL2hxf
pRowqW3tq9R8BSw5DQOEv2U/VNPuMV496hoiH7pWFUDB474ScGAgb+bhCDmob49t
I10I7QXwqzkZSappTnsYHZksioMhKmdm31xwk3pSSPcW5JTOS+aFDTs42IHNxp4y
Oa0GTYaGHy64TexnHuNSrUmGDvw4rFCkBmxkQow2lME41OY4E4/5rtPlCmbVmD1b
LINLdr+6CmSVVRR4lkq8raeqbj0n9w+aTQsBkB/8bVwx3d/rT6HwtQGH2k2biflT
+LxtXTYnuaOwBQxOXhIYnoUgYJTksGeEEBpWjn1MC2aP+Lvct8LoBE5hzYi9Od7J
MMz4LEpemkrlcenBEocdrykMFtRWXXjY17gzvz+/xL8ppIiTM2zrLYLPJ4H5msQ5
mxrFLsJzT97ZfV4VKoXYV5c86wB15EEn85vkU71lKdobv1tmU6IA4wVAr5zpqMXq
WI3JmBkp5ojqpw50HmFU/Q3R2uPEClyNNrhsO4sB3+WH2guBuyhp7csaLVcejHEc
1RXI6yo/24A33EHd7OXPOmlJ/pXpSQtY2K9iE29JYqiFvxRhf5sWxSSWP8QOMlFJ
067Z9xuY+ueaWmdT10XcKn4bihDM+1xyCWhCuGgHj32dJbKUdLCMTSktZNJME3UY
WmV32U2NUDuNgshYkavMu1mi0OX7RVKWmft7bdzOqR/IRVqaASN/4pz/MOI59dWp
M0BSRrvG5s5SDY6fUhYogPuDSIes28Dgr5xS3FrPVItIXu7lYT6Rwscy6tvUcdlx
cqZNpvCSklUWcbJoPtam5pY/+1zwOKgtsHs+08jQXaOXOcSV9xQA7MAX/n1/XJe8
ZXCQAs+D5TPEWH7t8KFWhTX6hSx4fUQwMx1xy/02uVNJBTNXqHKTHyuNORHkEofO
GeUPBdqznGXdo6MFl5r2PpnwfGZEIM1cAzNQvUCMqAG/9RKRLO9bL3COnTD8Oebu
gXnnxo7fsl70gvma3I0pLiH1x6rJ4A3iQrAZ9ekUuT32VEifCkoG0VEnT0NtLVzO
RX63bb4wwhrC8Mm5/zpHYF0DUwnsM1LfPxDDjs17UuqaFk4P3eBA080sbdek9z4h
Lzdq3ma9zR0e0S71mcBRbYeQHLB3bQMagNXmOBCC2bdeT3aReAkm4s7oeCY4dXsZ
Sy/HlSCAFDcJitIdp8q9tqVjbLFWEn84BRRpK3UiGNpdRqmGHlJBdCMD/+Ahz/rp
VE1J9cqroWxyRZXVj1ldGFmRA4BUE2IUrQk4zib4tTczE7N6IR1ObgXRULIYAz6W
ma/cjoMo6NNsxQ1c7ZRtSOSrj2g9+RDpFJYQwqb8eU8Ba7OffJ5m1ap4OWR2RIUM
hkbjR5CAbiscW0ID6ToGG7mpK5rWMRz10a+9uGYpNsi4w3InVIH28Y+UbWMgwJzO
ahq6dqtN+caywUHvjK6ScH2is6IxBcHFv/2nrHJ9VWKXfS2SXt39yn+mByCv6hHZ
X3/AV/Fqx4jUfEzahL/4UpGioJSfHzi2DoBm5vPTrWwFa+VQ3pDeox9J8sscBUYs
eLr5H1k+vpbqDunIQ0suoFK5uilVT9KCCs2f8yURmAg1mYt26+P2xM3GfgvAgAYO
U1ELEcc+f/3Lw4jvAtgxs6yt3wSuK7z/nKMoP0XRmQ5qwEDgYvrPyUoZJZ99Gtby
KfV6LR9edQNRbPhTaa50YUgjF8IvI/k08bKWpNOqQtWBS1WAKEIFjUHAShJQD6WX
LtBWp+SYSOHXqnj6/jwtycTxz273ZpbMTpKXQk0bwj1rcONyq5/IwBC/II8/IN9L
D5HyHKCp0SFjPMyvTZmmPA3/OIoCk6poWU2jfHRB0ipg8SSLJj0T1Tf3RdJ5JIvJ
sb2PvDuMNFYxVCGPJijIWq0SBEedVaPa1iarVkqzV2wNejvifZolrzPbSufXL+JQ
XZd3zqqlanW1U1NDUzVT+m6L8Yp82B1rv7ipGR2qlAK6lengOPhY3aDK/HOjLMV3
HGGppwiA8sOQ/ZS0+a+6/7csi0ZXr+doFrmy/vC+8wrF8As0GDpdPK2CE3tRt4Nc
J/G3y9/c7N1L1p9LYWURapFvs4ui9WrTKGVU92skffUs1Iy3PXyKoiUMmXcNEG4/
NtyO8v/lBdEpUhCtKTX8qtWUYGrEik5RFjD7XDHDrxVDPGlyxktfXHvqsQr0t179
rFIRxVAK/KygPZYuC3px8g+Rd5PhgPFW3VkbKA8Jmh2r+jG7RWWGei2PEqm7USTz
Tl5zSa3Thde+XoWCKVRRc4mj5Mvv835ja0c768wMm4aZOaA4zEuSJnxws5D5HG3w
+w7ScHaxvAh6XcPigz7synw9639bsqKpzuDGK4t77o0V+/soLPUpGJE8eyim5Out
Rjl0DtZ6wBtGpdfMt+uL217y5cSPGG/To27yrX0zB7ueAPZ3jKMEsWAsZo1Dmkfw
8kseofo+8SnFZxMq4Al9aep4hiVK/4ROT7C5pAxCJJKUPgCPdvycmlqkxfW0Xc21
Udbhge5PR0f8MPii69mlvhW+Xs5W4vVaoFwPDIk0zB6pn4jXDRZS4DFUYdH1wj25
SBT/6k1jU6Oen1EA5WNquh2PcADzre4D6GNEa6xkQWiqS5j346MndDmalhbwMBkm
WiCDka4NTvkz1BFQDwObbAa38gYKL4QykK1fmVNzNmldjKKq6hz4rAYGgO8DarHg
btOXusAnml/dxMa+BaPctw==
`protect END_PROTECTED
