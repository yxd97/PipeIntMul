`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3DgcChXYIP/Su39n3YBI6/41tImdNMGapigrPfFBnb3B2vlcSYwonn68cL68C7J
sIk39NvscpmDEjnkfQiXsuK1YF9nRZFgB3Ft89YAvY1yYV58uHdukPdwNh6u2Frh
81riL7yDnR3BVR6/UiI0noeGbEsShRw+jjGk7PyE5I01W7J1antFMECeSuSQrM/p
YZKp3yJIABtbXVScubeSr1GguNTIBYJYPNS+iUvKdAwDVyiQHFRa5T0KopwO+w+2
LOwg/XoEQUoKCPGURxtbzZEFA/TYejDequVxhza5I7DtV9hfLJ+VHwf1f3QrNeow
m/19WdoJcxhW6sfLpy1EORmcgzvBCHus1Ifwi7TPwKbCj+dBuL23tGBz9URh78qj
sksuYRFhTcRuSgGiO6ZWTNBSidyqiOKnbv+3xp+pYIzZcMbDi16FrwNH1pRVQnE/
gIHinCTzttjYHL7P/Y6ZnDLtlnylYQ6KAPXmWPA5mXhRITxT+gNnSMtq3AQfOD+p
TVKdwXZP5QVFKh+c46e5X46ptoj+BoXSjiaV8VUitpec23MV2EFnF/VsShisdu1j
4Pg323hmkqYz1TCAzhydMLW30D2e0E/6J0KnR3CtRVNFrH4KlpcZ841Hz3VGi4ph
CfHSV4cS2hwnavUO/tjJA8zvfdsCYXw+sAIGYMBEo/w=
`protect END_PROTECTED
