`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFp4ScLQEZeAtHV3hWZFiXT6EaTj7aTn7+tB7xspUdmi9sv/EAya8beMApQ0AXb2
GLdIQCHyv8wABPP9t0Qn7ycsUSsZBhNnxOWgSaxhrXzxcEur1spkRuQHMk9NFzWD
fsjig/SQzHZZ0tgiXsevqnRd1uuXItPaHYjav+ymzbOcqaUyCuadZLKa+k7QHYXi
uUOzcR3hwNe632dASPSqpeeuDczXohhlls+rROXABOl0dVdC/cY+8Wma51W7skgZ
xD6itfOK+PDtbasZAfJ5WsweMpsk3n77mYBk++YUhNUJLPWUXpLvAJu/XZ1r+pb0
W53O+N0os9klWloLRhK5xF7lsC6H8FgTZThd3nGSKyTQqBEeKjdQRDimlODTtvCl
hYLDCrTtt71VRR5sxKx9jrhuggwrE/uRT1CcbUO1KkM7Sfm7rfD0dO+q7hO2rCPa
YOG3EAyEayc3OZgp/NNdaO+/a6ySFOdXXCVuuw+rNGDslJeCaYQM+CiC52frICzv
vB8wLuc2b2cT+PLQAQl6kgjEg1zYUORM/1gEKqHg9BRG1p4U8eqMGvHCqNo5uXoy
uYqILwepys4Ywhp2vQSMbg==
`protect END_PROTECTED
