`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/ukxK8xeOxnRzknp4v5oPkEgWFcz/j2k+9Nr2XpJ7wVON6bWy6nuupMdiSog26q
gXxQwSd/14OiUjqJesNlH+gZuXzw5YCtAXRpdDFppU4WLH9FwjN/VU9q8fnFO9SZ
Icc7lZZfp4w15InIMnmVONrZKuNW5MnvunU/M++IwvPYAVunO4xK1VDZYiQEmtd4
9TsoG9daVe26pH+fG2D3vCOD0Vk/OmtMaDAeIWq9140jDQUOFoAeKnhhSTSOHblm
Ok26eI6XKC8P6XSfHxb+Zw==
`protect END_PROTECTED
