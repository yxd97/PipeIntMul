`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWFgCFSEGakVbdqwhsiEg9P0ugElo/ZcrKLk3s5pSrQ79TgmoC8Udn45+YUbszpA
Y7rsHrl+YpADdBNC43dX5XDbZ7/l3vau6LM9QyyC2OPhtp2AbDDBpZeRSGXWnKIM
FhngF3hvA6EJCxxEbtUAiscwn5YvIuLij1YkMh4FOr+VkNTriEBiZltIXZrUk7O8
QrbkHGdo9/HNIjjBuGb0c5EnaykzyO3Z/gp5pKb5QBB3B/jSEwZZV76fS1sW/Glz
Et6YDvtBGgAOmViaRGrR/VjsbYipkk7gYSssgElucENF2fzw56fDQTEq1gNhD7mY
9UH2yYkEHa6q18bFozs78p0i2sem2YJOaA5QK8jkbsH83PrvacNKD8KHrePkHakN
ZptlinKnmUQ2mOCsOIQOkC3ndV+rV4lDK0OfXPCq1mESL+rNCyijDR+4V+zVIsKd
ZYaw8UA0d5fSBVpDvupyJHrJnidRENFUeqVdb2ghaVokkRcRzM034Ru2I2Y+NCfG
jYFcxNswdFMD9rPoODk9v82NEtnZLPqq6OaIAQcTvVSPzD+A5bi9IjjIoXoTSC4g
//jPbcHTAiJYba46naQnESgzW8pC/lxRQr0J8FTmdDw/WpTECtZT18cayBUsRGu+
lxfvJde7wvqdDLlasqu2JN43SCsNcB4jRxno/gFOQxuQUszy5zoXrpsWIHgUi5T+
wBIOf3ElFCy3ygm38ifgGpV9ncKsYwqKzuTCCDmRUDxVqt4DQYtLvKj1UGldP2Gn
9wtXwOTdc7HsP2OmkAqnPUdEp267yqrVJJGKJ9ebsBWOaPYBAElLPWQ2vpiAvgmt
pFi1zLHzp+UyQj0+muyhG+66eh/yCh6AHYJJfBJpzP2LzpVduQaGhhP6iSboAHPO
Y83d54UMuKR46ZsZgFIqevL6Mqsx2C9fI31wFJnBvBnQZSzOA/+I+c8k11Owm3zr
wQnYAj3pwThZzrgfsd8dph8OY4xvQtJd/uN5LLiI9AucVNWyW5c4GO+kk867646o
WL0rP6KgZwv4hRMPHTHUykh1iiidmzwYeh08Df936dpIrLMcsKoMcuV8mBVS7kE1
OZKeVCV8rSoTl7+ndvDBGillPf3Q4VzgPdcghE6Jkt6F2VVE8LDb2/WzIhGDJ6F8
+bfEuFZ4YpUyMc4fKFscznTh9hnMXQpuD3uaVH+Zo3gDGkXn4mBB3cdb9io3WtzW
Q5I7JCOs2NrNsi31Lapc/cO/bpyQpBburAqO9saQtfpGu8Gpxkstf/xXGIInGYf2
9K7QCLEk7jZTFkJtOWB6WZ/iPPCeaGgPOFHlIHp2eRb/GL9KHDOTnK0QTXNzn2Jw
HrcH8ta7/urgMjWJuaXYCwZejQe1akpooONFMgwkuT2B/9xzNC3aCu9Ax2mN0dHW
BPJbT8yXolkc+MXTlzHcxY7w37l/XgjlQVPCjHCFKP6dSkSN+xpv2rw/h68gUIIa
rZ8gWLwS4elygED2W4J0QE68GN8fXlfENyB6+JFrScoAtv78V7d3b6dwxjk9v47V
DmYOUULW2f+pA9mE3UkVAVgVJnch3AbsI2+zVzIe2WPaFgFIOcQoA1zA04c1gyQs
xVmjxVHAZYld3+i8dc4rY47cu6hcDx9FSPXWhw0ufzDwF9iEAfp8hkyeodPhbTxy
bXEziDDrfYYO8S4Is1sKs0EnpwO6YTDkSGgL04aECZkagY/YQB62DGTlBK3s514K
o7FxcLatDKupBpBNPYHvzPZ90+Q3kyTC6L6r1GE05hpX1u052ZM0WRtZyZY6RA0m
gZpRMrdT/fVTmL7fgn92auumYaIPUXrxksRZiAvlTpkJkwHVcjHf0jXkdXCueAIm
T+6M7BVQiRzY+bkkiw6mYRz+NNYYGB1+YcyhDUuER5S1RxHz9+phV9dycJvg9q5l
DtKygRWkYQkEQjhczwUcQujKjUMm+0ApNM/A7inB2Kg+IyBEn3s451Jmh9xtO8CG
Xn+WQJFLJHHY9RBgtQH6YwBf9OToOjq/CQMQ2l1BohoOcVLTYAm9KUxLKHrqFp8P
HcRkJNVgV/1n7Aw8PhoxwOzy7LcCzZFVJ1XJON09ZPJWwsrRHaUjCSqRDtb2ezJz
xjC/YwJlLp7Jy4kfyV/diQXN80ygAqE990B0e8B8EQFAq+kk/5J1tHOouE3XPMXu
IEE7SIX3PqqA0YMOOVpj9nhCNF8wInKrpgx5ny/DgsgD5Na6RitFj3RF6UEhGYpM
7XkMG0kMlWJS2lfY2gkQ6broRmEtYRcyjCBHwEhhtkYwiGxMmcwkuikre/p12OsR
YqwN2GHSIRgi/3DtM47c1k0oIXILBOB5gvxWf1WupfO/TM2L7aPF/qnGwbjr6oPE
X+OsWrxTVSyFAClTqXZkb36rekJjagiXLJAsLCHWRX5+v7Q5QHXXBu+MZY6q60Yn
UHqEE5RHTRDu0Z148J7AUM+EK5SqaH2VeVque9OBv3SpgEhQ8BgfcwkaXRGihqlc
4h0Eafn2xHxpA8CXR3aC6w==
`protect END_PROTECTED
