`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Srri11rEaCRP3iDoFN8EovEkCy65QK4D6xA6kaljq4siJx66uCk2dcdJDHGjVBnJ
9bXQ2tA5l8N0wOjMWcW+f25P+8nPIdECv0WB1aA1mHshTOhie9ODS5+JiH0c/a7X
0JIS+eJl/H6dVuUbEFBkQ4rn2IbDGG6pGeg5Q7pRPBPHz2S351dquwCY24vMQerY
B4IOC1muzqX+bRMV7tTlTWFh6I8s9N2wJVuXqKb0VMMDf1Ag7rBtwV9RpqZLrfxR
51PIuuwAv/2zWkX7AoUF7v1V0V0U28wgB2NykB2SRMbTAXRdOPLiZqrLJZUbAYz6
1pJklm0lLR3nK622nQVDWwtzpgDA6uS4YGSELHOcL4wr0EtXA2dsDBvKIApBk9Kx
o5o2cGyu/FeCUKuhdZel0Q0WL6TT0QFPPsW/V4N11PlKntZyKA2bn+0lUp3pYA9m
YFkZsYEntAsYoAOWIgzQmWoB4s/jHrIZ57dx+fbf5i00gDjm9TofiQo8ut8Chiwv
/yFP11ewXwHSKvVRuBXShq2TBHHYVRrgtzVOpvfAt5IE4eJQZP1mjiT9/ha2ORZ9
7TsccnT4e1w34E1634z4Cg==
`protect END_PROTECTED
