`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oFer8jnlRZTl/XN+ke1Jb6yvNeHdFt6pAKD2OddQJa8Lrzk8+6B2s/W50QzB43Th
JGz/SeOL9+T+sQ1MtK5d/gVxjHb4SpE1N862SbBlBkMtpd9vNOvf2SQLEGNNUVDz
wYNmXWWjomJv6Jsfhwiy3e4/h1rszEg3puePqWNsp7i+qH1YdScdo0MS9I61FM54
AbVzS0t06MYKL1WYUswTdxFzrR7qA8Iz05zlFJPRyKZgZsaF+JtBhoU6Ge8faeq1
8zOHrCke05ZSDMmpDnBD+I1nvqgCRGI8Tgb7k2dgvNuWMSTtadSuI7nGnGXHd+CF
oTcns1hnYwxadJYaZgYoTsSuEMZjId1B52mjdFbtiJIH2pKWnAAgO2b/XO5CWHix
/mprs5MEk990OXzihLldjifCsP4UXxx0sPAjAAaW8FRqzWgLNnPfmKfPEJCr1Sks
o9ehZ0N97O+cJzfN19TLGGLt5FglS04yofeSUipM7TYBZdST+qyuHIvx5dD50E3A
l6ygV1vaizY1AOh6ZQmC4PP2OdDJlaZ9Kf9DdeYMnU89MkwSqdrxsq+H0JvPCir2
7y3TCowD49fGWAB+7qxe6KkReZPvLzO9qmq4sw8L/3VTJ4HJk3jW5qOElt4QacdH
GGwJUFT3m8WNkMJCqEkOcaIYkz5LFjPIvVq+M6D3ywFXTBw8Bx7+0k1xJnUV4Kcf
nPhIqUz2hMH3anIWJG4BxL2kUTVHyPr4KlhkL4W0KO4vKN6z8Q/hNxGXK3m4qNax
Wng+pL3QSeA0/Wa/PVzIr/5K4sCVhfNLL0PtC+Jaci74/VLy1zgcLN+RqGPAoxTf
lMHlsRVboqBwLst4mNcaZtHcYpqAPUoLxgUrZjb9+p1zoc4ZEoxbfsPI+QAVhAUw
KkhFD4Hkw5bh8mNrbc2H0vvaqM7tS+z1BOhzXin05WfYByg7o2bTtp7IqZ+MARiw
jA9josonnXNS2fDk0UJsgzdm3d3uYKDIocsDFMogR3hr/qt6WuX62jki5qgaHLBY
zxRlW9+R4MlolWGc8gZnoHYle/w8Aevb458kj1J2ElCXArqPMkMd9F5/35o0b7tU
aMFCqmocTpaB5krmfZ0jbOZhGCoIAlDBQXdHJgVf0aC02C/gPpXrEAbtt0Au3/Uk
BBMDdn9a2J+GVt4y2xFS1en4opsSFt0H/Agysul66MM=
`protect END_PROTECTED
