`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aepMa1Blo73zAVQK40w//YtC6kuBrCOJnDclbABH1Tkrx27IChZDLUUsHFHGSyfM
lRGv3b/IrKRqI3Ooh7okErkUcVmrWw7ggn1qSv/UltRxFaAK44cuLCx9g9hI6dcr
zUa3ymlo3fQpkGqlS/zOtyRTnvPT85XldBKip0IA7WfbmFeEr0rdLrKNyvHc6BZe
jaeMALYVGt+nuDEejoyt3J3+OBa5nFWaQwnVc0SANe5HgTha0wb7eAnPU8m8ZMhb
IaOasUgC+UWBTYGukJpaqBwobLZ4VivYlXAjhF9rK/2i1t/mReMDPacymw3l+WQj
`protect END_PROTECTED
