`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
blIHNe7ga9AhAw+KP96MD31hgIY7AGBbAIii9zupdPV+BJhY7KgKYdHjrTqHymGI
C9GF0HBntJmYc2RUVVKkDJ0udm0YUhyZTUqNfLNVksutdjpI/Bs1/GnfJUroXUsf
FZFMDYMVyzY7C/s8AFf36bkJ5RZmMXh+S861dJ5Rw0iSPYgMApC1zEqtAwY0uf2o
nn7+JeZJI6tK6NjfoR3UAdAb2axXDh0u6TLcfsMKpol6DmoBreKjj8F7+xBCAMoj
/EMzFfresBUCdG8PTy8yOS5ZwssSC7uruhVOvXk1/GyUjoqp/29WTvNsHkiYrwLd
a6fQrBNF15rfmQFeUoFy2dNmziwamifxjRyrQCVSMZU2xHygl2Km/4rpDTFb4DBU
XNOjadqh1xGBev6OPbFFqaKFbi/8+Dh9x6PII/W1XHh5+TZUQga5fmvbgp79nyrm
aJyv9h2GKJu0/DLV2G1GvQjei9uLErfmQ9utFP4nnEGUA2VMxVlBVvs6xhFvkvfY
khboof2ocUfzSGUQb9WUx8d2Y509xo4/nDjlaUwt2V1bKTKpqKcKZCjuUZistLFl
IlLKlhpCdbioPvidQAeufj140fLB772LiHWoCHXmTar8MOjUuil2rBj8v/GXr4eG
jwwK07jeb1Lv4YCsBzv2Ki3cQj5rWwdK8Aj7rdnovN99No0LNpLgcgIXMqpYYYok
9e1XkbiIP7xg7U7F/CWz6w==
`protect END_PROTECTED
