`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2iKTc8w5RBgB+qFxbHoSdon8xM9PX3EgFOu4kTTMwiBZNIenx8b7x/eMBsevmIrq
Lsoeg4NPboBzppgEqAM1fej4YAdvaC4hZEiZjNSCwGHUsre+szjGs9WhoKnLte+9
z7gT/Gs+6VDnqVd+/EJ80dECXa2zkIsQXKgeCvsMG1l4dauuoZfwryK6qnuAEQUN
uW6iWc26K6fOHRKxPWfkzg/O6gtsziEwtsfPOXHij1a6GqXoDZbX+kKmIsEnrn+N
aGBJdhh5yWgCOU+7lcRolCFr1u/Lu5P6nPJRopl/Cf02LG9BjbmvKfB/D1IEThSw
3DOf6MtL2E3VffyhyNb3/26J3osaZismq1//hvOTnAdTCsuJstnpAP4JUgYFsIqZ
CyBT/45VMq77hsaCkIfETLQ2QuzGkf5kLGhxrW7Urk/oY9EOSCjMApfYhQI5IkPN
bU7rQgFbeXFDKR/wHp7XGAYXluaapA3ltKOAUsuX1UAQkwngV2L8WWO5U+URqDxu
`protect END_PROTECTED
