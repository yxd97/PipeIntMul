`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nWNcG4r8HrQDZuqwzR+7avdOprZtwkThUAyknRx0RfZPveLFq9LLbqS8JKj0V/Ld
y6DMTl7cTh50X8D/56tJM9kV3RoV+s0mMeNWPS82saGHuiUDqoNsFlJMBZjMRUMz
lwuAh6GCEMkp++Dgvn2rAQYCrDKjep6QehZ5IsZGxPBEQATgn3EKOy8V1a3tPzxE
7gg/N75pQND1XEvI/p4C3TRBHSjETSRHqFf1/GMOjjTwA/jALcLrRzHjRV/GpwOe
K9l/5rSmtO5D0jOi6vo6uH4RKCHt4jEoOhK5S+ynm9P2PRkR06PFiZ1J+3cRouSe
0zvp5k5oF+IrY4Y55RpqJ3BqeJRdgn9um8n2rzUZfI1ZCQPvOhTtpZIO1iCgdPQ3
B0FAyEyiZEKlMyc2lUPc47prSnupVgULhGTmhgZY4UkpGBTgIrjUvJShwcyTC3Qc
Weql0CBLbfzm1p3hj6ebmbGtOuemP15GO2NEDZjdOCqelSY/Q9oiSE8kghatBESW
VR15vZI/xb9OCx7bZTVGF6BDgxT8Q9pDVe7DEbbfO8fcE3StW4Zw0+u7uJRIUEPD
`protect END_PROTECTED
