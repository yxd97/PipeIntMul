`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bstoT1l1OJEQH1BjK2gTVwyGlr5QxbfTjzYCJJq22km1r7xB+DswVvPICOZqvast
zvPGizT/iDsU1Q5MNS4gSkoCrQ1hbUAPrRnE7+7ayjSY7sPyOLAEqnyoWUnqUyAn
nBFyxOC7U/sospBZfkUnxO74l0NCKYX8/9TwN5VrB2luhyK8PQ+8b6PB650u25AT
Co4aeBXae/wtqFjf66jvgTf7oFA3xChwY8xjDWOkz/SLmBthE1vRtn7RU9ZKbGU6
NVh+Sx/uFObsGAd+unIYDz/c4KpoXYENSFyOwRNc8sCuZEy8yXy/puddmLwJ1+iK
578h139WZTu9RI+uys6XbNKMpyY4h/PzIcGxzKs0OMX760paor6VdljafnWu9rFR
936nreATTxKxeBgR/Q6tVoO68nfiAQZhCSFzzkbeZkKIYr7O8sSych2HksUOcJyK
cPEPFjH9B5LAX/MWXwCXUwXCxiiPFItakuQCRZy8RTlZYedjzS/x/3JgfrWdCVXE
UvwYEYMdkFrUfaSqU60X1Mtvzmjca53+XYCvK8Y3rydcGnH93drvoZU3KwWP11h9
cFG+3odp3OUeqaaLVlWDhAFrksHBo+Azdoix/mc7JjKlF0W8d1uNxaio2c38Z1z4
xgQpNaDmn6VWMAVgcgBWgg==
`protect END_PROTECTED
