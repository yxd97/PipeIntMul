`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HoEGfMpNkEmFq3avpsEyh2uuUHwnWRauHzBb6BgGr8IcPGkMB8miDXLOUKKd6Ge
eVpuY2da5L+SuMVy0b9fBhjI6F/+KOO7bzjhM57l/CPxD3SbRQsM77FueRVIfIRS
bWktbNyHoiOCxWEiMV8n5Oqeyjb3PLyqq6WxbfI1/burS9qx14ittJVgmz3XhaKY
RGbxpariQh2/jeXXtiq5BLhIkphdrSlw5jRBa92nzpdjyWBT2OwfTF1dDMBWfp7x
L1h7EwIxK/I5a9pmxL0eWrqGvE5nqWXYIYftK6mYiiKMwU/fC7tfI7clyn61E8Se
mVJ1mVdoe5NYjm3kFm7eQKeB3CwjzSx8i6pAzscGNWUEPoVpVx8Cp6gbbikVD2Xa
bezFHkwR37AjYx6QrnXYZHfyLDDEW+20qGrYvmD2gOounv3/ntsW/rsJcpojJoEG
8fpRTuFhuKSZ7jfgX6GMmCBy8fv4vH8DZelPycV3k4oXEj92ipo7BUwDypJme1hZ
I+5FtfNOWUEVhRsY+rzR+uha16AuZu/CBg5VFk1NsnevoR+NGY90SwOjiaR/uqB1
qadiAtdXLCI0DF5B5/sDeOYeqpSlVDHJKdXxaIB+8yOEubLIuomTAlh6PFvTIEv4
l3G0eF4uJWy7ZnpBjdetBwhiLR+6smgZk5GCN3N+Ph24XjAxIlYq2QqfbHHetq0v
n4NkRSpCdbw0SUGo3hmsL7cFODmhwfQvNm9ndgCxzB2RzqgMNWTr1NteKlHpRuxZ
/aGwnQRju0oF3wfFmniqeqOHM3NJqxIFiPPYjn/KMxexN9ocO6s9rtXxRTJhiANO
XzhLjMYtWK/xIgNaMiF8FHSGN9exm9nQC/QVifwEYvnGYR8dUbjo9+Q5pqqO/C9b
CmRnh1PVCHvdPqubTvi/mGjHQvMwrLDjH9UgGUvsmhyH5hff8BHCyg//dAMd/h+2
wxeCZSOyJSR3aUYKlAi4P5XjUitycH9FHbVYBNQeLCloS0qMYt48wYQ3j0HYlLHJ
QdB1aUkznbjtAO5Lp61fUPFKYo3eJlUqr8gkzEIotXTR7wrE9Vm5B0WxDmYrg/hh
RbJvFxL0786fCao72JqHpgc5ve8dUPXEsRdPVVW3Q3Z+9ggOHthrQP54K7XYAS6c
2gmJFx21sJPLH6TOpUc5hFO8leOKswZVviqMEY3T/0TjuDYEc3RqVq3PURjbcZNS
tYC9h9HXgcjsD6hpH2wPK12rWAZ6DROEUXq14vfV5D6Z+SSzU1qXu7h6HqB2AThA
yHe+sEzOSClMJOfUhquGMS8ptD0dm+PC141nqFe4Wfg7B9OptfgHWl6n/RsFOjtb
tA4Vs1EC9PfWZlACer/M8OxY4UZg6cPDkU94sWBtPatW6823obXteOGfKRCcbaFh
OfG92YVus2RqNO7l0NPrLMGMEa3PodZF/mawmcaaVfBu8NvySUstiB9hVgNVACPC
5psk5qb5ExcDMvy4rfcopeTRaWJf1L9WbGovNa8kOE+7OpXvbCiU5FpUFgMyTB2w
xx8W4RWHyfLAlRn586/km7m6xOrj7k/UgoLJSRVxwAeTVPX5UdiFibHbngTUcXt5
wDq7OcJe6NjMFNO/88w8hespqBAOkzTDJX0/YE5kAwAw7zTuWSo9rFuUi0vw413m
RXVZpwo0SqeBfFVu+HhvxpfWUZgLrGkefmcsAB1HFZSUs5wiPK5QgWlJt4O2vdZj
YGnLNnW8nCq51U11PLE+ABkJPYV2iCA7TOi0+y/8QpK3iIVH5xTxLLb/5lnCF58m
vhbt6r3IkGw3S7II6a5MKBZsbeA84ok0SKNeVkDY7khtECg/FxLpFVHZEO26eTsm
skfa3OhxD965bUbJEn8fj8esou9O7aGn1JSqXBOmeg45bbbkIfQ76xK8s2bSAKrD
W3A/LQZCiOwgdlbQVtYX0tmG774boXq/70UkC8sFXblhaZt98eVrp7ZavfIJGuKz
S3xOSzAZuJjC9P+NjdqP1Bo60OgIo+78PIViv0yTv8NitNqiprQ5yNNFtNDeydH+
djKSWNxwpM8S/XMQhXnuyxhns3wBWqtQacfHW3tS0mFG0uKZz3NpCrZpo/rFtkFD
UYWxMSIvlct084fQDyumn2Sp82AAl4YJrWHf70rKj+Hxlm+zPyKYY0Cuy+WdHzeJ
s9cXycgUDJcluJuPvRQx7v6SDteYRceqapAmdZOoneEN3TtaPod/oUo3MK0V5SdI
7XL0ZmPT1eaq+XUVId80AQJGnwhlWycP9VE4I74ikxg9tI3FP9USOcLqNl7Ifstf
zfF3H44s2QyAr1GuWPiujypTYtBj7O8uwihcLfDRMq3p4D8cGBEHQO4wbgMRbW3Y
Y5LHooSfEjotebcZ04x3bn8zWXpKHJtvXdByOpyUn0Uqq1BFRNwc2BjwleN2ai2L
MUPqO2Zf+dS1hRvKII8EUreUhgO3kXxirm7PLIQupVzwCD27Pbp6LIPur++cOPrK
teDgFOAvOZRXNrNbLwVPZMo3rdsiwpfJc49HFrP29BC34Gu9dX5TWUDESmOOsOEn
cKuq0RNNACSc0Sme7sgyOBpCKVfYWZhBBn6SwX1KyrxFtecNCMsoWPT44+th3jhJ
b9kmyzhCLjjoHCxIkf7Jokkkwu6V0NGUVPabomM2j7CUuNeL6Zwq3IPnMJRgneQY
UQRTt6/0RVHBL51KhsMq2jzgU5qKfQkfPhidccsrYc74teHmBKUbeZ71vu4u/l1K
RYGwpi8ifqI6rj2Ds/++KBeLG3ltK6j9B7VdVnPAwL9QuY8RM8/3q1DVfgsk/tKN
3e05tIk77yjXhQtCMhUaV4f1vMUT5Cjdt0rCeZqb8ysROhtIrNKxc5+D4O+Ye2LK
rWOwRlPXlfMpxLzjH0syn058KNWWdUCqDikvz4zR+L67K7faIWdb09WG7BjwAZcX
YMnpoZKrhsaUVHcDbBGZW82LEIMmLvC/CDZ6d1REHKUQRc8QuzqSDT0dF4Zj8xME
Txv1brE3zHrtl94vJMD37kJjcgTXDmMBFPqLLCsa6jR5mXhfoqRzT4lYHpMZntSI
+OuYx7ATQQG0SnNNvsMqe9j4bc8ePoJnmbDNtZK6/vdYNVTcbls2VQu+uV8Aq6d+
CplZSqR7s7lzYuV+PErdKSvR67If/f/AV2n12A452iuwYxJG9UlYSRZhUghs7ew1
QjcFUxYo6nCTNqBNyExXXAgBF9OjvBvM8qlD4AQMdsiyciLXBzo3hUL6lButR7to
Pv7lVV1wacLHhlLJem08VP8+AXsluLAD58p9XK4I83h/lqUP7+00hwtXMUaavhrs
3G2u5o0LRWtDHrlUqTG2lLks7UZfDX3oVN8ihInLqJnISwUWhQPu4QMA76DN0Ybc
7GuBG0KfOMMp4KmYeyil1a76Qhkag2bWgTJzBd+vkByE4HgCHc2RYIg3WWfDOWTT
U8KvZejKLILNa8nUqFH++rSe6ZNzjbVVkgTzBYQCAPF6KtejvZmey72CkdIt0LjM
erCuJ9QcLIkH6MdSmu8MRjlb/QwJ01n4C3Uedi/UxED0eA4v+FpienW1Be+41foN
SO5/+vFSJWpDI8Tfs71+fpudtBfqxe116Jo8hS1ea3c8aFH4uCFlphtokAur5kfz
JVMmFpcxIsaKW14luOSt6XIBgpQWMXnVc/kfB1QA8l69OW7IiDy1t00L/WW9m7Rl
K/Ex1+6kLgo/DHcJUFxDtZ6MqryfOX/3FmVheeBjwFhukXunr5C7b8gWcd4MvzAg
LP1rlutv/WCum5WuyqFEk/Dg5DHg7eDiHvBABsrCXdekKbeOZMptO+R8HRsKLJqz
nbYMTua6J9Rkcl2K9F+KYtdQwqAU2Fq+Vbkxwit535qJ9Wb3SdjQPdqNm8GFxXcQ
A0LrBrtemWoTHrSl36OjUIS1Dw7AtHbEUGzy/3O3+QTA0a30LXctLD0Ys7hnPouS
nDzN/7iTvcJ60TUfZBzxII4b5+Ba7dmqW5NQiXyvT18CdSqxmLBhTJcWuNqdzsF2
pFSe6Zm6Zq9fV09J/bOu0KIXBK808xIcrXqvsDugzIvAYih6hgeqXx5/mF/Ko3RB
veRyLcbMoKCMFLRY9uUoB3EP9nYCq+WRpyC0KORrdOa1RI1lhPsgzhiC6FkroOyB
dCTjIYc09Y1/cdL2+Vnku4Lfp+bLnmVEfwLz0lUFFAmuavavpWQLJsBXcAJu4ofH
loziepWf/66Vo8krqujyDmogVfPk/aSSgAdf3VDE+HP3dxqZ78qIOMaUcjL4UyoB
KaL/2DS1xcLOZ+QoiDXLWFKc1SWo6JVNggTjT9H8wQQtjzvOW95HzLbPfdqRyBOV
j2Qwujz+EJlNI2mRkgnk+4mahWKDVoFRiUfferMY5Fdq+1qiTPRSPVL6BeGVBFJd
sc0nyMfZ2PEvA+k65Y+6luUe02VbMJWfPXpaOQrkvKmJzThnEyWVBuB/+J53Fp2a
H6P3luOyzks64UKuOby6Bv4lX5a4EdZccSVsdVTLqrhOHGLgpEi2Nvkla5RZcpH0
JJ1xEpdnOit0S/T/lxAxldkh3jMsRnZ7Pf6LMf4updy1Glu9jeOnglFrJTIBGUeK
9ZoQ0bhSIyhSSAaDlb9orSGo3aykqu8qfZ38Xzyfc4aW7nppGko+gLG/WfyYazHe
O+mC7hyvjsssun+VLicJ1SFoaiou5GgWnAFvMpfO62wOGrhcBJkfispOD+WQK0qW
36uYRmpmb3CxGx32fL+TTEiB/RnsqG5HL2+UHUQMcmmknBC1l83eQQQPla6kfDUb
zPXmSo2sQ2FQOh9SQVrdTz3SxYiPkJkbh8/qIyVImr5DJwSWHYwAa0JMSv1Zbzqs
/kPk+75xtUfw6iHpdjqwXgmZolVLJcgXOZrMoR86hpdfFx6ZETg85IQbkJP9W50T
DO83I5E8yot9fhHKfd9ZQcc+XOt7DxjO6MSO/DfXaJc7SXSmdeqQFt1tMeDmxAah
2r5x3sI6f9c2z2iAWSYshrXtO9gUNfh8kK0N7zWZWF3Y16NVtmC//XGNReVflEI5
mszMvCMyqYeFfC2gRqgl7+L4ITighwpFyTVKcFP9r0fZHE2RKpTksjhZwqKrj8AP
P9zfGboyuZ4+OWNaPy7fFSDnbyloABrbiNSQxCY0DFUxYQP3Rf8RqlJPi7XP/AdO
Yau2VECWMzbMK+quk0zf87rE4FCELDa9VLLXv0TkcDgxyc+sIivC4UEfo9ql2sGR
dzI0JcajEkZ7DIJ/jp7gKvrXKEghIkuDfrnzJ8/8TcKvOqS9u0i2d2AUeoIhgV5R
xQD+6b40LkMmoz0b3oBuBS3G4NDwLTtk/DjVDCDZJOqyZQvfhZOVA3zfmRTFSl4b
bAiszlGdTrvZz9CBgm0j8G8TizTgOez6FZGv7oPDrvZc6luncLE87mM8w9SA2R8K
3eiQdqul+tXz4MmejxQOS2GFwVsV6aAvRQyhPHogMkTQF+yvQCbqp6NygoZDS9dI
PLVXLOF6qhiEn/DPiileumnv9pDhZzed8cgd6eo9m5tFd0ZPmW9MKralYtPIh5Tz
hJchCqi1RaIQQDDF3SSOJQ8q3eVhapWt7JjzQFMBim1MRqVyHMQpI6PzergMQ95q
pP6rVVF1xIfT/9Uk/05/kVGieI9HVOdaI7k4W7UNwMdhX7EfrohVieWGTSQyL5dV
YrtakBYmx/oi6iMm4w9CqIc6ZbWID6ZJvuILOkCXCDHn/mA1AF+3bWzmzSsJ6c33
ospMbnGiGKPKwiqUgobd4h94iZs4uKempLONizOxi2qE1i+K1qZpy9HG0tcg0N5l
4/KbVzRacrhhm+ICOBGaevJcX5KQfPuoM+uJY5TDIN3xmp5KqR2rIhier/O0kkoT
1k3Sw1pSDw9/8Ts2vIKD62Pm4PM793bYv+1msAupiDOYBqE7fDLn6LvI1XCS/942
QBOlGHPFsOsCPumKbZ8SBwZ3J+k8DjIQTVct4xw3FLLQjIZm8/VVc4J1q+pb/5Tq
dUPs+jWZsblt/BUgoHEDL4MFetNXMmeNXZ06vbWipOszW8HVrR/fquStI22/Q+Rl
3GyMF7qNJLmBpa9Fht2bU4igl7MCJyOX3Wk4doBkzVwxnh9KNs7AT7KqqdD0hj/q
TPu52fgI9/HqTI/ucBoQodtyDmUpXqxGhc8zNhRMiMBREMnhpK/L1yIiq0PrbC4u
NylVjdlC7/6ptEbRkuDrKkIXXlKPQo65zn9T9HSeZWAs/zzSXkwtdiyYCzPi5CFe
GBlh3wuxwrkj6V2R0TP7F25V1EXZ300l5DoXxTL2ONrDvPmUhSFroecjl1zu5vpb
j8uVFioQO8qyWMrfej6CR4kgMPb1GfYiadIhpzKKTIbk7TDm8lHpkkR7J6sCvzzV
4usgIAUXrTioz7ghmtXtKvnt0gCg6wA+L18dWQoUcxw4+SugBESp3y691bFcgeTk
qpabwFuuruvP/xTFlpbWLG8bhrly2Caq9il92e4SeOPI1jaw86jMhfzFmEoG4sM8
IAtDbwX71xZJzZWCdJY3LLIMDieI9AOo8AsqiqaAOovfEKmy+QAJfrzQRE2GV/53
Uq2wNzpsi16LPNJeXs6Gc7nyU51bJQ6iCUxWxZ0xDiBlyEOb3DW2hSA4uAzui4jd
vA8IhcUJvtO7w1zIuOe0iRjZHwi1dZlC7qJs4xZgYsK84benLWLbzS+yTYH8t2S0
BRsXiOAC/KYUn5LynSzmxaPsxUaL4ydYidhW/MSAL5SCEqLPsKHTszBEv1QtBKgR
urTUnAkAE4T5bWeOzosYxWEBmLBKf4K0YG+fNQmtGFuRc1uVnD8p2bUvUywLBBWB
1WX7Og8349AR8bDkBHCWpJfN8nr4A2wIJhCGH58Z38jWBM/usdBhvmyZjq6w086W
i7t26Jyy9RCLCz1JVzQVymD3uQsKQ1NUBBR5RKxfbawRViexXQM9jj7DufPB93dp
SamojAe1aJ0pSWRZWsPfTvD6qbJUbZhR9NlKEvSGOyo+DycmQDX6tNL1hrGUpU3D
IUNZNHVCFhofGv7XMXHNR1f5yVwv+SgS/MVDx4UNcyLvngSlTdswAA2QhBd+Eyee
UWh5hq8hDgXvJGXRyIPbZGB3NAw3q7PnQP0TdHSEhOSn+2GdV396ySmWtpZym9VP
QtmoMRGI0GJeDgSU799wMDeJ1PZKF+tG+Is3tBV0y16Tjskf+Re8lI2ESMiD7IRT
nxfE7hBgRknOFQhKfipyYVw9MCGx5gz04wEknJkxFqfPNPsnYwK7YBIoo1myKPcE
llscVxEHsEqGi4tlYBhvQLKIwjNRFWnEjDKcgmfcMicwYK+DxVfGujsVungcDDvJ
xPHyyHF36UiTBt2xk9LY5VpXB2wuAFcY7br+h/xaur+K1f5RENqQRoQsjzQo49DW
/rG7qZ7mR18LRXMZ0ITCLQ7GTpFkUXLkFvQEgcjN5rKpv/00o4q+3IJSNpIbQxGE
+mtKPyHuL8vQ0pT4XNawfH+k2zAOAG46FOjl73lGBalyfbSu6OPrRSO94WDiI3an
6Wj6e4z4jGo6lxJMf1sJbIG60zKJNVMEXfPc+SEhPAmnSCfqTK51uxCq3otHu9Le
Qy5zTtHhFwq0TBwQbD87ILXOTd5EDJBT989gVgMgB0cxQpMU1FrGolEXUru/1RFt
PxkCjisGebFeKiYQaRFoy/TxugPu58HFD7lNIlX4SPmJA1/81LWSyPz8B2niYXWt
HedFhVKNFv5HpatGT9ohazx6u1M975AFUXUbMsVFmoQiplgQj6FrjOiCZdmqk0Rp
qF5H18JObII9mOeSjvULxLvQUT8UNNLzfGEoCvn5PoaXggmVeykfYDHu8wGw+Qaf
tkU6effhPcc0se/jpdEnYgKDJYF/yXNavqU+cbdZAbNBssYDFGKKWVUGxgADMSe3
0bVHYTEArmuiM5qSVN/UdyB16P+VzBygQJaVYy8oSDnESYrs1qaUng1jbYXbxaoP
3ngAOWDRlaGe/Q86wMxR43iXCMlwazXAV4jV7L6G0BcRKrIsp6ecyZcLsCgsTWQ+
zKtAuJyANcNGhmM6+aneR5FhgxRP1eMT6VNXGAXwYEoPLn8yh1gTRpFqWLCB9Vua
j2vZ7M2Kf4cxNoJQ3X5cxEqqzbcB5PYblvJnQUgc0D7Fisr7/2QoyG7MPW/zkbOp
VLrUGvVql8xC7F09x77GrwV2zPAYHzAqXSfDXa2x2nAiuGWsCcPVx/R+ZDaIPwNo
kQJlbi7D7FC6axfuQ4TdgfhK3f3TNRMX0Op1CW1U50rxkHVofRz5e5tszrRQubf5
RXyeDtLiRAwDCUJ5+izgcO95R5thRrNqTOaOSOr3fFhvoglaPJC8rf5wPESXJK86
LveGBLB+KQ5c47idunEU7+6slNdTrLHBgfPlhgjc8ObewzyLeDKav1TJuND8IN/6
CBWO8Gmx656dlko7gQjDfjPeOop3R1qexsngtzGcolsh46AHAEf+iqS/RYeZwPIV
xFkOV74SpaNjEcVDZgMBgvAynY4XyNtu4STiihiyxE9B0jIr30Cm/yNg0/mqmpCn
MYQmnANHWmGiHqCtqEyxWuZVYPA/yiB/vFDig3GUjIw2jlKvQBI9wDNPVEJh17i/
Ye/HgRSybyOBBHxLQD/YPxkM86AgbxBTIg5+0QIcCxCvUJGwE+bSsiN7Qmvz7LR4
os5UrunX8I/49CUxgFiUpHQ+HvOBwDAZqf+hF4y/na8bFUrpvQXFHBIdw3yDB7bI
6QV49YOPhFY90hZLarGTmN3IPRLWwainPdPiS6aoGwo12oAYeNLQmKAQOFvJcL0s
YyYutx4dfXLkaZO3aXYmGWgUPpg9tNAEeM6FQfEqO+NVKAYRWhZeYaoYPuWvVvCP
xcWehVPiTvAK9sbIPj7o+LXh673PdKeX7UkSK6Uz164IHZn1h0NzBwDwRVI99WU+
tj6UOT/0hYfmtbMLELold23INGyjGDh+1WgX/oCSahdFeWaX+132AlGLwYhsdkHx
aa4hrrhwwEsUs/zb2UrnqW9fZ1q+gIRjCD7jFwnk5nnOfdcshnOX2vkFOMclo3Pj
c5IV4127cqThkqeEwPMzW3rfddekAVlNl3KH7kGIoarKde07b/xYZW5gkxZvi119
YFiMd0HMAEqx8pm7iERoGdMENZihnXIjITrRgYe9qkeHKy38xNvVwzmLvKPrRClO
WnKday23tcR3SDYPraIdY01oNA1jIVXUwdrUeRMFKZRvU/5NtY2Ood6l4KDC02e8
u0otgEwPCbh8dxs/mm3xIWi/XViUYqZ4SIV7Hfm+QB1RXN6Dby93brCVUIGOwMAD
2ICrcAdVwAJP4Vrz5kVu0gGI8fftRxBVi0/QNRFO8h/geq0QPZsZDIH+8J+uGHmh
YQrkbmkM978/09tkHDjYRBs5LmxSKDtH4SZmx7Zi0kouKkocEAC38vo6KqOWUeIT
KCIq7ZftsxyTVj0LaPqtiD1Q3hHXIBWevd3z3iHba2AAy509biPhDRivk44A0mA/
RAO0HIAPo5ym551wMdM2UTp1EzzPUD7G5YjEs4pBheYgCAKUCocqcW3xp7Cjj6CJ
pOeirOVbcGe85Uw9BQyvM4tiGsYjv3DOOzsBp7Y9LdyF/jQCW4doQqRFXI18u6sB
K4NAoDN1FXySr5zkGoUdGfDnmJOPA8EYM9+Es1AfRb3dEcT/H26kKLkXbIvSYV5V
I46ekcXATY/wXGIBiyg7s6X42N2gAlHydM4TB/6636pXpzYI+DEX9lMO4+IDREKn
BU9tkhfXMo0oWh6lxt017QaSaxGuKbOWGv66MnnVcN3Z4e51wzb0oEltLk1VZYJt
k/dop6NGNrbXZW6UcoiG4p9wBxrUNn+Q5EsSzyomRnGHw3hJsEts28FbUhEWHUzK
ajgRBXVFh4B5S613K4C7DU5VKcLrHsqDtrro8CKNWhZI+o7TjNIDLN2+Dv7FhntE
Z+uu7Mno0XlUF9XYX/vl0YAISsbW4BVIm5q6sgmD2dps7DmZXA+U5P1KFHxVRVVU
WOvinlxm+JcHFaWgLoT5yZtqEBDVKSuCeKdjSpp/3nZ163ncF4FEXpeOUecfP49K
IvisGG5tGDttoidRgRxOxxyYqxG0dAxwaZGGXIvKI4ulr/t0HBbNV9YFMZrTj3oG
WAG//yZXXNW4D3eTOD6vkVug2OcvSg0z1b8MvxRC7lyjNck7GKRTApzhsWZKyf0l
T5T6mQchFo9Oxfdufi9D5jYfUbztUEX6nYPbZzq9G6swHi9PBAA1edn01s/ea6hi
J7JVqCPysO0CQn6ZerItnLgfARLwBrQ18y5+2RoDaxWgxbUCUMvawopJrg8X4uaq
KfARvuRTea7QGphyI/KaJuVZBDP5Q2LFCf1ObPw+R9XmW4z4Wvg6/iRKyHm3ICRQ
Vhp4E3vthoSSMRv7QttePAFtDqYMBeE3zKZWuH89LXnHvImM7ktoBm3EkFq2oFJb
80LTx5cXE80SzDccJ5HLZaYpAhCKkLdUw9TC6tfph2wKQrk9XrjaGCzeeQfnyc+C
L0woJsg3NPVf0WvywxZtVpOeQL4I0J3SwDmMtHQR+PZSEOtBVWchrWYVOLUHDVjE
BO2oeFPmWX2kktA+zBNdbXvlUzcArEK/K+wk4s7L7pzTRls05S6DSRZOBnbVGdRr
g8/Q/qWHeb8zopvKJNiA8MoYnuYy3MV+S0zfWgJh+4mvv67JZIJiUSAQ1vXZnfJo
qYJ2CmDQ3jvBZBZIW7EncXNfQ88JrUURRh7BwJw8NWTRTIlbjqZ/Ky/zd2Jrv/W9
m3HnPmzoWQ1F4Ud4NmBbplaBmDolc1wtWjj0FfkXX5s0nWjhWqfkAMzvMwyABjYL
ivL3qz2PUPwWJOkKhLy6RUT86WqBR5f01CY0KMaUi0DtpHoKWK7ziCJ/X5a4sBtH
0lHhl91O2DlsW92zfsiI1qtqGIim7jO3sr7mQBC5LYLQhvx1dWoxHo1S5Aeyaz8p
2nPPz1hvqBloDjXefuecOXdLaXPhDQVEyUtRvBO2Qfz4D/OBByORfCeRStj44QxL
qghiRb3RJ0gU/d4slcGPRnKB71PcTyTjOZVgbcRNBzqzgv2hoQCB3cBAunw43nYy
sOM7WnWvtFFXDn8hkBSgBsB0a2tfoFCkS+AXxps7aUs5/Ez08vvEPraz7hPq16UQ
68iaaQQPwGqDcDrii1IG/hs8y19VdlVdOU9WJm2RIhZK/vRjlbqQ83S1hmWfXIj2
PlGV+166X79mZdhEvmHN2spXiItxeCOJvwpQm6NO397Z1d/58/6i5zPreSUHhz/C
CUsMrImO6UzBhLt4Hk8CDhiOv53rnCirYKaBUe8LuYbZcW21EsAFQ0rMd5tCod5y
8RSON48SxCInFAc6b0ayn+GOKlK0OhFA6KrEbi26u6yRLpEaFG0uqBQXJb3j/Uzt
1b3VtTAOjmzY/aZ92cLNeNuCRdX+S/C8vC1iNkbWQ8mJCeO2Mcv9FS/HWCz6FFyJ
fNjKMydv+zwaJSQBwCtApgmtP0Q1CFksxOMtcrIg3wHHBkWaxl3gflLDhCBjmKc+
GMvSl074+kAS8tovjFHBmbm0CbNF+n9bbTech9fshjBQlmsdjh59JERzd1coiTgk
7iax2/o48K+EJNLJX9BBgqrCPCxbIo88rvgwnPaijmEkNqETf68N8TKzy9ntR0zQ
hC9F30rzO8inv3N9ctIiexoZEEtBlE+ELZI5apzaYAqr67/CNirx7jcAEz8khMNZ
b3r9LwP9b75Lby2SRSvVYUvyffiqmPSRC7DDFinwO6O8DDurmFO6iWrkCQvmyVo7
W7OOy/+ClkXy/hBwQMDo+1mh0R2b0up+B5AdKUUnyMdRvaUlNgCKu5TlDfrxFgW7
6d1RIwwTk7ZY5UxZVgggxZzUPVHEoCbMc89s8/mke5a87ittMcQnl08YetnPrVRS
cxP4qUBv6i+2YWrNuKgcPe6OSD7nr3MeC4YIxqnIgQuSoVEieHv1aXhnPD4LV85O
MpASNym+HhQB+IA5QI3Rb5a65KlPKJo4pUP+NMtLAj/eGNJEQtwtLw2B4svxyJd/
F3P1GcZ5FLwviJEwNc4DbiDtPpRlPOu8zcjuaKniVqueo3Y3e1ss0k5R+ke2vCPi
hZJOyr6lmG8BvKJtBn/c3Eep2405TtfLeGcz4s1BjgNZn/vjGSKOaRS+BW5P9ZLW
pHz0AoBRKKiukerFtDL1BhTwTbDeBT5VE0Xk0HgIO8azF9CGXhfZuRo8uBHBcTi4
CSeI9IEDQ6veio7AfprGcGubGXCYCOeziVNHX20TRelITNjE4N5ooxqehYn0vqo4
wzsKYW8yvF1XZdIlB37s3WW+WsQUdqYLdhPzL1n/LjmVlqyK7XTfUAVQOc5u1tgV
4eiqwtiv8cexlN1jsgOSbGqt2jPO3/zBF3Y70btng3CRWNoy9tY4D10xqrQ9ROPz
IdRXPeF2z+uw9/HFecatBQO4UIn30mAfRF7VcYvwD7s4ZWPk0fiMPmGb8OjkIx0N
W6/gj+n8ywBIiNQgJIXA1d/Amk6AYtjg36cx7Z1rhhUR2Rq0sYnyQpca54qAOnES
M1oGh9KMw03pjd90eHN4dW/HTV74R3rVArV26VHN+zMSPw1HDH9WTdos8Akp0u2z
zuAHw0KxHU41cL3UfBy+AxxX/o7WOBw8ZlwRu++MjuZDl6GgpVuxW+EUknaQ+Ryn
GJCEljWRJ7bWlwGqBtoRTcVkxLRcL2NbUkPdPYONyLlS+/v9XQ7iPHHxqMn8MO0Z
mX4EVPoNAL6M21YDddGzk3DxYbpI732jDfQmSGFszmdLxun6rbWbyy4P634Lfq0Q
DYSDWAWvIScfzMaEqZY7d7EuoHV9vpwmGWLAg71V91uf1U+Sjj+r9sPYAq2ha6k6
nzeDfm6y2/hvXYy7CPwKP2amPkpev2IIYKE7C5MZS1SRvi0f3ooLVFWyDuwyCkH9
NLbtZ4+pp6TBz7s5ESZw3rtvlYpMOrrxt4dDARcHw2nve7jvo5r7nBuUwrY6fZw6
BgCHVtrblpl1q7JkKH3bTiMn0lWQmAtrs7Kk8mEJVL5VVDT88TvPLs9HYMPTkyDm
wfdEH9F/WK2dz1pGOjYbDyQLRG3cd6Sun9cjBdRsnucoR7tmu/Jl7BND/f7q6Y1o
b2wVAt+lS2VibRfZ3xAadp4Iy+bUmOBl8L8l1Yj2FrSVJ1hDKFLCL3GSVRDQGyut
Ta7lZFW3kH535D0RH5+onMVeDZVTD5G6ZsQv1yRmVE7AOraQeneQL202fyp9PN9K
30ByXmBHbaGxHeo5j6J/2w==
`protect END_PROTECTED
