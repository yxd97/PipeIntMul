`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTv3ZNfr8+zqtuoAUFgmbwjQZV5SJgXH5sMJ6Wae293WLrUUVDaWjJAFNo07PfGC
IUP53FtFuY6Y3JVd1oQuTsCO1rImRvca6J3ugz3GKgcitvItTWhg1ww7GljRjPGc
WXG5k1uA+bjDkJZ/mZq3pJ8BaiiZpTc6kKeeJa8d70lRTGYHH28VI96CCx8W1pkL
gZ224ANPoDC6YYIMjxYeFTHimSDikGixOLfhbcy81jkLeOoRniKMzyExG8znPAjT
xQAPFinkJu29tkeUMRcYEL9mBYa/pSrPWfQI6t/74LsbiOPAxBFh+7a1BEksnFxr
M2YSbuL2XYnIdDCop1ZZgcQ+bYxev0Sgf7O8oT3Rvgit4yAaleFMTeRa//lg6cCY
AzedLnu0kk683UouRe1G7zXTHsBXlJ/yzgqNWdyWblFRasn/56ARm4iLc7dGxDpk
ctSJHuxLOokSidePyCo9+T9FuqR3sXn3awhCEcJFVMmlJo6igG7GLv1r6AyLyo+7
nIT98C+ZUYGG7pZHkGey8lHhQ6gBjVf4g6vzsRhafWd9V8o2k1R/u/tlaYYXKN8V
A7utOlfuY7elAz+XEZt1k/L3hXRdZwY6uzMAdm1bySgMiwoKZzFzEzjRqe+htotS
+xyqaRBiFtUsLhpHKASMO4LpOle5CMgvuciMr/ImyHs2d/S+ArzT0mL75iLHjlpj
jk1ewVx6uuxSd02Kj3/cBjzkuk54uzN0SWH4ooNP3rJRIYGienKlGAJw8dLIOrQf
yjYPQYFHbUSkpkkr4UhHN9BwzNczycAsLH8K7JZsZA8CEBTNert50gPuWP7SqVgs
yKdsfnLA8Uqo9nQba0Km/ohJsocbJ5UrwCpotWwNXujLwQrqGwSl38RzXFypTGzT
2/fz/R1fTPqvR1uf7n3un9Laiaorq3GfGjpwSOsh4RG83B7b4Hetm++//IEW8xCi
`protect END_PROTECTED
