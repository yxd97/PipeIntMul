`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WuoMmrY7fm4VMzI6zEzwbwCfgisv9+vwh2w2DTg7yUuN0qt00l9wZSvLYWG56s2C
OYYtl3uX9GGvbngF7ljmFUyPt250wl5eLgJRTI/cMGxRPGwkE7yEX1z8EhUxdJfi
mi0qm5OwVGWxtNL+zGrxaD1U3liweNuV6plSl/WYPiI1lsEzXbkTnxK/FdXZ6uS6
WT0zUUkKFuWkm2/GBxV61ixSLMVUZIJArUkfDswt+pc9tOq9c5Skn1o/MDlDgVQW
Xl8GDqxIIf16UiHjTE1I9/I7VACptbzAJxIBHq1ZTPM8xF2DbpkUFJscGOeRSrnT
1Ry3HR8WnUcc2NoFERYx7VgSi20kskx07JE0s96bWCX/zYAV3IjHEIwLl9C9m1eo
8BwATTjR/Yq5MNC/dhqlaHGRZcVWRemsprzIrZEni1cO9R8CGohhrqx1Ep6BVxUN
ucp9t7N/uPP/ANnRHrlqGqZldQw4iY9i+14n+N1d/sFoy0XtEnXXEOTADhS7aLt3
k8FRAhIgy5ixp/VgNAwVoy285rnt7/OqQEDjXXFTeHMN24G4oI1upSsZ41aTWujF
WK092XrQxIE1OXC0JdketQw5GIeskD1/lKOMH3c2QUhAVeeBkVuB30nTAkUqT59M
VI/r4xQD/KVsMjx+xfrjpYSV0eha/5WAwt/Efoom8F792VWhfdcKemTa0y93r481
8f7ppFvDj+CUmZig6707Y8G5kNkPNeoqqEnPGZAms/EyqowU4OOZDbJKz4/cP47w
mvcIeixHxitukxuv0ayUS7ZFMP5DZw09TGWlEAG2Jw+UwMlqzSBC6va/nJgqBF91
TDSsHBNOnlR2IdO5Dd9X4sEnoPuudAb3g7gZxVICq1wsxT3Cs+A9/5oFMCVnLkpk
3mL06wU2U0Be7ccLBDL4Zw==
`protect END_PROTECTED
