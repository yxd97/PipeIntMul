library verilog;
use verilog.vl_types.all;
entity IBUF_CTT is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUF_CTT;
