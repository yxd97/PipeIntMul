`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yAb4rQ/3pV92Yc8M23wFgyK2vMCR21IK+7WMMDW+CwGmfdwkTmhf7yKAifdvut+
suG50UOifX4CMopTTiBeB0LdlHvyH48Y76fU2D3qZ10RDfZpOCl+EV3r+R/1jcUa
mI7Qw0ASpmEce34yGI1r0ryUKFZOYAU032f8d4WHGlwxXdPgGaPAYxG6387jKTDE
Gljf04Z038nqHUc4rZ5ZQhKV1eYCfjNw4VGJsjaegr250UjbeaRvWwMPMC7cq9D6
TMjtK6T0Mw+kWp3udcyTrpXmvblAJyRyeeHGAc1C0ts=
`protect END_PROTECTED
