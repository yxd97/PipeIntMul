`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggoGQgVek+SDLysUGf1Y8XNw3wHcH891roxfHLp2dmF4BSywZPHdqtbnVtB/DPkS
0GwgjceKLLjKQlzjLTOQYVXYed8RUZSATWd2ic8ddqp/M8HAiE/APOr+GnAcW97K
bcGzxxtbS2VB3HArbFmhk7SLWVsW00VvXpKotXHOqvh5L0l6cMDiPfcRNj+LytqL
sgEX6uatOHeNmwDiMU2gGqJB71e11aIFhzjgjhmtmqKhDjoWNM2xJ85HeESDBNpb
q7oO625aSPp7jmmbd84TW0OBgLbccxCEJPmvNYD0QiTLLOjHJjEmZqG6KoKHw+VS
IJALPjWoLJpYlkGQ4i7i0w==
`protect END_PROTECTED
