`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fPT/N1eyJwle4DHFQ7t7WkhQIUpKfrlDxbZVP5tCZYvpcsJLl1GrTZKtGC3+/rp
a/rIfX71NeqPV0yKhiwg81e3X9S+6K1hdqQpvs3WSyrnWe1G8MzEq2xlKkR+/RYV
3Jl61P0gOIMwMmLRlLChmi+NjlPbQdkfngDWWPBpBL9XG8NxWx7FssdKh7AA48bP
W4ysBAZu8EN/CyFYnnEW8ZDErI4mAjaDSiydemD53ptvT9KN9GcfozrIZIZqYlif
xGHAI6b7k5mOX6AfZRVpx3Z98u4zUkCaHoVeGhHkjSxFtKOfw9FpUirE/EBHw4pB
lqs46i9qFMvGSsQ8dJnpDmHEP8PSDrq0fQlARy23jFEkL0CaxebCQyePWZNNI9qM
tvUXNwFav58TrSUME17gfri7FNAD/ZC/1qMXvMRjlQ6GD24pa6qs9CJu0GXRkMSg
`protect END_PROTECTED
