`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JdSgOD/PCHATEZOzSaGJOB+rPEfndhQrylp+FsPDZGEUTZH42IcoUXjDxzePHAE2
aEnCQmchukSoeRVwQo8W7JE9AIxpZ5HGlz3xNY3iCyL0nScOqfBCRyRxpDWZh3Eq
FaTUOGCt7gKZMtWCM88amKb/OyYkLcQ1S0Rez70zpfTfLztGmcodE3cbQxQKidrz
wOCu5tSiTzXj8Y0Be0V9l4z/XfohucjjJhdmDrkAMrdjDQc3gTmsrEIDsjyQpagc
6I1Ak1tHe4HJC3zGA0lS4dztd9hKYpBd46U12saMtIt9tyG1D+R4fUdG5WYWe+OE
mYp3dsX1LkPSmWs5GmSDQn6OLQGdzPSn2bc/lm6LBnNIIE3orXoGE1cL0RdFN3As
`protect END_PROTECTED
