`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sSA3Mb3trU36mkuecDyWa+DIRtCBN5tBV07/zg/qOlxs3AeAnpEFjPiFAmUZ6BXv
1mA4YRyMyqUqx6rIxxtCbjocsNfwJ1WikK9+qe4kr8pP0LHlBgmSUHmiSliEGLbZ
AOYXjARFkI2w7PD02kkRpopEBOlvE+xKqajTJ/yLwPhkMs/XIKeD1OCUJmaeZktV
SUFzBldXtz3k+ITSCphs5NjRwKjYgSU+ISF9Mfl2fNzBRhlxrvJ+6jCyYFT+BQzi
IHAiOM1j9yv6yme/7RINBxlKSVXgCpTMNLlDfB0whqh1NehGRrOrHCJ1QwtVySYg
b6oZ13Z4ibnifbzx5k3MrGydd7zUUpexGBgLyvnP6JayJmBc7194pKRrcvOlNIck
`protect END_PROTECTED
