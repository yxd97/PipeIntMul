`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fF9sTfxLBkwJK/2Z5pRN9GvCljALD999fAhahT7S1GuuhdJ5j+33b2pst3EUPcSo
P2ZU0YZcLNGg0nZFEZrRcVHcyfRHQEBnJBTK9s0Ow+/pUQ/X+xmU2uUEO8tCGnmz
xLhCtko7ogJM8GbjIbABhXSwzE7sOzVfPFlg2vmX4m++1WtXAR415ZXW1Ox0o94x
rpuJHlTfOIzznV9J8tpPXORXl3MbC6n0YZsxKXYJkWPzKtxGqm7c+FdkWDJ3m8c9
UGPJEIJLfrSsMjMm+1Gx/lP3ORs7U9DuCDXEeTcu083GPVBz8jIND6bMarj7DpRE
U8+zAT6Co3VcvQYorQt1yTb3mPg0nPn49yOuy3ezJuTP7WElRTiD6MibnbfuT1yD
6/+ovncM+UAB2dFXLgKO+kcfqs22xwWJ9oxklNAsBMHHibuN5QtzEjJCo7RCtavy
An0pS12gYjgyZnph7287+j4akyPc/7Sqjk6jJwvMslwSy9K283fvDEdSGyUhsdkb
E1b0LXSmpwu5x6U4VoitMA==
`protect END_PROTECTED
