`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EaHvbzIWMkheD1i11zaCGYIKT1t0t89ruBYzGVK7M+kCdiJkXgR2FSWobdQlXWDc
n/wAy2VMSFHoWhZuO2B4sdNKZd1wusRoDz9oX4BdPk8heAvounAdREledbh04Nt9
o7RW/IGyk8xwIPz6YjPQTaUp1GILVVfT9TsTthzCr1i552Gk8HHmzgRGkjUDuNbI
UvFZKUQ/L3pnWTBpfF/zRqp/MZB3XJ9tRF0cQFbvOCiey//M5/zSBBo7S1BiAY7R
ZRWDtbiQnUTub7XZErSotPGhmSpluT2D0IiATC3tkgptNW76mXSjh4AzG0nvswps
Mk0jR2U3NbfpyPBZ6F7mk5tGPDwztwzoZ+zRhLVMjQZj40QhdP7qdotW8EB+RWfV
BUWP/leS9Q9sAKt442/iLftSaVf3J8nwKsI0cg/W6zGbsG03Uw1OdfdV1UMa1Ytu
yc0x9EnuW7zr6o1bOkRyxAIJdmOVECm7ui4ZStR/zy7EVaXsA6LQqUNDPffnCdez
lYEpq4xxL7XVzDvHS78tEhJSQe/MCVapuvd3sxRcWRIZ8Qg6k6ENdfzwydXkzjmg
TN/Bi5+untCKxULVeMhKx8vt5fINQ6SPuR5oiwClznbK9O7JzhWsbdswKm1NHd84
0CcfdcmFsC7adG5ylaFFpS6xIy4EV4EBZCQn42ge1tzR3vLZYPN+esiUbN8KKMKh
ExreKQJGkMiWMaUcAlf741j6zKf1Xr64LbxwZPabG7GVjTKcd6T1lgK+HFj3eLHy
f4H18VvQeTN1stMIb44BT0kBvnN2zFtAj3S9OwYU6zQQv8eGwX4Mkhi3tKR35Oqk
xT8cj+BkyO7mYuUMZvbJo49r4ob2P6HWeXYkuFIaSlNnp4/dW39XzUiDV08UQrYR
YBAnDvBP8ERxDb6TaRRTFpfzBA/f5Q5UNsK7MBhc89q0j18XLzd+QvKtm1Pudscw
83670dxj9gUWFwq6mkwiNXkHyh2zbq7Jv5Ti/cYRadms4Ll3Dh+1D/BjNIscGte8
WBL5p19x06ME6oC8XDQrm4n3MJkLwuIXCXTyRpBcdXQI8meA7B/OI8YLQyrUgKLT
8XHZVokiGph7OpQyro4Iti6mqYhthXjOUifbuCkjeHCF4AV8KaX8Tfv0aStFk4QT
gZZlGAHkNV9W5HSlIq4NpbU0HT8L76vB25M8TLxKZh33qcLP/yLKW/HQXSicjiag
yS+Bz+NMsBhpo+10gXuoDixAKomJSXbpd8QO61ldxok/uCSc6h4lF17zuvnvNUb5
X+7lTmzzCWMZ+pa5VslBn4l4TRH+BToQZ802NdjpFlG0y/utAqBbtwACYKkPzvCX
S2bdQJbWS83WJcR4UfSa4T+U2HlNfY8ThIerPmDbDofuJgU48rp1VelcHEnKPTy8
jm+N5w8U4Uf0T6veZ65vxLNyq5Y8pJC8lxo2g9snHm7VQJONtBTY/c6qjxnzGPKx
fh9fSWYlmhJ17mnJHu7Hq4CvOge194nsKGmVckoUUZ+wj5hDJzBgvPHSewwPXa7y
5yzMxmRZ3lCs3YTw0CVEiI6LcVpiRdw684Qo4O+a//wPCwvdxI9PVJQllBeP1WrU
3Ldu1N3FuqJUdy86kIC0G45zEGemaDWMt0C1vHmuwEEFj80aGp2cjLrIAIUBOzj5
PjMDS722dspnJMmpT6ybYfv0eEoF8aq3wSPOxWBcrKZk/nQ2mhE6TG02ESTS2UeR
1I86u6nr1QCwBNrXNL5VUPnOPfkgEb7hSMAdxqp2UPsM8yDu49+GyAuW1fANiGGD
zNBNBtmfJAYGe1QSKgwagdO6kwMvHGF6bxbJdO4rkVD4bRN4A5P9flGYp9CJ2kLw
Ynhj5OptCxjJVuNFdDF9/aEuuzJHiDnLxTR3guXr/M2KIzoOkCEnk+V4OzJoooWS
+OLXw8hSVz/5H6Jc5BL2Lq6LzrPsNOKebcjbt78OIPNjLTw/orml3CNAdkwi1gzU
I6dLY3309Q7lrPOc0c2XmHN1wXpo3IE0taExGE564o0=
`protect END_PROTECTED
