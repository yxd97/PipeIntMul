`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C+BAKbdmah+JQU+3CpU/nHIVAaegq1AZuPhef0gYbQzB6xLzoXlQjeITfx+t0Lam
EOJn3xa2Zglgts2UedNmx4f2wR25dgBMRsJpw5HSTq1UH9ts36vPAJBgzh1H0ynn
MzmzECkdS4KQvptXMF9UV1T/nBX0eCGFX6a4Hb8HwfZo6kw8RaP0/6pNCxNN1MVJ
tjY21V22KwxIxwR2I6epO1wrWmy9BB0yC8NWo7hcl433XPXja27PvxDd75sBEoVE
l5nfN/Z8xIcD1zQAjxyN/uJdqpd8P78dk4lPHNXEiQatahlNk2xZizbJ7IXJ/vJz
8OOUC6q55KvOThasC6tChkMlb8Elc5sOM3txYnBKoaGqgXr/hjKauqYBef+8FwNa
Wvz6kskdRbqfLWZalNIt6j5OhYYep3ZSSv68AOFwJC7ZOB5Rga1HuTC235D2M1Zk
5RelULw5y/dnvyoSb2XmP8KHITZJhNAQNegYLsXGrXMzC/+sbZ9hJxAgs2689J+w
5t+yF3UErM4e0yoqDpjnKII/ZVuNTszE+qCwyEU0jTuxvzbohAVKRA+xK2YOeA88
jgI0PLX9/XsOgVwKlp9SwgOXW0NM3CiJDGVICjVqplE8Gf0jsCrBLlQqPx5O3wBR
dfL/vfPMXJaouejfzpl9DTCRroTZtiUBV2aAXP802iB3CPaD21bKBs4i8gsUfCig
FVJe4gXrsQSR3QcKI8zgXzJOpsUTYemYesNtcbubLLHT5XpsMEcnt0zVob5oPCA0
Q1Lv3PoeeyURYZEzSybZCDm6ex1/8GyJ1B4FzhY31t+i88Y53nNkolboD+tr7JvU
0zSfE8KX6/RprRDD5TotkUiuqp+R43nWiHFgaRBzAF9p5ixVq48cxPmHFpPcoQyc
w0PHxatnBY4O1GN3a/slNXjS/iRXeK4lp4vZAARUzkv5i2GQWQJ4+w2KbRpZNA5V
c5qZDp/YvcTZYORJB4dLS2QiFpDV1asZv3DFFeTsbKvuZ5N68JRbUBqxU2RuwJT3
eXd6KIR5KvsalVzCuNlOwmPYwacaVslE7smaRhRGX1GupUwbzKN+hTv4aVqFQqqH
Wj0OL3StM6pnCbxRAnqOASsN7IkQNF0+/bE9QRi3L6eHwaJdD4DEUXMapcP3V9GP
`protect END_PROTECTED
