`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1n18uE7iRZ7cfHuWPp/tYy7wDW1pCpo854d5VTCyWKAm3rj9Ibmke6I7JanHX9u5
+6SfbPGSjbtri9ltuhbnQMmsfdhpRgQwq2JMgg3PROnh9JlE5cZz72r1Yy3Y+878
WpkqG/FW438cdqCio7faaNavSA8DdgmtcR/ql/Iey5ViR5icJOAi9RX91bc7rFhi
ofvvPiSsg1N3+tpaK6vB//M1e+YYWY6H/PE48PgRCDDUkvmoygqxzEIoLuUL3+Mt
GuOuRzkueReh5CKy5CBYM1Tkx1iV8JqbjimBiuEWcqViJCivsylYxi2u1vEjC31x
LbZRbIR1zUxOhnxifIqFmIlQ8iDBKCRsl5WB7rJi+IUPBwjJGuF/zcEeUT63fmsI
tbrUtlyeqNLHpryB6okgs1ytTW40NNduXmCJauAicgU7AHifl/uLxvrl5XxNaUkv
af9T314n8MmT0LfF4/rm0eFdnkYOrQWeVeOrT7rUaByYBZyYa897LwBeSFIaZYSS
88RHt1iafBMx+LVdYy1WuE576/aatQkrUkNLXWf4TVtnW1Tg1EtpLlLzJIYEUpOq
cEdv54jtGy81PBxjGVPb943huOQalcyPbA9lnr9upw/vICIsC2jcmMdTN2NynqF5
/jqPYoxyb7RxBLvnkqVLrsn5hoxtJutIcfLCs/CRgysJFoDR7qBzFBBylLoZW89i
SzdntEus64uxHXxOfBHyG1HO9O6VYm1dYG9r9UDYwIB1NiCN1RUDcZ1Y0Rq1V0XG
7PDH2LOTaZLjjuhrZp8MrA5mPq5f1aSMYtsldQqYE+1/hRBnHHByeG/Dan5xd/en
vpw/wbBWugDRCVv9IVNr46oaOp2aDU2HvG+/rRs907USU1AuTSeeonmIJuM0aMSG
loxE32xaW4c3GkT8iBpy0TZIZmjw77Z30ND3CJWsq1R9fsTo3dyw/U+4d2m+jd+5
`protect END_PROTECTED
