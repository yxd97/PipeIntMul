`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KV3TH5gA1hkogN58Ap4f8kkrd6yIFOzkapVgyFnAom0ADBZkpFCTSlqy2rBVrir7
ka0lCNGoimSa8Myc2HsKuHtDR9RywwqxR8eC6U1uxFFxdakMFnhryL/WcWD+3lJs
ugz4OuTPn/spfTyBoLOVl91g0NLH7o3awrWQAYks2vjo1lDqeaUGPB1bxebmOAI7
9pOWwaJb3qwFkbK8EBzYD/UTPLq3jgepsGRNDqoyhAQjbxPptTsPsxewXPUe1ob4
Dluz0mInfoCoysudQ5Ucg4pon6N5VHSr+jmTCzblPphC9H34r83tsik0EX+7frnd
CKIz13L8zNhc0oLoV60y12RZiECBwD2LFfPMXfbWe10=
`protect END_PROTECTED
