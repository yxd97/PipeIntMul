`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgmDrNzchU8ftifXhgPWHHfzXBpVGuoRNrGm/cS8dBIFO5n4wDtyvkPf6QxcqufE
oGZAmCcMdYAGT400GoUfurRf9L9teo50CViLYJzcpOZEKmlDs+47x0Btvt3tjoPV
uEX2mMB3KBhvZW/BXU3Ig3ws5Q+oEI7no8rB7kkkmUEINRb3wYMFjKxU5sfVurJb
pGcUx0oSp+jvKT1TZbZdmk65QGx+JkkEQbqpNIEfbg9alGwoaDdw5z5VjepGLXdw
XvZLNxbbz25kLcxaTpwCQIxBSbbyOIiRsmzm8PUmqcaTciDBwmCtLTjuJPIMA8ae
l5FVGkFULhscU7fLEGxT9JW+4ORxXl47p/PE/EayQWubiVRnHw8w/Sh3Hdq4E4Ny
SXtw23nA+nSjgWbH6aDaYay0QXyYxi2iV5mWmyPRZEQh5u/2nlr7dzVGBxS2c5tP
IYlHZ8ONljJmgkXQZ57KZMcXx0sP4yQ72G8auheI59E2CZE3pIFJhC7DSmIG3tbX
axZx+T26PAMs3VXMfT0bAG4aOaQWWB3SyVE5EKf7b1VDOPh63mkl0d07oNiCRFSn
CWR9JoMl+kWbQpSfb5ezMBKIIaK0ysujs9p8WJQfaL/mbHekueexlsIngYBnO+xN
ykhHe9X3kNqh+dLI+Jpo6w==
`protect END_PROTECTED
