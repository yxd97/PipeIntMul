`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33g0XcCXgcFB6A+o0LonLZFl39lWXFtNoiL9OPxZM4y5A6tvu4HvzD4lhkw6M41W
ZikKImaNtiTcU5VacWKPTGIOyOmPGLnPXGRvbjQl/c1JAGdB+wkdnhkE3N6Bjzqd
7fXQJCOouNGkXi5YUqBY9DtGPzbtpsOE5cdk1ET4XHP/VaE9JdIPKU2i632iFno0
e010p8x1aRwhC5XjM8rahD5eLJyRtwAvP8gDWLEsDXUeKy4PFFQzbOfCp7mlf5Bl
jy5yCHQPRWecB856B1CQaHdRxgcXViohtXeLnoisgFSQKYVvxlJnFOHqDhzEVfhp
i++f+9tQsJAcoomNNMCuVVenGKXb1cu0XVHbXqCROkoLt7stlHQdEtmb/zpwvbKJ
RDw34fcaqCzDxIN2MYR/CDSRCEHtPN7B90O+yo1X+NpIQWT6Q9vrbbsZeSan3Y2s
ynwZ7ymUenLuYXPO6Vny4batGDZ0RwSrhQDrjFyMT+E=
`protect END_PROTECTED
