`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Q8K4XfCRXwdnjR7E0bP46seWDOQokHPMowavOk6chkS097vt00iJLjKnjLY8o16
ceR9yOEzNES1cMyOWvXY7R9FGN5g1NDOPkDmYXXDvLjvcxPnbmvD/yM+8gJG1dlh
n4JxOW8NDLR8GmeJr8PrkerZ5nbb1QANtV5/NUzW8Fm9hHIMVP3BuJn4yDMkhNfE
oU7Q8WSnyDS29gxV8JVnfnbU+fzlsxDNEFuynJk+2FrTczfUdO16KH0Ke7zhNaCw
pT0M+0cIfX96naqKCBMDbQ5D+eVeHAcF7yNXf6/1yPUb1aeXh6rvfKX2s2N2hA73
XJ3F1BHhylqigkLTw1YQhg==
`protect END_PROTECTED
