`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFT/CoIPKWdeYZa4oPLv7YCyPCQcER9m+RFDvnFuIemt5/L/Ly0I5tc9IjzWcFP8
D7IoXzRya0begKy5O8Rz7/4StL2ib0Aanpa0/JlcR35tj+YSsoGHOb6XtkUE4dPJ
KLqALATBlJ1KAiv9teawmzJIJ5t6He8ovcZeZ8zPmiJJVc81nacgEU7M63E66159
ADfgOiYI2cZG4s3GjXu2SfX6ILu6JTtIMmmx38uReGhqq+sp3iEfEj4yVz+OKSsl
Hs4mP/PiiP5uE5bSRfFkmjVUA8q7P2ZSs+HCWBqjpYou7fZuR8OhW760r4+ee9IV
XFvCeOJzJIsTBNGEGxjyGOgi8v1ECAESufKz5ucm1tmlr7+xqgBNCH9ZWN6BWJFq
rwpFyzK1OwvEjReNZ3iDe6MbjYTeNSedNQt6yrEi1ccjDnOOgkkXv3MuYEuR66Fj
24hh08ER/GCUWCtM49ZaKsPQTTrN9xMVfnKlqHmpMXX47XA6zhbdoFJGIohEGCU8
v8/3GB7DIZNjmZbIjV9Nmowecx8IjPTjAvOt70mgbMpSLtY/gBrs8TmxK5HiGFuu
fnW5j9wXvf/lAJP+f3gbnMH5NceuiA0OuaIB363DojS5F9NdSBUuLuAOPIq6NL9H
c1XA91j3aKpnQSRLB4SJoe5Jgxxk0iPrsWPZK5+epTlL1AAOR/11iHndTZFl7+IX
2suNsXOcqEXkGUzjiYZ/ok8Uvqz7/5BJV5wB0J7Tl3VM9ppovU0PaQ+d3Hk+dmOX
/9RY0iY5Kqa/doqfYqDV2pJERzBYOeAftxRADXSG0UysicleuE0TGn22/jRKitzC
S8OzP96waxcWjN7OnHlJzRjXlJwwT4f17OCjEzuJ202yX9pCcqvJPjXAjDPERTZa
hsB1ZEIFRCsovnVVWDKBVBoJMtv86PWvMIywFoIhEDbf3v5b+Wgv7bDcVtvTF7dL
VmO4gb5aPY60eWwfR2MX/RKS9A0PC/MGtihwAlWjk6/CtXeQKJNEi4ykrUTDbtmz
PEEY0OSDzr70OLqDHs8feSsszDM5l2iMJsBGxsF3AvzAGsyVTdoAlMUL91BHnsqh
P/wNUY/HW+SVGslSt0TauJ3rP1dqaR35wl0qKOqei09cB2EMZgNbWGHh2pt27Tqi
oIcHSoA797nCSO5CUQUcV9Y3zzi3bg8R4mFOh2GyC2mQJdvVo1xsmjSkqLIcEJQN
`protect END_PROTECTED
