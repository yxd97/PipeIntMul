`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p583FnH83IJ1Dw1piOYplCYWhfiRS9Wi5YZOs4SAVDaNWASW9CPtGjfZj5SfS5YC
aEjzDFyrm7aHBW8o5qlmpkeOy0guuOpseDj4wqOc9fnDOiFO2RDd23S01yReWN41
A1S+pbj/XerwN+bRVrwWbO+5Oyz+b47SCQTsyPYVhexH6bRAH7pbfmAesAEjzW2R
9KA5cspxXprzE8I5S7A6lR8W9AvwmMZ3SEjahDwmkBY2+8ovppk5CMo+2qE8XEvS
77rDiar3qa0O98an29MNC4va4rQhDFqyNJEt2ZZoh/4Bk7EeoMgPMXkWOwfYscEt
4est/WoPjPL71LJNV7bYfBU4tHMVTNd3fuu6iCBM9inudmw8ZvgvfmxhOcvwM5CA
zyQdQYENqjb9z+mvYBdaB7V1BpsP/9s5NkiV8pbgF1G8jyPPfa733l9LIUETVHDu
usYR/uD1nVf2oInZw0Ni6gp53pi20Xjxv/ba8RSNfjS39JiaSeJI4Th99oJIY4nW
I4GAdGj36P4TlgUR45f5EyquA6FhUAY1+56UVLnFcFua9QCiX3Rlam7Ihk3K18hM
CT+Fhn4W1GxyPlWMjK6Fbj5GKB4nDIWSAn6kZ7rbcC0LO8irmHcTbAd+3h07UUsM
9cr/ODiEGghY2QlDFb/VIajomn9UExEmSJg5veQcG5mHvyk7cguWVIkRhNJEaCua
McHgsp9BhH6p4dVsHqYwQu1M/ddto+wFOjl2HpBT0VNvhL0nCV4TTHrHmMIaNbn0
hfFEiofIidnTWIOEKJROdmL0RZqPLddI8UUSWeGb/UeXp985jyPyYlrpZ8TaT8TS
pltanJu3Ixr+MmIAdBnHdSGYmNSCiY6QMerm3qTZdwkga+XLZEwnRVmpqx1gwGDw
5WCX9rjPLqtvu5y1SAPqfwcSMeWyjUAnmnbSqAE5jw7w51R39rR31ozgYzSNNVKE
+xKF1gnz/G6SxOGGvDzjK9aaqm6Yrr4R/Lpk+FGJXWEk27f3LmF+y7G+qHJNeXHd
998+CK7JOcIyooKRDwE3Q5PFb9ry7hT8pYWA0MpeH8TVjUFhhBG3bAum0aXn2ul3
MUcf0Tf2TWvjBfmeXLjR/UGRnGw/Ihp/DE6jFl6PGZSU7tZqnZaq5InkyVAoc9C6
k6mBr7yRiWoxn658s1D9hZELeNbpRgPTee7vumWrAjnvdH/+rTb2v1YFmZSEMupb
A2o5MWK9He9ToCUnBAw+QBXaxb7n1Ofl95BlYu7cq5UGWCZiZ5VXxYLH6AAfzRyg
f00cIUy1g8oMpTFZZ2haYeDp7obuJiafGUOZcacpMArilceFAaWuDOxg4+hoidyf
QqEQkW60UtCX7ZsESokXpfd3rZ65L3PwNat+b+wCG+1RWy052/UL/1DdOXh5qmhG
Nyura+xwrsOVRP2pi3DKB4PPtIw6Dl9PxhC0gxQMpPbuejD/teM6GXzJwcnEKjPy
Mfw6ueRfr0uyg4DSoVfIYZvnh7qHuhwRB6oOozKOJHnv+7kUvLxx9EA+lGzAmrpp
jrjsFshxmK1kAsqKTgljtjrnCgA+rK0dgVjqm8SjUcHLJJTAE6TUsxPsokTlpARu
R6QFXYoaFB6U4gZF/pX6oDK2HWpBYYpIrK0r+Gq8N+Gw1chH3yII/rJ4vgxp/KVE
y6nf+EfCSOxX8g5cc2HaFTFfuSkPc+X4L767gR60JHH3O+y6SaMcJ6XlrGdWB/t+
hZLK8SD6r75xoTPN+PW9+1U6lxGCnnwo86iU9gQsV0JOWBm8+3as6Y9kr50jZT1o
c9o7BmFQOj5Ur1lzBw/RNsE0ghHw5+MjxvHoPVh/09hOj/KuhD8NmCVCD8T64LJK
hfGE/7xQtNwGyQHa7e2o+GvV6TmJ5mbauM9oIc0yD3wMBg6NCl7fI5yaUm/lvzTM
6WOo4QBb2kmzuGWkw49Fsx+/zJn8lDlXleX4CbA5RXDEgzXqxEvRzUdkllPZPUdV
B2yFB1AXvExRK101IAsSBv+XNxo/dqD4hnkVAP+UV7qU3A9nUrNisanVCjfOH/k4
m0nKK+ltlABiZorCAElI+06hjxoGhtk0HWI6WwlUoAKvYJCtc3IM5Mr4lY53Zx/z
U+E7m60y3QwzU7RM0Ea5Dpgp+xPyT7arihkSO6cejzkuz4qPQvZpu7eP7dvmz+Lf
aF1HNo00Ewn9vL3WDuDsQ7rPOelAgaJnDmUhJdW1jNoyKHx79nQJb2HQ/58Sr5wN
nyyPnzEUr4g7IAuA8mH3aZEvRDwyKbJTG/sMK5Lta/RS4oKqPMj2R4o915Zs+1A8
Euli2zC2GFw1LxKamwQGCw6DTsUsSNFKJXoF7XgY/tt/seRl5gwglgF8pmJDArti
iOUheFa+Ly2iljvpKBcQ3PP4LD7yNXILL++tuNYgY3O6yl/3RSjeOdpqOhOphIJP
4miWEBCXEAFptCzphov9kWv7C5sUdkzJkz9YC11Tj5huYseOfVdGKicHS0IaG9iC
T1aow85qBlgb4EODptmqcPNSrckC0kp5705lsp6axVuVWfLse2zAS4aXTEuXORGw
jYPmLvN08l0eKbVTalSNgpm1Jq49e8TOASy5wo4t8WI6h0MSUOr/USaOPNChA78l
zAtCfELJpB/V4GtVLkrqv0Hj/t1BpPKc5hBZPukTpX68L0wunCiSYTSfgVdSGtMw
uuOIXFrC6MypCj3oebKcLjvaMSGDomwDCuRQU4v0wumSdkn5sbkVYvY/Q/ZAtwxs
hNCnB5lNXbF4qogd0FXl1zxIk+aN3AmnkS/ZURe5onvfDscjMETkLahtZWY4ORxj
PmGjWukrDeWmbAQ7skMJqBsA0uO6lIEQgs0Jf4vUqyV/EhUUZ8gkqZvgn1V+lAr/
wG/cYWm5pxJh/RlAgS+VQuATi33FrEFPiGTKjSI74xSrZl6j6LBo8zWcH0piiw+3
SyGBnbWXk1AT4u3vQwjiE9uptXR8qfH58PReKTa38oudC76ZsYgbm9bMOuEI7jgW
PtfZfKsVoewz+HDOAh0+HpWZ23+1NrABFQIDma4uYWv6MjCmoiIuQKI8GEfPBX5X
moEll5eU3jb+7Tq0jE7Ggj26dS4ZAfmb3mYMR0P0OCbvfx7LNPToZr30X3qG9IDZ
GF2EslMO2+9T8dcIq653Yf4x7LzKg4WMXxaqdYm1L3IP9kKBfN2rNHj+xOo98GNJ
qwTr8X9oUy0lIWrK2PZO/w64ZIaJkPvPvJ/IiwpUrZxoMz3uD7Z6Wo14iV5ke7+J
4WndNjNqsD8DTqgVNyEsJv9mZpczn5dU5oqODssimnGvVIo22jYLBHKb2pWHAtxr
jPzXmSeXBPHdZfkMACYsVOL5IBvfpNvqWAoXvkfYLnRJzVzZTY13LL+sRd8MWnjN
byy8aDZW5uGtPZ4UyLwMpjre1LUHaC7OK/0PlVled7u98PhZuSDxc8c9WX+Y91Li
orMFhpnaHzeTStAUv7g6y2ExwYI3ON82zmCELJuTWWMaXEmnEghtjQ05G6b9vVha
InePxp9oaUX41C1V4OaA4IIDCpa9h362GwV+a3LMQM9J6NlPtGpesjk8Bn67pIug
keiLU66RMd2mxtkwhuUfXldA8PZACjsCU8aYu2D5phCLYuHfiiIpXhW/RhuOs0Ep
LBrmdc32HAlCx4IJHuB2WXTTsG9EZKzNYbf92B4mw3nvbt+x/Ax+iaBdLDxTdXpV
mqNjOvZcRUVte2EGCv1WrYeL6TtrVXGM8Dir+PQDDMDjkCabynEHL4o5gB6/+k3k
`protect END_PROTECTED
