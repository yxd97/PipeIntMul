`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZfDxzFcWkw2npJdnfGB/o2YTVp/cNxPBOuUnHaftCOBnL60Y4WH4kXYtjWtEFAj
AJOZ3egtVASRgg82cvisQWVjTJ3PtiEZcY8eZOwUd4hsCYZ2Ja/5UeQTKsRNS0gP
87uwwC111k/WRdeEq8/+ofr/gbyIUknn3FlGap+O/JMs3rmaSRs3i+uJjlIOOmfy
rv4JQpYrubBiPLAPf0DOVRT+cAgw9o0MfQLkpLSCXDE/DXcgjXyo35hZYGvfal8K
cKu/wLa8lqdwItTDrxIBBz13Idw6ZVrM4I4kV7Rl+r1DzkKCZviqxhm2eRcXLEMx
6Eg2rZ6LMfHzu+7v8RkGqw==
`protect END_PROTECTED
