`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/TIvwSZrvnhvA5ewnakiS2bNrxKDrH5X83cBTdDpraGi9qkO/+TT9osVHExFVmNe
H03CtSd0Mr10RZaBrndEsLjZ96BKY9+hoYG0k3o5//R/mIZbZq0VfiYVTQ9zgSnM
GWWPBfgpjs24Lo9NSZxvsleC1BsnwtMozhNZ8yPWBVyRX9yJ1ByEu8ifKrv/pIBC
Oele+URPJuKE0caqQ4t5xahnVgeJXi2oMAis1AP+WxKoFms97vjZrZ00s/ZA0O0U
lrikRVdxGHoSKo9oT7vGdwget4X8fQ1gUkATqVrtZF+umBkCOVMI0ewNn0s0Hj85
y3ky2TCDfF3Wih5TrVaqxLcchDgp4+7TmEkwgJYvhADbCqb3KSZi1NDxZcX9a7Dt
tuuOh6kyVGcGLULXPtWoHnm3DgqAukx3kn7ZibIEX4rbUP0xpK8JfRFKyBGgZoP7
aM+cQivcseKgpvrByE4cnohPfhOf+yPXq+ScRjFtBaUCXNLxLLhl75rLktN51lL/
`protect END_PROTECTED
