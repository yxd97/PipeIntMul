`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7RlE2oEhaEw8KiqBUTcAiSIhWD6z2CIvlkm1Wfzvbnps1XY63mZEbqv8Cpp/MWG
QWLak0bNCO/aQGsngTpMQ/yOdO0oAM2X3YCjPY2snA1SFYJSnrtGY4EMnV/BFHWo
e02NCkl3co1/UDlZAnOzZp3G0qsysXjqWj2g+b1eeMTojqqU2ISCAawPNhnuGxgZ
1sR7+xQrjrZ4dRYmKGpwt7R5ofGlxqHvzpQFv2h9J61rkxNeEEwYIA5JhucRftle
qOr33dDWg7qzDA4oMeFmIrhUeHzqygiXuK/UCT/Drlgfugj1ZDPBNs22X1qRM3O+
M96BVoFXOTHjAqpEd+NaNPNTHXtSK71QDFqUqwwYSolF5YWs3tyD40+bH7jORstX
A4s6+euGKz2wT65f6zAwppzPoT8e7lpqLfrvjE4BUfaowNA0jED783077pLEE1qy
UkWV8Lpgb4/wZEFbIDOAtyKdiZntONlW69VPQ9WBOi4=
`protect END_PROTECTED
