`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+wt+J13+Htb/f80WzMXHwLki+fxluAlnd4YzWOzb/2M/0pwAVNQipuQRzjX7xmSZ
sYc8DaFVlZp/oxlSS/wox+gEjljzEPxhNyFArE1JXpRe9wvsaqknNtsLMI9GXPnh
TkGKBdLwkmyFKYUiqdxTdCZVkdUzdAxj3eFg5W2qNKGPhImZSW8/D8USnZMwZTZK
1Doji+ulWDEDmvE+Ei9+1oBDEka+VaohefrlIOU8iSNT+E/SnrYU79ema3V9I8Xu
WRwFVD7vIiOTIv4DvQQc5v3fUf4i06G7uqt9zpHNS9ZJmX2r0xnW4RNouhaNxEYb
`protect END_PROTECTED
