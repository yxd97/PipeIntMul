`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EfNwkSiikwf0wgpRGz1HdnnZOz+h1vKYZXEys2Qfb9+ct6bYCUFURnk8uZFC0EEn
f5j5efsGCdqpjU7aUkWBbiR+noR6sQQB9eym7YC2JonEspqo7cLBhcBonlKb0H8/
pRXli+l1FB425DZ2wUxCP8ABCFm7WEwKjAbvvF9y2ryc2TwCOxtQa05BzTsCjMcw
TYC5ijC0WefYml7WdHCckEemXkIuvuiFX5DEuzXR589Sq8r7I66cqLGG5+vy9eOY
YaT7HwyAjyu058bizQU6Ur3cEWw/4fF4DKRFmMtK6FjKggq6b62m6AgW3w2vt3EA
THCqGH1UJPHmt6Qm0rJPo9sEuUjfSP+AzivrkWoUzHw3BCPcDLO7ZEvrEY0oNgmA
/+eoHCeOsGzO/FjTW1VMeRWNr/poZAaVhFxnTfV4dSM=
`protect END_PROTECTED
