`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISehCEWnb8a4tJCpteDusPiaLGvFJCWlnnXZmu3rAEZX24WPj3myW/92CybXHnP1
6WLMdahuxr41UrmIQVnLTLavSRv2SF+IOqlQcqz4KnWAgirsrl+OcC1CVXseHeaz
21uB50+mJ2GPvP5oCSceJKCxYSEBpUKgEaCZiyWsX8hSjC+eFnI1fdQ9lUZ+s7Nc
CykOqFpZ160QdES3EoA8umOiwlnG7hdwe2LVjPyWQ0iYkNQJPQad03ARj1hEjn7B
CpcCBFU9/6VjbtyXLoB6/OSWhNOBTB543IjmRnx1I2piXiUAq0uScAE/SNidKh31
F/j+DtkwDzU2TP/qg6RuaG2uHC0G6oo2ekmcWqAaBfoPOEqXPzkSxw+4TQso7uf9
3KeC3kpLMgaH70qbuDv3km1Gm+HXcvWW9XzkT6uGo1HCNgRArY203aFfdDBK3TrD
uhZiXbOZpJeTLPUIAY9/WWsTDlYQxwaKk7eLCOPARD7g7AZYClsxcFtIEnT40hQE
f0alLKU5gdxsRs0SpiXFcElO/+Sijov+qdF3xnLoRMBL3NQG9oBlXJNetlLmqkg0
yjCEgYwurQb1FUC5nIJ8Fbr6fXVpfN4Cei6GUxKy5oGzjtqy0wfDnvLtXk2r/Rpi
/T9f+EyvKt8BntNRpLcbmuTdpP+kM2nEJVXcvFhYGRBhr4T9pyERAgYOqCiGeEYr
2Kvgin+j+DAqis5K8hsmahE9Nk0+U7VOzxTAajZjLovLhEEz3oJa+GeYxuEn77Jz
sDIfa3Ve6pgidH+m6aVgQl0Udzvuc6CvZEF5PiobnS/HJNzaPzOkjngHv2KBU4Q7
bYSHTBDfhWhnaQoPIE5Sopks6vQZNHIVGlxvbpyC/SYttTiUCrgcP8dynSI7kXHP
TpZ0Gfm+PUzJ4ltz+vstK8u6J/oqMXrELkJC6dL+q1PUoms5E0Uhuh+w1F0Crgxa
fyzfoAs+C5X6azY3ho95gdduumd5Jy1+F/13Ns9RLEXIrktwl92m3kp4d7lEbaFR
QzR6cifmufBVOAI3qQl/NtH0RK38srccN0lLLO/dxebLY39IOiIB9H+OCOaT3Pgc
olH4ZVJ23LK83/fIp34e7u3aAeN2r1Tax9Cgy/kbs58mZefnkoycPP4ybGTaKb4u
tPE4imwdSAVeYWQwMLJ6nGpb0fYIdybdY44SruB+YH5zCfTNd8YZwVOj0s5WH4oJ
TSMaqON+9VTFYjM9rIKXB/PTlxXKrMopndKY5bzHasJ2c0tYST8PIunbxnWrEbXR
ovilzaqBMeHVTCmS24Jam1bMOCwtM8DXbbKULtLuvJbZ4dcTK6lcmfYSNyndkUl0
5URScwzwXO0DgaUl6OO5gZjS2ykC+7Bnw4IUT3T58yW5SuYFklMP8LZpBbKz8V7T
Lvdrk6oiWtc8bRJYm1zSbwRQQhUsehTrqyj2rr7H9U+Pysr5YLe+Xlum2UZhkMWL
FZk0xzZjbcTI0FlVoq4Wx1St0pX2VBkDwAeULXNOPTt8dZTrR7a/eujyywindO0N
D5cvHSqW0Dwi7XEDE4ip4A9tmZk4n9C01N6yuGD/2KMZv4PpSrbEQrgMz67/s06r
SzAtqmmv0bpD9ypzzjeosBYpJuXzxiGKazuZPiLeGL/pvPw19+huTjGYPGILydD8
HoVaBesZlKFgrhm4jW59ezdAoqbb3fH3k8Osx+m0a8eii8N8mwyRuBWjTs1MUh8c
y8LB4s3NV0tEP917z5NyrwD4J66OQ4tNcMa1oF+lpMWpXZQpEdxEUN2umD8QQBbx
4ZViLmdgT+ov1HO/tabXtJm2+TVAjYPf94dAL6ySvOwKXguD37U7nuggcdHNY/1A
fY5ymjs8xVwwUzBmtXZshYBuG9uV3UKWzkvZn6piTXa3QHfHa/ss8Xbj1uEVmY7c
5Cl4Y/LXDn5NaGGdlD7GyqYayEkpmkHJ5ZZ5LzX486k7wRU95z2XKWvMbfdTd4Qd
lgfb/kjzF1yJYSBqYavGnET/orGk0lEqSZQ9LfJfnUihB/XondANdJI8ZxN5maEO
PtkDOkNllYwik34dgl5AcZpa2L6bHtrmPMn4Lo+acxgEYn8HDvGJxX+/p/aZjw2R
ZfOXV+pb/T9Azet13iJWbcdEwVarT2K1xQoqwG1w5xNRT00zDDdd8qZOBr23oSUG
65jFR4+pOfKENBC2TYS5ftDRCaSl2OfjGelWTQx8oXpPimtIG/hXhrtuIZAon0r2
PVIzutx3blvHdmDITbJlKwGrRB6F1GPZp7jYyRcVAPnQVZy1dz+BOoaO4+mOLeq4
V3KVIxXgqtzA/lQDy2DmKbcLWQAKNWzOZ/AGOlBiBI4cuZtnHm34Y/dILQpbiPHQ
/PV687jyBBBloTLpAyCk6hrpcgSc8npOEs4wb7Ifds7ENkhgLKzpZ8n4uXyG+dCu
K0sj/PGPhx9dpvmulD7aipUyfJIuap+eozky6CZZtI8JqUafZ2rAtv2ZY0LzUs1B
0AdskRwUJ7A8mMv3P8MebYaffXQ0c5IvK68CAL6x25sSfDLpZglY0PwDseuXBkYv
1SrklTehCFkfPmrSzbkdoaukCwsAPwiOzkx9hK6GchR44AxYFTVIYw3IFsQmfeeP
dp12kauQ/06q5iEFcxRsCpEaApfEaoOIQ9fFCngcX1d3JOPSwmf8Vn1WYa0qDftE
qoiaAsM83A9Gk0jCUQB2qn8C48nn07JDMiKSfHdyov1mOsI7u9QZAHKrB8bPVk9r
+zhhP7c3lwkKi6Z+p9EGmjXXv4DeZUYykoBP+0YN3MeaL6JUg7SiMWIpWhykpJNs
T3JmrdwQf4y/HcWaICEiH5awkE38Wn4mHtMvVJ7J3x3IYOE2o/Oz5DuLrjlqaPMg
z2gqyq4gXSEG2wO61gO+zVeXBg62IvaAgSDJZgGesCgQj+RgyUlhTPEWa9Y08V6V
5d68JWzT4YdvihI9YolL1jNol4FlLUzfrzVAm4Bnp4vHmHqxhr3erA6i5oy8U+EM
TeAjSk90gp64qSIH1kMKTk4tSbfa5j+az3vNWrT4O52AYvVwx2EUnZmOIi8JxWy6
5gvmDgr+6+mYBo+ypBbCUkjtE00llPHA14YcdpVliLlNMZt+loHkUciVDV4XfyqJ
Z9eBpd79sVtVD033caM6cMSVg7MXWEJpzvAcfZ6nV1mIdz0ufur2uL/jk8cERP5c
esPcO/Ig1eY65LaY7W9Tx3Quqbvx1t/eMLv0T0R0+lgrfXm/lCLP3QZBRk31qDko
EHneKOz4I50YLb/6vebux4Pizgy2mxAf+ISw2WLSuizl2Xsid1M6wVN8ZnsujZRC
6Yymbgw/c/6GuxsyVDtqCdwqTE+6x3oZW/2z+MRVJfhIqsesP+R+GjIl/T4b5LM6
FG5Ji9686X8ixjbwQ67afvG8lqy5xVwXptiqRiXdbHeEl+rBFwxGlG5ebf+p+NQZ
xs45786PCm9uTWPRV3FiFFU60ljhMxWyh8ZmmFk+HahmyjhD2JfO05ZV7zxeRInd
WvlOn/EvMSMeNWStQp8HFjhDnUcr5rYgObgit++uSGOqoU9bmP6tW1ij4JdHsTUm
Q+2nPCGeKjgGVueXBxbbdgIyuUpS0Or02k9q4U9qEG+qNO5UzH55UsTFa8NzgsIt
HlouvvYEvPCP5s1xoTSVz4rXvzNb85PJEUJ2jC73VA2z7J5/JrZVCOvNTa803uiF
r29m+sh8A49qVLDeOEnx+lJJj9by7GB7eMO+iv77zfqiCZ1Jiy/I1LOpZ1TJZ7f0
yI//usSA2LpH/N8F8Y3Aa7SOW/8Kqipr8bzLgg8iMErzR9bvMtRkVZnpZFW6WF5+
QgWLmI4w8UsJOMN+DrnVZcbCalVOnbOuFwjwgLQRymkXMc2Tfdn1fuyKYsAqEB8V
nX2jSApaN4rmQ7XfD8D6RuTCdHTwGlZjFJbnhAeZDuf5kvn77aqkpnRjkzt+SBGU
/xVPmqsopHKBjfEe0zuv6EeC6hWeGSe3+V96hKYEWScncpW8FzCds5hQSMNkiifj
agsKaGTx3HaJwEZqM5/ZNeCF6GGo+0FrEeaSSOAH14iFXA3sgcN5a3j9q3Ivudxx
IErtfMkcWi8WNBxnfDKs0+5iJrkYxvmZh8khfBIMLlTK5kvOhghhXR60ALefQ/6X
TGYOakKeuBSf3uwxHKFEr02n8RNHSfjkOpr/0qB/rlvz+AKTG/JOrxQWcXhc9+6i
lmcJy9s+ytKbo+yCA6UdzcEtYH6LFbCKj2t4J+RskqRGA8+tyk3B+gMCYBt/QdQQ
cLdP+WS4RL9tGjukiaDLAj/y+99Vxqd00Srkutkg36wqher/plWugDFmBXnztsbz
nY6zDZLSnvxZoAs9S32QBSgA/Q4X8Z/+RX29bt2hNfuoVUMw1IOcwjIsmC9oVcMp
aqwDnMDxiGEFCEe5mTX9vaS5ugsm9EGjgybnTXrmzupziTcU88sxRE2ysUi/j+4/
2qlGHl64tkItFClLwcNGEC5oFKdKHkn+a131ZpBAKzWqMi3VF6Qhmrr3Z0nS39ym
k6yJYe+bfVGcxrkAB1uDUB2iByzTU1U8RdeUe4u8y9hOEl+yhylk3+a2sB0Rrs5o
Ris2XCcENxJSWXJzOyZ5BIS8ukiQlzE7Wmq1z3MN3jueNgBZbNBS+1l2rbBtTjb2
QPExsKvao1e2sKXL9kk8grRhBsO2ZVuvz75PQ700fhSdvoV0P7T1rYib1/AZlPR/
KLcW/xHkjV78d5wHmO+wYo5xF2sD3aIfXh9LMJsjTNgFDk9a1eJWID3m6jIuSBbp
ob8BJm7WrC/zq6mow2iJ69W+lx4sC3kMuR+H9aE8K2NeZCYE0R1tXPRliAPniwH4
zUMvs0t5y8I0ep4Bp4B2hfsqJIWkdQGvsAbnE9XUxQcEEEI3aweZWcR+N6mIi06+
VyYiiLoX6hxsDl303DBnDX6bRbHxz4xa+GnGSaAHK7BEghS7PuWLTpRk87qre9Zx
DDphCSsulv6k4oWz59RLkF3JtY2K+GnZKUmbLsvR1RA9+ku+POXGFbMxF8Sjh2Nt
SuGlTjgqB/XVFwpODwJsSIZ33jDA45YXJyl9W1pzOoaGpMXOk21YcGP2cY/xUuqa
FypjsD4EFMu4YRdaelvqAH8oSGSZCLpISSa4EG/9LRUxyDLHEPRdVTP4eVRnMGde
yEEg7HulH4DevWl37R1wZeGW73SQUHuMhE6wKIVrHhCQf8SRaJafDRFQB+wXd7mb
yB0Fbv6Y9gmClQybnWskTQ+Q9EnJMcs0aM936npoz1wpFVM7wP6p82Ku9BV9VN8H
ylc2eBvR5YaQi0l1K+C2gi/tJpyPUZM0yXfPeyOdJyVfntCCtsxhTZlo0XhwsQKV
HxJOdCukjZW3IQEojvjjsS1v2s3VMdy4RkK7Rr63eKPQjkkRmM+fQiv2NPez6cIM
1pETpYopcT9JNKvXzsiQhc3maPg1t81aug8C0DPU/BsNPUf4SFMpr1t5TqSYoA14
K2T9e9ca/iOjj/h/jMkTkPAg9bkLhP1uOctPXDbG13TqrjYrl2AOqEJKlvWwPRQv
b2/qrrq8n0DyDj4xgi2bo/VfWQlVTHPosVNEApfkFg3l/AcBuL5md8IPSJHHIDmT
/KTGQbKbOOit+MLqutzBKVFzjlhX9HYoA00HaZ7T9Uy8dATu2RaFQupNEh6kgXex
MXlC7Ow51ib5YcIzVxn66qlyh+rKRyibjIs9FTGsq5gHX7wd9cMu9VwF+ZZTJxkW
fPShzf4Y5fEO+OfAJepxTKIBczrMX8tNmOVwqgGPdcWGXqyzc6yTpPhn6NpOWs6S
qw840Rb2zbA5j8RfC8rttyueqEOcPPhNsCMG1up6m1+TnmKA/TyGoXLCZFwEwk6C
jjzy7kx5/QWmZZIsjDXdJg/DtA2BANFSnWqHvfO3T1W8IOuuf2uvwb90FXVUvjtq
2uDdAwiHy4tLZDtQ5F2QEdmr5lLpfmShmG1OPkgcUwbU7X/dka4ZDAge2x7cEBKg
mFeBSh9WFQq7rorRGz7A9Phn8rXknEa1pK0wmFUcjqQtOEv3ISrX+//zzkzd1HCX
LVaEYpnmOr1NeoD+aTI0UzEr2Q+4cFRTY6D2US1KWLPYUG+GZ6dJi1ZotRkLwKpS
8E/rZT66+Fzi2LYmk/lCChh+WuafL+Txy248EB8/4GyMJXECo2BD8pDfykm9Ovwp
bHghUs3vwy1I/ivPu/gobvbyuGbG+0iOqJ1CqLmxZZjdItFisP6/bnXEjq9e7bPi
qFVeV9gCvy7FybClEBe88mOghGNhDS3uAwObGObfT5ruOetOJyIvyAKAm5a+57x7
wapUK1PFisuSq4kRn//5KIAQ/xY9lzNO1OpeqfPK5IAsjH2C//hTg57TrDmVCUll
/0AXg8R6zitBqPALVd17QSx02/cNqe0UKHd0ZWoe9VUDF2zE61rIiNyyOXwbXAGU
BrFd3dzZvirS8Q5A+r9K/ULWn8LfXPTHSadTwVZW+CcJ4TqybTNFJhOGe2QOd1uM
Xd24obrtrukbtlvAF6GFYS8QOVnUtKbGKeFSAcfDXAGKUA1clWaMTPiU+gMV2/fj
iM6mz7bmfSvCoUgNqtJJejrbghn4nWXyJSmeL0V0kNTHE4BohLBHoNTRCh846bx9
4KBWWtS8vd8Ti0N+ph9HSw1Yvns1aAdX8ORkTrOJ48Da9pVfHfRQYZ+VqilxsFGH
LwFS/5/kFX2qb7b+fRKXOhmlueRjGA5pAsZjWAubixfQ3BghpFEkQNuU/yEee50N
s5sIWgaaRStmpPMDTPlss+vxUp9bNXKPhylJa/f625QC8U27eVubHQiD9w68H1LG
hA8tDA3UfOSakesuBRvVoRMWBjzMpFuLLM0JB2i5dtf8CEmsCnL7ZugLkIUCh50m
oMuV4Uy4UPaTUf5RCIAd4Wk+te/qGmedFRLSBv3CZb9pXIDww5WMhVCK1HvvLgkY
51Wfhx4vTCi8mxuUHGGrhD0qp72YDXwsh4pCZyumqXWdMrJeMBpaw8nDaIC0QRSm
AY75FTf0bMnHwnEJ9Yy84d88MblxL+G0blTu1PXuu5TdUoD17GT2DC1eJ4iIiYHz
9zO8wCoaw5oIOIlKBg70NrHbgZqT4QgXzFVOpilBqINt+DS7lkvvMl6gFiaRXeIw
i6PFMd/l8sQwV1Rl1pyGmloNz1acdHJrAbJ7vpMTpZl9pYzcNf3Lkh4FomKTV542
mAGd35TPaKlElFXvqRGMzi9FsUraRb5ar5HhdsogsFaogr1Olql9MDNtoQyc7qTL
XFPyGfoNmuxUHk+Bo9J88SLQ+XDIOHhSrQunh/LJ/P46IeViiSmLj2E5S4PnZnOW
vCIui1CaOW6P7gHclD3amJ+oui30RACZd+acC7Bcv7EETppAOAYuOlOsY7IrwDel
Jm/6wZ+WoE2vq71cVHHagR8Mn7awhzjWwUkrneBz4tIAWUvdl+pKIgsNFRdR2jAo
vyLMcC/I9OS70bnCYasPuuglVHA7sRBOIoff4+n/kGXUXeEXHvQ9M/Q/tBDwjSSa
a29TpwTAvkex5mW9dozqKmNuX8sgksHZnzhimXA4YRu9XqNldmDMqUEQ/b6M2YMH
WfOh2D/p1lc2Plu9z8M26s7GncwzUh5BBmZN3vmpOKHQFDYWCjZX1xSVlA77ZWcm
qgzx4I5Yvh3FQ6pE32kTn2OwcJLj1jgZqf3NgrEvbZ2gON61zi36pjbAQRUtDz3V
APgguDfT4BfiKUKYRv78cuF4mLKVpjk6p2lSO+T1vInhNZ2tlKF9uhRhJGG3Y9Ui
nt4kyS87xTdNc2Al80ldRBnDA7TbxiD/U2iZl4DH5Ex4+E/j5Nhw8G7SVYj66bWx
bMm3Dn7wHQmgYaq9Ofd5hUmn3cFaBNlEcI8lDpz3P5u97SqNqAIK3MhfMsusxnsG
JRBfCq/GktL1Nd0HqNYXtwj154ULDLRBql8YRqRiOut3bpytnFNiFLYmCZNZaS36
mUHyCv+MPKSbqOXEwgh0oq6j91ocPgUG/h1bTBLnRQmgy7t0iGI8j+GBxmwX7u6T
69v2h3xHlbSD4p2YRDM/ATwQMQei0mY84Nd+xP7xzbbg0wLkOz5pPjbUwibh7tVm
FytEyTjq2QYm7t8qQVW8UcyukV4x7vCfLovQNz74sMC3AyaIYDBAfbzijFmV/Uke
VGv0not5tTS+mkh8vYFzb998xi1TNRRLjcQoBwkD2F4/Br3AcLPk+9dcgGWD6bIC
uKwEO+kZf1aSv6KrNVI99bQ/20+aSsTpwNUknCJjpI7R6hHcgxeBdRkohwvRt6g7
sh7r6AI1CRBhbHD1XpvHnxr+OigtmyCrLMcSOPcolNXzvn1QNN7H/9aM3rX1S0/1
i3HVXi0JtDu/Cj/QnrE04FflAsMqKGbDldwIGVGzAd+24kxab6A5dEs5UbHHJwE8
tI0yiPtJHyhsuHsOxZFAyhRrQk97E3Hsl31+JtaEWYK4nHZBo3GMJFBndcEdaVYe
IXqyjegMMSZT651z0BUgWNCKRvhulBN3sb0R0ylZ5m15FFHHQ9RdEb01b4gF3ab2
zos2Fh4AjV2LMUg2R6ZJIFYYzIDKTSQ88DXoXyKuJDqD33vjHSEm3elcUN4pUJzZ
gNlcTy+rXXU6FWWd4xPLUY9VuO+z/PILJPPsgJ4uffWtSkjCezMos/ICdPt6qzf2
PBB0ZuTHtHgn1LvC1NjUXuhwnGz6yKPb6UhnSJsjH4/NJf7B0idEq8tyI3eCw6r2
p6qAi6p6l8VuFmqcnWl3wldVBPu647z4G7TLxIdiyBQkwH9VkEZUNxCj2LjAWJn1
ouqATATzAp3ng/DaB1Lp2M8fcAuxG6zC2lUSLNH60fkW2P2TKwK8wUuP2scDhxFn
viTWhu87dIgGM7EOOVrh6mCtfvNr19ZIDQg3kiMtGFJe2Thx5nZ4662kRbupK8Yr
nyIrevvVRkftYU17wqw6D5wL1ZPNMEU75ZOb3LVzRj2MdJQC7paCN9xPdVu82J4U
xMkBtklKXdkBVttmFG5RViYV98Cn2+PTs9P8G11BcYA4Sgu75tT9iByIiEgXBG55
rxewjLc6Do+1+7BbHLbhkbpOSe+Q3xHKHuKEICRvfOLXiNdPfANpNkvICgSVevAw
b6Vlm2Z+uSSwNZPegU/sLPM7sJt+GE6BFWbrWzM3SiWscns8vxF9F+BU31mSwvD/
QZ4TaOicxKtmEggFgc2MeaMy2Ka5q84HeKjf+IiIP2t0NUb5/iu7M4pkO5rANiYQ
fQ4piI5Mfoo+PATv68AS1x658IRIpA0RHRHZKgtWTo6vYvn1eJ2m1qDktAG6nrQ/
HtuTqwb+baepxkFB1Dvnm9yEqYDdBEYLUh8j9KpUKblDMIIY/rvcCgcpszLvbJOV
8vCZXS0SBgSoTa2YSlS5UVS0PT3MuqlQihhkcn5r+Mvr7huDRG12imVoNF70ZyEM
vK2I7fXnpgjbclaforjvhkqzDT+HHMJxZLXYNgsB99bIHkdySMD7ELFvyYNA/ohQ
Fzok5Q8DEZMDP0EbFhYuc0iRdcmTfkntlman+shxJtSMdootXzlSSHCdklybtPyR
PMfeYsh0pzFCv41Y6/56VMpgHvK0gCgw8wt06HnNxPvSQxRpMfrytrrftHgXF50Y
Xse0b65EJjq/p+PIwPGQSvdxjEWTHIFP0KGgmzcX1sVxAwtRNKLo+xh4abw76nl6
j7nRFb2ICJMA7zAEh8KhTr4i3/Jpxo+nOicJuAeVpZ3V2qrDGfJtT/qOTXjf4zGH
F8jiQHqSwu/p8rF1yfX40X7piyX/rp6D/k/m/aukZs174odJhJSN/Dz19pi94vim
v7sDF1j62NsH2sm3VuYvMOsfzA3g6J/ZRyQwXRVie5ZaVWpOIQfIz2elpvJrCsfu
Kv3MrUErOaLwUvvuJ3k6Hi1NEf1gicO9v7HLk3UkzlOJl9Ht9B21y47DEFkDJ9Gp
z5ZviDrDWIKhuqpWKnD1B6FKuw5nhCi9Wt1P5dvoEMYN+hcm08Y80bFhrKw0upKJ
AGxGSOgD2XLphhGmzaislC3StbGDYOAD+fwfUu8ec9My5mPw9ZikoNddWd51MQ4g
37CfCYvhx9awD4ZF0YMuJfnVscvNFGr30ZMaaiyAFXfWbvxaskz+ygxiPPDGTfY5
FwVTsMDh87B1hdFGNR0e/baAlo07NTvtiT98DDn29c0U2ctJA0HjMAMeV8A9FOn9
Q6zYp+xvpSoSssIWnC0msKUnaC8SJo4iA83KVNZs8qeqheMAdnFibbFBq2YhmNzr
wUjT/hC3KJvIRi9dyT5uAOBwdrv5oH/QWYVvxCTSrSXMqTpIE6SUDMv59SVC3rbS
LuDMgJUpkWI+MenG/SUj5QgO3poS3LBI2fXny6O4JoZ/DZ9gq7Gy1tx++5CkEqVR
EOSkdPSJclapVTyu1P5vhwt16Ib0fVON4SzO4fsyHM7AY0hPdJ1+A6GAJJVtj+8A
0/THWCCkUuepJooTIldwIrA0D3KIHdHc4QAByJ8t9jCh17EJozY2HX5a0mddFziW
fb5N73KzC0fzg7htNt/HRmNXrP26Y7PYUIrITE3YimTSRv9F4mV8vMtqccg+eSVj
KZEwGu76D1MSbAkWuESVlki7MEiJQideqgl5aoAoFssDFutiQx0RPPHt5MQZgJzS
X1swKdk/dhjBN/laB35QQPNfhztGewNbgvqnZjySYVtIE7hvplbsvONOYLIai9xq
BMmp1VNG8liUy8OLiV0XqvAIuQ60LpbtSNEaqB2ha/Y9zRFuLE3TyqeGXhPT+7rs
ae1xaIBUEqEgXqiXx7hMCe04Hv0zhs14Vlo4BlrB5H4/6qCizKjcFuuNNZH3+j4a
sFvB0kFqlMuLdno0/b1pEib2GxEj3E63X5UccemomS7odUC0Z6VFgXrXQGsc6OwV
zK4X54ijNpLMSC+QCDyJEKJOPFPHDPiLEI2IrWYqCiY31oRZxvYoHWHDyuNFBOu4
V5xxLXCz2SZBSy6dLknfH+t6GJFB4B6oXBEXpxm0g78xj1VmMEqhdrU+LjZpHBoH
5NelMhniHTICNlNFBXODuT2PK4SMG93zuj8HXtjdmYa3rsaq2o0Zlw2SfdIKKmnW
eN2TYwNlbwf2G1coHw/DeybrO+QeSFw+FkpWpTBtUvEjY8+1PrnJ63a5k3YKABgA
SnqCFvKQXmNdTVNTxFe7/T+EwcGx+6bEdgFGeD2Sw/+Wd3Y7x0WSrueS138sStN2
6OUl/yaTVLPMhYpNFUlb/3GqUwaaylhj24UkNS+cq4QXCaQLPu1aKfQkIudYFcZr
ZOqVjTTEbxaHVn6mvJwkvPTwXaUsRwx7BvPxhZtZ96q5+tjnNSmuUoui7XFdR/qs
2U1KrZYcsIk0FS1Tuq9jbZofSONBvWlCk2npExquIK0pMcIzuYItBYwyswRDCuNL
4n5YondwpQNjcntLB2npBr5RC0p5RarABt0IgTh2mXQQM7KskTWkq4ukX6tgn7QU
x+fhHRUsYysg4wLE7cQFqU3n+UG1iDiFNf1JCmOTZ95H0ztXfR1M0PGflUtGnQfF
wbqDM/aR5HeOsfnOQuTgqDhneitmELnw2R8988gg1ijQeQPmBX/uRW+dc3saDbSY
ggjdtJ8nT3t5vwu/IvFGEXErjBxgtwTiHwywCRIBSTyuk6UiEGYZ50gU9EE41AuH
vc6ExOZUrJOyWEoYhrK1QWHGCweiyaIcQXgMoi1azJQa7sazf3HI3IjkmFq64IaS
EmP4OQ1sY/lxBv925LyWj0I0AfhP7KFz1F3qdJtP2esC5ezQPqA74OZhTdGbeTmK
ih3lXRwGqovooLz/3uXrlJHkqShIlHvppf3ZkJ3ImqrJvtlcIdouu0hSRQ5NeoW6
095gqTBr41cuCTSa0DYJu4pBM/LMfMzIW7RIKUtRV5EEqD/NicZeYhEe5uwunNaZ
hI9NcDwyoqywLunmlqYeCDjZtP7Wo2QjEsJAhN9C9QUYva2NPsVK2wKEtFqkRMQg
RWNqXSkGVTcwirjatF4CMleo0BYYfJ0RiARlQTv7JW1IuC21QdEmupQEdFPxyjyL
ZC/FZCZaZ4/t56sZu6hSfAMmQKBVDtzPcsEL36R4fwrkcCr6BXzhmFre6BMnnJ3J
TrtMYkcPuUAtq5pJ5JGlQDGVVLbfCvzRjhPO9fOe940uqIePWm5XIWM+fgtukbV9
lLTEPQsRrEpmVnaf39KVOYROT06EvYzcKiyC0n+rmFO12qj0hecwSiWkbx3yeJrQ
ywwvHPHJv5sg477IXjJlvyYmwWovwoLjoU1POj4AB3I6wsxMSxApc21wG3mgMOfx
6wgOtuh/zG46GkW2PNID/0Xcrz+nAeHhSID3D7GVh3VFGBa5FF79BPRRXbvy01oN
Pr5f7qy4MtDayaEfE+/vggoPz+bBF6/HDEwv/Vnq07h3mMsJ+XW/6UwVuEv9N5yu
ShEYiIGypPfqux7OjAiJB6XvWuUj4qQ+Qyqz5GSjBDntHoaJ2rqtUW8Y9EVjpAsf
oh5+fumROPZf4CMtNdJhUTFKblC4q32MZPTUiMd7ToUx3lkxIVeRZ1PUrlselD+C
aAJot8wD8JIdxqgZQVdauhbt8TMi5Ihu2jJnBTrNerQjKk9Atpj6jARB2F7J9sKD
6QaLO0sWettBLe1J/fNHoqJP9sEotpVS1MkHjCTE+gnev7Z3eQ5X98XDz8rejsTK
4UPaeldVlc9hdiM4yqt1ljhFIo1J9nLc6pAWP3Sq591k51rKFbfhhWbp3QIYC9vb
T9mEZHLASgNuDpZEyeX9opsldb31aB9gB619GSCj4p27QjvyDetlvspkXw4cnHLn
Fr8Zx8KjVQwencUk8Gfq9N5MQFR390e2jSmK5gA2SqXPkCDq2toj5C6REz2UG9MA
BsRNkROHHdEvQS9cQ5ElSnpypSJIsje4ox9R6u5hLKbIc87E7Lsaw7QiDoCaYGDH
vwUvjyW4xX77J7545AT2KFcuJfJLdZLyAWYxRH26+AMD5BmDaYqFQXEAKnFMlO+p
hEeqbpHKqEYJIa8eKlFxcK2rJ3R2OrFT0XsddRZThcuFvlNhg+wNg3dGum/l31b4
HqHtmukX2X2ezhHwmVEbH+UV8rQkO3Hi50rV6pVowp9yZ+HHF4Ij3vY+wPqHmSHf
l4AGzZMLlGFV1t12BNJla2e7oyd9SeESJnNPNbJMM85NtMBQrxkEADeX244n2MAB
i7cZVbhIOynaPM3uspkrKOeT82SVazOiSb6eUPO6PDHbUHGIG9hlYqKiTRpqxsNX
e+svAus9myYtRCKyF/w0odgcShVQ86Getst724loJiQ6JmdMjXuWq07yGb/RlaSn
Szh9+OnvAbXw5e3+dbHyXu0LLcX1LmlNcVjfPsQV7LCBqnVahgM+sTFSB+PuZnYi
Y26kMFgq54sC2smnFWtlez5yICCz5EftkDIkXBcYt8pjk2EinDthXN799Adv5SAV
roOV92+cKGrlN3nyZ0DUSGixIcpHR0CojJoxv6k8s9vxobSoTidRH39QE86X3RDx
q+IVE9vh/Q9v3SCe5DirDLn7sdSv8Aku0S24VVrAJU7+hT0r8ZLoWyXkSrGvfJL1
PBLUEeUfzsZ2hgAkAksPU5A339l+eCwLc8wkZomvgpAKMrnbiw1m3jvPtwK/Hz4l
stLvAUgKe954A5cPhS8SnEj6xb98w3ZTVh23bV6MhP2017utf9sq5qjeB/nZ1hhN
UUeL+UzK79EdrzPq9ferb95Z9y/92JoRwY3atjegP+8TsjQDB1KYvqevMBHU1eRo
gSw6TwbYqTDdr2hR4k64eLQU7JSzApk1xQiIe1ymXl5nMUB+jWlxOue9SYOVH+OM
toC7qYTaJ1vLNJC36UYD/VcUtwqTT2NA9jOhAxGCHFmUckiQaiIqEmcHVcGhA1xN
Yzelj0uVbae6vuRg5DXAheQASRohhjEBeuOps07GkLFbUjOl+mL4/TuYMxzaOAgk
5b7BXm0vCRbkMBaVg0P7sxHWgeuPw42StbTWqILpP99eCFjNBDSoOMuzu19nMH4d
arYMiAistFI+ln9Pd0Sfa2uXKOIfbdfoTazHpERhxOdnib5sL6uCHlICpqSyKhiR
3R7f12fE0rFYo8cZqPrJsLxRmYL/rTltsue1bnNejSlX2Rm+kOdn9xQ54jkobXZr
RZ9qAYTa9smo7hYFFUquXMg9DeY3vqKlMfn3YAH3HZ7c3MHJb/1vjcRozuKGQmDI
xSWWiSQSxXJfw9u2QCqI+q/2FQZvjbQBfIDYwMsW5Wz9Uu4S5GdzeGlBkIoUTyhY
JjARgAOYg9Wh83vi+cR9kLSvzC9EfUhkNzXxHkxT/Oy0nL2Id1Y+ig16IoQ7GODv
EFHaGdL7aOSZpEaxrE9Vsctz7qK473FAp70gjr4E7Vk1ub0e9wvyNuS2e8qCmfNG
W0Yc56BEQ53cTm8CAYy+VrAMvvdrpeRqXQDTTkUOmgnIV2cZ4+qFfuYbqQGMUuDY
qu3HeFIugSqZZF89BiiYpvkQt9IaZzTKX3S7EZ4dBxnQHMo8ywI/qJBDDnrI+u4I
C4JGZKA0zXP/8T/e7Xeoe7NuP0sIlahHtrNwdfsI3Qpt7so3lKRVdDDSnLKBLhFc
Pai0bnh0U2Sw3a7NfkPfVB4sjkX4erSh/vPY303KXcbp1M4h+JzrJvdOQbklAOuv
4TVxemSKaONKou8NMxokpTrERskAn+sMwp5yUe6urtoDBgE2iR+nCUqX12J1Apav
qXANNBePwbB7zuBt0T67xHq3IotPcoE4bJ8k2saIxQ8ayYCljc4oJ3FNK6J/jNZZ
++NlM8N4nFj+VzyfdbLmUF2hZwlAoZRBJKd0477+jfyC5patw9wQyPLWLYtBjGQv
qflBuuh+65zNjVt98jNwMVfhcB4UJaNR40NLfocomxcF/WV7n6lC0xJckmZAISRm
XhgtD6UTDfgYL9YuzkqH5hY7yRK9Xty5U+WZDS4SZocylHytKfydYPSP6vzAdCkm
4oBDS+TuXlSpq4kEk1ktAutFp8rxnFzF7y4jV4NqumbfN2NUwjsDKdsRTPSf5C4b
uRi4IRQrIuuKwOnAFU84olK2CHMg7pimIrUHNKddyTNSenWuzeaYb9s5Hx3pV8Yh
SeqoxDPDYPgTuxNCN4ZV5V9YIx7ebgPCEbJ5TwJIO3fCO7ywSkpzNz3Af+Q2tTQa
K6xVMrhYssYp0jZKZkpHKKWsw1iuOvN0xA287FEDKIhVI72FAOwUjs8Ay7fETDnB
aj41R0yQNrfSS+ExQx3Y7L7FYFeIZYhNHnThajjrCV3pHQSiv3HbY/ybabDD1ILb
MdPwqqzGwC2xgAHUXUWGS0/+yyp66Yxj2UBEDbLoTbxCrSBbxMieOQcwGDV7jqoy
tYSscQ0f60dns5N0H+Ln0/v6r3Hc2KMsp/VhssPgCzh2H1KN/5u2EYVCX/s075UB
1ubi3KVtB/HQ2TAqaKE4KH+Z9Onr4V5qC9o/xsW/LEQlhXkFnKfg4vd3CaLfcPtO
/azyNaVERChWLFyQNewHfCoXKICHRfr9nVeKFXCKYdV6aq4HOQU4jfLqamJuV1TG
t6RdI6l3x2zzWfPX8TqHU1ymLpN0deXs+2xWWZzScqpGbVOWKsxJJmLYI3u2jGDy
fH+8QdIYngOeTEMl2+R4FabfDkaexZHMihY3565KZHlLnYsCyjz3CvmfVP3mUCUL
J2gz9EgBLwqEVsMQxWhXwGw8pqvmrHehtOot04qmL65AF90tngM9WuJ13vWzw69Z
jhv/VUtt2B6ec42WbYCIiiMf6DI+rCgCJBPk+xz7drKjQmxmO3DNt0n0ODSVtm0n
aRTNIpWM+8WI0Jd6SimGY6MwsS28XTe7tFBAwiyXHBDo5Pjn5a7cpD3ETmGk82w7
yPg78uKFDolI3qHkZcFnS7Ar+EVXCFQBdCoQG0eGTaHbVx6TOcPNKq7RK2qnvv31
P1ClccnrcQKc0gm4BkYpmzrxWr/yzJ9IsDufj3CLgBE0L8IbnEL5pL+zGGT/rrkM
5eabpdpo9y3AVNiVspwaogmylg1xjA4Mt3xblkISZcmq7IdaEhnZfLdVvw86Hqsu
zx2f2uJrMxBKJBqCnEMlzahd6x6CdvI9MYKEOeGq3Dgv/487yAijrU5eojbUcRD1
dtgHZL0m6iTJYS3SJNuTYAwDdJ6F7Z+CXndkC7BU/ZF60cvjwr71RYQTkBBfu0zF
qpD9jGSLHPUb4kBucEFwuHQm2wD5y2w6GLFXr48B9PFDA3aGdQDAyHV4L/8g/jc+
dZG1DMaeElgGJF+d4pTiofK1ayzvebXXG2rS2z+qtIWFbpJSBipbBqGEGJYUFtdi
vSD7ioq9gkvKI8u9id1jZiQAMshj5cI8hMyGW+lzIu+PTBKsGY4vr2oJH3nPzgXr
L3Gj91xKBy0cTMKdZ8uH3ucnaKK9YF/PNZXjrxLje8SjpmhwaVBuHycbmIpBdfy8
zC8Msir8s76Bkl0G/u2ywr8QpajJC/sy9wE3G47kbHE7vMirEt1Xoq03l4Fn8kok
MZxzC0F56n/SrZowfM3V23wyjXPJHbBex3xGEnuUo3GJ1pZb65FBsl62xDUYbo/b
YLOoDMauhObdXPX0Vh1YxqbsvGLtCUeucacYmwPSNBXjPAR2FE0HidPnf43Lfdeh
BeByoUSbviuIWSl7yan/ySAEWUX0Po8r6I6Ec+2PR143HQaOdn33ovPBngY3u5MO
NzJ2dXTcYswQFOfczUhwL7mD2NLH/LZr4GPNkmYKRxsT0O7kc3SFyLP0LrEkuoZO
0Q+xt/+SatTlHweifBNjp8uqunFsDBJQyO0/xlcvb1guO/gEUQmfLwLski71KcVc
jbGbW5gXeoZAl+Hbr9mMRfeI1rAhq7Tl5LoTbtX+6biUA/YIPqeggcn8X8uzk5dG
yGnkS8I25xpo4stfrYDMnQ4NyxkIRllshVErNjFJF6bU8t/RJjtY/uZcn+cVdVhm
IKIT+ixiicZIN1lnw3AcZPtp3sDMb1/O4BjYHTyJGATapM+AmwUNzC+s5vWCTysj
cl8ZdoOWzO6TVHdlIvVwzVZ3WbFVwEoyGASm9MIitdFV7cXebfhvXpB/yoLYysUh
6GYmxUkEBqJdtlbIcXhkqzt7PI5DQJA/bDOMD5529rdRo+7Pl/kkSIIJ2I5CIeFO
Kp49c2pkly2t6n3qFFXke36hPgGD4DcZusOo6yYDT9gu0ktglgIk+oUA+to+keK3
My6UUXdeUffcH2gT/Aixp/FKfvEzVeYr07agxDOkAC5UcPqQCNx6oBAoy2/KOjCU
O20UW7Tn6x40Hw5tNYdX+tUhjvrU04nq+hWrcJvsCSQwWSJG4ov7tMWRFS/Z46EX
5uxEMzh+/qcBmowkGsMSucnv7+dpTteVBdjlO6ItY6IBY0J7oN+vVAkjFxk3/hs9
973CMex6noaVGK94gz3CA4stIU3nGHwEh04KP27A1WcBPO1/SWJnGGQgnhbS/RZS
tj4FT/VSBqlvS1NixT+9MRpBDrKKsgpadoEzOgz8fVr2mfTHew00425IKYiD2tAF
rAUqIvSaL2Po2n0f8PswO9DpGaYkiTa0z2AkbAOcksx0cnC/0Istj4Qxvqh//dvA
TEVqhpTLa6hQzjjSBgZNAWFcHrRdsQ/gqr1L1E+CuJz588y0WslYAvr57tPyJISS
uDLWuqYJEWBV/NkaTxV7frpl6SuZDdnvVd+5HQL5jdvvvvuTF6X/hZdrS4YtBPIs
fNNW5HFRn7/W5YEEcDT4q/NamtPeJFWvE2ObN+Kqt/BOPJHbH+3jBu9vOVbhL7XO
KycOZdfCf5EE/wG+UVmcMUHCfxQVP1TharBPIiVYsa5N8qVC7cy+4PVO1kupWy+w
NlkjVyGD/sPyMsOdhmWgrb76ICriHG+0/B3LCvBQQeP8bUErgfNI8DTa3SvRb7bg
hm1xxJsSDKcHsx2XpTnTL/k+sRDQSKaRUo61v03uBA4hK5vWp1LGvMLgsRvK+E/m
oKYPrGjgWI1KSqJmw7kdTJFAeeOY7QeVh+we66hZj2vJwl2Hl0+s7pWAMKQKEQGq
Slj1ULuTVjVuKE/9oA23UOlWkO73eeWVOVbOlZ+H6YwJ9br4NEqwCJund7ISL1Sq
9WBa1U1sF/DOUIgh1EymVrRBiGc/7RErKpPCS1bipLrpsSsq0PB5lLK8tDBPhHpP
zDn48s4kqslCFO/p+Ik3oyaMD5xnVwmjNyQlslSf3hxNrzbKgKtLhsStXtZ7LEz/
6neTHTUC478w0nIAPVxtOQHRv3ternb4zn6nw5O01sxT9kFa6dW8G06wSKlMIylr
clnmt4CAwW64Llrm9LXIidHCYusb3Gb+99FS1xnA8bHHcJz1UvFN2Wq1EYfpxZ7H
m3hslo0+XknN6jw2mukSo8nCCLvIA/PyBp2gJBwGiSJbyoPY9iUFNArJTDqHmL5Q
fwIfMVBvMHH5D742MRbm+wWCeYT3TcAsqSJIwq89LSRpI3ZcrKzI0w1J7LqFR0RW
l7k6S/AxH2P6x3Wmm2R6eIba2IpDrObaFS7Ou2EgGUcjasuiQViEtnBW4FcgvZVN
fLdu4hsQQgKIc62Eh2HsbIvU90yMQg+qR+yugZPre4CYyOIamRa211H0tJu7S2c7
B3xiKj1HJnbt4k1SHjLN0GpGuGdVBW3KbB65rvoOkNG8LjWJshFQDZOrFUfJ0fup
DLt0Smr7bRoV48FohFmR4JZ4rPgtfLJSh7OAnc1Zou3kK6PPHu6qhvzc7hr2EWjA
KVUUbpRapiLWbPNwt9prPhRq5zaygeyd/Tdgn7uFtEpGVfuqXMl7D+tHfTxKZiQ1
LZ/X0kWSZMXRynMQ63MUp52EjSbXwJwOaio3upasHm6LmFOYWMymEf/n3sCJd3j8
wcPL+6bDiRMQlQ7NdVePUw3D/dttPW/vFO3gJoD4v5bmnbE40p/n7felpHs1apCD
dsxPHc3zDgOHgR8T1ndQuGLPByLCwztm+RXy8H8/Ckg5qSNSe1LMX6T05NnycszI
tp6/5Y/w5LJ3Pldn4zwN4augfKTYGvfNfZXJzH99ukjds5ISFqMVwmI6IuGXPADH
qVzyX818qkmF+xT7Q0pIkrSknzhMrIup7jJIIjOGsIshZNXF18J9m/msu/nReYqx
JJopmLjXyzhK3oOCkD8aGgOxqo9z5LC4onYc0zwSUIBCwfF30VWKJKUTF+2hCH0d
2C01lkJvpzts/GfU4ewOWN1Xylj7JT1NAr6CmmnYY0bZnIb0sGa93GZryc8in0HH
fJ3ig61dcIgHstTqyDQy5hHS0+KV9iYDBt/MLfS6kw6t0XyW/sNkz8JDl5G3Aupf
nMhV7BudyPneL6oPw4b3p9sdiUG6KkCEKZtFaIrNSATHWZBWT2Ag7mnWaUFIM2VQ
yHU9KbaqcZex7OxhNBM3SapHtb6Mm2ZVqVAuS7UtKgX7H5NAL9dqvmBIxzPosb5K
EGETqNXl3irPAPFJZi6KOQtVZsdxew0rZiS59tfCY3fbOEeJIu1KXXZXZNmF2RPx
P64v7e7P8GJ+xZCv3bhoDnHADHSWkHuDZ0z6973iga5nAkMbmaQtQFK+fHuf5oqr
nxmdY2vYmpCr+n1mzYscbqsHIt08FRPXtSPDrSGxMfbxrItmTEjaPj6z8X91suI1
+/SvWNkETh4kqufpCJQNB9/LTuVb7SofFDYMUOeJLcV9cLP/W0w+JyzoYCTeCfYC
UYAyVD9DkI+u6pUirZNfJ/2Lpj+ax4TKT8xEiQAeFKgues4ps5L6hWpSo7KoHO3z
dHNbQsci9xRsmkGgs3kPeRgc7Z/mfPRE2Uc4/LegBZIQwTX7wFz7qIb1EUq2FuPN
a+XUHQecoVOgtKnPsl6wOK871PSQXVAdHqgSW6M01iBe6EKY4RMz06sn4R4MAv/X
TInf3uCymEgVAMvf6OQq9J5HLMTrt6kopduMoYsBESHyezdfgopljNpa7Ay1i7a/
DZidEJnvmbFzfhsBWYPa9SYpRjH2BG8CRIMhET7jrxgRRBb+Q6r2xUf5jt5SyYws
/+eaoNyRRFvKpKw5mNXHZp1DXnKqEcixppSA3kvrXtDuw33ATk0XRAZa3VJSWn2G
nJYTog7+zOYs1lKm6QpUim1PLzlFkpg1IadwM8rJzgJE+kQWGUfVa7wT17Gud4BC
mlHMESenLL3AizZsgCmnLERQgWXy3sdBsTZ2iKVPCzMTUddiUnvqkSLu6y6IMHwm
inrU/YdR6n6bn6d7cCmhcvJnXXG7fKUmQUZmN8DkItgN5MqefMXR/WExRtx1OJFZ
H3jOQH9Cob3XNHsHSRtm2IQtUKGioEl6iIZ4Pqt+sHacKn8ECwTxOw9k1fZXL8/U
kvTBb55n2YZeOXTiETpJVVlxpLoN5udqi3znypiHCYPwhHPrZblwQ9vEj27+WX56
HZukyVsapD00nnLeopT+B2y1SHw1Q49Qnn0IAKbAqGxi7oU9HFYFYh2ocU+eKoVT
yenG+ATosUP+fCCGmtFLDJ01+XoKGvXGFZhe2euvgqtrigLZt0bBgXXUEgEPIa7a
uzARPY2UCmzjWr9FWXTwfqqhfxX+xiqh6XSXLNihL4zQ5VTDWbFXB1w5+axj+hdd
A2gKObuUrrMnv2icKESuGLL2XF8LsU6y+6lU1V/CGvi0wnl3euKlEAzgEKP0EIX0
DPe5NTV0dtWK20UuvUW9e06qN+nDdkPYGO970sNCC36GZhfYgUEZV/ADmwRLzwbF
IWYYscHw7kmDO4b1hi9S7iSAxyvuDW24GTJ4am9uSuu1TG/5ASnXiDOx1H3sbR+b
QKO8kE0KkTAqpYm1xErFojlLbH70ffl31JAxhX0iJecqeI+1e5OXcPwdOtDOabh5
jU8cyCR4zqfgjWKd76C8y9By8P+7mZc8niPQnKOjelmEWyNygOfgYVN5bFlzuR9y
qCh1X3v8AgMYqXCqeC3PD4H3gWt7CP8AyjJ28KGskWi40x3RaidpUeOl147lNDEX
x+B3/WtQJ0v8jrUUaN7AxtpPI+UUhL8qTp7LQyzpCxWakLWID5/0WwgmAUQ0sbLJ
V5ZNIBMr+YO0BDJ4VyISO+Ff7+mwh2r56rHDImyaLRq0cQRGjCQbE7jFKUDXMl4A
JR9/W7gTPhDAu+h8leW64i8gya44ZpotA9LVb0j2C8H9UIJI7Kn++dktF8by97Qw
ZFNNnMaEaLtbUU+I+SS67sRIagAxZ4u0wp2/BKyfvcK5EBO6PvuiPE6/eTZMRHe0
XS1SExhmsygXPLqZSQBZjHsBSqwAqRNHWFakzOzdYUiWl0JRbvExChThYdV3sMpR
W1RxtIj5fjNHm8c8+Eg0aLH5zaMf66uRFl4/Z6cSoBc/G3Hqs4aGbqaqUGeZFN19
Vjxk2bS2TMi7g1IVZiUeUJdUZgc41kU4GmUb7uGQE7odg3KXJh2hG7GGDhlE6cS5
2ZHr6PpHbXdD+8VnK3pPcT/05bpFi7I80a+iH5aNlbbBvHClu/e9cPhHgGA9J4hz
e+FeK7JZ5SOhPHETBgb8LJjKboMfN/1tBzCMjFVE2Y3EMm2kizp+ONeuC3sTg7PI
lHkmGYbtly+lk5E5Zsqy+LWkbTye1OR1zYgL5Tb067L9ydZB61h3UiwAD0yDet7/
1251b42gNt+r27sanIFOb7/ZryNN26bOzIFfGqqnbyXJAPTTXqQjJ7Fw+hCx9o+z
Dk3wV6yePqhhiYzLuckl5J+sdWqMR+fIlJjabe28DwocfjTcKV1tJXJ6BzuytcZX
NjSG3uymJ8tZdokjH77paGTZZZvVnnaup9fjUMoF6G0wFAzeEbu0h5FkH7U8Pn9L
XL/8z0RKThTbDRtXl+COgM5/SxKeIJGZGi7r8rFEdej4qb49Uy1bYueJ5ZobDcYe
bN9n1fox2dXIrkbz4rAteL9x6qCigiNsngpMxYY1ans9DdMlJdT4Np4p6lzakg2Y
+aDoDixYrG2PLwg01N/bhAR8QGNEeBZ0ridUtCdLr/ReI/tJWKy2elyUR4JMbj0G
UaDDS46PrtjUPuwlpuSVH13f7akWVyZJ7n//2jWbZYSeFIYigi8GKB3ZBUqO8IEl
b3MhpWMZ0ZiQItO4/jLftoL4mBJweHP5/nmQrSlsSw5qKarvUa+II4CLczfK0k+v
3JduEObNAQvhmjxFAlg4Eq2Ejhe8ItqsnVo/MegzSViblITHHqYfetU5QsrqvgsR
oyHGEDJH0EaZrlnoBaqV9yJd0fmqz9LWhUi/kUxPi6o7j+YR3N0cKndy7tB8Fhmj
pUeVl3RrIdTaN47YiL3SeE+sts/4k1ESrAKtmffTXWdoGopZ5iG0pTtlpcT60BI3
SAQV9qLRPSdrjKSXMaigf4AeF/mdhMHJJVT/B9WrwrQ+bABfZTl9MrTfSAG6VqrV
QnhwTrfErhe14CzFn9KtNzG8p2XUi+OxdRrKRiv/PuV3CH3B2+2pvKeS/aygPD7g
pWaqyZFynp4/g8okBQOqTr/3RzKicf5csbsjarT2z6+4wJuMCmVf1fPWWjZR2D3H
rzo3dKCGJncqe033dlD+kIbKj0So4NiJKfUL6oY4L1tbZUwKsVtl8P4m3P1ekEOF
QldGSBGAMflY2n/zukCA+ejhZEMdP/hvK3UynvPb+Q6hXUo3Dmkr9bCAdMH62v/2
2nV8CfRDTlLjQLJcuFv9VNeh8eqgP/q1YltTdpMpmLINH4VaTS/hNi5h0FGCNu8m
i/sMJBGna94Qz3tRV4J5j2ucULPibWHzZotzfeZoeiED3cciKkGNKp51a2wxdwy2
3YykhcfXScVaqG7WVho9S4uxcaYs7wMezyKbGilLT4nawpSVlPUxurgaI6N1MyJL
vUWq3ulD3atNf9bgbDZwlD6Fun0LPNVBpyiqlt8UrlgB3DN8DPQpiKo4TFKpS8FH
ok74gUh+eY8sTSB7V+9Bt1H6Nt64De1z+9TUoY8Cspn8jLZ9V0OHrlhAwszacmiY
O8PufoNFBYksOL5c5n9Zu8t18G+ekwifMo1/uTy65vVwlAwPoN/MgBJgvwwdYMOL
4wt0QDQktvLpOXVyFsK8YS4ChCRn2Q/Oc0BxxbC7OhNaVpeJim7YLpp+pPZ1cIvH
mrRzpjD6bxBJFqoIefs8woZFsvzJx2wWji1kcrJePq1SLCJhHv4afiQZL/iKMZLT
5L+QCPdtZLFNpooJ0uNlIB6j+LglPJv+VL9ORR/2y1QYHnMikpOg0y1pKSESm66h
q/Whe97Mx3ZuiwsYOt63i//Hjh1zz6lcUp8oQM1ezjEhiKI4bs2CUAAxfmb8WZrS
HSTXkweoQexpL6L4X128pSE7DYpt/smRqMLRtFZVLojr/lw/Ej9TWDQaEV3VBnUZ
karLMwMKQxoRx8O0qGoa3ZidvY44/m3eh1+XUah2dyYfVikuADi6DGMwjrXb3G7Q
D1zR78zOuGgS6IJm7CHYNTVYF70q8VmSXRaUlk52YY7I7dZjrNoRBGi6bdM/+OSs
sGj9rYmKvfngTf+10OGXfFtxK7oJmpMpzS5aYz0/27YcOaw7sG24BURHBq+fiIBu
f+g0J9wzk7njJQZanMepGLSdnOi8Z1ha7QLHA5aRwfM3dVkj8w6CnN0t3gIemduZ
y6s2IFqwaGuWIUJGqO8jqdcbymrtpvnia1LptwRo1l45GS9RfgVia0R9IpEcDaxK
bzL8qfRelDLaOiMemha30kxyj60GAnzTWm0aoSmxiCAay5m85p91bA16no2pPPTZ
aazzB4gXC27hgHTaNT5eNNrQ0NSPpeReJFH+Lqx8Gsi8VUy9vJgx+dvcnGJAvop2
ENTqDr7l8PPL1ARNIiCB3s/2SrfBTQfwMzEjVQBWQIpbYEj+nebCVenMbYBtK+WE
SEZ6vp9lrd1suajjtlq0N882Y0n8+c4x3yOS4mTPjLfDnElAeAQFDjwm8KAbyPE/
tXtwBj25bTAyP9CBv4aZ7iHC5kH/9iwvFVS/iFyjnPr/+LngLaeyvTjv2lsMhl9+
Jil2payldzM83uT8shp8pwt1O2+EUQMafQvK5nMRivhu8WItWrpoyuBen4WUeeq7
J6S0fvPoQN/qKPqL7GhF43oBTUmJMoSeIm7wVbEvRu9ZWhzxWuDLBxVe/Zpa1pnP
o5ZUJ4+auKx7qhxMEB+RAjo8PJJl57JqxqIH6FKubAxqYfz1o/77IEhy+1kV8ZAP
xNc8eghWmzC+YCO1GrMjLBOLWwJ3w+F5d/oQxnFT5XT7OS9afqwhmkCNIqG4skO5
dHk461E8FHd85Wz2C7TfF3nbvvRszdE2NCr2PltohG8j3P0ruWPXRihs8if6L5LD
tRhM8Mh8DHP1ooos5BWF2ZxymdDbfJ321sFmZeo8PqD/yeFdfEAGPpltkagYHp0a
POe/70bop+NDOBmESRY59PEbltVm061SR+e5AQHIwoKlhqCVZmbOEke7MBrQiWYP
TXwQbPyu5Os9GAe6GxqgaQThoA5cRpFj9PC8FzLOpbNAdTsE/EHjeV9T/xcXpkZf
iWSYZiawW31vgGh19W8/FS/oq5joUf0lW2vzBWkiUuqbjb31yDS1NH11F0GGDY7t
M7z6+tMXqwz3EBPFoEnqiScQVdBXFvrz+34/JDcltjeUk+84tJuWkJbtsYT1bYqM
wloTn868nA+WOvUAukR10qKBMO73TG0KSV1LQvMHciGlpSH/eVARlRvzt4X0eE86
V0Aka8+063mGQZjeyD/kPQYRiF7saqZtNF/tgQbpiPg96Jmhx13b6JZyQGLBYjIh
udP8T7KVmCoUqSkKBZV252PBdHw0XAUIrcAEay3LMor5XFIT8FBeDS3oT2SJWA9f
O3A4vKVQdLt/juwrZZUdQ8DGjk+nGUaGL3QdtffUhgNlJSQWl5pKitb26eGRgpAY
kIKuymDuA1Kspl0kx/uymCZBTx+X7gfSE7zypTuv1bMGAFcSsSFCI5TkvcjROkDA
0NIibq583qTGaBn+yC8vud4kmxy5i7nT5mpykD8QkNnP5WbbFQ3/WAebyanx+U9D
biVg+jXKNo6m6uavgcTAAm/mJF+iCwBGkD289sgRswurtMjROwxGT7JwnARqjpQ7
+qc5Qn/DCvRkGZErwXqyV/VwWgqVN4psSkfVO9FTz490bSBLtxXgim4bik4pJk99
FUE97GraKPVM4KjHsiiB4bwRA4kPPER4z/c0AuqtH/rBb7r/urxYxK1wtinL0Fm+
WSn6g+aZxNJ+GvUkPyn2eAszUrjj1vAlUnk6V92wL9SUs2tOPfNJPVcMI3CZdku+
wSKF1++iAqZ8MNXJXR35m8t5Gl13fWQ5OdoA3jAi991GWMmugSzUVA7wSt0HoS6p
5FC/YNLpFHUQNL/u/BJWa8H8obpKZ/4u3W9Z8fS/rZxhe5y7PUVDggUDfIpzFRi7
IYThoz6Q03FLKMPiJCfmmgJd6y2S2zq3WBbBU+z2YmMVVhkO56dDWfbL94udRQxl
WyWsuyllwBHHvOHzEO7ldGpOhDEXQLIWvND7XxwtzIhcUiBAqn5oo7MncZtKMNeh
E37BNwj0y0RMTfpyq/F1IzEc4hV4sopOXdVNXf7Vt9eY2m9ckc6RI3jdCv0NQ0ma
Gr6a5oCmZTpeqpbkmdX0aj7BdV/Y2OLNHNtU2saPDp6dTiqaKSAO2Sj7tg5RLQBU
2dqGayUVKcpHpnro1x5yCn4Md9w9uRTzk7gIvrY+r+tumCU/fBBq03NWnvJyx4K+
WPpUft1MSQQqxQjPXX+4VoflnADDO0988VEVnfJQSpLq00dqYF2CFsR9N1wnXJpg
bNto59LAq2q4qEWWp8HaKmQ4+SI9QMSWUku4qZEtRa5+dIVYdXM9HwzXDUCpI/09
/RKOKbMD6d07pWBfE046v5NAeHO0vkBYag9woETDb3gqmR2iUiZ+oZpJhUTubPvY
0vgNl9rjKmBb0C5C2KelREEeUF8lbPxEjqKRpVLkGC0z6AL7Lu3Ke/WE3xAeBdkt
fXhFAe+hsmMIG/BlR7MNlLGud6yWUF0cRkDvVyLltTXYYLPL+mdsbYYA6NIYlB4a
QNqnmLJA+POd4BnVPBVUSWER6ddHCeihHLDzW8vMkorByharVTOHbrBcApkosYzY
EOPDCExVYTUhxd9FNat/lGa5xvsegaMhrLcDqyTV2ZsGLx7v8TM/rwx04+rEe48Y
LKBc6mjqwj4fIUL43jguaF60aKfTwUjzIkCXbFIYfLGvFbmPBlnrnbPZx/WplzQi
RP1xctFSk5s+UNrSVde/BzRL0J45Ghq5PkpofML6xysYHtIssqJqG4Cd7rgAs+0K
Wz0B6vDuNfQzTL3sMNbQaWqA7vr+gZS+P5fxgyoyLXo8I76C5Ls069pQyvogwz2b
RHLRHp7y0PmduIkscEI2PSS9HHSSz73mRVoxUbJBl/zsBmfmR+XERUBIszQDKsDd
B9khwwSX7dtod5Yg9nHpMxXRxdCzSmEHhDDKXTwIbqA1N0tmla1x/9POg16ESY3b
Wit6sjwnz0biCosYBKwyFWUb5Xy6iAwJwiz3rY1OEGF/PT5s5BmP+bOMXq9EfdVc
cZrP2d5saa3G5DIr1+fVFhZAzlfmdpLF3l2Y3R+1VnVBRE4Glg7uZVpenKVGbf9w
53LxQXo6Eel3cmwp7MmO/ZAalMPZqWdsUZlsWmgmZ9ae2E1nY0YCTgTgmGK8dt5K
jh9Gk/S9/8HaS4oIzlUtL1grn45qX09fRkzHsnvGde4Tj4R6lNSd4YpZrVcB+iHl
Bnxp3GhGyx+tJlY1oh7HgiCcHHjFPNt/FcH0y88FYg9gADTcZBFXvnN8WHXImaBo
l/xd8jAvBdwvjOfA+H2b6Dy4k14robkifKJ5LyjXCuIljqlSeMUuUJtR90SzdzGa
1qXFZp7pXtpQSPcpNuP9L8iQFfxiFn9SxtrBW6BePf2aJdSVTKLj4kTv9LylUs+3
7bIGMz5i4XSrSPHXDS0pH6waz95kAajcxkTqNC/h+6k1Nv0OXLZJq4SGIMD+DkHe
KfQt2WoAAwBxlmRJT5omltytw73JnHoqfQusre6lj4xk3Web0lQgsOV/0zOd+w4W
zXizrcPz3ZahEkJC8d+KuLLB3+445+YMWvr9g1w1xNmeLhOvlQYYWnxD+4J/ooQx
bmdlgUlns2UphKWy0DCoxj47kdYOm+I/OWtN/P2eVzhhGwaSpBlUYS7Nza/ZtE3c
XPthxKOKdHy+/VWTxtUXEIXU67B6FnbbRBb2YNbERp/fxkIwjanYS3uBQvfx3g6K
JQtP6WEJ6mbiqcMwJ+998Mew6uIVjRROLwcVYnRKFVNzMiLYMFkigWpSH7wcaOhE
+cTvh+/8bw+sEjbYUtm/aDLY2KhTxxXrjiuHCG4xitViJx3fA+pnqFq9KUJvuop1
7VHcGCyI5ta+RqeZR9z38GlHZVtWBRZexs5lTPEEJONvLIFUghr+54OJT1+cnlvQ
65gR27P2rGcqjrLd1iKECpcn8y+6oWF32kmQsjbmQBiWM3WYCRhG4qiRiVXkLBZ1
h5L3esbw2nVd/WgHgsw/4QXntVOXMuhN0HWb/3qzo22/aJ+y9NjdsQVIBQYvjmvv
idOthNLpr78Ng+9Oo96L3qhlXnJgsI/HIKxBsTuM1mrgK0//AaRJatgDNMk3EVjf
PagpF8mFd7kiBzcQqAAYAF7zc1WZa/oLW6+8yC+hqs8=
`protect END_PROTECTED
