`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SgXN8lhKRddOg7Sca50nVd0/257WAyfKko0AschddJ18L9/DSUw6nTfD5vN3RxvQ
0g3FdtedvV8JTS8MRsavrK9PXSGA5aGtqEi2BorDMeRMh6Zq9PHwHBE+fCdn6OBo
/thAB10hKbo61yNVEEJD6S84MaB4WDxmWN0nHGA0JgO6oVTa2hJ2phslgjpsXij3
S9u5mA98KQgkwx4MIZgJyX5lt1vef46RiXH7hE1kP05jTpKq0v/oMjyoosj7nV4v
QOrBSaaq1aiPxGhV8ePbLoaEUTwd4f3UuFJBP9c2j4m3Z+CitLKIyfu33k82yjKo
iZaGjXYnjKeX5lGWSiqEub2MpNvDcRX+Rcs8mcI4GuuWAQ/lJ2JV52ayC9TFqBv2
r7+GOtkYihFITK9XTAIF6UTNuE++4cBRfY9n09uzhTcCITQ+i6YTLr2eNZ1kT4ZN
uMFUTYh55+zSEMzduGkfPDXCFRgIhA254UCqiyXe/HAdAKBN+ah8AVnp7knOoQYB
CUSbt2ZP6QmsN8EhKBbobL7tt0eNqWNyw7Iyn0bcTes+lolNJjsMQpff79nl1NA6
TPOqcalcMc9pGX649s5gwXVulDqwv9YaVBtf+f7I+PW32DuiaPSpuz4FFCgPeqUm
67mVS9OCkJVLdhmNMNsCmCEK1RIzqJk3lv8M5MWIZI8THFIjD910dJqmGwnsP58N
adqeDSJB2qbiRipU7wZsyEZ+XaRhjoVaZQBX8CAcwzkl6EHYrv2B5JaUrwW8NwIL
6DAdKazX6MBRGYcTw1fYbP3WPB7nkfHxmQ5w+TaAruKY6nqHac32qn8kTOQ/SKaA
zL8L3fsC6fkzxJqHh7zBEsl7U/OhcF1sg8oGd2SklycRIB4jPEWngajUvAmAP8/m
89iSP1qSFrGNBgcSBaLLIMNIr+x/e+pF7ICCq2k7HMQyFVnH7t0yFd9txIp5vkCp
2Q2WThHy/k7FlWH9+JJyQN8jmlauPGibVASOdzZ+mhwd7bCbI0IUH+BIy8L0eznp
FLL5qaGz5L4FUATIVICAtVA3fB5PEfjpZS18FXrmbDTjioToER9eDKPsCmwGZ2M8
i5z5equ033oWH9Optd5VBH9E2YDSZ0MBrGdZs1N3O0sLA2UQVDvfUS3hdBARfMTI
dOXLkssyvaCTuc/Jh/bfSg==
`protect END_PROTECTED
