`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pK6ob1uyNy1ZXyQbQEOFTalIaONamxgFnoGP0/2AU69NMPR3r9Y6F+Zxm2dLnODM
nnxHQHjjhxYbyFFp0Hxk/j0kTw2ChxFFnt5iFu0AjDl9h47eVuw+5NzUjdh/nIqO
OWXV/dwxn9dbDHuSb4tgKa8xKHUtiG+UjacMvLCUZ3pZ0usZYciNiJ8gxLwRMJY+
vBn3ngyhICZDwqcCM3qFVejvAHA7MPgkMSk1ee2ySLwZXT+oQeTG0RXiGrSQpo41
8tWKWh/CkhFFEzBZq6GNztbXxR4PjOliaHdumkig43q+aswGZulX3MNb988w2wrq
XtqrT3Ec+nHaoi23Q/88f5Gn0jgKmPhdDFEVGh/9KVUlIGdj+WdcE5gb+JCIMUMt
XtZRUQ4lot6syQeT8n6ONcBJipZhtVvR3kcmpCmOdpZDaxqia5S528FbO9VWFV4V
BoK39TxnXF5XD9vkCq/ioKsyGd8IFBMNKf9kzYh5W0lnkeorJ3KSpOTjwo8v00au
RI2LwYowXvr/HUh/5jjpDXK3BY9rcsl97CAmnQGAl/WmFhS1PYkYwZxMONHUfZ9x
+hvImsbEO6/HyQSQEC9q9A+gvhl/4Aer2oxz9zQX2C4ExoWnQN4pqV5OWN/8ockL
2dW2rfUPVCR56CxdFLt6YTvK2/GCS5cD9qOmrNQY+rI=
`protect END_PROTECTED
