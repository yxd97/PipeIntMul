`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rXZe4lhhAr3sz1O3LWJM9xeHn1SvgcBE2TEtv6HWZu0tRCeJKZ856kuNJ0qDb58o
xzxoQe8l+fCGUOTe1vxiOEL04ubb6ZT3xuvniGwCUycKLG26HLAcs46euhv4+1RD
wny+FTuuTAMS8ok828ViqRyOuStqPnQDS54Omkb2FjUDL3Kf91myvnlgwqpASzYN
37zqkZSIM+pdnG9e2/2B3+gDYpzM8RXld1/lk545SddMfH0/QB+C9CKg6h1NnEbV
TT7iOqLRgFdZ7brl6BWW3znxzYDizWtTpdUQHuiu+ec=
`protect END_PROTECTED
