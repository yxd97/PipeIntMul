`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
itC4DgFfZ1Uc/ZgYT6UlsbZuz2QAujZoayzKaTa6DxdTSqhVdCFJ03EVfyErJ3hJ
PLpKW9GSwpjUkRRPxi58DdfLThCUpec4umdpPqIDPYLWOInAN9zXYlz6ZfQrK+Qy
gpLAwNgHq+jwNE/EMvCqgwbgkB9nAFPB02Cig3N2kMgnXgfF6kILUCj7If0GeUHC
59loM7SJNTa+TDQcTOy2EBobhlnGtNifVtUQG7YiUuzlcSEY0LyCke+xPfyRqcZV
tmV52T0+UlhJGpOf9WGu793DIz2IruL8VImbt0iYMCJS4MPC6XWX5Xig48UxF8RM
cnbDoiEd+LnPslZ3xPQRoBQpZckKkprVodJm+RYUaCO3j75WMWsVfuJ4CuWS/EtN
J1KDtH66Zeq8+njUKW2le7YlrPkfD8k2+npohaR5LoFjEdk0ow2SZooh7nmHyQiy
CZ2JjZWTK6h1jfCXv/v0lFbhdA98onuKGIcwbL8pItcsBsGno1Oj10m5iZmt/2LM
vrSJVkn7IpjGq3xlNQHWzVv4F+Q4bWtUDQ1PXHECr18=
`protect END_PROTECTED
