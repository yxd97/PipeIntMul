`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uxf+IHBL1ikb+qk5WtBWOx6I8/cudxlFwp36XgynID2UeJiyyy+6RbbUqJZh8ri3
6RGgqo3iP/9HPOuO2VHVGS7qHvp00BvenjFRMeANtvmIioxHYVYSzHwGnDkpcCbb
q17Tc3JbrcO1I9FIEQ1cJbOnRlEShSjOYrTQJe4h9ExIGRqSPCk2ObP1Yv2M7pAN
chvJX1lBjKOBr93FiEHvu2DkHhUMLuRynJEGq+21WQKWg71WwSrN4lbOmo0woFCZ
ikK+80CFOAqLrguHUVzeGhTEgHqBNayv4460T0ckyjuDprBk/DC8FMTnNitsXyDc
e1bnEP3sX7STDFcGuRcG3cFi2PzG+E3pFcWQWBGRasz79qnxkXiNM0IPD1+sV7wq
BnLlKvHJX6rddA0pnhbUEPiULQMulgLIlHVZflIu5Fy53EkqTtKBaQuyykBmHoCQ
lwaqdXjct2CoNu+2i7l3Ez4FzrW2SkDSCwxmWS/0iF6Gs4AlkgR36i5XhFJonocA
vZfDDVVIlV1Mqn9QC033EasWXtBAjUrYnV6ZXjHtWPKMZBEAkFKs+IKMBk3MZzUL
aJrAw2n4qcTSz69zL/DzwPklMKU6DDGmDJCd7Ze1lypEejnChudzAbY3QfYa2cth
INxZB1Iya7S7grM2Fq7H5rBuaQVaDTUfzJYISQvDVB8xxevhHF36yBc0VOAq+i08
r1kOHiC4IU/MtecjNSwvffgt1QtaaohKPi9omFcFUcFmvqUH/bjs61xEJC3DADiN
iNfCrEtgiEj+oc7/HuK8KDvlUyP9SM6nkTsV3NKfY3LCg7vtmws/9dUIyDXLqMeA
aFHDqqhaNHY0wjXCfkVVAIKR4mMZkxgXpN4DxqLDEndy+kpR12DTUvtqCm+87iIb
3pMaLvdzVQ71C231aqT73zpXdst0Vw6wDs0CLgNv7OPxux8slqgcfIu08PKNhXII
Jcrs0yR6hXZCFkS2qOMuyYrpVBvFn1B65bXoy3TympxzX1XjD+uc0N6+fiIQA8kz
d6Iy9ApafQ35Ia4XUXS1fy3KzYWvUbLTwwAu1IHiLNd7OoGzeSzi5a4YjBktVxww
hy/HNcFSlHRH6hQONVE0eOGGrTtFKrDHfiL0/WKIEl860VN6WCtLN6mhg/KHOyFV
NKBHKVQnqGGiNbOe9gxJXyrK+xeoBNdaPXlUXe3GK/ZrpFR0hs4R2zujZ32f94RI
ZDz9ajgg5sGF51qGju5Cv3M2ofWFEgPJRwqtukWTyIHyf8pKITqoLW4+fOubTW83
1CLwMZ8GK2sx+gThCYyElJl8KJbRyrSt24lrzceUHxXrBHmNHOgwIatqhmNldDQ5
jK4YYZT+OU9YgauLpycnaISLL8Nk+I21z44CJnXKH/ya9Kid0FXHCMze9g6skXrv
2kqZq6GJPIRjg/0gztiQcx5D6hg+OyaL9A9sxe0SjNLChwF+1ZdQnoEE4G0BuJmS
EhFUJQJ4zbsn3GPNMv+RTbXA9mfCT2RfMwEzUQEX1ns47PYmK3ewzH5h4hbbDfT/
6W6Yz+HTC85b3yglGo5gFcGQ81YICallRLJxBaLZZrhkoAZKeTzIjI6uitpQzIZv
TU8+w5qZmuHrCLqcRre7+Jvh2AqeHSaiiH/P/VKjtu5TwxvtrEdJdRl0HWgyGqRG
bC/YtqXD0H0npVn72I7VGzD06qi0OZEVVvFLZN0mbJSWen/j5EQyTg6+Ia+mLhGJ
kHlmNlytEhbV6eYtSnkPrqtozPCKVH9xbXUJbK/V6cPgrmZup4VC9mV/NT3KF9Bn
KeYw/UsysoPt3XTbzN6J7VwgmtULs+ZYdeUPVAQsbfLA7vhjg16RP8CBPVs+gjqP
Z+tLBNXtFhMxq07gU2qdXGTrRVAKhTjHwvzGtclHFOhpPSLKKPWQFuNRCIPw0LVH
xMhf6kXhRq9F1wWAe2IXkJ4dWZBsnW1iOFqcuCkYvH23CSTMQLDGVZM9A9zhODYE
Q9QEUFiP9JLuefItbIGV8JK4kj5mYaX6s5cYwXC+qLZM9j3gbVAZywEI16XxCn0x
sWFIZ6g34ir+lGfaH3m9b+cy//s74zILNeTxa83Vm8xzPjTRqnEIJWwC+mA6kOXs
mEhLD7sUdfBYWyeeljH6HcPM9lrWhSnj7oYl/YTw8gwFdR8egj2lI+H2JUj6giSn
DdM6QYQM5ERPN3gGdfBZcKl+3bu1fQD1JBT59/w+zZcHB1r2v+iU03aE0pxPJpyr
U/6YBba6xnUqXSuIbcNEaaSLpS3jlbFofMHxTJBJItxyESZM64xCwja5FuvAeOOB
Qxht5duMDCgI5xFSJnER85xjsu/RfkesB8bUQy+SBExeJc9vnynzN3RrtbPPCeAe
eLP5uRvV+W+mOSfpnr/2lAc3vaNadAPrdHfCvqIMrhTQWAOCvqcGfrZSY5Y7hHNT
4BTDCF8zhooVZUFLqhwJmCdSuZN0n7OfGNY+ds27ojy7jqhu4uehP/xP8vKh3cB0
MriXIzXURdegwuZuhPQz4z6sMteLtoeL0gf1QEWisxR7p3IlrO3TABKFNnZ6a9yy
IDfUOsqQ42nFyUjXmHjuYb1U+jtnmUsFasRyiS1qtEjfvqawslZUWcZVPUio5jLe
22ZLRLCoHyOPdSZqlqsx6ycLUNZtiAXvNW9Z3o0xYUDqZ514/2Fg9XGB+PmnwQuU
TJRO9v1ZPluPY58BWq7nTE9AaxCfUKafuNDnto+hv6Us9Xq/N1jtg4cZgETN9/Kb
k8x6+pbCFdXU9HuxtE9UG7PvjWEvRBjV7i57ukwUcjde7MAoVAQ6FvlCC7ih1Bg3
5OL1g6VyfI2gRFjaD2ujTZdzrhBjRtdYS3nJHtl+79fx9whqhEHO65RKxbrzdjhV
xcb/4hQELcGL23SN3eemrjTNFkablH3mu7z3E6d3vefitE0988taz0qAYCxh8cP2
w6aCdxJpKiC/z+PoMxcjcKvQDbzIDlxN9UUxJN8FG4RiVZt69fXc5JdlfZ8yVH9Z
0ee7G6VuDOqP4+HY70PVh8ubH64Ze1IbJIgEwVdhbwXXymNcBzELVZHUaXSDvuy6
0squ1F1SWH6M1VG6YyqEbpculxYU1EQqxMYZfviTAsIPAPeq1HHBQ0JseiDKuvGs
6jwqt+G/9lBfwuo1dqdWi/pSNOgLTSJzdwmuB3Z0ag70piNNnCVIgBY3tIz/7jlq
npQ6ptSf4y8sETUziwJtPYpFfLDFwaQt4HJdtgnN4LPXSWoHj2oyAv8vTCDvRzG/
in2JJ2EY9EHSuinZR+6c0OuVGyCOehLpWJJX3aglNKVQy0jfYljkdvKNfmFVZS82
pGKPrDs7uLpEHq9tfpnuOO6WYj9W9uWLZm4jECWBYUUC3xCewp/LYgoEs+ZmfaeI
7jyb3vbT/65KJVNLYtQf1TyD+s5PkZDJW2krZSIhukekSuuUmsXsTDqNxoXWfAKV
mckNI15ddBg8s86op9qStjdOvy7fkeWZJkpkain2UPyDE65Ji+jTfUPJheBjiYH5
RyF+8FQjm8YVslozyQTMBqO0q6ypvsz7WVvI1ixNUaxzJUnJebKjNsBDlBlN01PW
mF6EJuBPcuoJ+ZXk8obE/9X0Pm31RrhVsv8wbFzzyrgNpIrHKqPEsszFiiRipp33
2uDbXnxdOWkCQarQeIG3nAAs+xJ04iPaAKAieqi5C6UwOk7e2F6OHyeYsIXOZ0LR
b3cgjP4WJtzWPhirV9Ob2RdEM6XYoWOIoJbemUQNraR1tPunv3PbJt5cdDKWUB/x
CbGVSXHgzvSM4we7UtTNMieemgTYLxXjWIuYq8VW+REvOILsavkqDGV6bUp/2RTX
g2Zgu7wbOb5xgDY+YJtEmYtIj9pGnu7mb6vY8ACm+7ffw/pe54xjaFmvapYUNIED
SwV5dxXR6GuuEuutLkq3szlXF5qKrW1VkpnGHsrqpW5dfpA8/k04hEX7FR/NLmN1
jw12Mu50ZC6qzDYPS8bIpAapQG1f8l/SxGaJaOnUjxhAE7qN+3cm8uuSALMU1Gbh
CgXku7JAbasAirdKQss8ldQ4aB+L8SHxSrlgBAr/xFqLRB08ABj/vPwmR/bpBJh8
6MlT/2baNlweszzLUNsOHWV9ktDH8BMX6I5FHnBmnYMdTmFDAFa8heKFG3Hn/csY
nDfoErCKJ4VjvocRBZ/7N8JeoZeqOkGU8UCiNlIpj8fQcnS+LZ2SeA+r6GhpcncS
UHy1OlIJ7pQlvHBX5OVu9N/EOKV1RQkuyW33zxsmKHudZ8VZBj0ZUIqNAWXjLVJ3
5a8X5Bg00BoJV4HwvOwn4wyk5udQI1hyD45O6e5Um0De9M8vKOB2cpvLjaLabyij
mdNQ+rznjgHtpv3Lt3/zVh6gD3yBPPRV1rQ8DKj27nSLbX2qONCdOTacTVN4+a/p
Xa572fct0XtZM4Ghvzd7+//HP/w5CRS+GhXmnJiPgexBSrLJ+dwOCrP4uCrnyzDV
9+dqrEBh4jiH7vFXsedBP0br4TTP+hNjZhIydQ86d1XC74CvscreA7Jst4afMKxj
ASYJ0UfR7V9sYTHSxnfKSq96myT/m2zzpd+8wgrzDZRLJ4OvjVM9XNiGzdjFBu11
C60ILODOg5lMrTsMWZGLxd4M+uC2IW5XS15N+lgka8d4y7qfmi35aNstJEzn9k94
+bN86uGQ5xWXXGoz4LJ8wt397QN4sGDDWrJrveIxaEZLAW7Fcz9Ca0uqYUXJtmY8
WdUXwkKM+0HKN8ObMGK4u9TFch3tCcG0y0Pir+BcbBPq3nf+D2Eh28Rjd56mC5ou
wlY5KmQV6fV/Q2wFFTF2H8CSvvwYFr7KEOtjK8cCdJps0Q7idH93mIoQgWaYfSx0
9QM3hSkJwVj89FtFN0oIv7CYE4K1+GAJcwyX39pjcJMLHQpiDBASFxrhxgys399J
AFrrWV16fqabFiD778KXMoPDDBsD89KRptYWZpYqw9HT55jV6kJqVEpL9I7x0Je/
+sQL0DJ9U5mo7KcEJ6VlBpLat0S4Msa9z5+szvgwFINhFmBm1Z5FLD6i72Dly2s3
hSCPl5d+UjnquRsPsLGUJBrDYM2jQo94C7FaPM6s9QFPut2Adh3ieqxt+1m78tOD
XWzy1T49fUxbjTRWAf/UiRgJ6rPr5OJCPBvvZ4lxJ4/5mNM/OHpp1sh/sMhF7cPw
blexnepNlcq1w+NfhbRoibWsXpnw7mPqbgJjXzb2Pv6mHVVKou0NeLZuVZVOVAa0
RE4k7VWNkzI9bo2f0Lpfd/qAeU6iIOpcyHlpAGdIs4xqByx5oadxJ3x8NrNT/UsR
TW4wuTMp1q7RiSyZ9cYdkqEMP3PlsbJDRnvYPRvOWmR3REiuyR3jsnwbH3W8k+er
3X5ekNCymVPSv+RlAk44HPob8GcMNQNEYpOvYjGPJPtU7at9Vj0pCrI21yWToXsT
SdtRY/GddTQRtt0ZL/xmzu9ExFDgcTyIDj2Zqj757l7O1SFx374Alf2gZIOeRs6P
4J7HEB5Bol1bCgkREr27LIGWhS+0p4h9LEY7yIQT6jq0wdFK3Nsh2Ds+1Uv2Jzzx
MYd53Y8O7a2VG6DucDLbjwq2wJ+EdCvyYAbFXTmUkbjMQh6HKZb9acXUvP1Zh63O
fIkVPkFAz8yySpcUx3fTRjopysS5GtJWvR9UGgwD4QOQcGPg+JJp1U0ijgxiLg0w
nR1fYQEskACSY2FO+jXHqemkCTQAJ0FfjSrXRVFWIfPLF83NvphHQ1hv97gIzK3M
+DWnAYeh7h9OuF1Au9cQlIp9QGXgKWr+BJCmBOwZLKa8s8nntBQogOH4/uxl6BAg
eUn2lX2LJZRU0+5FFyoFGPNgMnyNSf3iE+wHt33yYf+XcoDJ4M07Lke35UL0WjB3
VRolUMGiQ0KVySbnvSQt4romGNvr//mw47yyi2CmigPV9mk2xQ7tOtE+9LexJmIF
0wAXDGSXBFtGygXSH3ovaBSSaBdS+G/bFz1W5M1v7hDjr9s+TC26OIVilPgsiasA
djopI1pYLXNzLZNBTgQEdmvAOfu9vbvkDwdxmub52tvf//OxhcF3tjHwcH5crNTs
sU3nqOqpc3JBcBi0EQPCXyG9Ak+qNx6ACUnZ4RLp6h8TnogUvQ0MQRraCRVcuAQ/
+U0ITwZ0MdDMAlG3Tx1AWz53WZz0CCLpzqkjU7Vae9WlDNLKzvqDGvUcd/w+gP7u
bSOojqLc5PvDSIiMz8Cd2mFJsPg3iLtn7daaoS9v3NcgN8s4WBjOQNik8f4iI/eG
zRM6pYpiwyB/H3k0AYe6idQl0D00JnpRLh25AQny+3um4cmZMm8lv95CwScabRRm
Yt3KpX4oylqjB3e0mDkWfVOAIwfQh98plkeFuwBwzMknr7IdsZQCHbNjBkclqQVk
BOsjxSY79kQTEPxiPkYCrkto/DzG0ZxYWY9TrvopYSrcbbkYTTg3ZxctdL6D3nj4
0jzoMMSjAYMomDxM2CsUR5eXnasKvh1tBg1Zjs4BA3P7d9kaUaW5Yem6FmstEIxG
D6qSKGC6wV65WRMYb81x8Q+y+m1kADlWHtviEdUZN39gO4CVNUHpuhrP5Y5CfMDX
LkUbLgxLBtYJMRVQCgwNOMVnQLRWKjwHTL/9r3MmkhdrUN1MhIR4pL7yVgs3Lpp0
u2TEqVGsYvhXQaqomD3PSg==
`protect END_PROTECTED
