`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EmLsPRsrTjzg4gye+mEKqPbW8Ssy87V1swdhTwrK2IfRfJzeKk7Ocn295xTdmFfD
Hne9Z/uq3PAihpeThh7DCbXXfcLP1lpPnpzZ+RCvqjrU+XDaYv7Gr7+X/CI8G7kY
IgsKT9YT59fBeVojk+853v/umVEM2fOrEu8NBlNZxjiS/J3Pdm7LO7WzGWhF6+tH
63N7CHou6IpUPJ7RA1MkjbHgx2YXR9z75nRAUCKmIPpNx/uGMJW32g0XnvkSQc2c
a7hquuaP+9bfx/x6Dywf5A39OUOcNmdxhy55s+Q/lBydjY26QQUlwlMeXndHtHKr
q6pw9DNKrfctHILSGAAxU3vYcKU3caluAu89N+fgF52kFj5v8ETrHH5Ql79lk2LV
Du2vIksWQu2dLgywWlI0McljJS0a5c7xEo/zzC9Le6y/g5BRO370JUQoS1iTlpOx
8FqXnivSxKcsNSRe2l2k7bJFw7JqjAw+gbIee6iHZc7SfUSbSrxdHPQcCRN0Fr8X
FtxCRZoi4ZHSD65iRS8NqOwHik6i1SRezULEXqp0ggdHOw611IUbGs1DcWWItHM5
3crZlNY9d88NilFONCRyji52GE4b2L2rsj4Wue5thszNa+IkldjIU6UkPHN4cKwx
JMP5ORBfDMfu+2g4ghBYwEszKWq9Cseoc+JL02HcEtsshoi+dyBdFa8wciVrB310
H7fm3U+L93goGdL6PNzF7AWZOaybmhmVj58lCQAG1W6/GAuErAk2tcm6iN3P7ruN
hdKqO5kl7548v8H3fpe9B6rc+fj/82A6kMel6OAUGM/+u9ANUSi7pysrdljudNit
p8X5qsNomG4MQ5WR6h+hycuSCKxEv9p0EYj9mmzmk8go7FS7CXlYnk8APpWiJ6U2
2gcF+rxh1oVd6nQS+mLkEUW6UP91OalmriQtNnrpELBRMyV9CDbhqEo3yAYD1J7j
uePaM4eI6U/6MqnQ8siTrHW3L0LRlBZJr/UErgi3fO7u9nQcEmwKVTzKI7/BXrBB
AyITqBvmw9uNsO8A4ciAQZJso5iULI6z8yikCXGciCCt5xzm09eh8ieO24nqoLke
z/JF3x4ns4t6Tcm0wxzLXqCswLHg1mTsc07wZ+whbjyqiTgH1sNBjG1rIwgk3fhE
jifUDhO+REw5Sv9XrauCsuPPKEANrBhMNrHAiK4GI+utnk0WGUe8pxnlJtlp/Rs4
6FyaPSNXClDQu0KtLEFSPYeSr/LbenxcKfQ1t+Yk3dT3+7tG7IPc/1lH64a2plW2
51L/ku+gOb/1CmhqvuG8Tk3xaHq3UL5mU3MBBWjMK3vyfQ3k16c6d2oFuo59k19A
fysD8tOeWnhgZH/YsGF8FtBCb4ugfQkrObn4l2MPcwGkTFXSVPpZNrCZJD19C5/9
yRBR9nzpjQWMihpmRgwILqOr6YX1ymoKHGztcx20VPN8FwKl4SXSPnhnxLQBKBdi
Iggs6Vh9i3A9PUt41qY0m+dI4q7ViDsFS3FwoPp8Cgw/weBhBKwOyOGTDq94T7vF
Bh82UjHc+nCFEJDIUcvnZHL6beLtKiS2NPoUcdHe/ZAlmakBHdbCjZtRkigVOmsT
7hcUQ8ObBmO9iPwWshVUdQxTRdHjR2uVgWEJUUahOT8FReo2OQ6Yh3NIX85h02ja
8iDLnhWuhFsiyAGIu4xbRhdKjgeFO95gAlLf8pmQdnN79KPu6N99kBmgKA1DIi+u
sKS21X49nVtCu0qMpl8JGgGElwsish9IjVhaaCzx2P/eljkrxwMgKC9xt2pURsrG
3Vse3LGGIn6XjGqoiZPXTqycicsUIiSu7+aSf2X6fZqWiZb+01dJj5dNoi+dxuLh
/8oQCQ81vbViq+1TV0lR7gXIRwsgKAJELSddCp4rhHUxS+0kmTOy7gX0vJ3chXB/
hWEGa4yJYbeClXzNWBgK6llDV12Hzk1zjUShr7ALJfuV0xhJOiFwcmsX4mnWnc38
BamG8yUZsIaSZ5UasYta0NCW6YYqzVxsdGG52wDRS4ja5WhfyTxwnl6FyAuxhBFY
TU9oZDXWAO1fwASpVgGNfoWzkPa/zig5B6UklJq8Euw4MYVSBhnfPsYtqHrzdJYU
RVMtaOXaNYaUI/4sYRuAZlssVX3pBjPttCEmcZ5B18dZqlyI/w4jNydMzcJKZSMz
k0nEsIGuUJM3akXYYWD1TeCwD4mImyH9l+D7TicT5JiVu5mYPjHJ+LMInPOJeCXn
sdY+OtXydl02dciOnUUFL66DblvZykGOHtehIsLHR43mXnDWDlxP45iOrhqVK8gq
03eqAl0thBk+QqZklAx4KEc/YJuFsJ2p5OlmHcM85zVwsfqtaxE1wdnWWOyR030K
Ic5V1JcsZfOA651Dq1RtuVnoHgXnPaIOtdBHLwyAFnkURfuudss6xZoiFPPhWVmv
Q1q6uF0W4umSgzcuWTipw0w4uX4FScDGboHsi3bd5USJ9ggkequHb+jmD0VABiwa
qQxDmJc3lYiOg/ZbCberUJLcL9NJE6ajFc4wyA5wKBUXdn/oK7TyZJrvDJE6NtRq
N6crRXr5sg2oQQiAGvzD80frupmvow9tP8ykTSS6GlOzZS64PPvBKc957CnvmiC9
Z2FVX3Rw07+u0/bPbynIZJS5gWn+GrTPO6wa52MQlh1gO5fb0wxsZTlQqDS8LnmP
2iiSls5HZxW4kmdITa88JkAoZB/9Th6mse3cBdjedwvZGIETmPQ7n1NQSJSuFdTE
kTSMcc7kF8FHi2zTBVP98J4vuBnoEsZmbNtBzaU8qWhF5QKfldUVfEZaJS7aR6lY
sdJ9q6P9mz0hFU5hnCD8JC6Ndkrum4b/HQmbTzDdREO8vSkAyBigQ1cOhtDabDPN
fbQCsCRS5H4kmF6cjRFC89tZxdRify8x5X25iLs6/j2VFhXMUadUBvOnTwK+dD/e
n49UfSf010Z37aUe0wzSagM3SPQX5KteJYdSgJOJ94lRK/SMGjuUyJrvaf/FY662
+jBr8YtVXOj1cHOAtRK9g5XtmmeGU2EfbFIqLfzE4MCPGwOLIwISEQwlxGABlZin
//y/AhqfOy9iYYlnEXkPFgLsO/63yhpIqMohlJfpDprBbzGqYyQWA4q/404ostfT
pD8PtaVoh1RVsvuk52CVcAJDhSGpd5VdljlMNcfAF+8+vHehm2OoCaLGScnTJPw4
Wsv8/HZCK3x7igTiWgr+oVGNRPR/lMpVNKYWtIj2FtITqli/M++D3n5D+TNYz53v
ZZawyJoPJnjajZVMa2xxHuulABP0tZ9yW0/iVW1YJ8YzJP4TSSySM/yogwGxMfUF
6vPsy1kqhKIJmU21rslVhQjR7NUn1Gv0bicG9OBg99dGJVDwGjKcC1ODiVwZni+1
wE38qlxeCwgqylOrsyqeosecrlMh/UueCVh3AUoW5h30gZbtf7XsydpSnklmqWKB
x8GNBCQPfWetrEA69PQcG9fp37rks+TXqzMlEnFXDTPpfnejgpXEtHegSXbzSF9u
wjPa6/VJlODfiJBQ3QoP63faqFwST5A76ni3+0r7YaLcOrWiyeb1X67Wsd0G7vdD
zOANOKXjqQ0J74ebWT1m3vWMGZSvySKkcZkgK8cFtskI9YDVY2kRPhdCZT/y1nrI
gyfTYAJOMNIBGEVsjpvEEITm97oVGuDtMw/rNWi13tRNCTrw7udRIGXH0J5iiWGV
rGHm6SOkARKiLYwj+PR+hXJapKOc3rOILmOMoM53vsbij6Ra1e2mcV4WDV4E1JpW
ITQVSKoqFLOGcBiUGeeI2jT00FdLpdNFHtZGHUydAoKWgF+CfJ09iEEpQMqs7jeb
v8L8RBaU7fpn19oA5zyRT1kkj26XG+Gx/t0wz8RcfNMwFNtptE47pz8+b1x3LbZ5
gZT/zYMMIPzt/4hYWLqoTfy3Az18iKWQuaSNtN3+oA2srXoR5kX0I4P4m7smIPwP
Bg+NRCGfax585c2WgMXQkpLq7HG5XeTck8TOU/rDx+8=
`protect END_PROTECTED
