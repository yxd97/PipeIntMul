`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIIBWzgzo5s8IFNT7AETS2/6V5wtAaP9MkTJat+MxLsk+uZVthJGYfcSAerFKkUe
cdd1pFm3NQbHD5tzQ9/MynCDwziopatF4Pe7XgJMpHp869PleNHLG1NrNUR7Hasd
pQgzImNq/W8WrsD7rXf0+74Sy8zi9So/E04PZCGUR88Z+zej+RAfyNQqyRugVlW8
6nKIfQizwPIr7lCzyc2FL32cfdZeoEVAo7N9ovcyuoQO5Drng1JT7BIpzxhdKixi
SxUiK/F+kghAtYX6zo335YqmKyV4dxshNdXL+PJfVIVJzoaK/Jcako1FeyW22NjG
qYmhIsOreyrXFYlPDqcAQkmOnO+NRriuJjWV5GNPPVylz4rsX3K0WA0xn9Y3mWDa
D9pUn8jPk5TvUSqcoAuz2ONUOR4T6x6RHdH7Mq+daQZwjGFxRgC7NlbJOT/zxYmL
0zrtCnsBe0U9NzF2H7li9mYULZWJEGNqt0DKJgsmtzbH1KGucuOWAvVvh+qijHiV
2qRcJbt32LMyF5TTdVQ2SBowyNfGU66x+jx5AjScw5ehQHXE7u8s3k3rBCuIVuWJ
xWxuPSb2qoN2K/dLADabA1lf2CYoGd98V2XC1LYFO80420UJwcy/5N05BLYG/mMY
aeLZOwu/pcciwcS5a5uoaUG1AZsmCJhelTVR7r/K7umbn03qJYFdybzmEwzHK74k
O3fPl1nsiL/gLTCyqOpN/UidpzCorMyoFG2BGtzdDdwx5Bn+KDvaFnQYpvavX6Sv
BpkIEhvjgiWBAW6uP9E8RPM7xJ5+N+MmKztigBxCgQfX7zXQM8t0b/8iK/ITZHI5
vjy/97iE2aOt/G9BqLpeRrfwSCXjjZRc27bCOa76tagAZXtVykCF+LohxgH+iYVA
nv4yLoAEw+ZJ6+Iv2zmc8s93Y1WqAYkhqXcd7LA/1cnlN5YMx0E+wd8nDpz6GpUi
EAwQGvZDWEBXPr47Dgm4zweTksJk1oTOgtDt5mYfiNDlQGn3ZF53/97VHDNWPEYl
avj0vlRY0eVLUqyin8ByVr5ZoKmH7XxBsp0NpUYGLglFvrw6Gtyl2VqnW7AqzeI7
ye6qv4P+VgnIPRVcSZYxa4NAg1MF8vNpqXOKjFQ9yG2i0GSbWoSM3hcNVA5k4vFw
YiZYMr42+voZix2q+3kVS9cxo4Ll9+h2arPtLYlPWB5JQQuhl0tgjoTa8HaG0EX5
CONuGJmJj4y9gF08RF+geL0gORdJnhy2Dp372xuSk7WWK6gQbasr3zf10R/yNuli
HcJzF/w8BWUh/iJVtODRwgfckiMIsi2AGXb9G1Fv/qo38Wvt7qlQOJ5xaKNqKPKo
Y5a5AegwxB2RSPIPfhvqdxzRBFy4u0uMhn5m+372LSFwp5YO56thDffFmfTkrCk7
bIo4HYK9mfmMtDKymckI97k8hdBcMBhYW1HxZrruD/c2R/v8jsUdCxb2KnVPwDw5
9o6+j7m194O62gTn3zsdfu4U7mCAHCAbGIlY0XGtbuVWNcrExtG2Jkry6SDLeK/f
nezZx3nKzsojxFvtdd4e4FL1ldWSJeCgN2RRGxf5X0aeehPzUOWxnuUJi/Cvai8U
yPNIC2BlsL4Cm8n1twCkNHzQJEv27JFeU+0U6n6tSXVSV2eYzQJXdL7gMM/WczMx
xL4nhHFgjCWzoVQ+GAK/JijZjkHNkCmH6c2s2b36bwcGujyTIFwkOOXAVX19cRwN
Eheh+1VOs+AuWFNxGi7m9PP4WOYU2NZKFQd1XJbj7LtfWNdDJQexsZhgMXhJ1RVZ
pu0xodv+MFRV9pwX5saVmQuZEdxfoQKPtc/XDrMXzO9TeR4dp5x9OgQlPf/JJj+i
yve6wcXd0jvG6xdUVLSQKzR5LuqFojQE9j+wi6tINty1E5TMA+r52fmVyHpRaXKa
hCZL35dkveeKC/5h42JAJlOxH/UIDuCSXH8E/7rqyQnewANIQd8SJLErEwBYu5ot
0EhRDPk4ZwjZMEceFxWjgb2+mMHOPQR1AqhLKKtm0c78C3LO3aJ9KLHRTM7g5ilQ
j93xu0tbstAXsflfr/1B/fhBLmb2R/7sZKV3pzJ7zWnsz/R/dW3ZN1SaVL2zT1CU
8qAKYMAJ/PoNIA1ioft9StByWkFKJvHkSfuTrwZSFnQ=
`protect END_PROTECTED
