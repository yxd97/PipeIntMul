`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lS0Ln4eUTOkDOd9FTB2TRn8bDqpd5yyU4auwJj+pp0DmSpwZQNrnqaJgGWMYO1/3
bMZUg84WP1e9tOuxU6INPdkT0zkv+XxhB29zIkIFBTN2xGb2DAUfYP3a06BZphCC
7bsvx9UMBhEa87OWduyMFSeujZBejQ6OKaeUUZrkStw1GuOXgQ5TUSzu1gBVQizx
6TBq7sU2pDeK74gC67XUFvyNfqxk/pOM0qt2WmAYmovPrZ7MWRCEOXFWmaMxiRbR
K/Xc08MJ3Bv8NZyI+rz0BK8sbO0DJjPQ3GyORkgMq0eAvxLe20CKMbNdrkjO6Rv5
XX6uMbBm1CcTj0+FwByqB6PQ7VHVFGPWO1IKs6Ea4/4S6urXUBuBMnOBA942Onf8
mro+S3oMycdtqoUQ1sVGtVkf+05B/UAAh5tKgcOfQjntX54/8CC5zn7+wdtWGkWM
ucbJA2Dptb9TF8EtAVroFsaxOgmqX+fqjWHnO3IaXbejNPLa7W5vHbfu076M8nO9
22IrKsuOnX9UwPKFbzsNnI+Ybf9MaJSC5TgOqnpsuzO4lxtCQB7FtW7DRpnePZQ1
gT/nAOtL11iggI9ytt0ARE14MiOnUGt4klrQejrOSuw8KUduXrEV5mrk/9P3/PPW
LtPkGpVxGqLKMHKRHIV6tTIQ+2FznTBCyEY505+6hqb1Tw7pscbg5HtklNhUWax/
FR/egT1ZI0T5QjcgHOWaXPE0JSM24JMCwsecMGlJo5XyEG48yKcP5H/NCMhq92FZ
gSE+tGBNpficGEkbJnINCHuX43IfBRIQiM+SRWHJA2Tk3oWRbbnO2KVmRiNjCbWQ
i3mUwRfv76csmRVd/livBwDLFuJHapbBoztNwmFFbxU14iCntSPy/rOJ3Dz/NR7v
PTvXAuHh/YYpJFWhiaSrXvmEu8zjZ7J4OoDGVko6zYBwCVy7SBC+7BKfxcWnAwMF
XbYmnjtqqbSmeRKwL+5Utarim1wIyclVMMYyOjSNkM+N4+15w8CHS+2Kfmr4DHsa
6xVh93dKMyr9bKzmc/qhCzombu4XNXdVBDPdNBpgVUV0QIbUYijdxG9pARstPbGY
ts7VCDBibLvb1s8FSK9uQJi6pm6YgKDdty1jNb2ggzYlkejQI/ghUnK30ccqfdMD
uQpTQEIzuYOmBPnhZzzcZcRftsabIxbRibvhS9itoL1xPSN6jrpW4fup36EyYivX
CmxHs54SI5TjX9KLs8KGm4UZCbsMMqncA2U7Tu0N7O7A8AMTucT2IcVSDVubghr9
/nwa0EuSg3+pEutRTxOGUasTy6i48/AH9tMsMGfHe8Jd+OsFymPirqeCUM0PZHJ3
aYeZJqV1U3botG0TcE7InweRyclbCIBrMNUADkTXkykWyAmaxwOVSDk+53Qsop47
OKxyhvjoqzzgx8c8eJa2wkAj9y0z+DdYiM91anbVvGrkgB9AgyhFv2DYzo7pBOgW
x1qhf+AIIar8URl4e7s1CGQh2noOS7yQde0SNPX3dbX8bvHUw3ADUYt/0urTXEQ5
7q/l9e6uhwVU9nlPHko3gVTZsp50/3ZqvK8HNxJuuMe3tx774rMqBhijZZ75fYFg
pRwQeQuN4Spy0YVlRbU6iA==
`protect END_PROTECTED
