`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/0xD5uu4LZwLXQP1tpTIRmBYUS+3eSTlcgv1dLeCxzibvlWQ8tL7jzIm0GEuHydB
GIBt6nCVgZr+DvRHy5C0y5MrRl6Dh1LE0cJ5rKDaJiOkBoh/JY9MKQ4N+cMGGAR0
Jf2lEtlcVyBqYUJXKYZrPuQ+3WKz78e2z68GNq5afAHtZZHuqaifUhXmNID4amrE
XWFRcKWhOVD3eOiVrUD7/06kRNTZP5L5j312ET5s/T34sBFk201OI8qbTfUtHmS2
uIFDMMpKxvmYCYtziF98bs/PKPFT706rNhhv3mkeMOw=
`protect END_PROTECTED
