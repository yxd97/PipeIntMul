`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QkCtikn3Cvp9pCLL5RAxoOt6uWbl5oJCxboq0E51nPL9NYeN45O27PtqorMWp7hc
Aks2AoUx8np1dVl4OXBF8qhDcnc2EWoRWDLWywnpEhVyoLLna0QMiX5mAfMQQv6w
9VMUiy8NZ79mxg7PMBbLA7/zqieXMEq58VfF7YLn9f/Jpsm0s5snkJdWa5v9CYKf
0Hw6uzS11z4axzgApiFAcZQwJrQnf2jB4OTMi7arnyXnMpWM8ceg2gEJjxcnNd6T
BAlGwQNaWGvb8o6ffoLLwtukkOmJTiKZ54DGd4lBWIe+xF7PdTI132pfPH7vLbT5
RbCJM4chjMaMP2WU+DHyQuVZfVp83N62Frpeo94fAQ2pAtusbKb5cSBzZ4wOBGVW
d48jy3BzkuoRu3sGVM3smPc6Ishp2tL5+BoshVr1cwmdxPFPyB3djOp5XaIAvqRY
v6XaYedWqEfqUBVIN+cMoDRJCkYIXFgeFRoLq+wCrYqzYLUNEt3U3/A7Jhni5q5n
9Kr6l9fUX9xgwmHqDpgb4GaTCcOI3MX8RazaIeHiA/AI7CI09COEkK8RJUqVMTDC
Eh51uYfsAyZ+veRj+h2N0g==
`protect END_PROTECTED
