`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d+vK6y7kR0LxOqEH0z7gN8MzJbLXxuE/IQcU13yXqVDEpEfjiBdfCkhYqXbMGUjy
yQiglMMv2I7OA4QhsAxdABVemY/sxf9ODkkUEA90bXWmSWcR9kDzoR8sTGz2OWkk
1JzZE6rcZsOTDAK4kGYy9fIQW6gdqAJeRGMJWfJajQ5JwfVgCVMSRh5Hwm5ZgB5F
+/8gbXI8eXH4RhLsn2fGlV5xVgakKkeJkaIjaaAbp37YLu3Q8JrwyE8FzEWSslyU
pGw9ZOKb3qe4TTEuP0zsNZmS/jf6PPzxGVa0JHelntVrrNvWBSZj7qGwZm8NbNWW
7w+hiIQaJHcPBFDhLxYzsO4sbE5/P52kBZauyUlEWQ7Y1xg8UmBRSF83XRcbI5KG
edJdQmirppgzrtnbZBQ7RYXmycWLYkUhgcmvgC7ZEx/trgni9hGYmjRdLy5Yt5BT
P+vDKzNFUOE7TnfTOrT1yQ==
`protect END_PROTECTED
