`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6gslER/xeGvA/2YUpGxqPEdrxLUv9eIkF52QfgIRNujMLDFW0Usy3qWzRDh8FJkp
lLTGtK8nJCy7aZV7LnWPLQu2hCESUGZErRtm0PW11NZBb6/RX+pvjHOEw2pRWYgl
bKMWGhGF3FPVQG7TGLQ2f7p9Ssp9noN2gj06lxthTdUFRx9mDURVTyOVAAJ+Of7X
BK9TH1xnJpWOrB8nmAxE8DLT5abDB1iO0OP8R41eGELXXA1XxX/MMps0T9Da25vd
HP8CLnxKmL8Lk4nvAeKHXWIM8VJxHX5W3fwKrX/GBWLkLVoF87vcmJO9b8V4plTq
Agcrk943elXGEvQDwtxamGZrvEbEFs6JwPsjwCUMCt+V7Oy/3MXQ6OBevllArrex
xoMcfIuI0Kwxe7Ue2GS7FX020cKxRkAM+12CLdRONfEJqfzoq0a5U9Kp6BC1RpxO
8tnEsA9d0SGpiSbo0x6dqPYTiDpeow1SOZflyLy1PspYyC4t/iekv4M5oRBFaoO5
HG1qR8AyKL/MEXLeW/95frRc+qMvrWpawCrzf+MBLJC2If2iXWTsAV0VVPdc6CQ6
c4ZoHts9uWemIYi/XFda7BPMjRxCWh16dxxzswNGQEzH4cpB1vJllCIGoRpKOI4W
RSVXyXyIFh5xthNJ0eAeWLbqlfjhrx8vb+ZyFzxJBHX/ReIjdX62GTWK0p8xwaYH
Nun5AQFsvBzmLRjCVzhmcn87knt5BYZQWzpkEIGDBRwAIO/+XLEaMCbYdZNXOS2L
r5vqS+SMNHyP/EksmE3eljgrBx9pNLP7ApvjG55eS/dTISQQ0X0QcDkCwhkLDx45
Rn/dtJB/7marZiia8QqBOoIX3wS8LUoIMm69acyDvjnM8bcEsDXjHG/LzginjqcR
i4/nmfxPJZZghLkC6w4V8vwuy1okbLJi3aRWq5U3Fbo=
`protect END_PROTECTED
