`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VK4sO5m1fekjmbZZj1BWdXhvR2hDevYpdLo0BgG85VQ7TMAE2vQwhcKohZrq90My
KBpVSTSQe89MqayugFeO3k2iUahf51S7puZEOgxWaoDe1cT0wTMjXAmmqiz5oTZn
ijE4ODrSUNjmqPRIh0Z5mHRUC+O1g8sSKT4IWdUlexCkh0hhcdx4PeJsk//sALMZ
N6S1gPJuxFWorNUCRaHVeyfpFvSqFe8KGzKSW+S0BtuOvvbpWRANMHzOHJCUDh0D
nyxa4nfxDPlTKgc+LvmhU1YmY1+r47SqGNzy5YaUrCnwC+Qj7jOZvyKCO1z04ADn
`protect END_PROTECTED
