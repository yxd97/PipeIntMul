`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jlaw37gmRVLtSnOuDlOpTLQBYFMEOvaZXNN73F6GAFaZ6Ya9EOwywc2o/H+MEXLQ
r/0GyVbwnqrnEyo8bro1+Fdgff2R+YQJKKT9JZpmiws9WY598grWpOpvTM/EqyBk
YELByntPIKz3+/+ocmLnUpQQNIB/oscWe85xPmfRceRVP3f6S5GhXDRJOCyE/aTh
Jkwc8LD3mbAY/NQ1nIl+9cOe6WFkaHCs9YvWQFhS2qglMqRdr7KfWsP3vE+Y+iHP
xVGumx5lKD+O/ZrezIkfIB5ie+gzUNM+RClZSkF5Uw1npEcdQjwswzpRzvl3igfL
qWN4qeUrj8jqzvbs7s4vgyH9PctMFoQGlZRRaaXEmXw3y7y4MuzeeP0v65OAVfIb
jylLL+if9iXvmuUl01fQzMhJLr722vDRgz7sT619ivr9DJuX8YPzCt2P53EuKgmN
Gfsxm2mMwKKlab0VkQ4DTQOlwjjP/Z4BVypFz6Wd/fM3Q0I7hdp7D7kYAAHnqznO
SLBg4Wz/lWjh9b3rq5BJO1VNtsC1n9cEDas5f+Yvxnws0YGClZdXG+tUHkqQ6X8b
O5jchqgaBoBGPpSOoniBmbqm7qkCwpLGsUE+t3TSDLQ=
`protect END_PROTECTED
