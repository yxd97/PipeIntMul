`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4dAr1zFbPPud4fFh2/mxK+RDtr9B9AICztJkHGgBLNBI1sGEZ8XsiLdwKIhfgCRu
BXsr6aP2cpcZaCF8Zw659kDWwRlSoQBI7uTJCeH1F7zgz0g+IO9x4gaPFIIeVFMM
c15pXRL1m1+4TTSaQvGZ2VZudNte/v49z1/9WNloGFlGUXNpKIXinnewp/uvpyxN
m0pO4Hy55qT9U8nQelIahEUer0bR38rsrr4KJynBX+6uyJrC1PSoqsWPxQx+otAf
NcFr41r8dGSws0t/O6YV7BayaWOgEYo2I22mf5P2fCJjddtYCQOZR7rAeRzFYB+N
03TixQo6TWXdYJWReoD4kEaWHxCewXXKE7LUkGR4dy+XLHQZAWEav0YgvlcYJQXr
UusIz8SWYNssfKJ1T4QOR8wp/fNoasYTlsT5QpypclZ9m5afZc+y2QEqihG3tViH
uSHoBIXqkhNjFtQqbjU97A==
`protect END_PROTECTED
