`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LHSUJRcMbK+WRR52puAC2bfB1K4UTwLAFoRwxDOSX/xCY2/cD4vPTnUsiqkjsVM+
w/fspfeovtgSW2LJ+2f+ZWdElSfMeskP+l3fnbj8RGPhW705JGZiKTiqZ72uxGTz
K3HfoNhv/w3AvAlVs37K2MP+D5UKl46tUtLUcFVLvHNhD8vRKcrn+5iJzYYolz4W
Yw91GvVjj6QugUDebgn7yQwNCgMZy9l9VqXIcvOAWz5Tfs+8UUksyAfGQ1xRROjQ
JTMJBKcoayuDzhMMlc++tkrtBOzqIN4loN0v1gqqFbx79m9XA5mdJOPUc/GzF7XJ
SquzWZm6tqO53kg95MpTjy0E3B3h/3kSwxEIWHRtj5HST4dtdaQWtYmzSfYBCAbk
HxutN7yfaYv4sWA56HLkXW6Ag4Av3uZbWgnsRvTIGj+tIwLFO7WWaPK6yM6vXTsZ
0vORfUZNTZ8qXYpX84WJ541Fl71e2KN/k0It/wVs4dDwWC/SMx2W2Kibe5MMqcmI
ikONaK4F5SuL1IFx/xpCIH//wevIkPkSz+N/ZYB2D9dd9kXeJBeRNgMC0eYBAe7a
NSDaWmzLmr0KSUnDViK95UeJegmOdHXmdeqGq/gAtSJqL4JZHMPtF6wxE2KGfy0P
FPs9MhSShk7N1mHO0LxFuLPR4NHeKeUn8u2mIeDgbVOoW6jicHvnb35nugnhHaXD
5JlYHjzkbFz7NgETyxNIeMmzP5bhCOc6xNln1QEP/HKUZb3yzGJkCr1SIijzv9Zn
+UeAWKqTyThoAv34IGpVlojdIII2L/LQiM+lCOaQFCeJ6WCgEWoCo/Qv2bHUowv2
cgiMYk6vcB3UL/sPI+N3hPfaVlzj9tcw44jrPW5BOQSo4sx+RRBOn4T4uN0kTb7p
+g0/e6xttseBYOpSyevqIw==
`protect END_PROTECTED
