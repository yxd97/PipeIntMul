`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AyQWr8NHJFqRFhjycYJ7uOhDi1Yx2MJOeWB7XjozKlAY5tjze52Iv1F2ssJjQmzI
jc7n68FF/NsqK93eF+HsacN7UarETt2cvo3R1wImy7qdStHhFE6JvBnQRycXPMGN
5gD2+1ujrhpIjgrtKEvh9IU4UmWU0XvOvj1K15yy6NJ4BYxHL1TI3+NFEbGJ1Wgo
aHeTCbwhDgucHjKdg8FmaEqbWucHDfdS0Jx2P5xCdplqc2eDEva/b7YEyoDO6o+l
RWNXOUg7IVzA/hhMAywp5YSmrVRtbC9JgYgBDHz0JQYtiVNIisSOY72O4asFcFIO
kj5LXXYKZGssWeg9eY0i0KSuJZK8G52Wny3xwkd7Ig6QAolXcBg6aUEyMCtUJCW8
4KpLgkpUpNUdJSGTso9sLkofndeXbaj8fo5xwjcDSSk=
`protect END_PROTECTED
