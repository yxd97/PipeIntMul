`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6gV0glK2JmvN7WCbJnZlaNoHRk06au4nMgtkvE8lSjfVoJ8eghBAaqcoThiq9aGL
KZqjD7JW1IW5AHVPLht3vrWlItn4fNb9xHu0A0P9U2jg9+9ZfZ9X22uNEMzG0mSe
Lkn5kD4hbyYJMDT9OvoW5Lcf550RLENW5qA9JJCjjUDTA5uf1Zw9Io28vnBx65nj
rKI7N+BgFOjBKk6acsgg1ifLlQZ5QGJwSpEWzdLEOpvbONzZPO9yYWd5yg8jGQVl
FpgaBwQ5SAGzq+BDqiiZ0wkF6JUlwRY/I4J6a8po7eqcJcNUih32dngRKb+YVKjW
XZMLUNOnn5i23EJoUKMTESRmtTNt9KPGnyjDt3lN6HUpessM088C8w2LhD3P3Ca/
oslYiFipIhF5Yb9J3TPNxD2Pf2E/3I06vzoJ776QUhXsKjYcCzcjaPVOTkp9nG4T
BuqfkgraghttTOgS77oFesHvO08I3JSvz2sE5GutStrVksy7lsDs52YjA3RpbILQ
U1j52yBCP9Yo3NrP2XO2FXyQxuXZHVoWOI5q09zndm+eU224TxywccZV2IBK/mje
tSdHiOTJxCmLm2wOZ7WxGQyvhaW7QUEauPJHWQJKUlI=
`protect END_PROTECTED
