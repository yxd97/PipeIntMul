`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7S9nPuCPnF19umA4G3L4iyrbC5Zts/l7GMKfofgKGkGnNJqjKmuyPCY9SpmefiS
ZNpagut8KprA+VKRTIaNhgE0KIi7l2/lCLTb82HZFDdezc/lrhWNq0U/sU16Kd/L
yUHPbGmTNVE+oBaBizvsxpBWONoKzUpAUY6s3UW2Wuf4jrqwD2rOkCDh2Pr1E3IK
rDXdFN8G7GSZYSsKlSqY/bFFGLWzTgnIK6WOR0QIIfUG1o4OuMPtJEV6QU5gZvyr
HWPaFGNppNOJin33TFqsqVSF56lz1V87vx9OOVs5d21f5iLsWLPX9lkOHFQ2cYDV
clV9NQ3SjoZJeAXHMuSYsloL80YI+1dR1yyRSWKfnqr54KFBiPF3+89+3SJfp+RK
CGLEhP4lCy9U2r9B8hGWaBvKA1v6s1mL5H4/1UTG5iBEchBYObbyEnWyl3t3OhVv
XPVZ1dIno2bOCfYRfznX0joUXCopQ8LuCKnkN5qcl5ioABB7S6HkeYctfg8mAW4E
eMfGsRYF+tXs/qgPRA2UnicuUznaROQ16DVetUA6tliy6YYNksrs2lB/CNaTtmg6
6HoFU5Tqk7wAMjAKKbCi+8wCKQ1/gSyVKxJFqYPaC6WbrXzJ9QwonkP1/muutGDz
0bVb69/nMu3YdgaOFy5z/3/pBOGm2id2CIm0EZzp3GIrWDX+AXjMkXeAQ44w1ZrR
su7nd0w4FFV580XDUg4Euzrzrt6u2qhU/9Wv9ga6M5+Y+7GaEYlNFNsLIsGnZsdY
flRNjbJijudg/dYRslNp/yaDK2G1QVhK967MrTctLntJxyIZRhs6UT0N+Z3bl2ZC
GJIwBFKSOzpOAj7rAIhm+3OPItgnvyR9hui5nVp9UFptM3tkeIZxZYPJGTfDYZ9m
3J5YbHjpk4jtIWDR2xTue7+jjtvs49/z8ss0O4cpKcnfRJmpFSx0N1+gRvaIUmCd
3l9yz+RTyGAt+2xIol7eOaLp0GNmm4M9da7/3iHL8iQCLG93B5z1gDNOWxaiTXlT
vBN+jFyPs8pwTtr0CibBtdSaicNSopQViJQmv84yNWGkJlm0Dw5mHsGRoW41PQ+q
eAhDr+jJUbfypRvlPsYNQ4LyioebcwxMLacyu7qYk/vLIA1BljitpGqgMV+aUG+k
aD7h1yNykWR5oO0Hl8jOKLo9UMpe0VpXDRhbW2Gou164rwj2YwxleZJkbzaqRvZl
AY63ZYvREVjLkawntwE2O52F2rORPnV35IMlbSLeDDH/fWiy41SOYdGFJM3St3qd
pWdFeqmT+3HeTpgalfAZ/9sx/1q+eCldCaJ7rmkvNr8eddMb+fbXYEvnNvymQMHK
zcpHVFoKLsZN8QNdh0CWSTAR/6f5Dtnd/y9X9XFm9oQuYR/J5ZAOvIGSYObGtFhQ
WqfsQiAzrIwFsvn+Voe4zALjAw7LjlP+K5+bRiBqBphTDFp+/B6aUnk1elgLljbN
Q60LHxxuinIi/q51pID8DnYzwqvUyfHeb7fpuvRDVQKpnNNw6i7rO4ylVy2Gpqjj
WWJCm7yA50E283KMJZCI3AdnH6U9D5cE4X45GJX2BDzKQ80Y0vGGeEzsJmFnP65h
gRp+Q80/Y1rV8bOWEm2w4OKAxSGLbqv6WtBSjLbuSbK5YSj40PjJZbH59U6kQPLj
on1se4Q3a2yQeSr2XKLYns1G6eC/q0tQD0/KsPFwiASYJZYkoe+R1YrfpEiaAcu9
pZ9qJ9Y72iVaeKbja1fS7Z1BjC3yDaYp2ahlvM3IACNrVGd0+g82/EiiSd5tVsuX
j/0e7YOc4BVpz2bnfPMNvUnW4vs8Y7nMqJWoQpSjApuZoqMIXmTJ7xTijI65asZH
8pZqYgoEMpsQBcGSnOJHB8oWfazFWoqQKqOM+4WpCILUPN5paHDU02RKlrMf2Ys/
rdA0RptbcPzW/woFMSBktwGnxk2cpjZ87AxxFw9xGeKsVoXkQFjNkh394EU2EOnU
RH2Ul2S/PaVvGPscuJ3IjdUGVkhDxV8gx1VXkqlPPSRnubw/YUMYkZ03YfbSTd4m
k4Yu+B+C/VKBgzy7U0lha9iexAlT2+c9iUTEs3o2gYSF+J2VrKraNK5Rb2NSrWAc
3INmb2/EoqGSRvSMNCIxtsdN/UVWpZ+byzEcmD9vA+D6j6EpE/gohxTnJDDkHKQn
1dWg7kbldnwZ/0Ry8r0l+/vvNFtY8bSWtfnRg7z4wz1VTRt4/mr3bkxeIe2+ukCu
oxswghYKLtXFgYBrP/Co+QKYoklUb62tpRfxi0mkTCfV3UBZ7EYr+x+h+7tNsj8s
13Y0qsenxOyoSZi9mIf3ZKfmqH/jKHY4asGnlEIdKCYcz1WzONtsmeoIdYsvGv4k
X4FEqe7mcPE9xEGr/wbs8MgVqx7Gx2ggoCwnqNDxg2FzlBBbKa4YnlpuJgo/oO2y
`protect END_PROTECTED
