`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SSE1gMq1mWTJZm/AiGfIInKLydqjM3hV8S7/3yjT441oq9qefWbWT7o+LYc5Wqq8
vi4Lt6XczUHBlg41l2nEkrbIZt2YLFDgFnCBokF+dx47s4GJi0lt1QUkjTB75r4u
4NQmsK6fZSc3p8WOZppq2A8XjLRKp1otSf6k0DEisXNO03F4F9vbGuWG3inQk5Cl
D3GVps8YbxETELO4TGpcqNLwjM8GYtvt25ZcC9kTVsQgETMUeOCY+JcFIWJRkPrV
oiP7lkeZahAw99KL4rwjL+oAxy/d1wCSqSWXJ6d3CmvvIbk+M8uCSXAqZbI/kysE
00ljgzt6V0n1Tmrs7Y94YTvJDoeRqfz05to9vexsRaU4DyHXoNeI/YSm8v39KYOQ
`protect END_PROTECTED
