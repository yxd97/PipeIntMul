`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UDjGX3qXjZI1s+14Nbv41G80xnFKZioAXTQnh5Fyg0JiQBowQZxcA2uEKLqfiu0m
j/z69J4VLcgSl9rYoWvy5uFIa59ppV1o1oIZ+MPeycrYVTYLveJFxJwZdA4VWnvx
yrygOAJ0r7mbl56MKTWoj24RyWXcu6HBAksizwYeabVg7Ram1PoankeHvZdaBo8p
S8iGZdpNjDLH9d+zu06j1nhcBJ3wu/CB8F23dB0HjDbwGBAbAIS01L6dR9xkiT87
o1zC7m4QZya7sJcJtGjShg==
`protect END_PROTECTED
