`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9okg9puu+vKZNltz3Kf104SW4Ed6fqyouFkImsfmfPg/Vg9UZsyFODhiujByTD2P
rXzsyIWj63HinUA1PHznBPElorTOUbpedMTJ3LU3udrGHBIYzO/bQCklWz7RhKQN
XaZSc4zpkvkfIxeOvVR3GO2ovYfHowtpDanpYpwGZHTQbP0gCVaE0Dq5KRSY5SNv
nDqCPK/hvpUt7JuT7ph2a4s6VnyBiiSrxcCppKe8p8YDBiqkvlkjMsQJQDl2p+dy
zADTudqX8ZsOqdIIxJwO2UycJDbyCQwBsRsSqcXQBByosfYTIIgns9FjaYpNZLii
Ya9c6R+ZJfySDVLkDoNjOSTwTIBsl8mJVrc4pBNoWI33ZxL1Ien/za4Vwy1BijZm
LsVm6jgImrwkJOn+1PLlknNN62/JJ1+4lMlntfHxVS+TpFE0q5SfS2MwRbKyHkpE
kyTTtM0a8Gc0cEe4Rjrp8qpCMzYyCuneQGmvweFwKcxb/e+E+l9e6uwqPmEhf9dv
+sz2G/0BgijaH8Npyd/Ifn//Z+UX/dzkiSNHQtxPdiyl8nyhxS1yVE+dCmreH4rD
fW51KHg6zwY7js3KkTWSJzAZ80azviAgFshofbB7qOUF+bzsHALOfHQLQh6QGSKD
GDyoDp6AeYoGovL3tC0wg4NTW1yfEydgh47dynhIKm7TkgKof9LT0+yzun+rAi6k
iJcp9/bOYO7QxxDMXtYEChVYrjl1Buc3E5zmjwJCxHurWnljlCdoQSVT37b/idIF
UY00/Tpt4F9Ta6RcsY7zophaM5uCXOxdSGYTaB8K53xheUXFfAOF0IiKjsihkh6P
2itVqsyFBXBQjNhjG4OhC9/gPC+MbENdyzAgvYb8i+ewfGrPDXr48yZkv+i+H+D+
8Yk0b7xMYSpumQxfsnYcsCl0Z1xmQtZ/IIZADDMq94zW0sYyiDpNDYI05+urDzHc
4HNe8gxcXh/DeLG8oft5T8qXWIbKlEU4pml6YTyNmnyaOU1Z2Hm1US7ukmXj2kyd
Pj6VFYIDAZnd1ynCb88clcTAFKJCU2Vp12yZZ/9P8UbdCsV92UcO44r3keWRbJY8
F0+XErUTj0PnuF9YTE/rBgyORSYnLTApQ5VQfgdfnY20Jf1TVDr6iVf5EkvajFly
zjp1LaatKXgvcYlm2LAecr6xQwJzXLRFNduszXtmyGwRJzx6N9XVhaKC6nz+KoTv
+zAaPgjGl/Seo6mEN9FHJYRzM3BEGuwqcVku67HhjYvR+ksb0rAhNfsXScW97BP7
DpRo89BNW9S/2R9tHHQazVQ5GJ+l8268wC2IiTb1y05sKyoS2jRfBlSDHPONU0ew
ty3mA1kNTFh9DsmRTadIG5gebApc6VjxjjtzkycvD1xnjhC3/kYOlA+L7/TjHd6r
fd2rN3csJ5/T7m36WaWd1IXokDHEk1JKRkXvH5xMjIkVIpCTtyJoiL9n+7QcBScz
E28daC4n63Q1ZGkQbE8raDRL41hg9Fd0Fw21MGmKUdV6meKfRPWZSK91MwjtZFUa
cvruFN/cjghcF4t03SYvYVTbrPRxxiCoWYlcZegNxXXAqcPgHaROY37R7UlRN2Bh
msQVSc+NNDvIwDwcO1qqBcSVTo+7MUrNccUqavOo25C2p7tPCu1EfMi9Jhfn3l69
DOfjpWPjhkAq01VSjMj7Gx6ATvWC+asJFyB0iwH/7K5rNel2xkMBOQmnx5YzCorv
kL1N+llFhX+wq5up5vdw1cezrTv902eeVYDEXgHHV7un7PbT4ZtpTdSOsoFa44W+
1lFyRNP3XOqqjiDcmxmk/TxG7BFgQ5FFBENK92SLJWsGcINs9H0oXmvAn1ZrTQ9K
Lmu2hToyGHpHsRh/PM31WKH7qjAWL0W+iAfgS06uATkIrrh6fdnN3XNUsj8HO+H6
yE8oCj3rTbg1DwlrynVHRTuUVfbsixkMPcIkrXsqHgjVnKspk08OSHnF9emmn1SJ
i9t98g2d74xz7ag9XeOWRdGKJJNYYKoIBwO1uBRvfUGwCdlcPHOfe4G7KJ+Gxq8P
vqYQBojsT/Gb3wlV8Qrpg0Yuo0SGtCdKtPrdiK35DKtCdp++zO6pT35/KweFd1K6
`protect END_PROTECTED
