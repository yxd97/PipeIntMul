`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hM5bvjRKOImy1j+Z6tS8PKKfnlStR3yFtu+vcOEyoWdR1WZ5695OcyZaIOnmpcBm
1el6C5V59lP5Z6VGg8p9cs9eMvt0WD1764VOKs+bm0ILbToHZMV3/gTsVAhASSbO
QHlb56QMqRxZZtq/yJdCwk/MIyRDUKIlj7dIzSHUcJhS/oAw3AUNaHpckRzwtMdd
SZswWdPIgMyqEaCvhSQWx7X07zSHwoCpgeDltrdXJnw3ph72Tb6IOTC4Z2QkN08s
U/PLH6GV47IWN04RIsBvUNs17U9kiFdhdrdsyyJ/dYmaxLTW9gcfzbjoVuh2kgP1
UUatWSe1flPQzLp6jVBwKxKKrfA3W27dmMUIOU7K0W3OzmmSUD22lLUDDGh5An1d
Er4OjQ9VnX4MUigySOwgqMpzX4x3g3cp0AsU8oyTYyGYEvz4+WljUA7qmvRgryvo
3hzXoajdnYDnCyFSUdLv0UeV6DV8DH/TOr1sP0PRUozYFO040EcQg0yOgZGCIish
chgJi+zfUEob7kL5EJWlgyEBXFSFS2NWopwQsh+uivzQF0GY8CCsIaK1EHMEaKdd
8q+i85OJLhz86lTzGIRAcjNCcvnpm55DhxGjytDdzM6zcT4PxaueTMlDTPzTEZxx
wPl5RWHbeFcU+9zMbYMF87tq5ZYM193xlcfYdF5HRTiXbpGucuIyM0zkkbtd7aTq
Dij+Gd/TBR+7m0Lx+zrrhpqXSKVupsLhddcHntPbfEX/528dQuY8qX0tInitV9YC
UYce5nxivGbzG0hr+tcZ7cmOhSbxdJdkKb9ZeSi54C9iOVB1fsijYr6Dh5ATQFH+
WqGXoQa3e6SpwlnkrhrenmFnuIgGSiQMnlNZkte6hvWbt7K6YqaY8vyVk4pygPfr
A4xAWXkdTPjRRfsMVfUpuPbHX0cWvFRIU2mj6Wp+LKyqDrYTgoM/Sctq3QTw3yJa
oGMRW75vLU+GgHeEQD1Y3dwLfzkvf9UbnGUK2uQ7Vf14/wOw9CWHZqGtLaiedNWu
Xhjs1/b64ZHHsTlKrxJ6shgcydTjPbIYIFJqxOPEx0F5GYQylHbrMV2y0mMCW38H
As7bTEQwUpkxZV5ZqvhHFuYjZw7l7sJHK3sEAasWM9rgVFHE9Y28rstpTCEp28Dy
M3XjRXTBlNS0qyiZGaBFKbYoHwxN/Oo/uOBIwhtP9RwVO6/ZhbBqhhjKn7M2GG6x
k+sVg1TUznbAUg/APv8SZ8zh8xM7HBCf9s9B3kSbrmKBYONKYYb+b23rmpUJNH+x
zT/12sHiT8mcROv+mrvu2iiSZxolbSZNuAiKV2Cr5fQo4L+HOSdkLWuSb0UU5fPk
wNnFWSZ3x6IxPVWfShP4LzWS93C1U9hzcLUDD3CAXuEm2+PwNQSP+Ao7L9BqPr81
7vL5Jh8tbdfEQK44lcwd499y7hFwlmftPv3jDl9p4x/k34NmGcAJymzwnpPvfpWn
5ZJT962cBCbGJDh0dGz0TwdFAvf1+KFkyUGjAmPDrdHwtQVpNPHkjVHcO2L5OIN1
pVpVSguEygBA+IZtQEovCqrNBfUOaC5Wk/LatMiGdnHDTKLelYvETeTZiXbZ49g+
rA6YsDfiOokxC0sIN+cry5rzVE+XC5F7Hg38eDz/ydEEWub0sbw4V3EphKeOXUWh
0Z7euygliRGM+cF1MGx8Ek9D00SuzBoNr2gFr0DjLzd4vPR7fd0LXTwryMSW/YZ9
OHQ9WqkThxJTZfPkfbOzq2LferxnfYYQN/F95PgAx0kG40zrjirvUMtLYmfLu0kx
yYeSF2crAdcnRPOQtXDSCIFmzERGB+sdsgC8HB8ovvTCpP1qjp0GS15fOM8Q2QZq
cmilunGW+yuzvC+uI9Gs3p1X1oY9bDiW4zraWgRT3CEHgJpc6Q/ZRq9qy6lC9Cmb
J+WBgDNqmRKV3YunrspbWDeRcGNjf5q7qizR3HvEsq1L8PJwf9xEEdSppzx6Umcn
EiIcKSg3yktc4tqdS9sf2MJwBAPYw/NL3tCyNLVhdZBXf43Xo1Eme9E83W+Ryl7V
wOK4C0ZbwvlzQgdRSMAylc9l3/BQpQVgHBaBzUC/BTPEd6rmANhWzpi9U8cUqAm9
YXkcHq9XULrSFY97YtPbjJs7opHlGluvaDDT7BkCHTgpKCJWV/t6itubBuSEbXda
xhLBeAnnHOejByXEtNubmx0W42C3JKeaLJ74Zyyx+xEwHd2CELJZ8WXieFrwbzHM
ZhXLhjVwqFLPTVayn9dmqWQhdpeD38KzfDKBgaL7I0+GdrrUPLMG5xJQ9vaqxc+c
N/iilIDj32mWvITUjjx/iZCWHHE48YM9hWis49jutlwHxKHRX+wFVo1I/PxdVF3/
XXnayvML9J5eYqr8SPHBFM7HFm+Yh8pS0bgt79aMvf50QINHgtxDov1U4PSO14N7
Cp9RCFb9l0lQCL4V3oVRTVnUv8QHmGasyN70Km8X0EPdRoHrFonL/YhuKUAgo98r
Qwjo9zwT0FJWAjD0jdTx5GpGqVLqqeGL96Szdv01xgTOR2PqL5TIDX69a5rVs7i+
SWHOBlXx+KYgVIs7aBj2NWeBTQbWEIYbi9HzvvTG8SSCyw4pKU/elmTK8xwE8aAw
YbOXHV4rj3pmUvM/8fBrTK7/w9zZxbLnL7CaKTlPO78+bl3riNe4eD0tOeM0shhQ
fY9S193xoIr7JlRYaEvrS6DPeFXpBm1TtEU7b+pBPE/gKBFURzX3ohQBcELfyPgz
ZdpSf2aFiwEvWiBlDdAG0/xQQVe1tbSkGvA31TESZEQNRWFX5Duon4Uy59KtQAj4
3QUwEmMxtYOwFKZGg0FQth2EcCj6/bL5QEj0XpU5rAGAwZ7ygDH5G79fSI74ANOQ
UGpou9L1t6mYXNavRrDNYGCOkG0B5uJkkrhOHEBc00N6WwCADt2NKlwFbbmLKkXH
rqH/6fjdPYpxwfLrzKjnaxylmIj/64j/r5m2mPphdY2+48fVPGfVJC94bYpsHyca
DSdyXGfG7TzuCo5+BZ59kl/vPNsa2YhkLB4o58zA/Bw/wNaqJDHH/T7qwKhegR8n
eABsiggXVYqIaA253TRNy3kQG7wg6hqduUsZcrAff5oz9DzF4A7mIjctq+j6Aequ
KT2wH8TUZ2QPh5n6OxNOMv4U+ki3+m6vHn3JkDBBVpXX+Qd9EzMISbY1tjqCu4Og
x8+zmrKvOgykF3KMThCb+HaJHZ71YLYe3IVnjluQ5rgvgVwT6B6fQCtxWaVOQUFw
r9q+EWiNKSrsz53T2k/vs2f1JJkO5GLbVZLp97t71yV7sO59Jb1RPvfDWD6Xwpgk
Er9c/YoDEidAaZXy1pPXo2Uu+qTitTiYp6wH6YUSTR9pMwao2M7zcXHb9PxmBC+I
MHtGSuEE228MZTN4rZSYa28VZ81UIQaERyobUGwLwMCjeiHEIcVFXcby4IRm1JGU
gMRSaY3d6iNqYOfwwJqv5wsuaK4djGU8g/v2e6krtmn1EenKnnRKg9OIFoJSV7F8
E8ThhaXXzU1MKSePwzNseMyVL3Hf4ld250KT0thWPaRMS4qaRE8skhb0zZmGZdpk
FLF9dSBigOxsUqx6zSl/R7QehovK2im56iAUZzE3QD0KG1vpQlfbjN41l50NqMK+
ZaMmHRyn9qMlxLIfR5XTnGfbpmQXJXnk8qo+qpNqtmMTc4mZ9Pzwnzrpw6jbU3HC
vSOQrxg+Jh0eBiby9PaddaAaXo3mMh3YOUFTmhmbprUB5cQDzuBloSpT2m8PnBFC
50xPihyUxDF54UMSyj4U9sv0wxSZUhjAPYeSAh9Dlg7debEmr0axieG1rWgmNFGH
a389FU1SiIrhpJFUjFhewKDKyk5X9XWC4/vODhOwnBauJ9jILtsq/Hv1NI3rhgIU
Vk7reByTbRcGPbUttYtSb0C1Uaa9yHkTLo61d7HBBBV4VQj/cX+wx8TsZ7L3TtpK
qRo5JFN2cR3gQ2qiZQU6cFqS2alZ0eDnCpZvxNnsQmxVZ65PA9IXpRmSQ3LfqMn9
bnJyxIpDfPgsiUrTbnkgU0JFYsbUzIaAh7Psk3dA0jN9oKNLHXUMBB+FBNpP37XS
flk/FNqDtx+UOsvNDqAv5AMya4/tls+vmCe1u6PRbGfuV1ID0F9V3IJWMLU1w+Nc
8840mBZ4jceOnda59G3rt8DNXAVoe9XOe2D2aIxF3CPkFyZc35fSeIgWxTA2eWeO
3O6a/EH2V69y6AdOjM5ec9OSvaXVEnyXkAMJQC+sDNgKShpDb5cnsvgxWl5zr6//
Z4hCndCUSD81FASvVNrRgVe4ghLN1aaeIVAyZSCMk7TcozqmInRWZSch5J+n96N9
8B3jFlwQ9UfXPuYJzorEqswf2mc9PLzISEvrng0TizrVjZKkWk1j5i8/IUBk5bbu
uYe0SXh+obHC3eVj4Kw5huDMQgJWyLHsPCWFFqxK3TlxriElyL/ZSgChe4XOAsWp
2aVnUUvhcXJ9EG5Yimk/wWPWhdXBdbJA5dQBJPlrX22X3mp6ph1P4uCFW53Rp0FM
ZGzUYvNt9FJTaaAD5WtNqsXMGK6HAG/aCRcInAAPkHKI4ewAMwfiIvi1/0/VBhEO
PqLHyMMYfsRfV6oDdZLMXPhhfAEYLJyLOSEBV9FZ4GVfqIE6SgphuInsi+nbtwFN
hu+g9jvPKa6PeK/Zd9TMPRBwwj1Z9zIqWdsSciTdlJpGQ0AvbdjsMvNpJzHFmluV
sjqEhcZEOm6B7A+7FvbgufHpFNUqUDn51u9P4+5S026hhfhInTPh5qxapondUx4V
l2OECaxxUjAMirgiIKWGPe/gKV3jD2vHcArBXGxWkhtwQBzzquPL9mQw2co1IHM9
7/QMmP4nOEwNIEhuH7hrex7t9SO8yycO6Ekg2jY8uT1zBkjnT0VMaxN4rI1fe0Yl
c/pa9rdN6Pt2CGyVWAadERCajA9yzRImXEAM7/r7zH5Q+kWn84zweVyCegPJMbHX
iULBokY150fDlJHCVk3xpjrL8KmyLhCxoRew8cH1KPcD/O5DOvxtZUMq+H/mL1Oz
6bb/ilMVCEXG6X9eElhPO2ZnhNkhir1S0+ghf43SfiVsQPBb9PhKbZkQJwTSK3tx
J6/DlGGK6KIM6nkErYwUAn3E+/4gREz5BM9W79A+6Il6AIHcz6RxVnlq80jvXCNq
4QPgDua9qt3ShM93HwXSiknyKE+j/+owyC7shql21PMgt/9+kyGc4uewJ9Zh+gtv
DeS+1BulYLLGWn9WJErXr6UQ4hxg7+hMaoVVk84gS9SCTsMxpKRx7Xe7O8hua63/
OZR6SqC5RuGqsWTwS/ls2gSWhMNTxOeh6oZyMZyX9aYPrIK11UjpnEE4UC+TORiJ
7smkzDID7XfcPK1oz7a5yWNcEOEqzGdeEnY8O1l6w5oSTOMFODxOxq2MR9r7VuVj
30MCrTgY5pNv3EHX5m7YNqrXiqdWxuVdAPxgZWNWU1NNLAIdN0dbmWwgvXDGp0O9
AtHEpfZCwX2xRv4yHki5jFnZ5riTtFlxmBULMhiNCjyxrMsbn0RzSDH5yBfHTUo+
6HbCqoH0E/8dmeYDoTzwFm/w7JtaJ7wf3yxbA/mQNjiiKGl8hFwyhWzq0qf0XXeJ
kOkSVgUs9MM39PAdTLlNSBhcyKrTghuf2CFBKdGGgM0LEPTo/37bcSUfwWF3EndZ
JsDbRefaZADZ5/mVruKx/EgAVbvMRA28e76TuSC0+yyyWGz0h5IKu2K9PjyykrO/
/b3CZf0Yy+zNwEXGqEYvwWygN/hbsTGOlOMSb0T/wN+DQ/+mM8QH30/dSq1IZ2JM
9R2FsEWeaE6pW4yOvp0EC/3U0amga23iA/TcYTui/KHLEs3YxCbEZ1xkwBP6gujj
A7WjkyEaVY+GobdjRZz7ykMPFWVFMvN5xi9opay65BqVf5yhBRbsOyaku1lxaF13
ywHsWs0Ypf0q/6/U0RJZqbiF/YJ2utwGfu9opM9zp8FeI751upExWPM6BXoDVhZ2
3labyPLEGdnIWb1VbVR9oP6w3OL/Itw2POqVaXwTitPdS4THgLjKu7eyg+jPBlsq
zMtB7mDwjGrFDGjpNDdOjYForwKVkxINXtg34I9NndNmTPmU/3bQiyVgwShoqraq
xt8iJG4taYvqCicqRaAGP+QZtn6H75llYRJ6PTjDZlhExS68kF5JYPSTQX1oc+pX
9WGNGoWE7c56sf/KW+i4c/khLipon8I+YYrI0gn70BJssj+9LK68ohZqIpEGOSYj
Ipn/Gw2nRjAdBmM2N9l8LAY4Z782QyjY2zhC+y+ZtOQQzpSMBjRMHB8AJX5mhEEY
38mN+9bi2fLlVaWBVfn1swS/2+dLUw3KnIG9/IDKl7lPKw+xD9iB9t2wYn36xyBd
ZoJRdJgzL0RlbKlcwrSpaRkOsUmLUTowHahAm3LaB3JLJ2ogWZA06xgL77Zn7Vc3
ZReCAz1qFXQhyQJ7tbc/jMs4QXh7J8PZqUQWA+ix+9aFgE5uznQH4Yxtm8w2rjwk
L4uyjisukNi8Je/Ia+JuQM8lSUIfDaiz0Zknt9KiPkaT5esAdPed9sRODmlQOD2Y
6V7CQenm08WEeOZ2J0E5htMPi4c6Hv6Agt207yVBwTeYMIx5aJPp0jG4/58IENFj
DpjeXIIyzHKTwNyuG8agKEaYQlZN45UCs72ZIbqoYQqrEqWExUHZrJtnlsEEFMET
6rsdzXTGXy3PdxOt3UCj1wHITmgPpJ3Lf+Kg9mDw/i3av5C7R/p+ZPMqnXIny3i2
gfnrksFWx2pFgTixXH2CDxzjFSsuffjtBhG/uy8PEeuOLrvm7uhWGx2+zTJVbqwc
DOVbKmE2T2RUGzrdI5ccSxCyYnu5jMgvi81p66FdEY88VWdI7gvAywjQ/U7rALUJ
KbbdGU1DDrZK+awj/seXbsfoaSNl7TR3u/yoatA9Q5DiYHqnezmGiOrckFh206zL
WLSp/OhmJCrqIsa0tMi7gANcswPCcnEofnY/oXIae0NRolJ7TjnusmgaGOMaaykQ
C6KidSG2fV1iI54+dQ4tbf1MHa0BLQSrmrmLv0Y05BX45XAYug4xFq5DkCN0g7tf
eBJP+/V0cd/ZWfwpiPE5xWExw62wdK3IWnsnmINylmnLrE14poLPff+PFcQStxyz
gXfT6lPxH8niYyNHmD3XpUo+p1ozupKrQdZfSEmdhxI05DE5eEXMBdooxBusukCj
zXmPckEWzjNj3O1AE6xM5jeqP//8sTexHwgWSbd4RCJnhKZczXUasbjG8D+DXq8n
VpAw66bHzFwe8szBQwFQ9osbpWIae2EfsobvR+92vBtwGtR1NCOIJqfFU5ufWZrN
aGAIhF/KJie0oRhuZpxKK4IRu6MrkxRsSQImRkrx2W3kDZKxs6ybAToocHTsmD1q
EiyW6O4NnyAthZSWzL/wprTKCp8Qk6Ca/KTxA5x+DNePfNFGgPf6hJtYWxPDXx1L
r+obsr438L3YkmD7ZGrdhYLvNl95fMD9Y7ScCF8lZYVl6g0kpLTR3eb6tXsUcx8x
nwXu1hj/KzDn3R1ZDM9PTQ2xUdQfedTZBO4l9rRpIbl0IlOK+tMSdYobfXZQIKHJ
xuJM9KjzMixahe6qjc4y9zX+aoNParaS2EmyHN1sW/1NRhPpwG0RHF/tY0sBwRul
vCKS4dxe6U2RasgNMbHD7I/tUe1cwefnfh8rKp9BzjXGUj4jwdt0ia9vNJ8cquqJ
LXH4CUNqrCsWhj0dHY3lqRmHU3KaxKb0kY/VPJr1RFORDSSEC9Qta642xwqdf+oM
J+48hUgd8oIma69avlr6vio2UfR6fFvoi6CTb39pn4Z713J/drQ3zjAhLw89N1yU
I4eKSMoFPo1yle3+HsraOggoSdEB42DMI7MAp4ItpxU3ep6cHWlkmXVfwmTC04Jz
oCvuZcMJXz+EgpLyH2H9UjBntSjzROJJ2wUP1y/Xtx7beSfa9J/VkPl8jvatOzTG
j73UfF++SolW2YcEMl++Ug5QnCJUGSFjGeKEHLnclVnqTac/T7RMyZWrNCum0Ytl
pJCiFEcuHYoI9+Du83/Ilme+nS7haHc2cEs6C2PbSOhC/hUsszy/oOi5IgpuSAYB
uVMQBIxutdY1ezM/W2jc2QhUUUNC5yVamf+ySB2R5GSSiWex4WqWd6W3yZVAkW6R
2sHsAtiKgYucTTKFdZdeSv+H2Kajj//ZsLnbhBQWnRDIaIwLFWX8NKZj3dNvpDl2
RqQViNDP+U462scPmKDiqDPq1J8yGC2I4SIDp1grBvEgcEiiSVosgmt0WAi0dG47
Gy00tOshMuKDb4CtiV9eHqzECq1LtS1TcqoLWEGP5iFg/DrFtB05EcudJJHn0d55
qhMRyEmHzaKxlDkH4m5uybK1hYe6qTc2ubo6X0wlRqjls/q49C4ZfeZPKxGbKeQk
P8FU9AMLo07LE84v2kJBYeHAcEsZ8in5N0f4hIhG0cR6pn4QmZsqrwKqwytRPsL7
TSwJ80B2Km7kZy/id65AJyPK3OsV6zVkTjK/7sHxBqBMrQPFzJo/RySgJCD5GQYJ
3tws7Ue7YMihmPUlwZ9jSAGOtm3xCRyLJhUFZnk9PyJ98XdwgxOv3Os3Pvly60+p
ybYbtPmx+wmPer2GBZ5ATHgaKGdyw4aKJ4/PUrQ90D8gIPWMxgEfgGnkHuZ7viHD
GLHis1+f5OdzOs+wWHgyYT+iUwhxNb1QXRvBcVo1TgRZchr3nQyq6AFF37V661ty
fakE4vPtVwrsDg/Mf2Qhk1fBX/tuUXi3rB9yQaxwYVvI0NIJrchoT2HCv015FvAu
foiROnBsL4ekODvjvGnXS+PJvAnQpBhnNR10Tjw7yImToMhLBgerBXvbAGncVrqp
+jyWSdFMHRz10CdHjHpdXXX5UmfAdTWM8PvpYulhNTGshYIaXZKgv9ZjhYWH6D9S
lzyD6F7nWTNBtKhEc3I1KN57tpAkkFsCaT/QiAWKG+o1tCq0Op8hwHRWdWygaT53
ABOctw4vE8/Y6I3lZxm85wLbROh0BvQsWP2AnoSVlkBbCNzwQPvO6x8YFN8whHHt
b6AxI1tidSmTyEJ6+EapJS49QfHso/V1iDAtICgvZAjSL32Naea9RCDvUMjDz7jx
nMk5vF4PvBYTtFAHPS8TKfdclqtZuonPGVw2ulpE29AOknyGe4Xw7qMYjb5LkbBC
vD7r8r9VKYC3b4mULLL69kJZ4J0ZDmOQnohsEgBU7vT2LxpE8n2BkFJAGqrtMzk/
E0oqt9kknbq9ex47dlcL/1pupyDWI46oYvUvsgbYelo8J9XVGKStiTsG8LH/lq6a
wNBfJsz7YhnJlJCcNeoXlfhG6rf79VE56ZC1PbG6Z20beYYOfFWqH4DzvA8gFbC0
cOmQ8OAAh8tk+0hkTzjJLtE9bIO7p7DopalzsGoEiB1OG81u0agVA12lK+dTLf/v
C0WSnF/Y/c/0REPSO72m5wzgL9zQeES/YnJVxnAgSp3AX735WCtonQjrYuEjOpLq
4z477Lp/S5KFii3E1e0ojcG5E4sHzYOKjw5RmGOjhrelmgSgyq3t4pH7PEDtnKCM
X8mOPzpjrHDKD2RRU0mvkT5lGbdKh8B3S8g+mkENnxfSLPXIKm20jJ+VL5QKEcB4
YfKJn0tVEYc5HKQTgp39nqH4wDjk5zHqCFH8cMfXpL7YE8IJSU1l1xd9QZr+lR6h
uBNIMQ9Ap0hWpTAk1Ppkj1WIedp5YKBi0YFLtmAkRqQVhubJ+lT07dU+8Q1MeVnK
b5qIsVAi+HL+43WvIb8kAElKvCojvgYdlddXKbb1yntLqbICjYxTkfqYHXxhBhwm
zXw6yFvY5PQHCBryKGe7NkS81Y3WpCJYNbvapc8E8AS8MiDbWXZG5CJ9N8hZnWYy
APH1xLo6hw0ONodP/AqAaCgagqwXEbBNTx9voL/lR1OhrDYewF3eCfBnvrM8KUa6
AM+J1Ecle0EcGOrwvJhT2atF/cKILa5N1/Emq0uSP1rQrdp10Nd34tlMWsprlPaz
/aLCCYQOAqgbyt9H+QVudUXulCAyOCy0HYJ3B0NgteFJr/u06Hz1Dgbp+2esLj+f
8yQQVUQRgJK07SrZsWIccNMQcqR0KIosPNour6+ysxqYYbJ9GXfg6NcdKGvrQ+ck
tyb75B9TKIsK37muiQIR0ID/twcdoSlFySPxL7rhSnnxcOjPH5G4XMtVSsKxCBJb
AEK3n6iMBE01MZ5USdFOS7LgIPCWiwDOvHypH9Xa1g55tmjsbOKUufkkaKv4mAzK
maRPLUIDgFGipeqJ9F+KmnIcfUz+3iU2G3RvgSfDiKmA+LsT8DvQAWIYCVTdacfc
ayhUNCxEM2uMwhMvwNUjjLDzteugG2KkcabBbVnOc23YjZoH7C42EcPerHUKft6r
7Zl7dV+cnFpA1rzwRGIthMvhG2o0mSHxQe7BJ3EqDzezHKdwLfTyxJX5/CAQQRTG
VyCHeSkDZQotsQ9VBXlYmM3Gq1ridsXPP5tbI9xLkkFpSx7yh2kerPsVuyV9mjpR
NZiiheOwFeuYdZLsiCMv4Tr6okHZpYAe8pZERMLr4gY78P2tfKjkSpNsGaEkv90B
kHerOfktyY25E4QUIC6k9li/7W6yKocDzIY4Wpra8i3cefoG/Pgiw6Y7QnXEhqcx
fKcmUg4Czzi/kOpfxsfMTr0b2hXT7KowV9qbNohUHz8bLUjmSMcIkleSIM9vRk05
V48tSnNguRcx+Y5XCEP76T7uZpK2NtEsUriRqn2isv+i2Y408YbFQjxWGaih0JeF
YmzRPxd6+2ja3TwAJCSqs4yjCGxLBl6SIX/WyMMF6rltz96re/i+pyMvXsM5JJtf
UQFO7HO1kQ4T4nAqrfG/FpOxveM/aDTylOe0fcwB9D51rJ+LzF2gxJphVx9DCzlJ
fjW26z30ZYqkbPpCV38uX8/kxbgjOAhIHLFb5kzdrpjjfMn7z6PhfUKM+VhpCw+3
rc+cO3ltrwcgWLJVBACTVZwUU31j3C44gjusHHNB3Mo=
`protect END_PROTECTED
