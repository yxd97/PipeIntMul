`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QlIr+U7Fx4PptvGGytynWqXRBnifYuaJjqSr3G0yMSIoMigyL4jaKF6hqZG6UMWo
FQncShdx4JORL6iEQ36KE9AWd6s8gd6HZHROXVqF66/NBs34t2JuxdE5CMR5ZfxA
c4YT5kiGR9SfwiNNzIqFI+CWaPO5OX+nO5bgKlv0ZVh6N0ViBfeCOiYwJkjnuExs
oRVvA81MPn24qDGd198u1VXtZyqpZE8RpKV2pIpkVrxYRBEm5CWL1xMGSjxlj7W3
3+K0+zvGhxs/yHjikHKY5A==
`protect END_PROTECTED
