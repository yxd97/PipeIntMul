`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gfEzErCWeoqM1KHxwJQwyzRjlGUdhLwDQ4iwm+kYYYAo1FA6qFmo2b4lnuDLXInI
afK90PHWZTBRGmszX4z1mfQCAJcE2bxX5fmJ/fZyBSFxcrXmrU0F/GlPLbQU6o8R
PBbSRQpctuyvtJbfDe1KXjl7caIVmOWaSSTa6XI5x0EJgUZ6+WmWq/P7cyaKtwXZ
GBgdNxd6O6HsB1a9Uf+MhKn20EBGZC0RJAFPe6AEdv9vskhKBWC8OnRqzItur82j
k2QFKU41g239VBjZoYUuCRsd5xa1dzWDBM88ZTIPqwbWVuW72aM5i4XT8sMwqhH9
XP1lsrgSD2GlV+SULQ27NaGZ/XQesjeKxjEn4RyM5mrN8c6Zt/Cpl8G2uvSRs8gR
F65I9EiLHdZiSXk9mVl4D14RoMMud7CMeG62FLMqtvN7Shx7YsZ+rZa2KL2IY+Ct
jchn66slZWojvSPl6luK2XZv3YwKa4+r4QD9aI5HgwNSo+Z1Uw8jIZhijZVn6NvZ
`protect END_PROTECTED
