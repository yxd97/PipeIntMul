`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RURfufpSkynAkDWLselUwiaBikWTX/l1CGRGXSew8Oi3/PlHuMEwlWl0RJuYce8W
i8yRuWQdGHHpgm3sWV+QS8mKSxyGvY8FbJ8/1iirwcbpaJL85RnNu7gTKR/jxu/d
xHq3nPPCWKpNSpS2Ojt3iax9SwyzXqPvv98g9lZy8Jtc15c6l2tchr0Bbuvz9Agv
wFHOEhCCn0y4TYKC9CJC2va0YMwNV3pYFR770GSuVvjUgTEli6ZtIoihPCx0yjIP
rPOtOt/N21lGRo4haYPzfrguVk084MG7EeK4XzmUe8tYjx0iPZzTUN+2KuMchWBL
xRkKVpaFatSGc3VKH03Gh7Z4w5zNUJwhdAN3Awv1O5L228Ypk9BZ0BdOVQK80Ipj
8mj0+UQILyhToT2/XgI3C02vab7m0Kt6JzEqRpgRMsyLximHBVbZF8HoJVysFMtG
FZgdHvOB3jCDdMPGOpX5QFuYLATfLbzdoB5slPH8WICM7G/bOt9IPzRFFZMVew16
xZIs0AB+3h6mJyaM364l4kuN0MfrsLU37vWsTzBhtvG4xBVCf3ficwBFqd9LENkb
bYTqBYWblHZIATGfFOfiylAbpOPjWteEqOkPucYIiSW6dPzMpGTBnsLvcazyPJhG
fEOglxJLzR7N1AGXG75O/Xn+SALBTia30r2dC4OylgUflb/IDhyTg2YU9yP+3uJY
KXoZdAAVbRqpaUHjDSvCohO+pAA7+Ij55zsK4e324vzmOxqpDhHRzOpBjw3392ji
/OKzbYfiHf5Np0Sda+Y/6ujUdZjdVXzG1nL72HaVjCxtu8jtYBqsga71D/rUviOi
FB2ibrENEw5vJif5LKBrBQNbZJL6289iTPa5BixjAOu76FhrEnZsyCM1rYFgQJ31
D8FfG8DWAxbgP46aslUUEeT+sl6YjodfZonES0BvJQID2TVWIf5dIE+IS7yrShjG
nQREMAeUWt1zRCxaIUBCXzDmZiBc59PZTn0BQPrDn4W3pNeq/DFftHzUX/OlIBc9
wWGSd4TquMe4pLNAdDL6LPHv+EUUZhv80vf1O57WXqwfkKu2BwJmE8WNkHLlmd8X
qkSYnW4OpHSio5xKduXSDGKhY8gIgcznQfqXfowz0hgaEzAZb867C3p7nIZQ0123
mVoDOkX5VoZEC+runFYZNYaTS+Mt3Yj67/Gq4VOuSPp2uizZJXyEbQQxv/ZdxXzn
rh97MvWAnCgJB1TrmWJkQdGnykyxr0kfxASlPHUJfk2OEUl/xV8NY0T8MOct6ulI
QeQHLiEXj4jrXY8lJiIXA77aeQC5LZqNJM+uVrfJ5UPmv4XJNrRm2BVQS1G+GSAC
A7XatXSOrH9zkDpq5wHuIYqNlHvHtbpSv/w86FD+DSxYn+k7hIb3yGn7+6Yxq58p
HHTOTKsl6WBS0a0pu5HWmH/OPX/TKbWUnN0+Wf+I/cVNY71dVR3xfOVsG5eDdcqF
EbZpeDKa2TA2wcZK8PUCH3n2Py3Cf5jlFE+Wa/dWs5FL5WPhPgQLuE1JbY4FZVdC
U4Zf2AP1jrZ4TajCw/hUGwmCIQH83UKXqbtcuSgOcFnK4iO/rh4PEGhL/Via66y7
OfYKjfVVvQBDHfWxvcBuNDb72NyBVAJ/pB/QhoDGHlIBhrDUfgb8ER32Sy3V53u0
TYgQb9URtmcwYLFm/858CYkk769DMilDAoKDEK6kuKdPBkQjSEVT3sKbyfp64xvW
PcMl+4SPlah5UDymTgfYxcLZYmAJ8j3ViZ4xolhyjQ38r3BPGF+NLxSPq6LkbS3J
A0Q5fszUsReanX6Dv2lr70Dm4OCgwmEEOua4eQHAquq99sF9TdjGRHu3ACGq0L99
+T+whgnygNdMbx/h/GnXCIQSN5U8FLF4h+kY6+WKy4n9LaizGBmIEvWHP1L8DMCD
l1NEWzym4lLckBOA6g50erq98gbjibsxb6GVEGcvVAmZSwOg5mFzz0zAcUHBtT6Y
IHmx1hE/1ggBYVmrCKUIzkYJ6NvTo5DtsgDZOuY6BzkOUicgbPDWslXAQXjD7ZA3
6qY6ji5V4sOLXB6FlOrsmjC6HfXdfjGeZe/Ub7gjtHep2gcUciAnm3adkY2kazuB
APFaCW6FbPpLsmq9OOW0AhDUqbBUyOp/xj7MIcDz/qXVZ5lhwtXFMD764BjCDe34
FZmapOTinBaOuR/bouPlcWt27SEZ5YR0BDOg4CgZzQJ6ryFVPZrLuGo8CMFiq9Xl
m+CSCX1bFP9uozVnUIbBdbbdWBCzbiQGnGZIBj6gy+49LONc+07rqAtZfCWkjXdH
J70nkx2BTnulYB5/4pQBkYXb9lT1hRTQW4Qau6ODw6vcNrR7yV0ZBTBaHIzZ0qWj
QGnOLrOIwTbbzKSE5tdIUd+kncS8csCmNC+qEDWpSLJ1RnQem6T93//hdXR40MXA
nj0f71jWL7x9x6ZbpXD/vXS270e3CgxZWDMuZqpwAmZNAsLvHXiusb/EnIwKeRFk
fmD2lCEyagUnlIYqHVPPsCRb4Qxy0HCaxcvU8RiPwzD3FZfxSdLcjXmCj/Xx4JSm
eciNKNI4F6TPMD9BGLQC3+Pbg4GAr4zY+6hjuxZ0hwnT+0kmdmIs7UnAMrwTXOpP
A2iK7Bp/bvDk9QvDjBcNl9K1RJaw5GcEfZDCaYRkxdnGaSxfYff0vxDeXTDnxv0G
1Ilp35z4wVjUzElSrmv5TjzYHiZLnuYGfz31k6AmW/ZtUByCeLgdDMI1y/lbOd7Y
0Urz6JN8WWbRpYoQ1eYbHU9kejuLPSQ6453mkqZPJYOiZGRk+4InHpdv2LSD5bqY
NoN0wwYAPvNkHTymEeOaCVyhGLHqESdAutQTzRgNATyPJWT8mtzVJZnxjKKucNWH
gx2COj1OkPuPAk/kz9fNDKvKW+DPREHc9y/jBYVkVCByu4696Yvvn8LGCYt56x+M
9eE/ejTYePeZ5EOfokcHNgfcV2J0XNyRQ2T2G8wQYJiETgOyxaw6B0So1HS61NBp
V7nDvGf46dHwOniAuUaHBEczEyJ+id7x0B7/OHdcp/QJGZdEUJOSq/ps0812iyGp
uUV07DCxhC7dACCzfGJaVLEqL+dcIEWQWsoBqTGR052QlrTtbvBr3YoHwso2U3Ea
FmtmYeaStsAQTW2SASjLjl2cFa5MLRyaV8kcJcB5eHKCWtI6D8U1i8VMVozaxRDn
sVNIi6iAhwBZHtQSisj9nP8/crBGN0x6KCpc6v8h+Vfq0pdW25EhH/X7+1Pjt26C
Uf4j1yYrnk29yFbRbt/ho9Pc/vD7KCSzU7adh0V8Ivcwi/BmdvU048YFC7QpB+Ii
LjLCTv33YwXkdm/DBKEr1Jsnp2jv+LbHVztYWn3Mnc9LRvoan036Qx040D+8LTw1
ogMrwFwzEQ4OXhpWSH3fZsTDJjMvokMfc1vOQ4D//rXyCoIm3bWW5AHcrBWiEyCP
U1sqAXBdsYgQ/C22M8/36yHNsmJUvflwtiOrQVoBPpT5jfVDPga5QLQtcfey47Yl
OIuopSobfS6ZbBk97tHqsljRnVpDxd1k9ayp5fpwJajqJvhFRuTCKCAkJ2L0uBNe
5UdWeO6c80J5P8gOO5jylzK6WETfIyVadUZUymFYRhhbhdxthNuRudwNWLY5c7Gc
UReEXxr2pFMvfl2/3cxc0Q6TAO1oTZPID5lPUwD7sXWSpZnZLvRw4BZXYylk8fW2
qrgOI0ywdhFhOojvmxTAimF2UOblJL3SN+Wbm0fnacYIb61kYmQk0eNtgdlympBU
ZK2j+uhXbEkIV1qFGqg1IJBZe48iLvCpXezPLN7rwUFUHdMVYxv+kvFrV1ycGUFl
0bfI/Y+Cwaz/6e7OtQ02/5lv1XxlY+MKemk2iECzM0gEsRTYyDF+XH+3HBu+HwRj
Xw4gE2xflyanzzCtrKcKfytw13fbLopNSgPdDQSRCxCGYLnvdByqHBMaZz3cnlpa
H7VQ7wJ7OKk926r8UrmILTcdSPerYa9sqe20HGv5BPVQ4aRwLmkulvpFcF3stS35
5Zex4PtVVfsIALbx2cfikQY1iEN56L2AxXkWpZPZLijeWGkT7WoWeaFpSC3UU61k
sAITuiOCPErEQEW045fBFBSOLJ4wZ6NxL8/ltxtrohTydtCxPGC57e2jXpoubwRq
RgzZPOfmt6ose60MrdVzHK4H/V/RepIu3zakaEwBoKY6pOxZrR2E/oEWBijp7CD4
apLtUzygC6oNgNzM4nKLVshAyHdmLY+uEv2eAbIYjvmgkVfL0vETYXKqY+mIvQjA
/zC5r/B7uASnGft3urscbPdN/lxfVYEORLlGIflGEbiAmuYs9MpwvJcfFqrXnMLS
W9M/wBtBWPxivr3mY9aw0Vcwen1RchDvlFs4PGw5fr0jIws0fGDl6ddbw5XFnjyq
WOa6+eO1jQt/aTjp7u969onk6dgA2ArJG/10y+KspOBeXB7IeETrKbuVUyXBC9p2
c4A7ft7ShphNAwjl01mZi9qtfqCM3NtIQNMqnVky0soF+O5/G53aoQ1uKfOWJ5SH
1vceiVHoEGCnXbncdp1SSqnTlIi4sdvQCyRK2BSlN2GdYs7Zl4owXMsPQuccGFws
jxkihLWOR3mMHO5ybDu4R7s4MnMyHU6bml9IPRydFC/8zjhOufzz6mZHCfOgodGy
PxLZd+LPd76es7iS7NvIQmmvbqnuzZImqv6lNQNFu7jDgze3jG2Q7qHfZFlQ4lJy
J9MU3UZ/GlcjX0oyvvdEvPxLhr51TURSvXt3oOZQ0z6cOOX1iSfl1FdWRyjIrbGd
ZKaqAsc/j6N40Q9KXHQsRPT1mM8iAbJ1f/AOlohKJsoygUBTopDKHw+khJKMOxqf
vw45b8STrN7WmTfzdAPncNCKw0lm7oWjAT8YxF5weq6S/FfnHHJ5SThIDsME16Tp
5XSyyn7DMbmMw/KB4YMgP9uDLWDLacMtst/JNhuBB8+zemMJg+NWXgtY6Z1ERkw0
d+7daaokO/HSb0q8ydUpWQwsMVP9LNNz42iBf83vDzchJbkIAou9coWz4N0ZXB3X
3Ku6TrCIQ9xNOqQnL7T1Oi8ZLmzhYpMDEooE/IsGjjbKITXUwjlB+YyCvJ/+8MYk
PJkZM22fie0hULtoAjeodxTse5Jc4BTUsj7gPKkACL/9m75I5XafeAFi/EXVY9H9
hRA/a8rQ4nhXHxavmmE8i+mtH/MSpBjC59EXW6aZN5iEViLHqq2fA2bj574Rl+4r
x15l7tsPNlND++rI/S+3AoOPFhGz3kH3QLlDfDBOQsyY+DkjPZlj3EFN0pNsU9px
b1i5oxUuS0xb5u+GRGX6Gv+ER6Rl2mvfjovgh2d3vVTEPidFCs4BESqnQ62QDSfL
6SJPSjXt1z8PyYN25gqb6G/zhq98gjWwk/tBy2PUxY1wNOQ+6zPq62i1xluTiuvA
CKL4hWLU77U6zOD4b94TkXoybmfJ2IzA3lVv26gPhPvoGCnugrdDmki5MuDK0YRd
Sr+FVizTdpksoOAnPSWGsYGbykQhdxlyyBYb37x6Mnlgjp8PkuNSOVgFvN2sAB8g
uko7Ng4sEAYWjvbPIedsDJ0w1BAeIdYOx13CBe9PNB11x9vo2a50X+KwhUpxZ/Mb
AfKlEjg3didjFErE3e53H6m0NfGKl8mqqrZod6m069LmEXx/sPq0mXZNaZmr9Ac/
ak4ziPStZWlHSfaFHk23ZHTfUwlB+3qiSA5pLfiUp6IKauvkNvKNL8DAkz8mKaWN
Bh0PffmD4MXgsXFZG6k22/K1tC/zA6lINdB/vqca5z4nwIvf2zGc/3C46au5nEqE
sxUcg4w55N7/ST5yKpV3KjQi3sYYORmFL4iWNj99N3Jvery3O6oY9OHH0kyPKN17
wYkzaZRPq3vRvaA5hcpdCNdfmmqt5F1KjEGc+LMPmiAclydNZ8DrDP3LJHX7cZPl
KgByzw74RWf8hrpU71ss19/wgs8lkeWN4W8ZJzBZ21/B0eWMOK/rsIbeMuAT/KTM
beMqhwPJ7NQShAzCZqS9a5o4izvKUtes3EVCKE1PQHoHZmVhFtHl6GKHvw6ShsO1
tVpVboB9gT0nubJKxSj9zodA/2C4AlVAakqMOLkx7neTsIhEscTswWeZsF+tnDDl
hnCMLFjRzKqjdhrVPS3NSd8dXDpqwERhWjadjjezeLfb4x0+yt4ppBD7P/AW9Tvt
azN5Tx3E479HIvNb/ce0T1zEEMF6/0JlqJ8gFE+jmt8Pi8FTWo0XJ1ZSsFwg6T/H
O5mwwFfTMF9N9uYwPKUiwDFvRA0/q5+UUiGvvxxEhfcRdCYmscUAu/sQ1jY1zfvI
xHy/gKPj6K83Yfz5b0Q0lHnyas0lp4sD3L+FFD6j1vbGoV1goyyotSVIGZ+1DsI+
4EuWu0wkRYjh74LC9/IDbkMGexQUMpYsA38drbEcXq/FySOiy4pg10YWn3Rkrry0
v/gwsxzP4yydeTGm0d14kgrfS2P4z7MCld2jGNA9ty2Wy+LbBA/pyioalOLwG1WL
pDvabP+1+hCCs2XufoJGrWRwi8K9sudCY/3bvXGgjXiAuhhV5oTMO30AeBjoYOX4
YPbexJ+0VLsnYj6OEwow8ptB2gyeraBKItACnuEXqPmDb611pR12DMMgC/lc9dDr
Q8rvWIRro3kUYrRkfkm70uj5oBmBZ3guOvrQ6piRpV582FYuc1HQ5QvcX9fV2s7g
wjO7wWZZYNiPexYo8sC8NwBapTLY+MN7kxG4UtWFT5PwRczfJFpoikluR19ojlat
rvrbnEULwa7h/+oY08G/ZQW4qPW/umsAyAcB0q2f5ecCIDrOTtu6+rrqixSZE/qS
eyemDWIq1RXBoSfnt1V1mRdS+4vuQY+82jRj1P3ZVGELbttmyK5gxzV2+wB43HSR
5AwTEf+XnRFtXTRwBbczvq9t6ZZkKnzIFfG0oyjr89eFgqHDUypPqlE3RvXPhf1d
b5Wa9Z1kCT4g8+FcJYMsMuzlqeYX599UkN7Mlq07evN0dNLiWSP80bnhwwWcQKLQ
SrYekOI/xPaUZylaEuB+ix6tHqaTI1EAb9mN+sSel7brg/91Ks3wCeLoCHTWigr5
9my2mYxNrueSaX/iA5zusokNj39kjAIczEiIQNqEP0LaQAv79Y5IA7LjcRYHEidw
CrGsdFapSXjERUS1Wi8oV9bQL19WNpiabcvh6cQnUPIazDkvdBlbhZwcpqYtrDJJ
BORvWo8CDWNQHnZ+boWX2A3vDlDjcVf6hBVEbAhwXSpa6zmEvj1+Aw28tAhku3EQ
NnyQpwLsqd/J2a4Bb7gC8vplrdOgkuW2F5+XHsytONAUxnLgK68NKEFVAYv3pJD3
lmlVlmOtntKSlkJARnM/8Edxn6U2TuBI4dcxKOVwGmU/xXYz3WZXHVhyUgTOHOUv
CIHluZYfdpAUBzCufXSk6qOTUtsLOuHwyrnMWsex4FX3or8r2CjWnDlbR551bHc9
2nj0oyMJ8kmScZGxnYSE00WCj+cDLYbP4OeCMJRpcwolZzI5vIDAayGnNfG2auNz
A6Mxv9mxTZnhY5hMPjdKyBOvf2GkBHuTatKfj1SIkd7bCXlpz67MAmaFP99ka3uo
S5MFyfD+8Smz7xYfiZZV7REKVPErJw+yi1BDnR8KeFX/XgICQRBo6Kr/0HLUliv4
2r0uru8gu6ec+2Ez0rmqcYb5scgSsd/bEy8IdbgLjN37vg3c7XjfkJECPCTDQBpp
CiSlBonixAPvSQvTYUfr3wyifQlJk4F6NF/v5eRwXa8LJVCRom6+u4g/72jJ6EWV
Apn0B9kJtE4tJIFON3tchxKQH67xMfmbIHRm5RdROHJNGMoep8kz/VKOnxFZCNy8
qEyMp3hXFsdAyDwvSpsf76inghFkeJQq6lpq6hSacqsfR2mV8Ro5Yl3IBBKDQE9m
g5HqbGtkAo/t5V0TwG0WZV0qQiTCYs07msdK2Czws9R6rReNZxCJrFyFmu549L11
hx2qvTmZWtTM4JeC9U8CLAtCtZ2yqocM0N3OwKcEMxgsI6FoN4NxBgHeV/t+18PH
3W4sBX5HFaMDlRGJL4pyNv9lnTlnkaT6pfgCv81/WAm5OCJuvMXzmHyUwBDPHY86
Nqt4KIH7gjnieqfl4epk9HQK7HFuavSm9+qk7HeLGIqR7hx+J6yghi/clj+nsP8m
D+V0Udn+h9lRCI9OKo+VlOOu/v8Y6Xe6d/plsEZormsS16H2fXGzpmMovCHj2JTL
A9XkX0y9ZiUewRHuMszoQWIDvu0tBgzSYXiTLGKMpUVpe/qNP5nC9AJ40P8MPIGn
ytPVwFwiWpvJEOo92Py5vdtfbMKJcqt7d1ySmgTKKhMUzSqoREkSG8XSzzAZj80q
pqTSXmIx9rUHJzY6V8eZU6FcIvi0N6bCBwd7wGeEv7t3r5Inre+DnIvDsSuweB1O
/7pRrYEjjvNcPRu5WAsaS7Jdw6ieLe6bmIn5T5Yv2ZuN/my5W5V3eGLnwGYeR/Z0
OAwhzDOAhVlpDXL/q9Lczp+nEfVMjnhF9bNKYGsqdut8H2U9rpdxBfpiw7WJNq87
HdPAWa8DOhG/HRnQU8QiNSDOl/AfvrKWJ8lHMK07WdgrDh3K0XgLcPp6HL/CMt6y
hIFr3nb6bhMctN293bFWstxQfTOCmvlYlCnzOtcyx++FA82xAAiJxNsnNQGDcX4s
qDQbYIRx0IUbmkJreatjXR2SFFPMFPKp8+0L9cVPvuISAkavWXxUDPXo03XCtL0L
Uu1fgtP7wI4JvTgklm9AS4L5eRXJT3JhNB0qo3mUtTbauZRMlYRN2dgKz1hmNY+2
DPnbcMZFRt7sk/zMZmD9KHXROqzQprZYc+zejHSvYvdIYUyak1ER+gN4GDCgwkjj
px0PoQN1HeQKNVyEkbt5Jfc+Pa1eMFWeqKKTeYVw/sbeOMeaB5rWry3LFqK5FUnd
9wUv3Z7d7aFPe2WVuyW/UE8VgxHfjEY+IOdkmgIefShM8Ir6M1pocEm53KDxjksW
Kcc89WzP55KPEBwB8QN2BFikS7sswAG8OtprESPjw5XMuZYBpuplRJ5Pny/OZexZ
9mpp3fpZ/uZP4W/AvjfJGlGPY08uelWs3Lmi9jmRbcH7Ih1H2sUp+InaeyG7Yu+h
hQc8dO4G+xohWowXmaOuIoVsGzOGGuj6lNrJyJKG4LQSA5a8sQqkS4AINnv39ZWF
iCvQ4cJ6tkMe/FjgKR2lKHImfzK0K1jizYvBpkbA5CCkrDfzS8vCfpoP6CxIXsz9
3HbQ2NpnTZ292eOGgDgaYh10NbGEp01RYDkM2j8IT7r8fbhjwCDH7BbMvl2QiFOf
FtoQx6ij+QmsTgy3+397K1WLY9DrgpOAuiaQkq+uh3Q1Lug9tlI4vIICvvmrAimE
DrZ4gtTybOPWTIMK0RO7BYm6li70B3luriYB2HpTlH2Lg3lgbT6tTS2UwCljNmXg
EaCNUXmJs7a5d8LOUPbBLZFEzfbn1T57op8eFMNpFZDWpsRJl3g+tM55qUfmE0vm
PyaJyEKnn7ERxtsjtghpUcR2XMJ0T5MkM/b6u7kwOKY9P35zr9gaNFwRc4oCXBET
lYfQhT+sdOZq3SuHlG9cOQzCy5+BTIDPRjqhDVpp7WGC4ljdK5oOjgqUb8eYkiX1
QeQW5kJW9buCiE1L6mt0E0XZ6RBtTcc6Q4RwRYCQ3t5w+7wFiZG800D7dpo5klEi
YE4gPipufmY495QA24MkMh0YJOvPvnb0Kt+yu/7Ts1IiIhzDjk1sI65Pj903suXd
U5Pr6YMe9m3UDBgpTstTm5i5B6Z6fwTGnXwPv+gXYqg9OjRruED1L4Kzc25pRnIg
bykcSLe+m7Z+JXMH26NrY+9zLrxIM3Rmx4D9Dzz55dnkLfEJlpMnAGJklM+RxrEV
fp96VwRCOZeeD/3xQgw2rcl74WZv9MKOGvAraRCVHApoTWaVIHZy53SzLP5D6riK
pYTUjYn2ahX6XjN50E8oZNMGfEH0kUVChWSyZl9R5tgi93lJ01FXa9Iwwzu8UCHP
LPkk1XtKdLE+byShoNdN3BrvHQztsTxjDDUe1Rd7n6cSLZDF3mXFIRAtoW4Jmrmz
RrUoOIG5dJeOOrWx/OCTrD+dx2qm1+7BsEa1urQvzdxvaQnjg5XUPmzEU+mkuzsa
SK4zIn2qrP4XjrPrkpgYuHWN/8uXyd+9IfPyBDe7AY5rY3ucNbYZidES2lqRBXNE
OBhTZ6faWzoh11sfN/DnFYGobCvxxdP3RdcdIBio+IjE6PkRmJeKAR28AVU6i+SE
fxlx20B2VhBL62qqpnpjvZnvKxJQXJMyRVPFY63z0ktU/jwt3p92TXzJGLFFjkNz
4lN8dM1xI0eC7N9EimmFYCjBRG6T5CTtup9fcSqXdKbXlsqokSQNdiPwwo10OKHX
5Vu6d1MP1MhgvkUySHBOuWKZU3ZHvfhCClJGQI3UKStiHPEVuOKoFtfT/HQ3o5Jw
PrV4ibhmwCMWUN3zB4GsbqMcoJ6dey+1uN/nwUL/a3mVXlp4CXFwzARa05728WNz
Ut0JDoio2+zeeEMohigf04aI3nbFxgdzdAvspkibSzq4l2tDmXPBcA097Jap1S4D
udnzg3SN54pBwM4n3VuuefdS/hKd5xnXCqQxBnLJ5mlDZ5H3kpMdq6nQwL4nuRF9
Pyyu1RucakD8oxjGuaF15qPKwb5lTqqGU7Xh2BHlRYtYYONwmV+nU4ecUYkmXlQO
9QiJF52eCRjgvjATalMrgnWdUBky+Y0Sm+RwYt2meS+BY5oFC58FrMkvQ7CDXR8v
EhYZZyokgq3EwRPxHfgHgbs/I7K9Nfs04xc9dmrYRharyHLnTkG6PbZfdOhICBNP
WY4y6JJHkD97AxxmEzBcYvXqGHVbM4wtCKDmb2ePepmw2X2KuiY2CBHU4s9lUOO1
kElwa3oGOjSPTQtz6QH+LlvyBLOflt01yiBEjXQOv6Us13/+IJv0/NorxXZBiAzq
KYT8XVx+3HEEsP6Zu/97Mz3GgdlyDTRHYqtkTm+B+ctRrTqkMywtTzHLQZMQZiJt
oKXk+/RCWb5KRpEOwRpK1jiCAvgyHDsqUAPGYAicj5zpVNnXXbGXhcIB47894Xjr
9e34Cfr2jiugFMmeRbZ3yVTqT9G8ZD4Z4V72fHZvhHDi/4bsjliLn2xUtKulKhMW
aIC6KJgQaHCTJBD3+EEWa6NnvU0huP4JZZKt2zmAxvhMrx1O2duB4hJDCrP5daCx
XUmWVKT9ZMeP6fTRJu+oc6exNG60Hy6Qzs8/EVAz9hXRpTKwjzIHSnKMFu88GxNH
5iwhPr2YlApKQiVtSDQe/twX9JmX7Y4YiZPKBWEJbY5IZbKl3DgbyBX4EtI4ZhVl
D2tWNK+khQW/iovUN0bUjUSG6Mm85ICS07sji9uTyqZ37iW7h2POA/HmH3T3LefK
i0GSA4eD246bp8XmAVTtZu5rA9rfbAjOBZInlNaca0zm+E12WqXOgYDDCxthzFIA
O1r4SRWQn0kyLzOo+wOcrbFjTQrbEks2fjPvcKqBO9b2ZA0riRTdkIAqb1JU0tbs
fAVB6XzipQIb+rdVQ9+FRS4d/yWTE6uKCqt82Qa7jyC5MfsSi2COX+9+cF5Wrl6m
H3yc1nzU3ckd5Edj9dQMdHnl6ueWcC1gfwJf32Hq5yWipneT+nfousQvHXjFfnGP
5gAiw162anZu/KYcFEAMTro/V6neOSlK04kC3CZ0P37OH0Pof5dJKUyGNL1LTWFC
PPXw/S32jdE+p66NA1TP+Y/Xp1u1ChTTDSCergN9qWRFGpCA2lXK2tbuU54cUwPx
hReCj6VDq7/GFqWiqFeOaYjKdCfKn+tmbEWWHH5I3v5mxo8xjJ0uy5bbbs3WkiIK
jjJ38Thhqn/YMKNrgtAoSL9mMh4FMFyHBhq5jXn8nl0rwZBZIpD/YifIa7QLGar6
th7+CMOen0TKWV2hbP1ZjDbOPdSEmqe2zslcvYNH2FsdCWA9jKhKh+3dMDCc06Cc
iUDFR+VP78tmcsgzUs4sGiXWs7y0U0ynURWujFE9a5jI4bDM0kiLkQoAqYn8DwIx
nkfsCrAUY6hSmr6uPqrdP8ZN0aS7N8mRZNeNdn+5wSi1JAbUA4EL3332aZ1ZgVqK
ugkYfkHDFfhFkTDr7TV/OVUQnJyqtktCk7JRD+izJuE9tbjxtsu5r8HYTRN3Gv6J
KCZIh+rWuF1xa2JNrWkfw9+QAlJlwoXIORM7RHkZ2oaObFcv3+Xh9pP6mG8bTfoa
ps+xhfgmymbMgwh53OiGz2FjvTcFcCxoizhi+hAIGQt3YC53BoXtFi6HnNt+SMxF
jisL5Aceocqd/A+rag4A5PhSQtISEBbi/fKDzO7AcFLuNwtmo2Bmnz+W1CYt13Qq
aLqeK4cl9Fkb340ITqkIOidQGQ3jgEu12NcwOppiYXnO2usfUqd/9OsnHNeM/wCH
uoHBIpznd+uS3EJa1OBri7poZIS4nZa+zGQQsUvm4ZF+7BPHUe6YnSoJsmO3aiqe
0uylKMvQl4uspo+69elSOOV2U1d9TScNT/z6jNMc5YmQmgNTv72yG3NPhkCN0ZWU
Ohrurp7G3WMuOV6/HmYsDj4HXJxcfbf9P1bM6ncKPsb7ju9PTc6SXVzlGThkux+N
3Z9ecZovrEPTeQDhF7hW9d5NeK8Z0JOJKgSMc1gTZH2qhu/PaluFK5XZ/JwAp+jQ
/Ygtfvq7pRhM1t0b4mJhNCuvqESs5tBtBrX/tJNxSoULhEd2yRAKSF7sq8I2Xr6p
NBzwsE845pk6KxPhVqy+EnPiBvNNo14FPq07RXRvFqas2y3Bdvc3JY8+BD396JH9
pJK93kPN846H3PCx53F6WBo9wTX8KZcQ/XY85np8msxxJyC37jYAVOWnMtkcx9xp
TZbl7beDCVT8FXH/Q+PI/2d6Yt41VV3IUx1y5a9D+Z/SXova7kXAZPvCqgzC/Pya
J200TQO1fHmj4hCYRYqpGPWErEzPEC/Tz1Qnuu3jkU4Rp3MCtSGGh46KgUF2udyL
ZswtQ93DgML8voPKAamZxa2UAIAovbM6EexPllPhUDh7LeCXVcFtRhYoYxzn/B+C
8RPpkmQMHuPIReg0xiutDwprLHWJp37vp4ybZQ6DH91AgX2TcEz3ebv41XdhpBrI
U9DFXBQ+WYkaq0zib6+iF8VCFEsroqdJ5zJIxVRRUWBtNNcrvDarL0aWsI41Lh9o
Sh9D50g6ws00kqtk0Boc9z15A+o9Fpvvqnk2aYp9hDAG2oyZMbRvS/kQeS2+xbZY
UcsgdMha+g8opMyeA6XbjtrPHhySVWpfgmjW5d7N3d1QnNBD+MtYHD+MY/RkVzQO
5kO2Sg5x/u5OzaLX3QiVSndUJmhhtFmNndqn7V9s8ck25HIc7m1qIgkirSnOj4rS
dLyCys+e8qPLXbL/TZTeX9nBa3WINFvqOBofdRnq65w4FlwwI5yC6VZcR6Y3cCnx
5nNYMssVT958RIRRxhIbH9Qr52tYWjqQFf5Xt99zlqScihB5I9licKGFTDKgpaWA
KDBZwGQ2QnqZVESSEOqOBcYhDa4ik5EQQFRhQoZwQbjoFgQh79zKyW+ZjAyutyKj
yZoGNqlrMCpgsFdeqI7sS504eJ8PPqI4H5i9Gk4HCajYOBvP2RgCwKGOV95IgbdZ
nRrONdGDVetKO8bsNu8l5lD+azAvQEkB3T+bNc4CbpF7NcrT9dh0hKLa/uUGZdg9
ILJx+jqkox+AaVC/rfPJY3qp38JFgB54I+Q99gM6kYjrIVD9sZ6Eu6eVxLv6n/h6
gMzPpyvmwHuFx/NoWHqkpIIjTJpE/YAL/tOQ4BlaAwBqttSlIcIHeKKMj3p0saUg
E0oc4cxxD4pqEOALSlrNLULmd6HLdnO31K/XSQRDi6jcB6WC97vMteFC6h0zWr0R
bahFHVwOEX8U6FEeqx52JZLaqVF9CgD2FR3uHDRQV+4tvDSkZckBm5xYD7YouPs3
OLr00OAR7VrTTkPVhqDhiDjPU6CyFhIo4bV5RLuX2SDsTq5spDVSa3aMEb456lsf
urhVu5LlgyDFgV+pW9xlUOpmRS2e+6as5L1gzNNXV9rPBh0oy8Ct0bJVtpdcsNAc
FREIBI31g1nIENN5ehiMZehcwsEJcPwu6xquzzhXnTGEyNy6GoLeK7Y7Oitj4ety
Cccn+v3z6nsU8r3RaRqyuVIYuRLavFB2h6GlSsJIeV5YkC5qTdToJP0OPo7T+WH6
wEtDLt9gQ04gzBpWa5ep+ZHUCnmNxieDN+iW5KDuBgeaZLDyz25Rc91d3oEvXI37
JYZSE6ucDeH5Y5CdN+XQnygtDlVVJrTLO0W+8sk6pzrD+nqfn6FBvhK4HrL4yajU
8hRfwWnSeHzWaVrn9VhJXhStbeXMj79q7rbk0gGZZ9gRkeWFv2xjwzXew7lxaI5m
rPiUdiVAMoPspxW6DaENn1/WZWiovwFlaADA9j2bmGQPQGjJsh8MRVfDTGHNfPl0
ARNgsKMglx6+1NsGRrhFg5Mdk8fZtTlwJMSR+WCTxEtElOwBBnSYJILh5+hj63Pz
fQTJvXGrjE3CmL7qAYH60mOvrfdB/h8Jy3cuhsCdMub+G9yqZfKBBvLVTWtJXngE
pY96UcmK2BmBB7RtbwmwFHlmdq9ln1+Nt2Xhl3jRjbSgbxf5sdoB4k8bt3ZmbC65
Cf+3vnsFBolgEsq+YnGiEnrSUFfESZmRO72om/wAT88hKwvkktmToDORhfkH3/ph
z2e9WKM82MJfNh80EicIiCpbp1metlJotgiOBik6W6tjmvd6Ns9UgSgvmiZ38LNA
KMerXOxSycZvMHhgErBLmY9mNtUKZMoafw0p3MtuS2kvSW8oXYxXn7UFwOtV9FC+
FGPpbW0bo6NbBsMyzt3XBZ7fTYLSYXZd6uEqGjRiNx/iUIRtFCxNI7aSdcCXjsLm
h67TI3lL1MzQn7fg5FhnCxmapYeB6sfDn1UDU+ky3dLpxuJhHzqWVt2gYqKd55oI
X9yN52D3qwmTFPGsj7H0Mepro6YSEIEiBqR0U6XEcEtaOWEoj8naNy1Jhwi7tNj9
3MtLh/Td63/HsGDWVvCnyQieiP2fcfIjYEDjbU77qccAcB0tpoBl1fmrINPCqa1f
E2H8uhq1A18/dp1DBCltlAXDq4m9+RKA2BoU1N38fj2yLSHa0n0H6XVs3zzNHxPr
MgxIZbMAR/yEMS49hk83q/KUOOJ2rpGiNEUrCq6/bskY1IIo4UDvxuf2zW0C5yGe
9OtZmXfy880gt0ekIH9uG3F4ouiqku70L3CWTAp7ipxtOuEV7jnl/+gumn+V9ZJy
Ik+Oh5sZD/UBCBNjQy1AugDMhPFVLrUvjC/jGp0g6vAbVg1NDe+hOysAyvsu8zl8
tSiDaaFV6TZhxVeGI2uFyxBGvUnIK7S/dMwyXaUuBc5M/ruuNCA9pwrjjtPBpggB
CofkD5ubgX9mvhBK/wv5hgfaR/w9NjV+bBugwCeFzW6Hp87S7/fsn47aA1mo+Z+t
5TIDDr78hPOuJ/AZ9S9BDtt9KtLQVWyKqD+jqJ/CE/XwpQCNkndysP8+CDNb8fnp
ste9DseSI/GsKpc1xNh8KLoRbyUigktO/nlOvL10mSn30KqrwqLk9NIKHQRPL0Fq
O9YeyCdSKlY5zvffmc/N1MuxpWd6x5Dtty9B28RCWxNjiQfOm/pz5VGZ2ESC66zQ
cUAXOF3KZqjIQy3fe31YjyJvdaoyS8sWd812gELS9mPnKxH9iM7eoCMTzk3j6lDV
Z7+E4dKnBJ7uWJx1JJ/sO1ygyBbf/v+95Lcy5l7we3h8CVvJRCTsNusRRSNRrM/m
jJsUW1vNxEMszIZjqFtP4dl6bU1rqjvLPZjexKXmk0CHFNeZr1RW2/zJBYZd4L+g
jf0NhM92a8t1Xdu6ORZ6izUoFi1GNaVZUXqOHpKJEy+ul6lbWJiUFf8SNERD7nSZ
+Fe+BxRnSz+W4aaawpsdrqIckCINnY3REh11W98akIrzMxVahxAgNk6CA0IpIWXW
6+CrrfzRyyzKsqK7Jr9BkWHUqibH6594SeUx32vT67z2rbjnbacFQEZuUpluIFle
CImAoxsxTWxjkvOKmD2wGB6xTNbiaQDCwaWYbpXZJPUp31Q92TGcKAkzoFd43m5y
JN6as0/UzW8KL/6ewBrTbxIOtJu33A4fBNZGScqlIV14fwnTUbjzqpGrYZ1ie8eT
8df8yrXKkPoWwFX+7+PmHQlitoUdkvOz/nmSNJQ7Uh6M1BwBsur6EkSmsarp0aGv
3B4/MerqhHd8fESYbsbgIb7/AYInmCvCMc0rOYjpFs4TkcwvndKdxJzs886z+Bwz
bP0j6TOaOFUU8Q2jFoHMoIqYpeA0wtepbJASgDgdzJbF108lPevzLb636tOaOhUr
/2jSzEQkMyu+3cr8p7lGRKqq9qD1PpO0IOwpl+rdo2UmRAlFKusw1jFeHbiZoqyV
7aFSWPMHjfQ/4f59VEWZmIqpoG9j6klwBvSohUUryyCWLSFfmTOTHmqnJkhQW7KC
Cw9/ggjpGITbDfnQll4xxM2iJ5E0zzbDz/d3lN326klR6NPGLZEHNA6JXC9i7YhP
z/JeEfZBbqBUnh6WQN3D9K0RMLlFjVPqXOaflHD9IviRK0vLm0qh4L4B/E46vB+Z
3xC6mn1aaMa2h5XwoDi5uqU3Re41eA9wt3xYBPjwyfrIUHcGXvfQoMH3xtz8BqEl
nz41oJZAxDlDWsp3hftIBiaefivARAmLCSsmfKUg+nP/BhtQrJVWEhdOUSIkHhTe
7GYTMO8dq7AAjbrzZYjVaeq0d1loVD6YcrbRID2ZUkiSFRKRawBSQO9rl5ho7FzU
jsJbCLdy9mG+W/Zt3143tLMvwwMO3nY8N7IKlWUFA8aIXspEN8VGLv4zoHe+KVns
stp39e25a/h5YTIpDzH0pW4+gwQKGeKkzOdL8cYBzeH1v6UVDY4wP7PAUL0ttkPn
ueNWd5gZKvM2HsiC60KyrgqdILYVlZOnFc+Wb7psklZQQQY72ZKYPKzLNCYFz+2V
BffeIQn/AY0S+ekf08kKxZQCTlbkQQ93Ujb1/soKM+CPnFkjUWIgeVeUXJPStTip
hH6QAAzVXDsFiCUb9SJUfXZgCuaWjMOXzmK7dZ0UzL6xVD8B7UVlX19mWgHDtUn+
Q5IbkRRc35CTbRdvlaCvr2nlqFF7CvM6rafoCpqtaIJGrL3ZSVMhcK8f2WDozJ7P
fYF8tHN7NqxQaj9LnvxM/HY8sHix2au0oldDZFi7FmA8gt7egVO9dn+aiaIbpR+0
fJ+GcimKX4P954mQM6ZrlVEwanVjkNJZtU4Z4UALeqkFAOjIEeSN38s1CBe7YRkd
MIJO2dRZ1JXlmch8ig8r2lLf2+GxiV6jzjFN6wAar6sSqx5lhNGTo+Yy5a+ucctn
qOJM7Lt2ygVl6Ij1xIF6tc40+iH9jmsDYVcIrgx0naOh9/aW4oR146WCFHFng7L5
gLO+sWcNCifx/tYdlwTLc8rrpm8btzdBUtqzax6VZv0laXwLmiMGaHUCI0FFxV/r
vcOfAXGz+7LXXuocFrShf1QVghpLTiy49X0ATFhY6DOl/ShnoIoMQPZmtk4ygbRf
a1x4+eFTR9Ih6qOh0NgMKgYXSGc8s4eL/uu1YvXsImhf20gPqRsng1UMVIiFKwTk
+0LfvPzwjFhWBWb1UTsbwLvt79WbqNdWNZxGDeGZWyMmWzI6U/ihgLiCx2vmeucy
+/93ACr9DiwfYwVNAbWSIOYy7ZdJU+8Wtq9w+58lsDnZ1oZQ4VbqbbNe9USqeD+D
HLL08grMqgYFSIU3DEw8N63i3hy3mVVZFYzzbZyY9ybTXKq9ak4E8pLPCEz0Z9oL
+CeW/DlyKKlyYsbX4lQxF/mxk3TwizuBwDb1Y8CwQVcIlFMhrVHpmkP8ED5mRbFG
x+y9bjT675wYxcEqVC97mK/z/RrUmcHPI9r1RWP8gI6FKJy7PDTNOkRL1V9nK25H
tyNsziTmOCQQ3RAmfJ8+4GLHcjIflNMxVYszNBEVCNwklGLeQVlSoNYm4ZvpFOp/
gNhQuzoJ+POeicEANGTNt/rm/uOQI4r5votDrpU16Ur7YOqf0dQxYzefqlr7HoG+
WsKQjojO19P5RDvYJmrUWlNkVn73nrcA7LgN7F9a18xlly8K+4ay6BF5CQ55btsK
eYuGuol1h04PyXgarXhI97RTDN0hB/alQeXAH4r8Q4PMrPE3g67Wu2aqoWY5B9Ch
+lo6xgAvP/ndN0R7ZKytJDAU3xJKFoR8e4k45kv1lBKlHVxIzTTK0BQRuLTywzj1
H+cab2vFK4nlkWRdVj9cggxI44y3EAf5nF18FOJH1zUbntWY0aHYP6ZGoSOgM9PR
UhwJgW+VYeXq7kVzhLZQn9nwtSBYb1KgRrXjtpleapfHzmGmyWj7av2Ahkt4gtcU
9RGFGiu1MnIs3bQT/BC1+qTzkqC9CC1N1cYWfgMG8XVVdxhNR+EToEMUs6dvDfYK
TZlY03SutyfRStqP4KvFp1WH1sFdnz2qdhIliPZiYJVlvUGhr3qRQ0mPWxpzuipl
/Z9etdc7Pj5cx3AAxsEFrnGJBY/+3eit4xiOpkCfsOplDVc4KuWJfY7C7f/JxOkf
jpgptjMFIUeKBMgFLoMSy7NWNK//Md5l1sQITrbNQH9+NKZP/MepCO1ZrrQx8jnZ
5tE+E1FKYM1+jS9p1WkIXZl/ZAW3wbtbAL4qRbErP/voQH1s7mGQh1ZSbKhxnCRc
eRTyEiVf4NBs5TZmGugobJ5FfkkcceZ9fA1Qr/bjzUNWzIibJN9Wb1bZfNxSRSzv
Ydr8cr0JnQ8cDCsXI1Llkmfoj5D5WUIj7je+UpQwmaORSCodk9DxSphfNWRZD85F
1S1Hw3x1QSAAYleXhz/wx1ZBKpzXLkKYi3U02BFlSvfT1m0BjfbVZftoq1uLC5st
EiOQjW7s3vHhfHD9jrcZ6uf792BY/4NGXuPo5dVnM1nFG4TjQzH4dd+IuoKsSX+d
f9i2gUKobZcT8PxuUhlpYmRD2NnVzrILwtWaO/Gxw+royNsTnvdRJvx7zXvJXL4H
UD98uTYA3uolTj6qjHdfUvURzEaNIYwut6vYPJjRK6E9j8c3wnVntsnN0wFx6BhV
O3/TLd5UrUmqZdRGYVffDZGX1R4r1dzP6lzARXt56pzvlUZxlpW8eMJXjf8MuX4+
iMfgsAnvu08WyewURpuxpbnUKHt/JWWIugVuclfsPkSKfArutLUsoI5d1y8KJTv9
KBtJ7YBeLSYAzARCxbj90CSJuiH+0ZEiaFXoR0jKEw3uyQbs15hh+b18QDJVy7uO
Rd7uihLL0IEPKtXbeBIRnY+y3YdqrDdkw0pFnpDzmawk+g6BSvq6sIxBozglXaC+
DUFfF5m+RXxB4w17uF9s1czoFIr9ECWax7jvL/AukM1z1B7s5pA7J3Hg024vDIhv
S1xH8SU4a7GDAwNmt7g6RL4dhwRq5Rjgtrt03RX8aghIwvKZr9M42M3q/XH4psw5
VPJwgngApux3qBZJz0zL6kp6fgcqdLFMfY0xCTg9t3ZE23Lm7VCHjE5N3h3buzFc
tVp/3tN5PH2e4SWT94TaXKLc93tJkK0U8qMGAZzpwufQU9hgVNDujEXEHsk3lIrU
o+tvw6dvMUl2nJKb5zWeCJifnoQzdOS49NSpltdnakMlYZP0azFsoTqUst+KMZUB
mn1I8CEZzytes8Jhc/FBD0dGvocFg3Tb11H7a9kuBzac1EcClx0yj/4SyD7YE0B5
uKkCPhzUYJBmUlbZbt6ry8Getp0t3xKN7rF5Zp5kF9r34Fg2fcbvtBja2n/TZ2zs
h2zEQLa4+1gTYZLcEVs3mZMHVgyAv1KRn8SpwYGf//Ep5qKBMpAmuKVu6C+smx4h
3dS+5RZsLrXQcp/vePLEBy+aTuSFbxTqS2aQMxNT3NCYQYyvnmNOG7ZaBg46qmKv
5Hxz0+TwMyckXCm/WZArAQrHkIHuS8ybInN9TnejeEFq5gwi8zjAcI8l/ROzDLsV
G5cLrtcTxY8o5kKCbLudWu2757MPNef1qToqRz2WF5wxQDbn0pl6BC3SXjHw9NJx
tyHrKCrKa5DcxYHLrzEFg5YXKV2taPp/SDG0alK0ty/549dhBrdKqDwFTjPLWCiV
RaQSWojKdFwMaNB/xBnV9giJE5Vsc9W8tIckfArXvt8KrZ+pjqdrvSwD1vvdJefi
CajAeAnaq2ejEiCNX+WnF9wsp6i4UxZj5WDkJIV7ESTTT+g6z8Zfx/IDCXG01PU2
jiWu9vaf9xhjCAS2mpfmg1pFbfM5rk9AzmJU589h7HI7MqlTMvlgycHGagQ0DpXP
hMhwEhTWNDH1BAcpQzefIG7ZLLSRdtxZV+EemYV6gjE1pACjHkw01DEaqao/pg+Z
8xvSW0HklAh0jm0Ip1d0jXEVVMD/4cyFwWgTS3gyHTkDQAiOl0b+ggxWj/5KbAyo
V85nxXF/lO4zFegys19Vn/iIf1gGU6pPgndW2pwEGfhXZX5aeM/mvGckAA92zk/S
g4piRZJTYkFEsMX5g314m1nhZawRnW+i5vtMSYEsiuThDIUN72sAtLGrrMKoME4X
GXxaqk/U3luSid46ptS3M6vy+DhCM70xkPj9NfWRPdGRGFRVTBQxVJdPsphOEY0t
SF8JpV1l2zZzkJMQGEUrP1E6nJtR8YuqsLuiFLqcQiRlDQ37eexxJY+TXINzvGoH
cwFEFISV+94S87oJTj5FuXNHCqhMB6tBESPfvkB25TyxOIGV15Vprs/Rf8+P2/tw
Ky7Uei+4BkkG+iGzhN9aEetoHDD0wCrCuK19Vaf+ozYZYfKXiazIFpK/u0h3kdF0
5qE6TtLigYSgnW12AmvYuu3f61ytbRxhsTRHw+UKYFLvHbvwf69aDct7tm9E/Fs2
ovflCms0/U1WBDwbonJjaFv6I6axtYRyHRctjHRJSQR8l5Ubwm6XnnFjmArE0XIb
zgL15UNtsXBV3Ob1xpwrWridZtCLaITfBsjhxYD5H7FFJkG8bVFUOVpXFONRv85i
4HzWAOird20+CCo4TM57VvTxouN52R+XYh69el6t8R4cnudSWTXGFr+i+ax3KNDU
YuWiHyu+pgjUDYNxhcjhk3iIZuE5bCk0Fs6Rvy2tqdE1vrnTCOWUJI0wsoBi/41W
fQLLFWNRydg+xLU5+/OVEdKaXfWI6X/bOjPCH31J15U2dkPeZ5HPFfaOGVaffSKv
uvtRHwoUVOQdxx7Fn/QaUQuu5ijy05JYhRy833czKT5oXrGJHrOi1RuRgPrYpgvS
/d0c98xpqy4Uvm07FX5f8gxzkE48AavXPrBoxG9uhMtmgTqgMwldHOyJXqozZ59K
UScatHXXpX6sYVDBsuZc0fs0fBpZLgaMw9iNGQB0SJzoAC0vEe1+DzpAvjlK4d0O
5F1QV20mLexK8U2QqPA6HaYL5mGs+L7tPiI8XAygD8VyQspZETDofisRunc71JEf
PPByg6C4QhL3/lGAupCg8GG1xmvTBId4bpTsjMdl7g8Wh+/1kk28e44/V0ucNVCC
SGdCz90X9c6/u+ZMvmVwqb/5tDL+sIJHfNqMknDaEf5sOmDJPmG6XgwLjKLD+08F
tJPR8fGPDWV8VSi/lsrWLoMeuS/3CESut3gMV7H66RykCN0KyAOwRUrvOgwDK7AM
LGe4WnTztqsIxWxe21IpBqJ6UX0ytnqQ3m4fFiIaYw6TDqUYFGjfnnya3fRGrKp9
HgdDdgsRKSuTBYq+hp8o5PzQWH9tf38jlNBV/P+e+UNLNuwU+ZSmzkQiEAActRNW
IBV++2VxY2nrD1J8SzUh6K6YxNL+ejNy8EN1peRTab6kb3PzmGInmqNix3ZC3xub
DOpF289/VlxVhnGbF+hlNX44DGfFlsOHvhEcepjynZ0p2n3Z39R1Aj8wKZknFiQk
pzlKtPNGmplSFCFfqvqXlxYPa+MJpNjisQFUtyFPl3FkU3gTSGnec/bWPaK0Ewc+
0LuX0+CyK+YulBq7MGyRkH+TB4p2A6x4Q0jc+9GGY4lAReBfvs+Yl84gQDz8PD+8
1GwQiY+3nHw5YkE3zjKhJhJBMw+YR1uN+P1bjmnDvNBqCLzZ3ePV60R3Ln9MmyIN
suMf5YsmLgBYa9denpheZ+2EP4pZYj5/MbO4yTrFElZxIskEvvEcDbLSxE77xmXF
mW1hLr6IvS3NN+JMlPKPLs99SIMdyEmYkomaY2cHE3hpdOK9gWEtYuY/kXY0Tlvs
5wW4XISjq83GCrdo1PIz73glb5do2PqLUpLxwrR/pShQ2XHs2Bipg5n6eu+TvwcS
21rVuJAiuXQltvDYCiGNfpHLo2/1yZMMK+HVqSNF1W2x4ML4jsVhy+f+p8L1iHnw
DnbETqpsKQLtPXQnk5zSUx4dHjdKhOEG3SNSoaDb9bcuLbEys8JWHut8rrMHd4vc
StD4sx4RUBLxyGw1Xgd1UGxgK6mKgz2OjXrnMxZDx7MeBg3hyCKroKxqaefkMT3R
1VMr8Ndp5Lsif+10c+H+cvAVNJ8QPNd3mctYazg188gGOEt8k41Qx/o1LYzBahZu
EDO4ou2ZfZho+zWF6Ea3+u84tzhG8dN9KJRAwpOsQ8o+DmUJ0cYKaJR1ZV7pNHwV
dy9d54HRjRd26xO14dRyCau3CzRHiVbGdcGPsWTBOxrFgotqNrBI+dWYCAvyfGWj
7NFjrxRJAGWeg6PZFf8orbCwGGamb1m2Ev6/QZQXh9RB5HeSbDw8X0ZxgKq9QOfP
7UYf0II16JSNP2dH8f7ol+E44HjV95grOnJ1WGrUu39rWSX6GjpTGudfsk3XNkzs
jrIECz5Piatvy+IyEUJgUbL84WIFDWMCQ2ZkQiX052txT5rSSidJfz0Mv2bTdQGQ
YioaZoWI0Zunr0aX7daXpbxfntCMSb/Qht/oa7YGTDh0/Zi/CFP87XqHMA2a+NOo
RrRgtpUNY/T68WqE6/F1dOxu0eWikX1klU+tFdPhz7o87thD5GtwB4Q4yhQE+4pp
0k8F4PlS/1MEMtw/U20bS1PLaEZyH8D55oMxtHCuVB3Ia/h4JhejZ0Yic4y0vZFt
NxTSzynOQ1yqNn7/0PdYBp+hOI+1jkJPxhh7eSh3xLwohNtprr2PCa1EhTi+oz6P
86p/zvA0mTT6lC37c9215tXvo1p+172lTL2CRQ5subA5YKo2LGluvJjjMSMdX+VI
Iy/tZqSrr7We/Hz/coKkGP0cMEdnUXl3wOCNlFJ95eLMJrBXueohCGW/AQqHzTaP
pJo2OB+5G9+GAGrkfIghkaob2y8k8v0Px1dHi+omExV56cqzFuRZvxJdg94vRdc6
Vinp2qS6tosy5VKJ+/XSdoEMipDQTyY7tK3fTC9Tg0kyucFMM0NAvDUyPhcbsfFV
ohjdd2QCf893CdV9yn3ILQOfBNPQyy2w/2r5lAa3uoA+m1voaGTLs6nBJ/IF8kTn
39KuQ9YzMX+ujUE/JuaQj6rbd8xh54n5LpwxzjHfg4cbsqnTd3JHYLborhmYY9b8
rsqz9nVrPuD+yhVmilLB0Wi33/0lftNW57y1hBSl4Q33+OJgfongO8FKWXRjuT1g
w8AimmWJMVPucBONM90RTaE43k5yiR26LUCmW+XYY+PxB7WMN/Q6t++VT3BsQZfL
8e99u3kkdAskTttLwR9LJYWWo9dRiRVs6FD+kSZhy3X/GpZ0F6ez8yl8if3DsVqr
nrkeAp93HdY82OBJtW2leqEKowniW3MTW2vnKKW2Qff8lHeTDRwa+rdlMU3rPraJ
rKTd7B9Fa2IkKQOYiDsioef940GYPf8VYpxvHPxa7EMdzy4xOQ5zvcA9JuMcSMLq
41KlDxXLrG8ONQggEdnvjM+M0dpTGtgo1G+6tOeOAaRNPzYWaQgqCK+rBkVFvFxo
fnaJmcC57KmaWFDQpgRciSIaPUVGZjEVBShuCZzH63uoMZX7VIgzFDwtPE0G2mcg
2jsYBvl/ZwMxWiiPKmSyY2snOzpeCvcj+wiEvT2QCIBGSQDHIeY70hhG8CK0Nfg9
jkJP3UnOqcngooFdR0rxcHGkLUa3TQFE33evamniPSzWozvjzm3XW4UZc271pNKh
+GmYtx2UCzGtK/FfzzpkUUG8pAVSVca/UFLL6JXxp3eC8hdcpXv4APNyNDEhGyvp
vPn9Xc7ICGXADhpFNaEXw295VzonJvaeUhhSvlsRnpsYyl9fhVfCOqVWajU4sG5J
UUN1/8DqWuVfAgKMFcfh7SNRF8QNNpNbAqDZB4o8RKEUp85Au5iCMUzSKGm1CmH2
SV/Qnwf4XwGwSnnczFXXko5ob5+XL8ct30h9sWdMMNDes33SiC39l9Blwj0ehNFm
B+wUYvGQHhIIHA4yxyi22kg2xxgwtPM6sEb7yGPG1By7cr4c2iIW7NcLWUG2MupU
ifTxhYRnCOqg/zvAE2g/j20TcRYnMWZY8hCk6xdH890YP6Cnp+agyDwCGvGyJPmL
hTs8ZH7fMA4AknTJEjoQh76uTSd6IPXqVcIzeCyufGMjZa2TYMAQDvm/+loPbFhT
41CQTzq9PljpfgogA4g8K5t7KVCcgEyHrFSsnJm9OuP/XfxzapFg141YhlN/oLrg
wsNzq9sK/8mVGCzT0fAGXug3RGp5qHbIMlbKYXyU+bXQRt+aL5glKjVP1f7pJct1
foycs3cS5zO5i4x6THOkaPURg4Rl27WMxZyHo96gf15PgOARDBS97v3YI9rX2fv+
01NC0Q4TFnLbkBHe03meOKUCUS9kfEcfsp+Pukyu9QGABSTCXIqJtRHICw9GAqM6
YjRgmp0xKUTxCP+/4imkexmyIDMSyqtE+URGDBwlks2EUZ+YsenDe+0JuJmZU0eH
1klq95zsYlOGAi9rcRYl4/5z02Jgu1JlP6Z/glrGdu0Jm9jB4jY+6R1s6plUR780
prVAwxM8ci5yXhCIx4Xi3fWbg1uiUgd7LB++GrpPzqSCzx7S/eJxt94e15bI41wA
fcxUIuVo//oq4gf86IqqIJzBKPATP/zrYjpq1O/mViPuLtoRHQAWBQhphzo9jucu
yy9cYg04PFnZg+g6A5p+UCWWUEC3wVQBHpQuJ2VQOw+stwacM1g9hMrvP3C2ZLU/
VXvp1LwjbGv0w+bGRCjGFviIoX3obCdxLglIOUxwOthRhZfVGyiIZmXUHmO60y1y
wnyBu6rF/62YYL+iF8ypmotn17h/oLWP7RF4++01LbFxy7S7/EPMqDGaYLdgb92X
M6VpEfHOxHNA5Gk9lZ8H9Fd8FzuMSAR9jZHbFova562vYqxUvKfnroOfMzMr9+fZ
3LrIE7++VMwmI5ifUplhBuNAuCXrEZwimz6hO8oFrOJWmw0Eba/7m1jQRxpv61FX
7zdNWojieY6MUUHaIbqCb+PLQlgcEW4jTyZnikojrs5yfcgsh+QDa9+KFlCcVEmc
rF/aRgDM7wV8wIhXhK/Ji8E3eDOUv8BInbLpq607rmiRielK0GHI1N4I9oPjRVcB
q0dmgmh0xqlbx6/FhygUPgu8qnD7KzP3dIkcLxT1umkzeTGhMiAFSORJ0y4cRpu0
VJ8hrgQ0MmPowroPEHks/MISfRNGwFwBphs2JhnF9EPbQrwEa4c7ryKz93P7/7nC
DuXQqxvSBywQp789e2i0lTkTZ76+eXQXznsEKjtCznxCnJOFqpCNJI+IYtiPvDTH
qxqyIXieQgdUohp2f6HzOYZS6I3+IZrU1/3iRFFmy6uLXRgcs7xSliM6UBwqMuRH
amWc4Rb5wV3nC5uFOagpPI87aoNA88/0fLF+fXQmPAK7MpYZMEBOgsFUbvpxSZez
28kv1Wis8wUlGT0Nzhk+oLs0bb8LgoIS6cpaXMYBSMZ8b68D8YTIQAcT1F4y2pLK
f24Je6TrPH7w8zC38nAJkOyXUERsTZvRQE54HHufaHSx5YthIZ1uYsThCuOGAYbT
etW95flYrXT0Keb6gncyg06NmEOdEh2eXHACW9aNo5hPHPkdHXRreQd9FnMiB7P+
Li+/4P0/v60CmcVIw40cXnZaQVTG5Fjl/N6dddiN2EDo5dC6NivjFnGSXNIN2scA
03iBS4yKq4Jtt+ILbve9qIy1HhfBG2PZ06Hlp520OAvwjwwyHduNUhEv22ScASEy
Kbs72I0KbyY1k8NjVRvtc/vGHdubGs6g/g1DByJ6IskjLrpgEaIvOdWaUPmV0tJf
7JwbLOjofWKngPlgg5Rv+QdpjL8gBkRMFoLm3QBWzer2marNR75TIp6QpNHE5eH6
ZgcpmzRyNfFqropUWFtZ9jxMWl+Xyf3a9DQrTDxKCFXY04QFr/8ixNzKzEQT3I23
+eo5u6vndLbUZc3ArT8BBLnCJ/sjT0browIlLkYrHpn1UCJpxgeCMwn204TPh9F6
lu6F+uLXUNjqE0bpCSzNNxQxpNbBujnnZMXkV6EMxytNvklJ5gH6WE+Av1RlWuCq
Yrh77XNVC5/NdfC7lVC/ujWv+It6LjPOWn0GpEjTlS1bXF8hyq+VaOS3n7fT4PLD
oOc8und7D2WboBWiOmlAJXJhS0JfJzePyZYdw1LCP5UtEo4z4R+/Or+l4dW0VtuL
tm0T850y8aJtoUUW9mU4jQDLCttqnjBUFSO9fU0aebBQ+/Yx4X8kl7G7WA8KJh9B
hizPoVca1taJOU+1BSP/BqDRAmv2AUHRTcwKc1qquSt228pOC/+6npdSCO9GWrLc
GJJc3ZeUWtZw2sZEzoBXB00WuVMXiAfwwJmHG6XP6xYyK9KeiTWq4Osj1efJu0dH
5Xs4RK0+BOst2epkwMhY9AMSwNM+hjYIPqQolgNk47cd9i9zs2u8SUWswC7wxJox
1tF6xAwDEvkP4cTvf1yueaD2crmfRgwLPe6Fnm3iccvke70WvISEuiGsgYm4sqei
A1FkJ2oBCzhDvfgNcUUf1L+F8tT6bildSaAqLucN9xpzdf1eJqeBrdgV4JetZH+k
PD54cJY6x91ksF8VxHOai/9dTiRoJ663dPdsAt7LZW9b7BMIWlF9DElkgZu5uYH6
TRF7tdhqwffwz2jIeo16+DtGNofjoNLFQTUNTIuW6WQ1SHfyD1ZiLmrb7VY6+wJP
J0nK1sP4XzGE3tMsy6q3e/kUR6zRK3VSiseqsQXBqz0E2aDNF4q/ITy31iedaPVK
Dgyxy+3F5IOcOVwaBeEdcqSkM+yljh3HJWBDChP5RC6akBh2+fvZfYiU+1nFtd09
PLwNm8d2Jq5qf5OIreq82wwa7ryf7Y+4kb2Sp9w6U9JIVXRijXIxysVkQ/jo54ei
/TKE5Q8P3GZ70MJF/YUNgppUYIlyJLuQNwOm7prSBY80xe2k1r2HJqTrFiPZbysp
osIeXXMjADQMOxMPW+edtgOHIkFUGW+hD7z3kzE8aex3m1UiofEFzrC81TRr6blH
czPFOGrPmAy7fzUxwWiTa7sLZ1hV6DS+DrlbFKmpo88sQTMOh2450cgxzL3/RaJs
HSPu0tu0ArbGaymQ2LxZgyDug/GQ6o7TGVqNdjZ29lbYAIPanBJ3KPriCMf6LK2y
9+fF/H4NxgwyroKUF8g8eiEYM4LwElgQjg4W1Gt6CJVOHmPE/s0AprPoPNjidfwS
P0TBvGjBO5QeDezPGFWW06RKR4gSOLWA/fEZxaD5va3oegyZCodVAMSWbkodypCr
dAYzWHtOKkpYKZUePNa08UlrbE3lmLUF96hQzQqWwOwtSROfoUPbTgrBxnWOX0dW
8xHF9wXNdiypS8DduboS5GHMPvA5bdPSoCLMWrOeWJLBqv+EbdJ/xrk8tPRVVpA1
C81JUR9+Dlo4Ov257Zjj1KA3LY1dhOYCO5VKNUxddpKHEz84AW6Dw43kY3lqfkgM
KKagBzkKKpMgM0uy1i40F6JHHjyOEaDbp1SM8qNzY7QwI+qDndc4PY23TNRGMFGp
FrViTfHGzKXy3HYNewTZGwDgBRw5I0iVjB3DUJyPuVPbIVmzJj12Ni223eNtmWlG
8Vz+M7g0W3h24p3VA22WHkDlZB5Uzw215ryciO6/BscDRig2yjZfC5CSLNClqRjG
z1jQJRpZsYGRxOOIAVY0I+SoSCm9VUGmOnXfosJkq33cDX1KSKRosbvbFPUx5WsC
mYpJhEMLxwpa9nNHQkE3HKHRlfz1mDDKQyUMw9I+8xjN6neQz3g2N3q1qly+0RhI
WnrhKbq8R1d/aO3MP2N9KQQ/3QC5rt/rGSL4in4hBjpqIIWFOAbZmY9IU5cA/1Vi
wBGSgWdNoawy2ZiIIc+oD8Lbec2rfIunCBb1E8xawr9XHehE7sjec3bHdrB+UADc
RiL4VHE1GpnD4mahnwOZBi3MU6w1QfRTYPDY2DmLznIKHH9TLwMd+MEhJ1biZ8cb
W8uA4s1/PHOiA18j/KmXn5TUWToDvKF17xLhlq8EcWGNZDmwHLSOeGx1gixLxS+8
CleuOPoijymbDUG7V7QTj2yPTQODyJOo26HsTxuLC5t/FHq+6O1aw5Z3feKmYFm/
qBLUcJguANa9/BlANYRplNiKKKB4VtKEue+52XytefQvRpUgXOmURAk2c0DD+EdJ
xm11vqcIbVzmqveKQDkhEQWtQSpS+Lbo3IVGCxng0E0ck4w2NmYMm5m4E5przOwy
5LozHyqH8tHKlOABRaBNRevIkak5m6QFv6N5Q+MFno+fKN0uGQSMR2VZC7xmccg2
55r6TlKGtNQ5tdqBdTjeDOa5GIQJCcvCm6m3zSiwjpFfZJvwfY6UVE81Zg9nX3Du
sL2xFCV07iU3nTfQaPv9QeJSnTih6Mc6l0XdHg8MOd/YW54ft7Ba8q0XP7WZBJJY
/EGpnM/7lyXAVmUxi2dFSKx7m8hN4erD3Yv9ANB+v3qwnqhFO4EmwFIo23JSNjUc
EHCR45N9dFw5qtOzG6IIy4weyP7vruTsNd1r7tROAyy1kw33jOPMtoRdHKZpdEio
MBzr7+vcetEOojn7ikkQ1OE9lDL5d7QjksUOYxnEzR5L3sOuwmnVWhdrCA86xBpz
0CEDuInxelv2N6N0ZZYca+ya22VFmwTWkhDjUi45klvPalEHwxFOzkoL7miTRrEH
TnpgjIsSdcOuM509h1Szy2Tx+Bq7kyss+XBCL//th7OzIIRUFokvs8NEzwDjXsk7
3dJEYBoUJLRYbA5eQRFYy2jN8VWUXaDAwad7koY0FwWdKlqPMyn/U6DBpRyJbGgq
BOSviG3ZqwtjevA8O4386rHdZPLksjNhbgSzNnAvhvBVmEIVyCNI+pcNiN+nUBFG
X7LCyWLCIqE8pEHdjvzCCOfHN07+slbSXXCa2VLxmlRAQTzzy8kdwcKZ1UQdgY2s
OaX6joX2+sflZ5wrzSv2zq4biuLyFv4sb4nmBg6P9WF+FUruVb/cakJq7tuv/pY0
/t8xIADQItT8uecZh/hsTTGKS5V7RnqJCV6AP3PcVjnqwoVdO1a0RmULUz4khB2A
BIHYj3zUYjN6jK0c3BAgZ0wGoX02RhxUBnoRybO5LxckZKOAg1+31IikA2g8YiJ4
WqoI/ZpKD/IQqkuCdp1yX3+rNlj7e+U9dW0t6BEs1Er3++/92eRMmBwj6r0TACkq
VsD0CVW1czzTXnVFz3lvxF1MsFrCbc3t8/q4jakOVAyJ9qUBjjNp9Ywm+dkjD6x+
7g1Gi+oTJ1PXpkfhfm9riebYy3EqzYRJuoV04My6FFTnyOE37lix2AnqGy8NdNBg
+9U2M6QswEFI6ilIfYYSbVlAxxeYzhmD6jea10KfOS+GRkMNhobq7Mgd48Uo9pb6
sCfUiWMh4RN+oBfpGv+GFPmdilMI9zaE04s5wpLKUomqSHILeMZSaMI9PJf8499d
paw/kaNcPNq6Dnj/+Fu56mBuD7kfPCsAnbDbtTDgRnozA0vTuVzirtkKqCsw/N/K
58Ys/l96/T+GoXW3IIuLCeWZ9QJ1/ewyzMCo2L2JUjEegPq15/e6VJ0y7nOpoeHl
2adaOq9I+1p6V8hxyuf6KOqPrqI+Juzd15M0HZwGTkjUTKBoypvC33EAqPvWxTTY
qMe4l5olvyppglntdWMnjUChm19l8DQDi/uwUuEfw94BD7VIzEIjPR50VYx6DMNt
6nyA0z2YTvjp4wiPVqMmpcv4VvMGYZcHUd5UiVaR4AQYtt6Juez71xJ8u2kXV4dm
Y8kt52hVvJaws+9S/RQXIli6TFpBJwVPO2Jvso/EU2S7DyIfXvuHaqlQDZ1HVrVg
v4kwga+/P3XFFKfOzc4p/XWMQR/XrvtX2UPZJbyzC9BtVcrby4dkTm8MQDyYLruG
2GpQEvZuNLNBKCyZjI/ke8k6ry5TGWcbCYmJAZ4Ogn5SIPiqXn8ZYLYRBNNK578f
mmUILsWF8PIhuIN8k+JXsDpcaM+lr8Y2aj8k8IzTcqSA4T0CvchdthV2TOPSlkvb
uLnuaPfvHSsROnn8ZjwiqtdeEfmwGDljE9r1CtO1+74cp4u2JgEefQENWW7KY9PH
Q9SrJd2ORh/n7webCluq9BpUwlyVeorTBz43KSn5u1z0TmDDo7qhKgrbvx1W09v6
EkYZFolOATBZSQ9vzi+2dOEGm3NNw2aDsEw5aWnTWQCApY1mZHElTQez5h2kg+Rh
9PcuEVxq/AShvtzatYYrdvcgHZcPFVrHauI16UspusbQBVjm0hQupss764uHpKp2
qYRcR8YisNHZ9v1gDq/szjBT3OroYOViq9gAXjNU4k7+zay/6IcBlMRhkdXqSKcr
NIMjEK1jFlaJiIlbA+sc+n0QY/fYMMxH2w8bOM4ZgOFYjZOSCsAyfyN1tvu9XCy6
3gwkgZh/ZZWMCXcywWUPVOvetBMRPoHd6nl+gd8Z8JbELs5B7eZs0/p1ZYksAgaq
tg0HtxiyjJjlOjdxbQOuaWk3rCPr6Nmuqs+SDfx3iDm6CwslN/pvaUxvgjUNohMS
bJ6yjiNzwDMbmVjwua3FewnQJJP4WFFsaMbz4BwdF7zjFdGNp0tJUGR6+Uk9gidW
EA+II4gvQsq5IjQOS2rCLcusvZUfwYERvwwK0JuwpybSaHcdmWcJenBOobdHYD1h
dV8N/TXDEWwn08fJuuE/jRlGdGnAV7eL6bFsjwfsJvtawoOHT7FLZMrpJO0Jxfk7
BGdKEQ+2L8xvToQduhGxgO/1ehIk9eIrO2hD/J9tnN++mRVicUFBL2slrvLAytYt
oYt4VtfNMgSGG148M9SZEYKOhypNxguU39KMnalsGkS6baxl4cR0ZAdhkr0hKgD6
iak427cxf3+0u0hLT35Oocui7b+df93F2EcvgyTRpE3rliWeI/5ai/iJktGsCOYX
EHKGb1F0PSm/bc1LPsLl0cVDbZBL7q8ZUrF7qxolkBRSyhyTqLA0RuTJ7D3pdj1F
anQF/yN8nrvoz0yYjuceIF1KUbwDcgQmn8UqFcTQIzS/OSpDGuMgRdtJnE6NpCtK
s189ZlRUMEKZlfB/yXsQy6dfiIpnlPJEsFocM27iJosI396ioHKHAT1QVLhj4A99
xnoGshWl/VFCdOTZ4elNRHafxZS/hWYrCR40/DwitMNDeKn7Di3vh9Ws5kyXulQX
6wqE3erzA0D4qEfaNrFnRsr7E6EYyROVts+jd68M5ccPXOFjlAt5PScgNbOxoGDW
+vIaNv87IMOZHS6lz1YzZ6eIV+O8fIKz4YZgyRYihgJcL3YpLa+KohJxkuAZMkQV
NWcAMZ6Jn95VB5n7l4U6MV5K9aH2gejuX9z2JiSP+MYgeXv/9ChIzIscLrLckvv0
GQnrj6sNaSymIvJO5jLNc5v+Z7MCieF0dMrwg0jDVgCuU7qZH1e0KI4tWCt/S32V
lmRcxxeP7pIu7zfaWCZ5WDcnfTi0qMSB6WhOuow3HL2J0aoKgyfFgI7s7iexfpp8
Wkg+Vg5lGW8BqSlQywzaiil15NNI0EuP1F1cEN6hN0ayinAwAcgR00I0k203MtId
GHgQqpPfVlTi9syB9pKffyv+1P2IwZn5UvWH3+dvZm7l40tPLzSBVis037xybnws
P3oBi0ASLPgtHjQxJTKRbyyiTu4FTiGn1nXpZk0hBu9afggSbaAkTrXMptg2hI+J
L3LjuPrh9LAG20zEq7zA8d3Iv8/KWpciFAkllom8MIl3LBxjIcC3CvHi8877Lo2E
jM6QSUsWm1nsTqOrpmO/ybfTpA4hFtLKP2/6ltvmoPVmSamznU+YubLEH2EnnLDJ
e565pNADJ/ph7yg7fz6/heWAKEq7IJqQn/3gQdb1i07KbZEVYUWEHP8lw3NEajRe
MOkru096YzRJKeF+7nG+9rtzk5M+QR22m+5VAfVYocMbbDWnUfk3Lky1epytp2ML
ioUW2mcNocQTXuvKUPKeYJa8Czods48E/3tdUisveLc6ehDINr1jTL8pJQ7siB/v
THT3XnT5wml2a4papuyltrbjzdAdIDGwUilOmr9N9UXYdbzhL5Mak+pneAOQ6sfy
G8876bWaKx1XNz2W091lxEM3jLpSrX/jy3P6mb76KaAd3iOUowvFgwZCr2dfEbWG
RVIuUJlk8ghwcvx0kp+O/PWbkGLZsmmDzNTLACKp6BcW5fEbJF8R4/jP4N9D2/Xp
5yJ6HkFJ0+9QjT75gBc8ENAOG28Qz3nnJ803RsItqbBqxS2mheFLqClzITvXg3uk
gIenjUBgxEflQ5uCQhl8jdPgDb/8nGCG87edHOxiAXEPN+8kVQKt7Lde+Iitvipk
ZzEiIz0PYvOfCDoh9rH6/IB83PX+Cr607xABHXkwpulq/0pCRLILH6MTx2reqXOK
eN88jsVI6pmBYjuKZw5XM6psJh9FEwaK9QwhUVnTYBVyI23KvmFCqvc/3JCyeH1D
CUy9Nq13jO11jtMAKmmuozgscwmsmnxv/9sXoNJDYCNCuykwxCDdEM+7K34p7O0x
wpwqlqJruuP1KwcKd7wM4v4FLPIsExgkyyzcypYvb3SX/ZO0o8perw0Q33dPDVPI
88eUKhyFQrrZfDLK7OhRqIQu6/rGvePHgNR91/yaBGu1ij/o+2DVfUA1J34K6dLw
txA3KPpkO+ysCcS5rjJ2JsB+2kCjThTuNDhCsXKtIcEElGE2kVfrpn5jS2ISkXca
lIHjuberiO4OaXuVAOdf2uA1WRew19hjI7hbQZUSz1tis//h6rp9hoLTp33xJ8H1
8JhTVx0sKhHa905FlShbw6CZd+hY5kQ7zRLTm01hOUzydgYJEvLIbwg8RuLhVuXx
JIZAtLmGcsHbOKJLZpzjNoKzWrnFSD9m6c6a6UtOH5VVwk19kIEXd2fLsKJ5/IWs
3yZLpaVIbwXpTU+/Fri5Wxi1/fmxW1wnfM91vUxw6lazX5wSRPcTfF6nffl+sJoJ
MqwZc36g5/IadlG5E4UYMI4LtKmFqqCZBLSANVz9gxu6f/fSM/d8K0cjZsCnxpIt
TarDWiFyzwi6+jmBG3lGM7WKJvGIFs2F9pcKma1MYToXGaKW2mTMhumHtT/kK1Zy
R92H/D/6QuL6Sr0cHPQAKFD+2UAwvWiwlPSJ/amQ1civgTTs3aX41wC1+YjbW+qq
1WJ3I7pCmAq2wQDV9fv9qAv6bw+2FfPYP1sZj+i79PjHgXGKHkOG8qpKdZ/obmJ0
ZqBnLCEPZL/9X8q9cFArbF1XeIIOXjxkOGwiX6gYypPPl4u2t82sQgeZeMAlGL4Q
Sj3fWmj9Kwmde5Sa8lwBuDYtQlpsPMntxexNDKf/z1Np9FhewYtgWiqzFJQgurR4
Ea2dNE9obF2hdwuSq4rrk4iHdw6hgxGkLBuWaX9fR2Mn1JgmFGKfc52MoCU51yDH
KuZZZpBFVPQc+/JRXfydpIrIbc7Q76HK2s+Bssgo/euiYCvWVGxBUZ6zPnf+iP5A
b8TuyYNTiJ9e5YSixBL2Is4B4kAeAiQMxPRy2jB2jUlKaa5zSl3yeULt+SRK6QEN
9YNFeUeBY0t1/UnX6ioHCTXx+TRCyP9hrwHZtdm+GAvu1WK+zBJe1/WVBrTabCyc
684DK6dUzmcjrK2bbU5hqd4DA/aTl5oGQDf2l0hiFCPhvA2cq/wN3s1zSDrmW0Dm
Oytj3SEX7slfxUjbHOLsFHjgLx9+YaCRS1b1TRbpZ07qjhaflsYga6pYglAGqGRs
DJEvdsDlv7GpwX+FPchQ7/mCJHu3FXGE7UQdESWn2q6s0+FrKMMDXqT6HiwzfdyC
LC2YA71gzw9o1uxzODYGOwWP1GW4fdtSmrg3JdvtWDA7c62RZYffE10ywRweiK39
U0Alt8sSLVpqshBNvCYX2nSGfBTBmeq7EwLkBA76AO71ljeHyJxhiP9sJUef97bf
Lr3bRX87QNzeosdIFntbHj0c7sqgynoMVJTx75kimSP+6tXlO4TwM5M7FfQhkDBu
b6LVlJFGr7QNhypg13uYpJV80jPklqep/cqKIwJ1Eq+xkgq6reHEtrRCk1LAdBF0
mbviuRpwIef4C3Iwbwms1fwWKBr2BoNNMhV9cHpOUWqG3XdEV9Aa+1EKoCFg52wg
IbKwpslPx3Dv7fSdZ5pdtL7Wb/rDoPvuBe09lN92CEvo4qX8Ro75BAECyz+W1yBZ
XPSo7gG4LmrFuVme8yY6bkJnUoBAVFhl1l6J4tEMe8LY8hMium0WMQ02LsnBcLFr
+jS2CWSnlMkjs4nPt5kkJcHILh4bhnspBYEeiXPoZyk1dvAAPSKLNNiRVqyTtsSk
mlCLkQ0oio3ez78jKzY30cMrd6P+ceNo24rRgAFQ44xBhBUxPvmovA4NdEj8GMTI
Gy0jEAEnFGdDAuestc8uvgPYoMk6IcimMBN5jdm4+RbGtupj3hczBukX7DAkntlz
oM+rcB1bTCjNjZRTNfqxkLdI9Lh+yL7eIhk3W83ghnAm6LDzVbmG3/M4kzFQ5VTL
jsdfdkFAV+WExesSZozatDWGvY68pHFtkx3PTnSypFzbJ3G2WfGHKJEOedE9xMy0
BBnWHWzi4+bT0tsb0Ws6OH1ij8xw/qCTQnUcjlWUCzXNCHNF0yDkn09yI3/+G06G
s78cwPOtZ54XqyHhTd2sx/Zqme/W7xZt0OlMd1czqF+L8AedILZqxkkhxBmq62bW
kTh8sZ+zH52quRyCVXmYizp4EuHLUJ4cW9vWGSwUcWrLtvzfnhYtGPmI8bBUeE3M
K82FdncQ+EJE0As+7Pa3EQsfYiuhGDspxV2wEe9csysTeMoVj9LzxC/9Fu8SPE4Y
FL5iE24mIzh/yl+iQRC0yhwo5kKBRp76i5AKBV6GNgJmJN+wWtZFHUF4eBTh03K1
2a3LTtIhmWWlTkEMrQy41Jag8KTMD9h0oMYpbt3Nj38V2syFLz4AIZ28NDx4W+wE
5UoESSTM2cCkCPVrpypxATXTN58p5Le5E76uDKcfVy5PXmiCStGN8/+mWcF/KDTI
PbIygVI/sj+d/kYz6zQebORXfYFNABu+aXcgLOmAhzhIDzqMfSRLwvJdQSu2EL48
veOUzA+eF/cHh54k/rBCOTssl31KRtlTfDXhG9FEhu/o1bXI+wj3gAWkoMzNfin8
J6daKaerBS1jPDSCYyxqMyopKl0vx6ILgFavvxXqnHhjkBBvnkBNhGtF6pcI9jh1
rYA7ZJW3OueU1Ba5V3KCoVUEEYR9wrFnMMS5J7xOTT//WDSqGgjxFt1sfUH7hnJ2
tDqQxCJNga4yrrsG0dxiOJYu6xR5Y0ySFiyE9muizrSA0Anbf1Q4BlgL5opUWUfb
WoIY/vE9clIt4JLOfpD2sz3jYnsq8Ye/9GmIy17eyGBHISjFRYt6PuUE1mnn0Z6b
Hsd8bSEO0tEqvDnMMuB1EJM+kEGRJCFm9NBynu0Qhj4QUTc/e2GkI8xnQ73GDYlu
OUEhA71BlMiKPBHMIAUXI4bPwryNuO21EFFxurOogajONciFdk4FFSdx35alQi5w
VFf7u5xMIvp5PFtuJEPJokfxS764ODsWJtdt8iFh6SGQWvqcyvQ8/9AhU3KTAy++
Jkxg/6BklIphXmyxT+PioQNVxnpjsDsTHVq/+m22srB5ldNPyXu41c7f1wkceX6R
xbNRDyjXUGcpTsk7vnHzPGXAqCeznwFliv9a2QRlvTs+uQCZit2VeB40vZzCQhkz
d/WLSj3KdSFMeptFXQMSn6wENlvrEDOIDyB7F1ih/8b7CqGOF22CdkwueGhduFXU
xxGyWXvrV3iU1v0QflMU4NXBdGDLh1n4jD0n5cmdjLWaJdHQzc+jNbbE1hL8rQeF
BsifNTba8Jdf3n8azBTFcRRnVIPYbcMA6xRHUFFHAGpLK68IfKlf/lgGz/9wp93x
qKQB3loWYkaQXz/M8tthoQqyTDU01md2MrHUTvGOZeAX9JV0by6WjNOMCn7n4KfJ
AbCBfqFnp57MRjUMsSgUus1E4RSegykXUZDmlE1mIHem59EuZ5zp+8Co99o3da54
1wpOiYTfPk4AVhCdzReL1IdNCQZZznzBcI5SE7wF2kecTTk++Y2Fy+vtq2omhUgR
x+lPWSSdHO165k6nsHASIXtsntK3HaT8+Zii5eQ3gVLrpYUDClT11ijBh0viL32z
KYsAtPqBvpi598DznsFbmifg1/9iUxLWCU4RztcY+E4JNf1DWVa2anO0jpyVbclq
lMJrLY+rpuVHCba849nFlMqzbfCip4PN4u9hj5LFSJYc8QoCjtxFf3Ps905xM2Md
K+l1RekBSibs5GkepEI5CCusjdFiyMsRIZX4xTlOvlhmj20viC9D0LH0KDMIiYjH
hrD0aRndNqhfc8gPkC+b9myMWo8gzPKgdUSHeG7T0SARwv4ydG0cjofRcPpXNjYN
LPASr8pVvx/cRu4zpX7DGIvtGxFGzhILcXV0AL6f+3cfgNWvPPPFm3snoryVaKq9
CL7fGccBH97gGzLQ4B9QgJlvX4+qptNABV6hMm8pPO3/J3zfZ6zp1qpGcpYDBAn2
CTCZTziuPL8Po8qDsHYQA3xGiFHoY8lAOjPHS+OS2Gfs22DrGK++kW2UkW9CbXsG
PChFcSoT6C/bkQyTnnpnIsSqMqaV43jYi7q+ZddEUHD6jK7IjWMLWXzTJbtxdBOs
BHHuspL36s6b2JsyV55q7ZmCM4vN9yttWwTsAAozNkrfc3f8X2jIIqRHis9w3PPz
uzPhNiwPzruxKUBfyAWYRBcnFLthpUqH55jqN6W1deavhbMR/jhNZ8MlT3Jl6g/l
yUM0nvtpCdymuYbAtCgSGhczi2o8T2SfzGuza58yHJE+XMoyv+n3GTZleasL2i5+
z/JMdoY+7BngbYvWH5eIMB5cel9fvz6Kb75+xl4KpjZr1CJXujxCSWkqnauWjwvo
Rbj1s6ZXrnAnCmqz6U9S2pmw/MlNNfj4BWwVxPBQIDHPAFrb++YJKn11alCS3a3K
w79T+N16feF2fNjE51JFD/1BN3J5PkBguSy/iqahs5fhZ+2t+VC/a83yCNwEsoXP
YL1I1SIWF0DP98GSjqyz134+QG/kMNF/az9IDKXQfyXJmw4zAxWol0b4uUT40H0p
SlUvk3H2TT5lLmBxbIzOmsUSLDKyJfpNwq2F7WL9JO7WHRaDrOGs1pKB5u6b42fR
TH+ZrIVZ6/wSlgZVIgib3OCmU7dHNlk5T2vzEA2VTro3D2zMCsJgnGQrw3FMavUK
4Kla6B2QNz+7tpa42aPfqaVzR9K8havTFHhOlVOf+7L1t1QR9P8BSfd9iHi7Z1cO
4IMc2rU2GNTElmVgAUtiSa6IL8v9fFkst7IwyPT+DwGz3lyoP4J6NzRPD8Fy4zyd
kg9fNJh8yPhkMqwvjqqnVbOq5jll6KqP1L2uXHMb70r5KlI3S2/59h6+y8tetSr5
5CU1FxHO1jtIGg5wX0lOkF/lgK5GiM2jdPGXPhjP4xynNlShGqOWyA1golvfQpVC
CHI4oh+XG6mJLmSZji75zC1XdrhQlZn+2c9nE1OCkkwK0eZVk7FaVxFCkXBI/7Td
oL2hRNfoyDQQIqrOtMmVQXKorfUzMnd3jBqW+oOQEq40N5Xz8fbpJ62CeHB2hzao
PivLMRHeyDBWL7AMv+aHPrvMBPXSh/HUu0J38pqK3+G579FECGgSM4kSRMTDgADP
geNDKhtc5qqoKZCayTmjQJXGj4j9guVNAJpTtykDqjk5pGhjuW7vVaCgHBK07ExA
faRNLJ0ge/Cr/Y7uRxiellzmsZoHQBy03mrT7qVK1/DYhQ0IIIsRVajRU93FV8xg
3kOo3o05LN7fDjwWQJkhhIw8OMImr3Z3siI2dZLypyOO2LIJl1hlxgahQ8wqOl7L
TSkMKF1w6KNBOrwkRBjQNaG0P9fcXyHKoybyBEEhNZAH7p9g6uB65Vjl7xUbV6cd
RaaUPAM2BeqQNdMd69LKo32/GbFQ0vwagk+90OENPB7ONVVWh+WyQ6F+ZmyEFTtZ
mxcCOMoO6Rpd/XHExxMZPzjNWmQ+xYmBCd0upsbiLjK0EkqJttQI7h9hhceCG9oI
IBq4duQPNIgUgXV4FcIj1h7c+3B9Ra25fHklLnReLL8faKEFn3CurG1s0UaXyLDc
kNnbH/T51q50LnXQ3rI+CpN6lFP7+sdfn2aa55T8a5uVn1t0K1wA9U51HtjrocKw
R/JKFxLwzpoqxu+KOr9pKf7zrNtjd281NwQPCOyjVfQC9LkoVA6icXMhQQzSF+QF
X/jKnttaz4ctKXNQcVlEabMrdNkOhmWh/7caWlO2Syi9H9FiqvDaCOJYPJFfs/I3
I0pg1ZdQSz0DmqKeAwPhrXp+oRaFRcuYXUiF7LIoOPg+LeNF/GzNEJ/xQTiKCpsG
a+OmSGf3iBOOzNDH5QCpcsWLl/XfGm1Cm/+KnyOWgZFONlLVjoET0ZqFOEFLJ+I/
i10NPMFDqk0CJOUY/B5S9wqZ2Uh5KqCfMl78dS4X6nG0DvlJJ/BrwGzbh9K568nG
/FFG6H7VOvVDFg2wTHlD43UptWoNuFImb30rAjUrt9ox5HVziCrJzyiOFhQgxv1R
UPoaYcyoCZBRAszUSfBBTmqpfIGk62JU/9W9cBnnvLp4pijafXJaxmkkTH4c3Vot
NU4okF65ZaZiwPmVY/RtrdZh10PVGYJUi1aAjg6AuKD9twU3S6nvEGQIdLb4AdC/
ZZ5TgjDMmfvE5xHI08cXzSH1YozA9b+Ej7EcCAC2WfGQRwuLwvfG072n28CMTyVx
7B73yxt0Oz5s5wtLbYM/ZnFADPXqqDmYoLjS54fuVr+H6MmeU29KjJ9s/p0T9iN2
LmlO1YsTtQIsAe9a66LRtGJsopOePZbEI9wjGIWw7ucDIW31jxZPYhbmxM6JJl4A
fxAXfAYkmORkPffpJ/Pv9aG/MaE1DPRWEceJVTaYGnBVWE9JLX/hY4pydqn0uYx2
iL+R6+ZLJZ9t0kdp05dPN4dplyuqWUwb3Gbn7GvjPKg8bJVZQELHX/erLSzM+Udg
A7ZxcqBJtMadfq9SvxwaO1IcQr8a3ZsiXdswUMHVEZR+4qASU3IXxV8nbrc5SC/B
aRT6VWVjvE01ESl6VOQRewbJLQ/GcdZVH/ufyMbGNoqII9+xtEkmw7aawzQF18gO
6/POdNSzH+VUJiprKz47o51FKyNa1Y7cju9tuoAq7RoPoxyGYyLz1zL/pWYkb8hm
Wc3bzasMS0LauhwtHfIOUjs1SYUr2RoTLxKhuThi0GqwQ2s+vfLi4iEyD1S4whS+
t4c9LEmp8YUnaRov8gr7br7uINnh1pUsktUECNGHZSJTMBjMJjE3s/rxsbViN/HU
rBI2fJii0KMvuUjyrGEVVNsvKqoM60NUwX3eoL5QIfdZlBl5YERDj3B3oiXuW6IQ
a/MtJtCjyd6/ZPY8FArSJ/o7zjFHoovSNLVqnhoJ/hrah3euyHDPLhKvGn01O+k8
LnTEkgew3MlORMkpJ29WYfPvsXFmhe/VzbuFOFki4PHHeVLnqb3mecoQUE90TH32
o5guvZ5v5hXqjzNYs2QWpGtcyQnZ1C6R9YpPZsKgH4acWnmtuT6jy9p11R17N8af
yTSzljKSufAj+MZL/QCpOwHrKS08MwFXEYEeGfCArHtQ6hKxmsksSglTKL/8sYAE
z/eMiaTenOgQCAr1BEBY7/EOMuctdwOQib5GgC64S1CF0NmOKYlRYevrdzLxJp21
FY2nX6GSaATiKBYrXe83Hsu8aXkkgLVojdozEkv7BXgBqHGWTlL9+PLmAyT3coA9
WQGy2dDSPq95oJu9EYAfL0buVZIDjeMd/YZGV4U+uFuk0KysHgY0SOqSPhAep9Pj
+ik0BoXYAFLgtaa9WM5FtblVIPyrzgI7ydSwsicNPGISdjHwe3c/H5UixSMwUXHt
k5R3hdwFs8ryfwGK9ucJI4UXeF8mG63niZFs045bnhscFnsJcW4AZ0VzvAEPwnAs
OmLLD/ZfoRNkWJ/xqu1QmPt+b14ypP+qMRedDuNfC5p8LeTKz5xtFhqctB/1gpM0
i/dPE+r2AiRm1afZXykznE2ClN4KneMxMipqt0APOp/ROpQ3hJMEfGMJLZAZdzb9
JZ9V9CCxSkLcKcZ6gQGyhwHk8qpR9ZY5f90UEJgVDVFoYHyIjZMQ6iprfEq0Zi23
obLzEJ4q4Gz2Utnsjm+jmLLhQiWQw1Dl8C+/UVG32gHhN4WuoMq+t7PWqvBIcCWM
YZjDIhq1EiGYHLbgbVLWpS0EjQCxidHaylCm9G4nhF33bgzKGK1PIGBfR0s+gUtO
V78m36O669LogXgtaZf8/HjaL2pbI/vOOiY3wsVSV60EqjDKb+9Ov7g/JNbYyQdv
7s9Y1/O84bbswF4IUVqcnwJ4xngZuXS8iNhJZYT3NFw2wHRIPWDWVyB9ud1m1u/l
iy1t3vmQwPkJ2AKIRWSa7nznfBZ9cJ5shjp1U5Fwa2WKjvP5t4ZasSk7tHE8VY/2
KRHcXmJgllFppQC9sL/v9nCfL4GEiGScCGHV3dbmEXGeE+n6LG+HsFq6mfK0+6cM
4W/WT7khiU4QSoVUrZvXVQzpMbFVQGS4URRgo1LQi+FlGRzz4YWbVKdDIcYAx6EC
tBe4lM7dCGqwaLbS+NOOSRp3dWdvdNFQmXxZ2xta8K5vZj3dQMEzE0qqq89a5U31
Pr2EMBwsTk7gV1tjUp3ut8+SlJ+BRTnRHpyzibhoYMTXRaq631dt4WC8AxtX9/bA
KbTm0PSo1u78fZyqk+kx1yR/drTR46Uuru1kTC62qq8y7I8GBn703ARb5Qjenqus
S4OKzaFiVBBU+Eg3CuhDdffeTJ3ocs38Q7dVAWDz9sU6OMtV2HQGJ4fjyGcRdOl3
tt+ZykOkVOtwLweKSQ7UhUfAhaUcQbKxB77t7B+l8dXZfcINXNjLtuw7c7W4fp3K
0T/ac8F4R+/lRO36jXBkJFhwKf2bElOZwzJmL5o+ra4a1kD1jxfEpj7ifB4zPswN
JvZXDsRZoKTCSOY+NR/tx0TIP6Ooay1E3KF2dLGnjiajzuqodgEzHJb4Dry9Epx8
ap0eIwAvGXpeuJktm6r9jUD/60CFJ+/czqkEJpYydzCmvjh3AIv8J5VhPBusNm1u
UbtyKLlHLovm1x/pOSvLe4cK2ELnj6fdUnRAFs9Lmfk+5kNEnkq/qF3rVgyKumuB
7JYAIn55l8EY2Pj8QxeCqGDPmhmlnK2MZvuizxgNbT5n0ckzNZ2nDlDGsBDAWzAo
8XMOnhb3J4pHArMBoQRLI+IEQThjpw6eY7mIZhLqfGD0FcgZLr3TC6V51EcEQt67
Q6ieGoq4Yo/2K/2bkYY6xyPkA21TU1opKDPNFg2Uq4h7StN95zkBCSnFn7lAuLI0
LUXQ4YPR5j3UNcVGhuEr6GPO8nWlwdFge6INnvFUnVAzDa3nYpjbP4kM1kjxgTJP
qFTG40rQsX3qsKVwUnXvCpZ3DCJazJx5jMvM6ie1iPS9uBsPuud5lmQafLGpSSV8
gLgjn1FXNAMI17T/TZpwj+hhbmn8wAJeR7IC7E5iwAwCcgxTAdwvo0xgSHVRFrsI
QvtlqQ5bhHWXp8A/H9+p9OMvj96uPUiLA1jyXDGKnqVqBUdCQOhNt50v7EWSbJHY
UzMzM+cuPYnD+pvrTYg8zwajsKe8qSDlkZ4kJkkOGbkfumlf4fWmu+iu5TqVA7XR
TbV3VWmyKWcdgr42Z2pcmF/ZDTtMvoboGALGgiRZY3l0S1c9S/1lmct7bsjNDWXM
yM411J4X/cItSbos0jfJFWM08QFAggzl1Bv7qvVJ+JPFlLJKeK/VG6rAOfSToZkG
vwk7Ghe2ZDU4ncK15pe43zDAGJ1lrmCkAhe480KP03UOI9r9bbRrXhR5DdnR1eKq
BzvqUbd1ZqsJcRjhkraCMcZFJgMEQRpsh2fbCTO8VtwdhdLtAua1UwIjFaK2ySYh
tF9GjpeFaOhGUJOGUszc+hIpZ5llQawQqfZYgyEcNjhuFkPnD9nP1hgJPIywPEVH
bbDyLBpaPtHvBZY2BAvnLhPOj+hpRH+Q5QZv7ZyTNGj1BuZ6TAZZwe1efF/Yy4dE
DKr8zOmD5NxRPrVwtRWWu49X58DaHsAwxMaT9rn1utpgE4qWdJcaA/WFz7bt5VWC
XSLi5hKqeq5TZ/V3OLF/NiRkbh73/hITqkXEC7fsHBiclz5QeRXxyGXMD+myBoMo
SQSEBo6NSpT+S5W97XSVi4auWUruIh9wvMJuUG0g2dqlCED/KvJ6kjGvMqNRLlUS
jqXZ/Gphp2nb5mu7ysV++XO8czaeksxPMEUvw5mD/rJoOU0mwqbZsONYWGzGv5Ke
sDxLPpcmpcITaD/zo8qDN65N/FOd9SPWG/HrY9t6XT4vSNOtSUum/aOJCYW0nQmd
LxEES8CEXuuxQXitK0hEqLXw+KN4+GCNdE0qRfvp7wFIIVJ/3ZxHC7FbdCqwx1hU
QdCvL6r8Prjf+BqpVz79p6nI7OxxDlpjMamztMcWNvGaycxZWYfkNVCNTjZZ6++9
KPw8XlFG/p+JfNdu4sCjh9Wcy+Sd0dCTpKcFuA5b0Mge94Nip7RN9fIIu6Q8RC5n
whTk5xavJByyJreweji/6l7+rTWUJP05SACGwXsP7CEOF472YEYVyXoXP5YTa46u
0Nr+9VolUeVBPEnSyAiLosa+3tixbqnQHREyChcP3vdNPCZ/sj/JNrxqvACfthEQ
o83urvR9S5L3jqATELMQsgHDMmtVTyU2vXjuenkTXsqZPkQD1jJxnAXc0XCn4rp9
aBiI9dcxvTbvOFzpnXYoA1GKasx1E07IBZfNVI4WWqqo7FBJhToKFhYYl677SMke
ozGoTir3nWf3xf5jW/IVx1EaMnSCD3cHGAIJomCUMUSOojn2BdvZv/N/vA1PWsKg
F5hnkLsS/MU+TfIamPmGQvgKJCyV5TkS0CHXN1pL+Y7HgVI9G8UUynObBtwQl2uI
wHXZzc0GqcNCPFvfBLO5Vr6wlmlFwxOxXOdYYOMV0t8bVeKOdxOz2MpNDvjYStbS
TgMQalI6My5+chbOEI5YYhGU0qWb6rKdqD2AnAVJy9zQQEmhbomMZZZ0kpGXz6q1
ZQGv3yldZag4BAe8SxMvqGbucezK47KkA/u+DhFgWGt59h0Vwf70MpIC1qC7gslr
OGyHTCYXEO9VP+NXEyX6QFC3lM4AODpaHF+HPrmzI1PnWaAYANjR7NB1UGyHhDCq
a3oEnaK+fsYh62j3ZTLVMozKOnIf841KmeOgu3B85x5ZqwbeATd/pOhQvlzXLoPH
iCDdG7O0J0KMaGZZrozu+yCdufBUmKR6tOZYPxPg71Q4MoFQvBHPjcItPVyzKwKV
CUNFYwTrPRx/VEKqsoAIv5htxgG9NHGw9KOTes8US8/5/pJKeXUAoTDJjROOTtbC
WKgw0PdYNTs/obZeBk5x1oeP+AsQKaNTmVK3Sggs0keYLdAY1PuZmedHkElp+rxr
MUI7i2fFKKWLPyXq0RpsOgUmfcDOAsq6Rn7uc+4wzM+rW+qWhdyexhc9tHM6l6ao
et+H8so4x31tTX7l+Ab8eW0YW4jY/ZMoMso2yRiHDMsEzQsKfAT9AsFafr3QCh9R
+rPXc/AIikIWigv6m4KIO67A9mX9oFV+Enf1FCn+/g5SLkcojZbL2VE8TJduHqGm
h0T4Ds65+ODmKaMs3MAWDmW/oxUaqVK1rAJR/iSDdqc4PNHWr5H+RV0xWgHthIHB
79WS/6vdkEjrcJ/QNiyB37AQHTG6SaZJs9YlaHav/sxxKGUfYH1SpiIPaVDMHAVO
ymWfkbVS1RWbHp6XCL1xiLMtI/CHKg929zGju2gz1vARoBjs1nQkcP7nE6gJV0n3
TOYl1AIEqW23nn1KnQCKWUatBoBjuXEXBkkLW3VrhrT3Vy4Qmxh30lMGLWUAd6MD
idSZ8tcCBoKNwrgikm6chb6TOGi0Z904ywqpy3zprsHCXLzxoOZf4KUDavOT1tsH
8TR/KYLr5aLFuEzyQBOj59dsTgnfKso6wCTtAxfPv/9FZE3WA/GDFamWQ2F+Y+m0
rzzgyPhN8+w3skGEtINfN6Mm3MdQIBdXToAVgxR5+PuUdUlyXCTpC1GD4AILIGqD
FVXn84GOQswEVpH6fxOFuNvcDu0gEFz3BJMgbDB3AVWwBFr5jiS8KLNigR9IBsVK
hWpVKKhXBZhFNujeBzHpjS++hkQSeBMRy6bXIdupWLgr1jUcYssEq6+NCOT9n9l8
rOw/2MiS95KMTZHNIs2W9OBUHhBKd3XO3FsBdPS712I6heU+D1MJrSE9W0iqos2H
jHwlTpgT0KPiMGwpbpdKdLnEMojYJRpnDHFyt+VvjjzmDcdktAXwYgND6edCMEJG
mB3d7gCi5RG/Jmomn9ZEJIsgqsSfAe9Ry6R5vLFnJQWcH6bmMQB4CpHqSPhpojij
L+2zOuAiv9FFArV0d633wcgmxay2jCJ+puAAcvCpqufFiPMR1+qcc2CFM1rWTUlm
5zQakXjWtgZo+JJE34H/9jBSRBpquA9W400aYIR5I8roZXobIdY0kROmwyYugqnt
MVMOGc2KP4ZNsWiG5L/KrgyqzYoNygGeN1jKDDr5YOe9JG8/7dEDqGb023De/E3h
rDWPdjXTgIxUaqwClMxUOWLhymztp7FvwPtaSpnyYFn3JniXVeyhp1PgYbHy32zB
3TSt20qokpZZB9TwrwwiMUw11fWs5dhgxTdSVonEDtBJsJk6CxokWgBOw1LjMxnG
fZla9F/4AR0HVn35i8kzMbRBjlialykiZ0YDvSkiB7Xw3/3R92wuEVE59uyuz8m5
YyZ5+jSNrdzM+f1RKv1eqOaL/5zS1OzUKetPW/tOhRg9NPFV+b4D2TASw5MVjg3j
AGgrtAeVN0l6XgvVRHbQrBrL10LIuhmbEWbd0/adgBLgj8BzXpuzBuDfnvydkMwk
9hD1++nTklLu1OL8ldXbF0Ur7EWpmPSiuY42VKf2lDYY+uy5iOlIUzR8BkD6uFKG
emqnZgHWQ7x77f9JP0ZM/R1jgbERQCVzF29bxMyQ3YvTrJ8peBp0YXRG+hIFYGsD
vDDafwFrqVPk30BQ9/tHAy9rypTb7PJ8YxuHYJiOcIU77gykAHKV/cDFoZjbzc4X
NCOPxD17qb3zm8pQjTUlRCL3x1284dXslw+Vra87imMorLLfRBcD4YWnZQPt+D9E
RmuRn1ADSVXO8ZW8g6fW49zYlOWUrVv47A4KyFMXtREdW0oD3aC8Yk2DoNDc7ajB
FeKx3dIxbnmY1Wc+8RlMVIQod9UN2mDuo8rh74AymWJu92ZiMa3ZmosLLctcpKKE
bosD39B2TYJ73lD6LSWsc4Oh615ZitxSX2jH6Yf54vjYqH6Oe7aHhPASZoKfwi6d
5ihxfR+HVFs/n7DSjYmcYsUEnovO6euiuGmAR6BwFF8loB0qyz+mTKxqi21dZiPk
sswvHkpSY0DwzqQcnxTXgqfdxV5U8AtUGmzEmWU9q9ZyX1p/8W9Rwf6cq/RYLbvf
/IeSV17rz4eabykEj5N7wofU0vtARiLGTUrqIVNTp+zS7mOoggMt4K9iyjmWwciM
HR4kmIngkeeM+rVHPfER1+dbxH9v+9Kj+HAzFVNZHfNwlA2UkM4kW6tmzw96OOye
s9qHGRIZ2LSerrcBXxs2P9WcQbm6e+yeQKxIYEWYgQozOXuYTlyRL1BJR8ImOjVt
pCthn8wTebdGw9U6ZuEoMlb45XXjvWCcKnLHcaWog9NXiB69MXgnJXr/R/T7Z4mM
ZagRfVmoaWztvGr1AI4A558aCMm0iiw0/K+9umJ4oLTYYBYotg6nEOl48qMmco/8
T0nL7YJNISvIpzkwaf3bDQ8p4TAXui3SFU/Z1dK0dZBznelqBEx5GNxneghetYsy
tJXxqIPU0IJCC8XqtaAU31qVRSZu1huioFcx1QZXu45o7u+hEGshSQjSzNqZDcGA
KNDzY6oAPm0uGGqwkEQ3MWMSbUoRa2rVXTM/SvzuyGWVlXsp9EqGV7IUKPB0hyph
RVCxM1wlSmJS4kJLRsTXcM8AJYaQHtc8NiDLt/a9LN7Eml5pj9V8UZbJ/ZTSE0F8
2R7MuQXayLFQewve4/i7qasG5hbsmXrt98kK6kGl96MvG0t0LJeLTsUfrNSOnB1S
Lcg7/jMJW/v/mHCYy7t+7WlX6/VUTBRZWf56ji8cav+2Vv9eXnNlf5QD8fGguDXZ
fwrnJQXv9zBT5e5Ukh93npXNoDIZUhWhx7zkgsVqNKFNN6OGcjAUgIpGG8AE7P4p
vEWDGkl+1zkif6mCpzgndchUWphABjT0FKpmUSGbDwunTf+aJVma6zqVgcmj0PGR
Fp/OmpeUaYtgfBp4XLXHEc4UwssHSpovWsm8/zHZDW6PQnmlH50BsC/8Ycgfq/4S
rKOqonhznGrZcjc3tKz0NA8EFBvtJdxNyELb7Y36SLzzlI3lCbuVPbp7NbJQDn/n
DsMUM/vjgXgNSiVFOhQXkuCb0ER55VVsVs7soD3LVvAwT0OlWX+iKWKQf0vM5ZrN
IhguDt7cMsWPtfWgRLwUNn9JoTMtTHqkhiXPha1HzZE6CqKph+OKZRfSMmPF+wR/
19zcY43aDfORyszGUjWXSIoDU+eOboYJNNQ31CKEnc+MebXnjUqyF6u+qXU6Xzsn
fFPDpyR9v05I2luRNQJz3ep+8egg8PjoSLNFoLeLodwLLhep1CgL9KsC6ufugx3I
Wljqq5NhlmE3A99rY9lcDPxByHAZRPC09M7Kyrq1zTUlpaaQE53UQ7rat8+ylAm/
AWu9uk0kn7pKrWFFFz6p9HuDnO3NMhjTjVqhd0dpufsSlCf5kPlUL/68g5DgWvV8
u1U8jRKe1oIWSqbYy38kGZ8eT814Pwj5AeQbbAoljePZW3vnu7gvQqpy5zpY3R3Y
qXayy3QeQVQ/OMaDY8yAscTTnuYnrvNAfKDednIsu5uxoTbNcVbBKxAlXSuNFSSq
kdUa838lzQe8MoanlSb3pRPbsnqvV/tMDIH92j27eCN7g7A57yh9tS1s0ZE5HTls
P/mpH3Xh+0SuDyFF/p+hHTBDBO19iQweo1s/rX51aBp6h4JsRZiIjAaMNKGRVLsy
frg1ATVnY+5Ur9rsKn/RuVmELqgFXn+bvgVRvhFUhOvZsNQnKEEzhR4fWoVrnDnz
4L0wuv1Pd+D6wQ0/byrv2ubLWPh4+Rqj8nQJpt6n4CiP58FYJh6E9Quiap1KzgqX
mebWru5u22RSfQty4nZh8HJW6Ckq5LTGWMYDn32NQJxZX7TMcWcQp7YWZFKjfHNv
9rUss+/8aDpKQd6kMW5lxVKNndnTEWNtoExbhGvooOUANo7lFjPykQRAo/3ICns0
a7quPary36G0I0oPTHm1Hp5LWdgp77asO2CS1O3cA0hExhvpZAAem1sEDy4pksjP
DU285hfw+dGtf/odCeBhx+DWpdg7/p4iQVI2rm3figlBf0vr+Wz5R9livzM3eK5L
t7ICa2JI6nr1/1SJyrDJxca8LMSxHEBbStpuVC2/m2qqvcZz3XMZnKsYS6zt/4wm
9LQWZkPjAQuzmZzXMjdEzoBTSekut/uWUjZjPtqXUwTdSuae3g5sxz/9ZJ73Pyqh
/f4ceZJYqkePtoDRueYQSuNVe1JQrm/lW4VGajUOaG71f9O7h8zM/yGCjY9U3lpc
u4XJt28MLeLF+/DiGfABP28rxXtzIBkr6BRZE/LNEZ5a0dDcevfxGs6hbJ2xGttp
WyrJJrXidD0AXJZ+bfLdQkD6HfkrfIKecDX3kEhRQD4CJRkjUzh+LOkoOViK2HoG
la0Hw47rizDrGbM8Q9cwSRjRDJNTJlDo8gTL7vDSMD2XphwJ5xGUCZSZh6B4THp6
/ZXZk70+89hTQzT2OjFCcsn5AW89o67tgC+/Yb6t3kUrDQop3FwgiLfDwono+3xl
U256kzCHtRy00Um8jt0rwaIuEZ6bN+TEW7cF/VLEgEcqNz/O8m9o6ecVNhcjRKJk
gxqY/XwQ53OX5bGxUnbJr+xpLEiEEuMLjROP8eN/PM0BTwA5CDAuWoK6WDWYG0tn
1Bv9zqFTyUW3tyPFCZcxiAYJaPi/5/Ijfhs58UNUjwaomH8uI7SjsEoaKyWhs1Ee
RExQYkNTRf8yDJw4FP36rkIKEtGES3C5u9H4Vc9H+dRIXDHE8di+guAvMgecbrUq
r4niXLB+hVeNbDVACJ/uBr+/TTEcibXAt2GiaSBUzezEmIvQFzW8S+oi9W6M7h08
hfbaZE5Fo087sHckuCTztKPlUhibEwtAB66yPgQP9u7SsEacAVgQyVBV9gdmDXUx
0kMDlxzlc/eJz5JGNr+vcXhnzLMSqHzmRxZtpJs+wsWMdkPCZq/VrGOc3jc14Uvl
7m5XfCe0NImFn6E1wlmUGIhJ75vhIgVEUi2W/YkBOYnOqKNGo8r/4DOgK2eArrUe
MrPSRgJlMfBPXsRht9cSD/WJoKq9a+lTliyDYZAvArk7YGtqiOhBoWb4i9Nl+Myo
fReOi6Y3cJPsrRXc6S6c7fiCUHhOreMnYrir1bWGSZaxCCYYcrst99DS4VfeNC3A
e1pywRhOCADFPJ7/9+eYxQNb7hBZ056InbchALRXABhr7l/J7oWCOeye4oSzdT38
C0M5mQcgaQmDNXMQ2A/l0B+u5/DG7o3BQv2brb5QpducLRu8MqXnnu/IxWiwHpsR
9PW4u+RjsznYV+xgHnH1sxN4SSFWU2oPheDLLNknFfN5t3jK8B80/J5jhbNpZgbF
tUeZdxbqaCF4eVdv5kaQu27eS9tI3y8Qn161ZFIAAzi3wZm7HMVuW0pHNsIU1x/T
FTw0rehnyd7X3921hkNOOozX3NXYdoHdDZ40ReHdS81Sqpce2+f9XsNoYcfwrzYa
fHrt08pxaJBIfSpH7ii6psWdx4LKFaBt3XUoe7XPL0zOY4qUd1NGMteXPOgkjKaA
VwKjN+ThegWj8eWB0u00OR1U85r2VUVVmobQRFzQJfo6SMlpUF2hj6IancCzd0EQ
0Xf/34FePThpZEY0r/cwtLYNsGM0JPJAHg3Nc1AJ/4Nm2x/rA/SYi75ir8v8FcFq
bsKCwxT8oW/5JsgQL8fGl02Hz8AX7Q7IsAOyV2vAl0ltUeusIZHXwiozzAqJyXPF
5FdW3K4M4wewJeoM3+m26XMfzOQLAj6pgCoFNVHl9H7wuCwHPHaowCGADEkKi7yh
falrZ8RyBxZxVvc7eK9nhUFOY/Pjc5Ow3W0j0yo1PYQZXNrCH/De/hEUDM+2L6lk
nS6CsYKwj9ki+EJPBh5e1uY3YXTLwnt72/YjjyIRfxsviBmTfLF9YJJNVBj4rhRQ
XN96ukKNEpJ3jIatv5WEYghTHgRQjO4AHUWPrRrI0NBwKRU0KdMF+5pGxjl/R1Mo
yPHiQjhDfdKeF+jPaiIQSsHhDHfXye+x5BF4MgrRLwo7ynjJWlZ9fnxLndv2NAQ4
G5ToYOV8dXtVLjJG0I3FXXi9mCiJW7KtSd3yjkX3WOAZKi0031IkCqbG5Hewe+a8
faj7/GF1YUcu2W/nwQcfng8kKoBrP5AbWR0/gdCUc32k/CoRcGj+63WU4TO20kPD
/7j3KVCvkLrGbN9TGEiBZ8oXpbe37ehywofvkuSdEfjkY/3Os4pVvWWwbsv7+Nog
94kCvyjzspVzw4gcmOpRZC1e7ixCDB3xMq5FNiy5gmyqNfTaG26acTPXHM7+mcNx
QDIyDgJX0nMi1aQZQQM1ixxqSLGgnsFMwXCvmU2ctnhd5+XAPBsB09RPpXQu0IEQ
FErTCc4aNFXsUrjSUJJXDc7A4M3GJhUIXQ3YgMxwTrzVMaMnIGaFBluRIRrYLYEx
G1kcAb8wgFo59lEelBdVXAwhPaHH2n/qjpI2uUfhvu/sSxXsbcg+3WuFColcLln8
A0S6WdSeVRyMLJ7VlWLyu+nLkfBJZQ5STw/wEmppcUv+IwXOXg3l6t8gUHzM4p/I
PbktY5yCo65Gd49X0Tju9r1/7inV/1fJBPVI+a+EyXcqkWk+sjWMw3yWrDBgIy36
vQr9pnBwKv2ZWlb6iN2JxnNthSn+I090LwXdJPyUNIt6JZN5aL7qoDAPR/8W/4VV
oCpmCR0tOKy3QPK7R5QnXfE210Aui0GZ0s8ZY8AHGdtBDs2Nhz7Lm6Fl8rxVRNp6
E3V0Ial+AtYertoFeiJ7wWVD6oOe7xwyusAY8CQy7uMQKoOAJrcWtED0re3vks7E
3mJpfMuLqzX5oeYcWKf6QEGP6N98z2r//2wgAFjlXQV9xNSRpUsHpnZapyjtM6aN
h2iG+2YudZ8Ht2PqUI3Kskc+VlSEssZHNDspcO7sCTSe1UTSKN0MXoMcPfR0ptKk
aelTGq8jJ46hCCN9DJknQC9Ut2Qhp/HRAh0d5IYnhqcLi1LL1TCiORLPXgpmpVGj
5cxoIXCevi+7x2/jdnyCmZKIPprfLhaPjWteHPgvPd5l9v3Qbr/6L5xNeCfcc7dO
zJccZnQmjstw16xqRZGOQCYetrVwVZT1eLZppnZhlPMEv/IKtfh/tLNRQHhe7IDQ
vIZ6/7wi4Roiyd/K/d0VTaqasKnZ8SYyryVEZbvSjg+m/Eh3eNs0jx2amIXjC2ge
JgWlRn6xMSCmBiFRPipjWaQryMnPIe+88dlaECZ6VlUUITbq3Sewrap9Ks4whbWl
+Yn3jlSgvD19QkN2Ksb68FDZqRdzY3M1fW9zFawMqE1Zf4SGq1ZgyXzMERju+fFS
+90h3KYWaL5C8TLbaZEtrAdURZTePpbDfxwob44AGagckVaTH2o96f22/JsgjBMK
oCNyyYprkyX37PtP+UYHgcCsogtJpOFF0+vtGKVil57YRgsHQaAw8AVoomFHYMTC
tx1j8kqRE9KtKV5p5ia77Q/QYtncSoEjBuuFtUeE3GVxlEyHEPGPXUPlsfob8POn
e1UGzSBNJANziJx520uAA06NzEbxp2vZVYl+n+NU27fNRnEpeL2TkdVUSTKmtpcV
ZbbzuMrn72P6YWQhisbQaOhJ+5HdWdLwS42kcRmJ2F/NGmZ2prnCiD83iNPFFkQM
NRe/XzTxEA9CnQrNgYNy9Y5FA3nrHcnmBQVq/PMOuRvI/to7PFpL0cVeFYKuvCjN
FoDWQ95WVeaIxU1Z3g3UO1Z3VUAy9A2P5goqhQf4qjMmRop1r8Oi0WOd5CuIC8vl
2uoeIFqW4BxGEMhbweA4hj+e1kdyPf9HVsnyFh9AkHyuyTQUZXF5qdLcZBboeUbR
coMAMUms5DmzRnTBnT6ZT0yhU/JVRSdXOqjtE71VpqiLe50ydvp0/SUJRtcfqvsl
ysUDF0wL7+0OFoEVq1A1m8NDjjVkZ72OozS1T3zYi4BfPKeGuiyHYJun0pQch177
5yzogD7RakFxqoSpTllRonVL8erh+/JGTrVyLula3I/c3pEXKVR1yVX+r/nz70cs
IWQUMBTGyekje1cNPpIzHudX6ZO4ZPkLOsOQRc5bcSaw9RKctxc5uEdhCGGni20O
t7/y4SjPYt1Pl/jhu/yZ0F/azEGP0KYIVN6Bi42AeZ5/ryRBSN3msh+TstS2VlqX
1kuNROa+Dlsel6eJlpMFdVHFCEpQDm6z9Q4je9X0lgOJcwPI8xjfq3Pkdf9uReio
COI9wJYs74Gy6juTD3+0RWZUCK/xgsorz+QQ+hyTm687B1cll9UsFEt1rcEP3qoH
cqTLXACmq5LYwiIUIZbRKT21pVDbaj2/T+jJNrajEIJyV0X+ENgtzzhPozRo5dye
9eg2czk/GUFgsnRC03uYWA/ZLaqsSNs845c04zNK9pVCuQDpGmbQ8iecIMq8K6AG
FvvAUI2Qr2tFMrRMa3MUUX7HSXhtuDJ2i2X0VfWvNkZn7xXkKsPFCT74EO+w/QGu
MjHOxEZXSZyptHyPihySMa6pyUqWjOOm8BqJEXmRSmLKlZ5e89ExXs8LVfBHRWqA
48clko3RXuG0upB6hzkpopMJOJIqndZMZOd0dqXOcnEj32q2D4XWL3N4uj/pOcMg
MfE5ypQiRQ+D43s/aSSBpJHq3JPhyfNQLJz9XRfjoA7/jc1H0fY0iicNNAVNg4Bc
f+yElsCGQRN0LSsjdbKSoBpGZ3JXRb6NZMmaqVjoHKtIQNq2atKQAb/WfD5pzUP0
lnz+xojHFiUOEA2jZ+4tNxiDIBiqBkY63BjXYViUdXhXTT/iDxQ9+gVSDm5DhGhF
rAQSi6ElwZ2h1F/0GvxgjjxwH0/R29nTeBu4DEHs6lacqPXwyhzGh7bMEHMNMjM1
9cxPf+SEuswUYUAf55EIWit7vc0pGqwP+1+zajRJU33Hb4xa+QsgG9e3IFnLwusV
hVP9HObrpFXUp9SXc0mqQBQ5ppGbN7g+NzNuF8AjGFw4pE0GYXq++B2ahWrUQYtA
oG/CsJQggy+NG/2I52pOmsALoqlZMj7RIjWjFU6NXztnnXhcDfqCms322/TWG8Ts
gcPTwtxVuzAC/K3M5mBoshEEsCQvmPTVRkL1RvV4oWfkAuLG2OlDDLaUa8IfMfTR
opOWyxxeDv1gmoqkjOFzjSnv1glWttpY29gQk205qSLcuBdSN1OYbknPOGBHn5mY
6x50cZYwxQGq+Yt4JGDpGDmH/9jh6KNY85d0cgxnjocaZflhuF9FTWiISxq1G+wm
lxr3QQGuToRJ2RcRTnwuqx+KE2T3wCSRNMPA52Tw4lHI2H3KfKAQUKUk5M+A78hn
jzRmKg1qYUmBpT3Nt24eYDCcjj+DVXCLbLLL6w5ZD0nt4BwYPc7fGuztr+TBAkxk
BoXXtEa3fUIZhkgo3C/JerXzPIeNk4p4iyXUC4UIGOURy7zHdB+GfNrKVY4IWqeo
aJXUi32ASDJinAsGWeskRlRoGp4WEDgPgxzt0+rMcz2MAIw9XDMAFMMfdAZUfO9Y
wSJcv7WIzrS8CSbLLOwzLauDCBPESG/pjc6X6M3Quv0p0zI64Y3kTkwWJzQ4Fkh8
rdGBsI56z5nYfTLk1zGBK8WnRhU+9EGX3itQ6e8lGJG/Z1zRgIrOU+ug1KAhIML2
07pupugs9P0jUCGeN74RewHddP9YvkowJ5C5BqEEnb/4zY1+IEaFHX7TtWnKj81s
952fSCQ9p8BWL/EB9CqfzrMLo9izgt07PF5S7KywQHevPJx4kJ0aC5KO+pq3+gGz
PzmQRifO2rQXjB9+5Di4s86JN/K/9y4V9k7q8LfB2CHO8d1THXSw2PqLo2NB1Ikj
is/jzvIrWAEaA9+aGOLy00Ud6pP9JvHXJKitc0detPeI+33V0Xt6hsOiOdQl+WqG
O2Ya50wBlHBECi+PwFPfL95x0Z4jrtbb97W9Ut9bd5TWVS+NWC7lyDTYNmzWCANe
CRVfNY1P6Njp0BWfLsEDVRrbJgYyrasn2VCF7ko91kKn963l0+edNjHUnq/7c/kI
0GIEFXW4+hpTNJ6qHkXHdKIJYZl6YlQXWkpOkpg5ZhqtoUpu1QRF8ljRdUR+dY5w
46MdT8rbxHXgTdFACsVLUBrPVtIdq5J5iu86DP9UV5p9KSHqRVgl9b3xxtHkeU0c
ZBtu4xEugDvNFULVVr02cyl5t/HGA3y/J3M87E5al5OR/KrCdK6MievXvOuwNaaq
f2zXpJjdj8/JMRP4HYbYndwunopxb7+ScHJPCs9f+oJUttMXgLLoCAHFyJRm/yTm
WPrruu8w9UPhZmD1qZk+/wD46gKxzt95xfsWH7fT9aBegcnAI8cbp4hgX1/EdEOk
xwpdbZRtP88WngHmDkcNB8hhrrGALN9JtzYtPxfS3ZMh68Ian8bOAxAzUze3Qxzs
Al1vD4vD8QfF5P2ZuFbXzSLXz0etvyVWOpj4PEbNGOdAievmYdyAqMt30PybYVvu
5BmBC9IeAqkMpL2FiEFEsWisxb1owr/G6T0koLIlWyAJlYEIP5RzcMB2XVDGJm49
uvzWY7RHKwuzo1h+/zCcgDl4BNm/kpqJkv5y+i9A2wUdAnw8fp3tA+aj2aNh9wjh
ikWBQjzVliCtPBivu88KWFL4YmVpID2oMGIU7kQS0HXOlmTEY9idWWaTyJinAtUj
G6ys9Dx7JCBmLdplvHUYTN1gRPlKWUgdg5VX9FGBBSgCqIveWBKabXrWtAi4LvFy
gKL2nJ7WaP1Zfe4KYPErqoblgSTtLHqB/xTYXHtoUBbb4cxr7H7HdwflOgV6ZXVB
dLJGERx7RP9h4KOhGCA3so+9Vbdy2bkjAdgVlR/cA4ixvRBlUJZy0QmEaS08xcWj
SdzU0WNGXfkGYm09RGYdaFsrKhu4PINT0BQ3msIrik+isRyeJ32kXRMcBSXa+ToW
ui+dGmSoc6jVSEGCSlGOUFJLJk5Xn4sBwxmOvLOTOb/D0t2qm8N7OMdpIL1VNWr0
3f0+1xEHMxdvX5kdU/Mn6AaVm3UmVf1eP8ZB3CKO1ECymnlOulV4/EXBaRekZiL7
jnLUiWA5KkrNrxMzFYdo9u7JkeybOOZRt7bMQ9iRBpHxlOBcsgZdgHWrVBjEiu5q
Io8hT7pkGV3vyyQ/yen5W6aykUcrbb1FLbWLIOtE0nqlo+WlpYJjd4CH7XKHyAE/
e2/DyGItilavxNv0+UJlNSgkB+gGA+xs0uJ90VdhYHkuN/eJnhf4tBFo0Ahf3IFi
Xx0BtaQTv50hVhPtZzWgKZb9UNvxn6Dv+Y+yRSWtOubPylUHjhviOVf7F2vVLXrm
rnVusUUwncKxUeeqvxZ09zI0uhsdc3fpQcjER1+P1MwE993FZ6eFe/NuQY++Na3d
9+hmHIFOWxG2A+ctjhSE0N2k0/8nzNNcaXDCOiK5nPgz0hVWMLD/cwcHnPvxnBgd
H8olZr58uirYEWfB1QZg6T377bEGlnqBoR3p8NnkqMRTVn53RHv+JxTW6afuXpFC
PhiQjAtbepBalIiUU0zsM38v3u4YfrUPaZQBk8q5gl8xhDX80GvKx5Nd0RhHmsV0
bsBiQX+smN2EPgiOY0pYS3KzRmMEw97kvImjT6qB2FqGx7evC4+VoZfIryausnrz
wCctprXs4DLLK1Luo6vjAvUVBrJAZtyGj7gYV+AaOMdHrPeSRuxsUFmfmqkkeaXL
2KDqB3+IOINtv+nceUW9+QIY+SoqXvzK6vU9vH8lmwTqlXvUS90iezuqYE98tYXa
XZglWo98IFOJEkKim14N8KDPpGsKITabwXKnHOJHemcHyBFJW9VPLoLG93K02zjF
tgr4v9x2E0jSfWOk8ZHIf0iZrbNUO3CwXuhVRJetouo/jfmBeR5IQXxOJRtp/kUK
CMZiVr9pt2BCJYWdQ+6QRc3I04mO5q16t0LmXC7DTK2Avqi5WCIOcRDKGv+HiZJ8
YkYCn3U+QG+Sh4PIG2OUZlrg21r+Sq+Q0YZsOItsPSQob5Mohsabx0U1UmZcDRx/
rSnrIyLvkYGG21qI8EaAdsqKez/BvZVS66bnlYT25aJkCFzipMNeQtrE2X/Q+R1L
VNLoaaEbA6eYV36NyH+N0oC63LB8bllq2kxL6RpkrH05bxw4QFVbCwZmxneYSQwB
NM7ziYFzSj567CdWImF3fe88cNGlUeE0ms3IJ4zQi3tPm35lLjlEKmP8xSRQhNka
yh5NY2CQ8WU7qdpCL8kQB5Xr4SvxFHDmVJ9U8d+mJa+90/mF6gj+0YCiWPbsJbZL
GhPZaioVcbwEUC1DsOaaBrP8H3GwrUZeZuM6MD8ZRfwBWXuVLjXF12oLLOfqe9Dh
W5qXXOEWNhwlEa9NA3HODf3bsVWzkdQzWV81qBXs4ORyfq3TrcseB324pgs3CBc8
5moui5IESOS6mnxsHlcIckIOtaVfWl9QRRvVdKktVFPSmLZ1xNM1Z29ZQA2Ool1j
tR+tMfVsR5YMN6IqPXkimdihwSZP1ODR6T6fIeWnKFUsRWybG2SYjonPRWTzPNtc
F2UBMrq8tq2UdFryanoJciVykugUKNv79d2juP2FtK6aDGGKb8fpt+UnGbNgtwsW
KYmNi/U6mDpF35FtFYHk3hLKfuLIBTbkINUxil4rMuTVjjBT840amcfujerSfxOx
6FDzR4y6jZeGGGHbTIsRREtpVPEOpFwsqmvmPG1CIfREZgx1jQpBWCO4mzxrIEhG
mKwA7yBq0b+VXvIOyB/6dCWxlwbOI2gBCwFCNeLFKr1av52RMKWRxArT8gKfHVY+
UX9VB2NLmB5eIovaoCXLRwbS2V+1sgyrlLF0WmxdRMvUMDaHf6ISHqw5ELl6t4KO
jMTmCnuu4qN/D3KfNmfmYCcVOnuhJS57KN/sovEm+atE4GdKtGprXjZNAV669cap
PX1K6DHSNuOlmkl8EvIKz8CSOgrwbsJ53+JmU+X/EUHpOJBtDK4PyK5hHkyeSHBP
3V+8duWXEhFXM49PIgdoIAdh/Hqyu9uExe7nmbOdSG3/QU1CFE3CcGPwyFS2jHmO
URwdphvVwwjRJJUZhjXFTI1EUqHn/9cUak1V2jipNrYGXPiKsAMZb4khGRRvcM/P
AcuE6yLDOi10x8nmMrAb5e9RZT7NWC1HJBHhTTMZ7RKiXTEAaqYWNOduHEm3ztRA
TZdGRcD/ZKHa8KnEXXSL2H2BAGGQaTcH+I7l6WwE30b5CKwEflMO/Ng4eW3fC7cX
JkZxQKxBb2hRN3U5pyYtgkIqx57NVUm97hhm+tOAqTAdqFlM/YIN2DBfQxilpAvP
MuS2tb8EXK6pfNEa7xQqieMQLer791+2n5ExYW3elmft4CFnC1pCNGD28z0OqQKr
rjxGnbD0W3OwPVbCBDdoNaU8FMYYLdPmx75YRw/8ocsEGf7d1RJEYxDANhOj4CUE
D6sAX+YF9Iqjzq5XljT0nExiPkEhfa+bsrAUPxJh8JloJ+XaUOvWw5PiSRP2VVvO
WK71IQjfpUyXg54K0qHrYL33ACcE7/IOgq5jzmmkagaunG6gZKsFi/O+N08aOaIQ
4kOaDkfumUpySemH+4UK2aOiRRxaIPvblsjN+ipmF5t/iyQ7Im+TpBqdVcufXSjq
cJCbNiFqTLUbo4o9x7FEYlc7Ml90oYoEnsXRjbfYzVnkqkImdmf3nFWe7Xxdn6b6
hQ/xcJKnC0hG7+nAVCerup1+Zea2geu6EgUEApJgahSBAYArrtdE6GXmgsQpDhyT
7gNbRW427fAUoVApaCK5TC9oq91NL9U8xPtotijBOEGPKGauc/AW9nBQCJh6LPaM
N8OZw+QMZOTQhAq9flJP6ES208SeA8lUTkt7iObCwfo+aKBF5NhoBKu4JvGtI1mh
fo+UlfC9MF17241Sz7DiMdSMqgEun829zPEarT/PyeZ8RGec5QjiMiWZUb4LBZ4t
Oec7REbWrJf6sqlQ9p/l0ceMq4hzIywz6NQ8WV1PSjyFG1IwNOqq3y7suJ623C9g
zMeUfAffNlZC/YSuzgVTv0B2OIUDOXuwZ5juaABtyTWTnCv+WmuiBQ1pX++/Bsj2
ahmVuiMzntK0tbc1H8GJdW1NqL+QeXhHTtqoFcBAyv9U0Sgc2C5X00ILWSrXf8uU
ZSGKV+ak1hPkrBaLBidYNbL/aLB0Rkt3W6u0qs5Q3yMHl1ibYhkAwi8cje+9aiv0
jq+Oizk7v2sQOsW51oMNoLo50AnKVOaamPg4b0HxbsUkAVglZPg2Qib9BHZdt/1Z
CX87pkmTd0Y7NEh6TWrvpK3HM8+bTw/63FP26KWxjM4BZH8P/TzHFhCFf+A6HKcw
QY7+UKtvwuxhQF9c+36GORcSIkR3Ar839TM3s9RA86FjArT7kr9ZIdvQRrQck0/A
5Z5VSipbplzLznLVkMldRxjZtmfa2JrnKwmxq+KbvW0rNZz3GKgFBaVnOOvlFVJs
1/KmUXoTtGDysC97yPzGij4U28sy58boDUGfkMJamZdtAils3JQD3WMIra3kYA7m
dDdaGleHs4lE7zNbcGFuCKAHwXYRPABat9pBSBGDUqi0z5rRdxm8pEZhs5pp36LQ
ZPhlmwRPk21ZAIRb3x0nXLIV/IP6d4rGtjQuh90ew87VmlFRoUxeTLZxKjXEjbMZ
9WesjdorJZorjxOqMowo4SCYbwWx9uYJNOTES0TN8JlOjNK5dgKE5PBcn0LNBFkz
BI8Ccseskxs+Dhx6etHMriaPTapQI6EolH7BKuFD3v02VQ6f5X2+emrL0n6SOEeB
XGVnPriQzwqiV9fohSgDB/gdSxyEHnMUi12XzmI2Tm7pE/if68267HUvVUUe+TcY
jwWJ5B7BFb9yTwhfnyZfUoyz4tTeT05dsFq7SN5laUxkiqZhw/44x1//pBr14FG1
P8TGWC+E9a36TSSnI1dz1Ibt27jiUSyHPHr16Q4PEn2KJhuNVvni2lKYQU2p2Ixf
tykRr2XeyCuUekSVmBs+JuG1lvE/gdOjuV9rPQLvJmEd1rU41jqHNG/rL4al8iQq
PLucgwat8RtNFpw8mWmrNO336dsV0FquVhZDj7+oDT3ayabwk2Ij2THZ5nhNy+d9
H6Auh9wZy8AEIHw9OsHCJertZOwpQCR7xxv89Sno4JDrsHRw/5FNF85vckSOu43g
mzpptFdqU4+U45V86lmIUtpVsvuGvzVfa24bSqgD2rvh7IJkGlCjrTmgzY/+ncSP
YS8k1yiVaC4+ndetAfEgTZgnVZOVZy7GOZV3bcokyDO3Q+ovW3Bhav5i9a/ZnrN1
xFJ3/DFIefHZ+ayBacpXyN2I14EYcKyq0t/fuXJfJwXaWqA4MaMVppbyUvZudYw6
Igbhd1QuYmt3OeyogUR2J8sBEjTXaOyM1UPlPy2Cd5GcGlwKakzermd5uZ+ga7gs
npx40ELW4+52XgdlsAis0kVzXaC4tzQDvlPElO7t4iIxba3B1cc0EM0yGi7xD/uG
nns/lImTFjkxb8/GW/Oz+wuQxNxBfxqtrg4PK9F9+D9LPLTHaCH1ZN7GaU5eMbar
G3B5Tiq3UAUhkmcAknxKnANx5eeJonpuRwG/i1hLnfNOaHLPK0NYmTkg6PQm0fwC
a1EFX4iVz85PyJ60FrXM195+hGwSXGh3FMKR7wqEn+eOhlkh+JiD1du7MR/tMI5Q
WGa6GbzAlcGnMn0x2amOn5TiYo0vzzXZFPGGz+eeqIOXQwLq6TOdmgVb3jMs7DC+
hjjIurUAPNuChW1OJ4Ym3yjMDsmfgDTO01eqy8fuVBtPANK/5hYlLKLhZxbw4QJJ
dAeF6KAQV6Whtl/Hb4BIFHe+M7klGRMioY1pyGqgwzi73rJc2EYQbdbKZAF/6xez
iC/0iB+T3NFCm1elkvZ8ZWG+1Ust3IMNoV6F8+oA1YFFAN2Ef+bb+MG4pvK2hjLr
VlclpxQI+t4xcD9/Fym4IzMqiJEEbgjEuA5Iz96gUdn/a8h8NZRQL4KTy3mQJgD8
JQc0mRu7DNR89/NLHqYzRysLXV7jJcjx54+5upmH8Y8JTANeRkGIYflPSH2yG2lD
kVqNbxU0r7cAqtHDSrjCyT/0mryLo3xtIbk6U3efEjIA239DFkeNKLrGh0l+WdeX
B8CZCK8g7KQme9+xHHMygGtz79W3nt3U7txUKkDYWmsMkdg6gAok9piukEoFXyEH
kL7pwtqrd2Mu1YUB+6RDa1qj8Q0jVhrLhg+CSdag/Umptb/1giWSdb7upgg1ohJu
t+eZF/xB8tWP6grkekYy22NEm2sqRMQHqKt5sLUoPr4a431bMQQCDnunSAt9xwcU
6p0H0Fnft6/TwrRM3BSOR91bU0hDjjiSXHLONoxy3+HT5MSJyPvDV52QbjynzcCX
/7Z6zgZBG1bCkMYi5khtplbcBgdKj9XwVwszxSeBDxrxI1zOyRpZxA5WCZaItb89
b+JftdV6MX63n9S53HGPLQMdQcFhMMXTeeETWylPAb7BsKKp7TW1ONku1QNdJUN+
v3s0ZTiZKHeOc67ocqDpK59/DC7i/1jf4rr3vmKlL2vo0TR8B4kBi7jp/Z8cuigt
e8Az8j09FVPnFn/C9GnmN4+HXxAOAvR/p/doGdo9B6XGTtWhC9jzop2st0wW+pbB
y8hX1z87RRPFaYJXFUXGDJWk5GKwVVcLJzj7ZkBSYsNPh5MZS2rX7vbh3x1X3S/E
oGNbeDcYOV/woDnJ0rcpxBuwSvxj3JFcYYJX6X2aV7WvApfI0W9nj/7YCAWISLL6
NGFAvUzemUgeVawoY+QDXAd43dmcfGB8UWca7r9k0UYkJCvBT362c/swFZlzwB6i
sOgHGuZcSDgJEGDzf6zf85hnc/zIP05+9i58C03zFcftATJjD5aO7A2SKLxCh94u
RIZnp9Ahprf/Hu92UE+NY4wc1G2chGcW57FkaFlx3xuCi+keFqNud3vo0T+OiY4x
8WoMkyxhG5eKTOmZM5FMIzUec9kyoBj71kBdrfaApJXO7kfuio1on8w2fon+sAFT
2LBBmvGt85jCA2EBDXIhk0Hagx2ULGtZDhvi6InwIVX7tcSS9XKJWwzrl55BPRzl
8UH3DpblDpM6VzguF2SghnQpR08Jxb2pF9RilhromEMBflG7JRAhBDMAUoiU1WFN
P0jYL6pnb7yKNug8Ea3KikJ54YS1B+M9vie0lS5mxrH4QdHp29CupJyJ3WBw6RLd
JwFFCgK3Adxq9RUYxUXMcoc9GPG+eCeZJdYoG2KsMipikenteH90kcRDjosBe4/O
7Aa789JKUqUw9/8vmXWoUgiL7+hAyOlFWSYCi4D1jkt5YCU34wU7q1yRyCHqr4Fc
Gmfu0DBYjpB5poJLOaeE7H1G+wMcr7v+HR2G+izgo5m1tmzTmJCRLYE3bYLWGdBe
mVxVvtNzShGR4Y41uywzxHAGmjX3eHEot+hWp8oC9FcHjbKXnEoqHWph3lSKpkx3
g27hJ+2D6Srw/8e0BT6YAMEt4AsxGpcx5cQ88+sUpFEe4AXPMf1Ik3dSwKD4z4kQ
T72XyeZF0bJEq2sT5N2bqO6YO+oWpifbe+H/Y2T7JRMxbz2OCxeufZmDLG8WJeof
1oYLU0xn4uyPPqEakB/xwPKFXTn/EdZN9mFq4OjJcH6c9uCtw5ck056ZvLgaOxZD
8emsLJWM5S3fF4WJhNVBQIzATjOzYKq9DDVsb881+NYenUYbsup9tt2mLxCYPdIu
CJTe9yZF+gKS25plOX8KlUPK2ZCfGMOqeFWHRjymIQnIwtdR2o1ToKd2Y0gpUyEW
XT+K+7MVIz+zL4LHjQHp1NcVKFEurIb7mC1z+QbpV7K7O5/IsSzDHw5Ogrup6BAd
IcdnDmtZq9KqrjfausqY8ZI219z8/CRcvPoGmnA0UiAToZcr4zVAz9FgVvu9cUhl
BfDgHpyuYR6G9DK5rFe3wdD3gZudRhqM2PHyVRohfE7HEI93Zdl5QSMgbwAuYQ6W
d5hAH3TjG+0oc6cIrtXMfACm0p4M7JOxmaAGYnSGlQaJrX7XtTsexcWwE9hkHsEY
UIyMYDD3+gZ+tUo1tqfiBjnDz09SvK+yMC/Wx7VB7Lz1x3Q5Zp9si1Gyb93cE65E
2HA77FkfhoiVjsXHixeHJO4i2YBCQeRG24Ao3fPTMB/3SnFk/bh6pCDTPLkdPtlp
xWq9TS8SdJPQKcyb6q9IaDa9WzCIwXADOG5wQiz57/ZhWpciCj01UezlvyW7yeKh
cp97q4gKLu9Y58Ah7dZcYuTl87lqJ493DSa7hTr6AsT5S3B67koD0XlYNbldiJyG
5itoaE+LFeCxqYlO2iAnBXdVWpcfnE6mzm3wF/DOFcJFyrKsJpQ/jljqVfxJbyY8
zV9JsBvqNbuDXlRjz/5AK7oWj7fUnEZPyRJRBOikhf8/kfP0b3lrcIGoqrK7S1Jc
xl28THMx+8BN8DLg6Q93qRSiOw+OoZP5LuviMT/KV8lOnbivgfru7uT/wK1zcAQA
Yr3ghXdBezS+aHsaXj0kBD00L7aPDd/Y71/vUs17e6Y0uRmmz9p+9ob0W6EL7OBs
idTR5xRgfOaxRG/4ER8XRHCLUZU1aY9XuxiVnoQva2xSkMHtZsxgqAuWDW3xvTNN
9Nb81E+tllLlgPceLgsSzuApYQwUlqn3si796ch83KFbEx+Xygbu5JAmJn4RVU7u
ETx/BCs4pB+UHyFWikjmPJwfbyGp09ySbfcJERxEsdZidCFoSN4qKXT5dVjxNcfG
3Hl/1pPPJl+7BTnkssPMG29kKqxgLPSy4VSQdxX0hCnXnuLwIfM2SYGzW13FTSp3
kIw1qw5N/b54NTtiV89lkv38pJ0u1kreikrINhBNZVN8r0h+ypfbKRr9KmsCxI3y
W4tW4JGYVwTXn1Ll2lqXynldPMzmQ8+9pDy3d+Y0AC4UKsOnM3yUamMFPIip5liJ
R40jSOJuVCDkNuhn7H3iqVyqCKumkxWgEclyQOuHrYTpmKjNVuSz4IVUj1Jcs4GV
bEInr+a8KiDBRuTvKXxom3DGKVLWLK0857mWKIF0Ic+1X01NE2eJuEcCqItaGkU6
WNHFVLrxPPUOmhmLDB9wFY12e77S++AmnOteuwO+ot9OjFG08KCm2A2Ep3DSL8J4
OkMqKXmhJdT4BdVhB4gSiA+0GqXitXgNJVzXas1DJwOZoUAE1TMV82fcwn87kRHQ
U6tcipCTVfmVfgpPLYJPkc5hVqmm0BYSQ1sT3ptgSLMmvT3gbWe5+0oJoklVId4j
5ldimV0KvOjd0oTNXbovaq6pRT95vJ5l9Mg8aCu72C7kifmDREdTpoxpiCf/59Xq
/ONVqEJlcXpVZjVwBOyHvz+HL85GwTqxjcQ9hOHc6yqBzSrkq2vztWcKPp4WvlHO
AnoE/QY9dTtBK7Ah62FHIBhBsKfHm40fcW+FyuxysE+Yu/FHkwYUdJkqJigWoGZ5
Mb/hWR9KC1OKJEG0fnBIwCqBoX+NSdRcY9GGnguj0Eofp6mAERlJl4TXcHNPC712
Wkwzf97MPMFl7xPQGlpG5xYPEyQ37ybOxyoc8IBnGkhwtHbPsdYIK4PtW9eifI59
o06/gvvi7RabjspBJn8apj+XdXEY7iJjULLj+cWnRNmtAcAW2q6VScnzi5o+N3HK
4VnWCfOtqcdCZD2Bi6+ozzI8Iz4/iEAS4FWKtKtJcg3FxSODWoseEhp56272UtD3
0kBQ6l+HseH96YOjD58wUtBMTssaezjU0xNWyDM8FMx4LJX/96VqDY1Fd474HEgO
ko25y9rW6H25JbC1GD/lB4pDuEkuQ5uCqCppgGNpQL7sGJWCmLWJOUkWbBqsmlQs
UxHOL4c98gtIh3y+rt/3s1iHgl6+dRjSoX9VTyLVNwlRvZBd8kMIxwY3LvHWa8/O
L4YDDyFaiyeQ0X6PBrcXokDoZXOHlNTIpxmXx+ajIj9Xr0Mz2n7kUMy0m8KWbVEg
eak+/X+WlYh+Yv0VYlNMXCGeVMNDimNO+Q984M1zsCXMOIY+yFnamfM4Y6iVN80z
/ipHL7T7uU2DVqrNED2PRCgOUYDoFWhWtx0MrfPiMhjhEnG2JunTNms4+fupcLr3
XATJYrOWAsr3FxKoIMFnNf1JdciAos7iGIiIgfg7z4KM6nCp5HJbNAutG4kTdKTV
noFesIiWaXlW2bQM7CC7UcUmjHozjjBf28wDSfXiB3F0NLbhIC1q9r5MJZ5+t6X6
DFUMkMLu1EiXHoqqDklXt2qMs4MCZnWDo6/IcrBBA4Ok7PSeMa/I3IvbSHHDnQuT
5Nv3CKvbB26dKRi8vBzsrNb3H47rOSjbosgUe/7qfmT/t3SyZXUerrhGzQAGSaiV
szmiE/Rw7YrfsDAKKLpQsdG0+pZJCURZPvY3D4Ifw5DisqbbnKj94OJAIUALWWEQ
UzmtB1GWq1wAp06+aR0DZ/CJOUP1MOROcLl3gx87NSKfXHF41TKugenW+gXE2C2l
aZ/7AUQl3DBERMOf4YkNxur8Kk9ba/+YYpL4PDLBU4ci/WayuD14G4Ls4sNGNevY
zvB+USFyFgVxU4YrCB2gBxwAkI86vNS79BesDIl7KHKX8+lZlGkjpJJ2yo8xx4Ik
fmZR1DFsP7Jc+IajHrudXhw+ksxVbvhtXfeNXK8eiDgHgrZWQEYjgN5kvbBnvNJd
632x+myMxsNVHHP775z8V0cTzypxTMRGoL+MRZAhOKYDep32I0TXwh0julEGaRg7
Ra9nIh/+Ncqy2ujYWqZED/FKEPxPPorX6vUjDqYTavVdCEuAauqgznVb9+hZoIeC
CvErHWlKNW5Tj2rK78s3qBBMXjIYv+jNxjRNXty1i1Q7JwyMBXaxHHLkI9Y1pEvv
KQLoJP1XIjsqFVn08GQUBl92Mi9YvDozdEHk9aiCOVUFXRHfr6yybntQzL5gc9d1
J1FgNsoPKm2inAVFdBG8W7W5kRRAkhS2geTYIwMDXaH6rVxFKbunIkVLKyQKaGqI
0LyzxwICeg1Fnz2zHM312qzrvAiGkuAizO69ZiciC50atCzsr+V8uouNg+WPgS4j
qOUcxRRuU07J4ClXcJcVBseXdMTrdOrfVWDTWgX08JdAjz61u3Xi+R5K69JSwZrs
iQxt8Q/zJvsuq467d1YAVH6xH8/1aYmXZuZHXpe2xL2iaVa1fxf2zMKfUgLPwcKl
2ALiC9Gs9lLii2y6DeR5wxrj90SkJEPweZFkw1nb2zGebR1fUW987CNkQUzG/7Gt
P2aPrRPr8VXAFGJOGoCq9ov6W6hCudAc1yCyNNIm8P1qLW7zQjnFRvSonszacLhR
s9L+9aRV881zp9Cpe9HCT2Fh7V6Gzm9MlW6EhH2dTqBYB549GXvc7R+4FRO925vL
vUzEJZLUl8jbvVkW7PW5bn9m0xuojrHzGI5M1Nh/PZz2uqGXJFpNqf2tZsC4J4oM
OU1mB+v7HtItyUZQC9sDh6u2zwym0LBE08ynEAlGIm9HKweLShBy3k/yPhp5UxR0
MtZpPMjXvXEbcigR7BYP1QXm/TmYBKbWVciz0/j/3rfu5JDJ+uGA0mEjIlk/xrRt
jn+L2q00KabbHe/MauUs5ijSrdkK0MvNvH/VabJ1+SK3mxml/z1DlCINpihxdMUo
pPhtRE5DO1SewnBm2I9sNzrrp5TybCcVRSTZvwn6kPXHAenEZsNc7Wi/PBn/+4er
hEFiTKooFyIoDn7IadcbjKx2Jq23LZ9UqSWqKa7gCfPEkYRKde0kOZ/hhRG87cjt
Adl1jtJ9Bl3jgXeubJd9+9N2sYK/TX13YYu2o+BR00ua/Wt4OQo46fHFEJ5DYQ/m
FZw7fUiv8WZsfD5pkNadFRvNc38L0jxuj7HYWMVrGgFjQerWXmDXGD9C9uBfbdbL
yH8h7pu402fs7sWOL1QYg77ETIDcK6y+KFpFBKvQgxc/nYjfqMsNLekhWBPTF9t2
cIOmd1RFxmoVyczB0VEdArQj4tLeNxurYlDr6It9/ed1XxjatNGunXbnB7PzyvfK
5KQJfBrxVrMrZEsVgWqqud4LlbUcHco+lSd1dIrWUqchG4A4a5AyuGyN48ixykTp
1uH1TtdO8OIAoVaT9JruH6UFGS9bASNN+qnob2giSHDfiw20e/aK5kdnDHthCVjz
rTj/YMhjXcGhxhlOzTev+Nu4syX0b1aXeDibVKhR8CG3rS2ZPuoqkLUraSD4Kiyr
NN7yy6ScAV4lpucAZI+55INIWK210uSqn5YhrTOZqKEPrp8qov58Qj1unAD2CNZw
ITD7vAPYLdJbFg4wgofaIcryZ1p9uGip27FOlrKz0bLeo51kNMTZ39D3B2zlepCB
q0XHuJ8Rj6NEpHbXzrnn4yp+DpjllGryiwQVoQHMEDgWWB41F7Nyr0s2Fj9YNfvF
Qd+qtQcjTmNume5RZDz8LUgFL1DZtTCCXLreliptwdrO90qkR9JnMWH2UVbpUuwO
wFf+irzYlqYZi4lgIGipZbV8FLzwoa1FEXGpbJv/E7D507GRe004w06UquLtNxl4
eWcxx8wevgcp1P9SaApRIz46/lIfU8AiPXSkEycCqnRD8fcNeQQCM3ptumfV4jrl
MA6fdfcqxp0yv7hgBIofiBRSxo/N5WQeELY0lqXSHKaxoJAslouOK2K9ZbLzuAGt
rwlV1w+2173eQzQnlZh0B0giC9Ylf4wCsT6eNJ/fFoDtWEPiZ+OlmWvy5GASorAO
vN2ocjREY2okPIAjl3YjR39fdlthN3bdQnGGdGmPAHXBHPvJMX2SJ4Ktz00KzooZ
FWs6z3yucHPw22ZGd0DgrezcH0aqf8k6Zoms0EVZHZ7/bMDQIPB7iGWjO7Qm5zS7
38KOkz+HavZtcEupCiOEQkBWx3YvtTpXgPy4lDgd7w3bIWRaBwcxxI5lyliraEfQ
c80oiTIy5LRTLEUQ1c2KktHC3Dtn0RnZXpWDD17WGm49pZE+HP4EmEQbWeUapk72
2JEPHdBkoBaXrBmWyscpXzUDWAy6/uK9K1oKA/OLZDhWXOYVuflmRcVSH3A9xLUr
T5g3rHhzr/cN1YLYhJc2p2JwYrC5IJJ+8zK8UA0YotxgWCeJDY0mDTEZ5HrQr1sA
vl/F54ngKeLeHJeUA/9JZZcHCcxByJkG/kaE5Muo6jOmod72RKmdyLpfHEA8O2MS
4iIMnDkMFU/7GKEnkY5km6TRwfz+uwNSEuXzFSqCmjeMDYXiCw8lEvKuhPczsPnl
5u6U+Q2xGlASZKlA/18qT7r9pfvnpU3eLDnWhDqhMuzy+ypXCUvYWrwXEKtFfc/c
0nQP2eHKdvZMCGkyFbn6D/XguLGEx3vHn8PNA50UOB/xUxvWu/YAQgy0JWTmgaxi
JGT0zNlSxX7jk5Jx2nSf1Wnj/79UkND7zU3UhQWShga2RmO5cetSYbpYXmHNM3o8
pdVpENUNvldh/lnga2E3ZTfdxHte5oij399C7F/opntuNWSuBx2aDUG/v9h9oWBk
AXUDxJhxNOOA/dtYaA41mw+9swGYoWXa3ubx6OVMn/t5f8rUDeVvWk0luvYubBWF
7cwEBcQfU5YRc3FGBZ8PDKRwRAb1x6OES7JcyT//QyohLANcgt2kjikSw9ptY/XV
q78sy9Ic8Pfig+0Y9iB5U3yW3UK9PkxqtYD37K2zN4pg3R+xmhZLsvG5LUW27kHy
Mvuozr7APmh8e6FndBQximUp/UQuynfRliDJMUYZUjfUtfxwVKGSkNSystqqK2JJ
WVFJxzZyOei/mSZ3dfJL49rV+3S/HBwY7g1IUiL7I6gp+kJruX5cJsyqe9DDQ/sZ
QyA3Hj1p16gmcg9CDdFD4lVM7HvWd3eHcrpmrPBM0CXl29yItwCAKEg5uUrxIU5X
gFxLnwcFDYmRKSW/sQHjIADeEVEQZqc/luLziaHIfxfyzBpiSiASBJHA6hrFeQ54
DRlslrSGpFMxMM6QD75OK3CZpOmJRvwUKHEFZZkIIkdt9JQzJ469xed3+GJgFcWv
HrSW+6TilF4ivouEYyWxUUp+MicY9nJ/aew4m5Kj3Abr6BEkkCxXPKm6Gk+Ldl8G
334Sqiyb1ZDX5qdjpF+8id++7L4b64AsKVylrueiQThOxM9AjQKA4EDKOecvnH8Q
ja8nywDm6lqgfatlPnW6u71lPHJNjQSiIcJODV5CaQaHLxWx/3aIc9zM5mPvzncU
rWzFAdL/eZnAEftAaEe2QJach4S7Vc7zKjZq4JiQ/COGHbHGYSYImDmTrgjsiPVv
1oOv8lYTLlPTnw+WVVHwUzAx9KFZaVBOUx0mNIfSOPgBGsuh3h3GNtxkPEmlfBFQ
EnUlcuXt8G4Se0vyNXRz78jUApMXuANe1Vanij5dIRnWv+O46MEm/0GgodfCe5Zu
3CEARvkadQ+Y2wbzMDMxxRhoaS1zl9irSMHTLDJV0fkWUSMD9LMZZRdno5UfdkKV
Z3SeZLhR9nnVxBuU+q9AqyAWpR3EiyMzO3LSrXJz4Dknoem4gYOsk1sjh8iWufyo
rLKMbymym+yPpnR+JC+5TPpl6ywXWeZimynVx8S19ZucvXWroTPqjVlageG7mn36
SIA8B0iWh7hTdK7PRc+RVhiuFsEuAZ5jNy4bQf4AM3dV8G7GEMh33uIZ85QwQWeE
TfR3SbgI6GroKGmO1SS4FliIs1gGdUjNXw7Jypnhn3gStJ1oOgDiNOhJ39QcEL1P
OUrPbNxEo8+gPWgjkH90MOpuMWyGf+omVFxELKa676cLKBlhxBIrInBKw/K1/TpP
q132JnG5KD3A7buxvSSYBli5FhnioyaqoWaVsfbq8vCWP1qKIRQMr51/aLa+2bEE
7+4eQllub5ZCC6vU/ettmS2l9qK07qGex5uIMj/4BhJ85obag2xsbX8cJFpM3OX1
zlZEJw2kfkjbrZzXdXxr7lHT0dvf5BnYmaPiTACHJFOYYg31T8sBMftYBoZw/qMV
q7WLsBflpTD9k0jo4PoigoqlU26nxneVHv++2yppQK9zh2BbpnMTJnv7CY49HUY6
uhLDelKWTr4FKfPJO4QvovS7XWVfJMple/KhuHxxECGex1lQeXEpe7nPH3YTcgkK
seUqy0HzX3LRR5MCJn2uzi4zxSWJfKrbniuB03Mn6+Y/nsX04Qb3XYnx0LlZ8KUk
TErmvKDg5h/8TfBuFIRjgEb/2DNp8IhpcsAu1kPtNZEh0IKNestJIpfIUyqDscXm
ix5aRG3gK75ck7exSYstu6SoXxva5byiPAvOlxT0InebAH9ihwG+GGA2dYY4WvNd
K1MydH6AnlmU9waH0gQXBEI/8yivFq18h9vU98MTMiiEfwoXhZCPYQJqRr6rb632
4JqTwqmMFD4CGnz32Fy1N6dBGAfOdkkmHc1mskqbbABgZzRmQvVHq8hUs6fN22PT
/OsUts+ZPmofm0YxPrCpjtxXysiNWFxy+1C0FW9dF6i49qeAqaOpKdDOfEGBfnpL
ShjrEseZtb7ZYMnzrXDhOzKEms69YuYlokn2YA8k1yqZ+CYFqrlUBpDpqNyZtFUc
SA1TFbI1jR2SvyxSE2vSZLzUR83ub8Ik0W3padxp/zV9s/6YbsxxaVIAcRTUSd9H
aVyVFDbGcI8hpWSUPze1TzbwT83qnMAvVEfR94NIoju/2l+PwePYK4153F3vpRNI
lT9cishtYTTA3wuQIyiIgoBBpJkK4Nqlt6senRxGfzn8IP2vAs5cDXvsnT9inq2K
6cJlhKKl8VSwdduts933hg+BVD8tNjfSzzgwwDpI+dj6RWlWQc9BxDWhvKeXaQSe
UuN/r7sYylq0QvjttbMCB5RQi/igFF8zAbu1vl0R1ajghUUvQ586igKDsuB4kIPn
HZIjs8P/yTAz3PDpjeCC6Atnq9qNgAreGHwlSQSUC0oZZK5f93xtzfnltgKlbuTp
V6HZ+O5QmUvkM0voKqK2vBBSBeUHAzq3ZGHlmnBijWRfzTdrkrdF4LLvKdFHEhak
OEVvgOi3n4xpcXTrg5o15TNj8ERvm6E1c2rF0mDN1gpJU8FU7Dr2s0dB/RzlSDEn
xX1P46wwm4Rq9wYIxoeqk2bvMBMgxwDe+ObbrMlh9mrhgYvdbbe3sXhKPh2qmmSv
n1XGmG1xWjUiNdqBEbkAG7mo6iB5z7r7JaScvu3gmD5Jkeqrq0p/dEsaWFUa0iS0
J9Bg6Bviudy5/QpBXvc7cv2WILSyYTBHU4YiHeHOc++D3tCHK00ichqfVn1eUS2u
R65hzwuXa8H6b+njn5z+iKyn7HvtlHSSTyryJWdcde7uPx/UFuXQVvT4sn3F83uf
bLX7/DwFLO9IBY+hWRZFrBSutcO3GeH1AFtA4nYx9pVY+Y4PlSJkfDWEPaI65T3M
3bylAbQYXLs51OqRzJj34iTkwxs7Fls9YgFJLYgdYdMAzdRKtByWn2rLfktEJVdq
dW1L95kaurMq/rXIdy/EDVeKoi1/ljUepfJU9opxNDNALunPxzHsVDlG8ePLQKB1
zTuK8H+M8k8kv5Av5QrUak+CHfSnGN7iwQEWTivzXrG0AYdLyYyW1Yh1FDOYFDVJ
cbXZk3rafIBjIWJAut87OBSVkMRI1iuYo+aYxswnKzf7RDw++3HTIPqWmbSd8Jh/
iy49TjY/ac7vewKNEyB6IZuA8Law6vvMi5sYK7wbdw7N4f7hT7LNeeSJAY00F9Po
fP5hXqr+gg7uxU711RG2gY3IYHSMHQ3NhcDaHmwZDepkz2aPRPLdMu7LAsazaOjm
Ukjur06CYUUmJn9HgoZ9kYAe/jSgmmLko/jOtpr1MAXk5VjhE/MePUtTdkgScqD/
1UD34j3pAZQ9+SxoMKr1QcZNGceEmDBZcz+Qa8KyecQr9EHq2N6KhPEyDHj+kt1C
6EPDpzf/B9a4xbcv+h8/LEmx+XoqEngSMGqcUkKCcMmIzeApHaAiFKfyud3CABrF
rEUIYJnk7rlaHgMmdd4mwbIm1r8MjNBLxU0Pej2F2M/NsPY/8iN+jAXT8MEkPBNJ
JSCg01KWpwQrcDyJLvFJSxYf3+6R/8vUYtq6KcHy77dT/NDmTMlfBT0H4SUESu0q
ReEHIcJk1b5o6lpbAwbBJOqwHMnpoYWnxivzRJl2IfFoYUV+nJoIzPbWehAL7np+
4XPCpoZWIbtoRpQLw5wsOLCsxiy8h7MszMV9rN9MZrUGqe2ilJxmS9RZ8yzA/WbN
nn6u/jqlmz7pbE3fXB7EJypbtZ64+mVN27Fa+4A3/G173CBipoejypRp/HrNGkon
lgWiCSNlHCz60JuILPeRkgy4OJF5AfLSi5dLZtoYt3faHf5/j/ylpUU0/FHf6kmY
eE/NnzvtKgxlye6a4CtsO9gL8nw6TSJbLhrIgnkVEBgzJk9zitaXJrXMYBRWSot/
HHsYNqgDyMqvgA9brvxnH+FkDQeEPxVAQu+Rfpao2AETk6VY8SvO8jQjffXC15NA
0c2VE9q7xtz4ytboLEajt9r9rLY7jza8Q/XABG6DUNjlk0RHVrKkWIkhXCHKtJEr
4+502DSNFHGP8/zJMI0GA07k2yxW90W3luapcx4ozsvcjIXF1cFS9lE8Gw7dqVAX
0MENsw5XJnUdBwvDcXrOMJWgcoV3ODBhtKcUldPVSQMVb+ByCuyZxxILH3VT+TkV
jVD5AB1TEPyrGw1OTLNeLgFEFGa75KBYJl8PxKKH91QHv5u8iWphOAHK2SrBdt+D
9rjwBtXcnMMTE7I7rkcZ4qCqO3lu+cRRhSxTGUevkDd22Fzsg0C4H7dSM+k5cMqj
cYkSsrOSt+7du8UM/vMBKuZVQr0oPIgTo14+K3JjVtoCEz6R7TU/mazzynlhCTOF
Ei6NzHkVOB1ZjHmnjN/jqOYxV7oSeRuFS63vCLpYcphJMW0umGdQT8BvrspE3oBv
iKpkI52tKkWYUR6l1qPSJfNR1fRMdggGJbAour9ECYkf54stKOzwsKmwXjNgz8sm
UUEymaVFNCnKQ58L13VPnLeQnj2x8PwRQfso+MpYZfMpQUYOV6Q47+BN8wJckGEc
nAF1gdl7V5xx0+/bvpjjFo4xwOvU5fsRDXBD5Brho0tGmZLzIW55aGOcADXZvrO6
1CGLq30QEihWcEMjAAJTu+sw4kMyx9n1ifADsSdE8qfVEge15mf8z7h2jYNuasaD
TlgpAxY+VYkPTCwCGuSefp3C+VeJ7zuYh5TtV/Z3q6p+WAorFM8+T24gYwRactPM
99k4nTEoe+N7pAGrxKVvF2/boOeHmzx+QP+123um9JchAIRZBAWOJSwT2ppnaxS1
+2q1Pjg0vFmMcbnKf2hrRCmmzrQQ/2vXn5FO8WKwXr753II9nouY/6o1wSMTvAET
iniK61dQFx6OoIiYiayeGPK0Br8RyL4Rox2XTQhVNpejceTtFx+1t9lf4VR9Qddq
nNrb8l4mv8HFCRzrx3ImUEajxZTGky14WmgFk7Gk7ODa9l94djeC2FjShpWuav8a
oWT2ic79pVjimtn8YHORwMRmj1VwSMjnh5yirzYSTiyKK0zKK1QBXMsN+doIVGs2
JzlgTbfGHW2PH2RjQC9QfbXSh6Jmb/XEiijbnw2/dBdxEsv7mh9VESYLXTXfIVJ9
i+mRcnBi6z7HjYXH415iato1qITo0GJa2jeIMJtYok0HXd/A5BVYBZKt2J+PVNmU
ML0aMgzL742MuvhwX22mGT7XK2DHjxW6+WsN2+GHPMVmhkGFIUwjt8iEpSHy75Eu
G2zSELcP0Zqx59F+cXJaADN4Gb62fu019xdNmyaHJ5AFy7zsfKnmJlrplR8kLhXl
c1NiDO7v3AwJlSOLu/h0LsScf0JbTT4IpxN1nEWqxlCaBiML/ntZKL2rULVBiWW/
lUThMi2lG9Nrwa43fF1Fu4eTCfREW1ywxEnCNGUejbqwDEZj/ibl4lczwuJUhsEA
oqmxTILHYoLdPTXCt3owpZreWUn299Nb1H9IjDiZZjzSnCYktfJb9puAsnqZpFV3
5pbaUkGgtm8oiF4GAMZryq/pTC+/88qWckJ6xoAlWTe8pKdvqJ3OUP0X9p6bhrtp
yVeFu2f4nkwDG5a0aZE3IfmoEx9r4JQWkjeXg58jQqXbw5F9LClU71LLFXXs/mk2
mc48LguzHUz/XHGUcx4W29ibYeoNOOQX0Jcdp7W768VPSa2nwHeao4Zg2xnArXgM
08gzZcpdHfCLnX5XEK1bV5gpaZ/FEEL5NbhKoaxRYkfT5lzujtrioDzrt5/kZFD2
HIU4wZivm0eggIqkARJugvZ/RB+LG9L7MHX38y1nkb3MDqNnpBjn1dpWEwphrQ+l
Mf1TLhUd/MhN3HG1g6FyPjBYF3AVK0IQZOqIdfIQTVpU2GXT3rLUJP8+c/YCmUK8
ZkOITkTLm+JBzGEjVzIRuUv7PWuK0u+uHKWNgFGfyTWSzfR22RYvBscufBrfbnvG
xDsBXIrLaA/KeA0BKfs/6RQqj3sEyFYZpAzaBWYfY3Y04sTPC+GiPFLPntzPKvxW
nxImZh75ei3Sb5sb1hh6nfcWRpcJEy1f4Cb2Q7+NR6AoNre5TZLuAaPh1z7YlaSt
lUwhEmsIYJ8iCD6uqaDBeBo5Z7WmOHBzw1YXXFBM/pHiwuuvMEfAdX1BEQt+nYRz
e1jmTiV4OoDtIahigcehonv59dzlqfAw/uPOh6NwbLrNHxlVWCmBp8atDcUqBS0W
ikLGWe4+yPVFfvwOx9Sxi8xPYuaSj1keUNyuUGQWY/FFIsOcst6gbKivFks8uJEo
AcU4sZtaLoqeSLvKXtVJSy34g8pKuWSO9G0nTfE8RyfbIPJ/vcWqoHWd0ke+iRW5
yumQHaDw6fdfl5viV0cZKRWPP+uKkYKidOvcrIRKM9gvxRxudqQvMFQKaGq6Us+1
eGuoiQGvGiQhkouJSNOc/bxENmXG7ZATkGJS5h4wBahOvpi17Wlh7CkKa6K74mdl
KI6eLz/G4ET1KdCS4LRnoGsXF5utfJssBWRtlQLtfZYq6P6VmPhWzynq9xcMJBQZ
W9Z0RJr/zmX/Ksxtl1l1zvmUqFTEXO4zW6clVYBpzu/fD0yOAuEGtK9HqAXDNeDQ
sTMcCQ8+gECDEUso/B0jqlyYkNiSSlldXbxEuL7mjcSC5cRYw+CEkkBCa0oPSxr4
R0JbQDctwJyR3gyrkAkKqUs59lCmLpF4NlHrAqtIv+nDaF0KymzJ1sodcUEFW9uo
7pScxnyNIs3LD9RGdCNIpG01olnYXxhu5rHxrIslt46/xaKRmixI4SbhDTX3bl3s
jXmYJDPI+Dnbg8RTMSIZ9nioaW/ptyQVQTLz1eFz03fchpmqQ6O155tHrai9zkwB
uCpIpZtyW9dAUE21iEDf+ptHJZFWeYNnLS5lVeYbXZC/1+aGTEjG8DEbI4mOidI/
qOfJeGeJhXYddkPnzGTwiVd3TDUMUrgE5odKpD2idWGkt6ghIQkH8oeeFvh06fVl
wEUsuFTageNt9H1zzTBeEsnPLioIMEuU2hwO4oErsNCrn535Lj967F8jQSUkuYZA
y18rqckb0MDOLnX4BB1dAzIpSYol2eAwKa5QXB6J/II6EswDMu/DAB2QekQbkFZ1
PVBgiDM9o5BCvwCK5j7JkZd6SuK7Jd1lMFWWp4++SL/onD7xEbMVfg2SO1QV2cgA
36o5SOSW9ZYQyR48bogShVFL2g5Fl+IiAn9SOuvqseLhg/z647E/C9TxODzrjaVE
iJWZLOd4vFimtjTnhjfPq0eHyKHeGNYOTnIFrrTNGBE47bjVxfo3w8eeLxLKM22d
1INSj0iWMEwkLUyTzDZiWI/1n8S9E020DVnaORMUP2iR7U24aZ4BejqonQicwEo5
GG8Ug0LCbmLWBa75wyq5NsZM1DjQktpW1gZurCj8c+Ml/h38TFY6d8jd3o1PRenY
2axQFY7U37cV9XVGbXEepUgteG32NEW59Ii/XDhLWzV8EoyTFUtc6pMZDurtHaGm
joRFBwtoukYJ8TR9gd6neFnF20mc+gQk7IQgAJ5ZVjy1CiE3UfexDds5ch+MTuc9
qk/+JzCH6siSLDHH7Rhee9FdAmDBIC+9M8XGGZngwZ1cRqi18eNI4E4klhx5Ukwo
66Tmjbid/6cWwhPX7PDfaNvBWif29Q4Tp55uCksvF844WR87TGqwChuu+hinlI52
twlN/BLmWtQbkUOUxIPCoSuYx37SiUSYRzYV9AgzEnFilmb2t4G91vt7eJKJP7yr
3HE+DsCXVzO37mJv6YPb8+NkpIEcEOb1aoilSigF3zT6mydRqV1hEhdCAW2yIH0N
3FjES8mY+z+SKnjRKK+/gvlNzS7NrCoqcsKD+4yCEnhQstuIlZ0egw9d166F1XeN
mqC2ulKVGlos+OoNpSyV3O5qV0pSmk3X5TfyH3pEKk6T2OSrmiasj+3w8PQSt23M
/LFSiLDVRwEkal1HBxuoDHK7mamkgzernSjmZ6UdgEUE5f1mNmqWrm2YeUsPhGsW
buR4Rsi6mN5x4ycJHV1OLaRfAcJmBV0Rt99m3GrS20nR9pUltre+YLTf9OpcPtbC
JmYq0S7RURL3EL95ENxKVkX/7kog10LNlT2XeCc2EVriaLNYllAlAz6q0+Hp1QC/
b2aXi+UKgOxE1SqOe6OK2GZ2w7T/9c2Sp+cGpte5FkpiMPqvKQop9EX6Y7yhjwT2
h6hL8TSbEnaYov2q8Wro5MTdAo3XpVOyqlvOpqr/VMAzrmL+Aoqmp/yaVVeRT2Kt
q0O1/8bViySV6B778rephjaO5/KFPXxRnk4/RTrSoPIPBb8VqX1G/SQPJhc+22tA
neHSa0Bewz2PuggqWOdW0ZRCu+FQJ+CxIwudM3psCilb/LXRl4+3cxSo1g5aJMKi
oYwmKzhw3bouAutwjS/FmOutOjEFZNWPDCp3Q6xEUTubfax6aV0b3W/XA5E056QI
GA+mlcaRicKPSaSKpaMlTOpANWOQt/3+tz5KKIaKSbwVffdg0kuUUXjbzwaBOXwt
1AT2+1XHHpHDVaqMB2glVesTvjozzWy2886ZycxK8vAQ8cFaTUHE2i9fi0xn4aDi
gAK+xBbPaXVOTtWzyCJkONQHe6m/fw36QSHgd3cPf7RdfFi9jVfcZEJdBLO4dLVX
Zxj6/GGOeiYs0OgSYpmfWm3DEabf7cYVLm1UP+7+Yodiwnmiembtxpc4nXBDwmaI
`protect END_PROTECTED
