`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3PJsqJCo8S0C+S+lLYQeNz24dUbKLPJRSgkXHX957uXYWkeF0tCORMrtFCrqMv/
7Yb1SQWSrHgo7cIw4m2pMrbGwvAu4/ekU9Y7KfG3Id4zDxg9iGrbANQYe1HH6GJ/
PXsItofEZbJ60e57apf5JHD/98J/V799bGfHblh/hyKhjoQIjsbAT4moPX5+5gUi
47kIeu4yX2nMMeuemv6WjfB1A/Jm7yXzGW16IZXX7yxsS40Q8jePaimvBIV4lsId
pqFnXTzjds0DFZ9GnHZur2BS+dtktyAxNMQFqRz4R/KVAq2XDYWlfZbkBhcDDCMc
b0581hECEGp21OwYefT5MDsefwMkZoJUaYC9FDFtYJBXioaPs5iQy2nzJBgbuOai
qkEZ+T5MlukXihE1qBdieOFNaI2vRp7hTzoS9L2s2TAr2YCR0NkN8L/w5sh+5DoF
+vVxiaRtcahLxSXkcsEUHeu2somd+IDyJXMvxMFv2PY7ahsdTxSNgsW8qvKoHb27
BQ0soxwcZU3zyZ//2jBEawY/U2ZnV3mkMLS9P62OmHjlSn60sHl04C5hkYm1czRB
zFcRd30bA3gP/a/IqwlUikv6cXVBwuvGefMxPLj3cAQuSFraaCoHvNzB5E2hDRHe
nubYzANh+7D/BjzoK98GuUvmhX4+t1ugTwWdt0dSoi0=
`protect END_PROTECTED
