`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihpdHhQTyXfJ7CcfIzUP4I17O1QM20cWm0gZfPIwHvWPimgqV2GLou1MT8o4/GyZ
sgQtyfG0DHVE4LiHywdy/j3wQw6wDbePW3ImYKskzhnKrjU3XZ5zWRl+3gD8ju0W
ywWFO5G2s1m03AhzBuZM0FAO74Ctnl83D4qK8dhC/VmDYVEAb++BSB2RL6Nf6NDD
bKL4V1jJ+7Ta719k9Vru80Txk8R7owDvTE6ud/v1kUIjotdU45a4Z14/uJepGccL
DcOsNvqTOBin2ABvqY42rqMCwydKcw1AWzCt3+ul+v9p9VNa6MsAIDbP/LuSqXTB
Dje5LmfH6aUL6FVdI0mil+K/XuZD2fcqF7NpNyb8yKxCqfW0B0MwkthXzIGnxsnp
Nsx0ZzLclVUp0deTtdrtQY21LRJZWCF5L4JaVY63qtUVNi/TDFFIxrtPeSR47E+M
HscNEFpJ8xXqNyXZAzhdRW50YXLb9tUsYuAEo0PT+FZzjBG4ggRVTqWYtcD+vKrr
TF7w1N01E4tMvI/ZNkPLHe+dJ5uVSg3K9k+lSEw3lWMleLhL79XoQOkbeCUu2XX5
Z6mns9jviSTT5z1nQ/xvMF1BrAeBbHwbbGZCagPdHrggDEbId/vnR6UBYW/RYYC3
mNU+BSMqGDmtYNJJZ4ptvVwcV/PXvkTiUdqyHtZ9iOMl5K0lUjGFseaC1J0IBx24
X/XBUzx4DNTF3mebpypR41D79lH8u7Bz4pyuyiKavpNYyL+IG0y2WcuqK+hSzEdL
kruSq4EtySkGzlz8ooiWXktkSMFGZAkRMoMLmd3Mo9Y=
`protect END_PROTECTED
