`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7sn6SSmmzImHwhxfqKjTxOwtq6CMqKJG1MthT7gqMWbLlgEVsw95BPlEgN7Gr3so
7BGXgLGENEcxBXmdQuUYjU5Nyf11CQVPYGOG5RQNMmLz0M4dZEo/rtKmzbwvhhlD
2WY6epO4WfV7Q2Q+nxc4GepJWBT/aIpsbQugyyvPMIeHdZPJF7GjNvKdL0tWu8cI
21LM5zUxNzke19NIx9C0H7ab7W/Q0CygzXg+03oNwyfhbwpMC8E24UdVlbJWa8hX
u/N8fSFkzwNuCBviHlc3FhWtu/zXJIC0DKmIzsLRl3r58ZG28Lb1DHYBdOpKXiv8
9zuF+iYOKRUfIqhbaSuSCr2YWgudmR2kD6J2/pMLqCUDSyxWMhWcwcg0jVu21JRl
X39fI0IvhSNXGQEzTNvbyYi/2opHoKXfXVH/wAVrfRm94DkqS5xqgliwRO9EBzXZ
`protect END_PROTECTED
