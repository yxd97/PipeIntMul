`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
806EMh5xU5DT8xG96Q6tcV6x7yItvB/QzolVLY+xBVU3FhkxQwr6nGb6/RchrVk6
lijfBpWE+/VPB5pWHx1v056omA/cYEJ3ByFaqBZoSkc3h5dkRPBivfqXSy0HTJzP
tHT7p4vnwrJXVgk8yKQE+ioV08/mGyF98zxHuJTNyo9+4gqYXfnoWq4LtJ5+PeNT
ElDaVSCO5XN52stC90fvesvdZOtDIh6gBViHHTfC9vT/d3tV/ZLlfrQamTy7y8k4
4qgKEwbJrH7UMi3ZwdiZipYlsQlxlPbYdsNTbd/Net8wLqnrhfZTBUCV+U9jh6cA
YWOWkdoqcv0tNnzBGkEbkEi8jl1ps4JTX+9s9IVX9YiYnuRY+vkFXL2/KvPGcoxi
OU3Wu/J4LXUEwlqGVm47dHpjk5CeQPeaCFva4RQSq5dBZPKO4R7hpF5xrfw2VVl+
CpV7HKlI2Nz/vU0padhRPH0M+g2zDGwGFZ90CLHdAWNjSUnZGAtAO5wx0IFsy75U
NtwxS1E2vysOkEsgAUbv6cwjEWN7iyEYlXFwbLMXWB4l97JrzL9a7RM+MUonT/yT
l2mbtLv6alJFqOTRKFTmeasFyrwNZXukLEnO3EzNUQEukOa8HjEg3lZnRdESGpnW
W3+m30yvrnGfip6jnnyMjvUoct2DS/w0suN7mKdQUBmaIUYE1vqLjUn6k2FRmNfM
1Q40hVmrzt9kBj4rbS0dfYg+JhZTYHPU0eRiB6skACM=
`protect END_PROTECTED
