`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iMDxwLnb0d7zFsQhEMGt5fApqxRqG9rsaUsN7D3yrh6XjOf1DIQVgoHGVHCNYkCN
kbjALm0e+g/unZnjpxR6lu9Gspi0vyQlICI6DwdxXMQ6q9+1M3hBOOyJsa55+NeS
KCrpq7Uz8btDIq9YoTKQE3F9zm/YhK7uiP1ykguVuodqCzB9RuEHOIX9C5DFGNRF
eieD1Uxn13O+94eQfE656KdgZ7pBEo7ZO+AvIXwHJfXEWt8KfizisZI23b/UtUcq
zqgFyU2kkhsq0vSLzGmW1arTnUTN1zRvwKggSJe9WnKiRLUkNXxVXUOX/f5jyGfA
RwgB7W6fI3cL5xQgwYlDdfOpZ/BE+zoQtO5XTXxK+H5QCk05L0aXioan3kzxIHAb
hAAm87QjveSeTvEjXd8o83A2K0oOOmiZD7ARoxanlLkk7aKe3dcMPAFWJunl4mz2
yKL+hOJHXhHU6M0yr07LTELgJLdalN7XbvbKq4AIO+ZVguokc4DJu5lWvDe6LJr0
+WoP70ylxoJCksLZHWOJ6PPoaChMke7DKqm5yav34NJU7+G8lex7Ra0wNQD2Xhvs
bug/3q728ZeTCGzpXrSfYLlslslR2CkFAdiAk1EF7C9sBCYhWK33Z3n9p0h43fUG
aTCfBXB9akdirKG/7nWUj4XF4qAMbSGLCOJBvN0+wS4oCfjnAXcDJXNaueB4S4XK
NVI+nW36GCsXplywUhvXVMSmOPYO2Jz34ViP1KArUiQ4JRTjhQOzelEC+fDTiU8V
SBZ6QozxK8lz25nCSHSOPiLrHzL86o/ZrsCL+vt9cderj4gyNPbE/eERnJ9B+Mx/
OllEmOvyCU4qOiGD8e6fQ7QMULDAcTrmSTeumyr11N7nW+g6bcIJeXzFr9DQxISx
Jaj0JlpI8NL/Fo0mrD/4CPkubj/OkkMtpZUXNYhkGttg61fT4vfqwqVOAy6z3pa3
`protect END_PROTECTED
