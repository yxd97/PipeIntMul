`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OzJjHVq0l4F4FDQqjj0hnY7Uk8cBPml3WLayF/qVmhUQGlye9GCJpGXhyOZjBFzE
anPTXMzbOkD2BDN1hFzusTXuY6ZELNjRfqaiOcIm/SmIa6LFjWL2b6x7aOWp53UU
3WTr5FVgektbQ7FtMfi9Ybz/cF41DDaTH7baqadVwf/v5cSP7qYxxbUxoGL80hIZ
LfGKLD/paiRCgfEFFesh9EkkVCe+ycEM45eBLG8otpLiXiw/+wds1+ZTF/e5RY3k
D89e2O7dW6qnm3O/xfBdUiQzDjr5uakuzzrX8X3CseF2RzlAj3u7YBKTQPbQOhSN
97Za0CxZZmZ51ESim0P/nQ3tzYWd9sct/8sIlAT5Su/JOTWvq7DGZ5FmG67PZOSw
KNU3jZ7LwNRFfPDO5f8FsVaPDK7jKLSzJupq4F36iN4UEGdnUqsnFqacga5A9tdZ
LE3gCObuLt42y2cErWkDMzipgeRErWC7Bul5IPlVPQRDaEYLQQGpfFeiI1u6kjiv
MA9Aly7+FjAFRHmBL5CHOobJl+FyEngSFVpUH0D320oHpVmB9jJTadBPCWSjIO7J
17rkN7tSeTomClIh8a0E471ZYFYGPSlocFsDLldT7qT9VNrt+4GzJACOb3XrAog3
jgler3ngbnXNGDoZ5iS8Eonq3mic6WrX2mbWEzIZhTnyVQT7ZcaWSk+ML9CV0f0B
1U2lDw9GJMO6kJbuTOf6Me1LrMeQW1OLTxae87RVMspAOoKh/xRS6UTaoAUnohDK
R15+hrSh1bQM/IOuYF2qn1yr0lnqPcwIDazzQsIiJDxz+xCkOVtRalcNli4GjYWT
4UJHOE6RbVJZ9eIsGESTfMNzNveGPVLCwlgaHV1COAnL0JlyQAV8dTvRNxBE/gGx
o9Ae0/lA3+wgzK//bOYAhc7szEuAuBWXOIhLebUyipZ3ehF1iKmDutkjlnhE7Yyf
wxQRF8TooHfhUh76tjbUjbqcb3F6e6dsWj0OpOw/k8iT1URg4WviyFSn5uKc5Lvr
`protect END_PROTECTED
