`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJis/fktBLIS11GySSW/PTo6o32oqb0Z/rV2vd9j1dg7xD9/DNUsS+3+0U7TjWGB
lkT9RMPNEBJMl8UWZ4G1OPRe4JM4wO3iHHelPN3G8nd4ArIDybU+qySoLGTDidVh
mWSZbibfiekrUAcaFAlcUTu8kyezdZUSidw1OOCRXFTOOQ77PbRwuRTnr0Y18Yb+
O5Bq8vXEfjfW8SLk/JXnvClmQ6+no0YoVf3/APRMTicZ/3D0zJqTsDUWvzR813Aa
lpydRm8uk8Vw7t0YHa/S2rO3LFqaKX7T21MAR5Zogs0OPBZ2BLejmBP0a0dgTGiB
rTF/Ene2UaRgcEcS79Tts3LvK7+OTaWThQEbSInvdifbc9gwVqOfQGzjFuJqhcIB
`protect END_PROTECTED
