`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3flIkJJM0RF17Tvfya47okdnPhx08HiMzHYnSMFdJ+CL2KCELkmZ3k6E9PFxrZiX
QFgjGckKAcDMtGWf5AVEHLi/8t74lqhFtQuNa3SrB+1aN5MMgXhaQTaWlsp7DhDe
4ltDk8hoIXuPBzc6pvjw2f6VYgFrkT0aFJBTm51e4AqL3kBf2gHD7kpZ76h1hZ6k
M+Yp0+oBW4uxyqLsEcPw5RxPKIgXtn9jG7+8ZgH0OdOEwBwkOIdxVxEdllUEeDCL
l1PnQgoAt4W97TmVAUT/fVqhnpQ3jXG6gc5/UHD0+eDAKfnkXcI7sxfjz4eAz8th
f1rpE2O6Y6XZC0um/fH2sI1hfLpGHaTk7i2+PJv1NKMTx/PxamY0iQ0nRyKvgGD1
5Y11WHwrP9E3onr8KI3z4zV8Tv6OTwUZa+82MKpiC5YbdroXEu/jfr2tq4TWIHQM
fTStCNxwgGhQt8ifmVosJWOerwQRtWcY9ERivVJWdkW/elcpZWDdcAw8zLt7GcBX
BSQUdeclwhlVjpb8Oi3T95hw5jW5DPabSYJXRHaexhP4Lqek/w2n2G++RS0/0AUk
+j+zO7rwC90YRLM3qsqMSaC66gUVB3ZjC1kqDCbNKixNiqVOOwds4VX2s8v40w5S
bKOpbr45bBYziFd+QINuQg==
`protect END_PROTECTED
