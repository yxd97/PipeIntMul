`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wS2zSq1MuO9s0D8ZGaATw0LyVj/RlyUrqVymspUQTU3WC4mV+SbTXW/+FSOt0JDs
lowwOwMOIKWhH+OJeN1mICRrZoLBWHNLZfnIQD0RcN13oeL89ugZ4u7Bd80wg0CX
8xfQiNtnzgEkNgWYnLLcl0+hu3PEyHSDZ524ptdURAaO19LlfCAycWO/L2XnpJ03
CF4nDmSBa64JVVZKjVDhMRcRDkSzbX33kXpHmCUKWrE8OPmC3+7O//5oJ73cHoCa
cAZSASNG5k5bANp5ijjV2Cy9r1iDBeHTNYRrdej16SGftvX30ZPyuFRHBhmLqhnS
Dw31vMuANSNHVoW7DfKgc1C/V5v9cQ76qepBHF3FXzfurz1Xq9E9a5H2yVLQO8MQ
Mq2KOwtgEv0Bx1TLW/wMrGvahS55y8eJQuXpLi0ImEngFdXcwIsc9UmWsfF6owSK
MWlNHKciEntqoxjVbLzNepAgzI/I0ozqf814DMUze8or4IUjyTEs+K/8WETkO28W
mkuy45kU4wwM+vpB8Mc4A3eLSOEvi6B4c20gd7cl6hLIa5HMNacJsbWWf3PwrLPB
q+4G0VyLfpCPGnoQEJ1g5Ad9P5LiaijxhNqQmAxQrvBAAxnpasWBpiYziigCd84V
sbj6vtfFjyAXrvU7/Z9BrQ==
`protect END_PROTECTED
