`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JlVG3nZY6zF/HqLifcPl/O+TQLPiZTfzqe06nv1ZPM/K1xlUFwQ8QBu574M84X0+
QSuctW1BciZVSn8wo2lX7LOckaMCwePlc+/VWlK702h4sKyTnh3uR5KoOwgmZAGL
xTNJ9MfnRFC2ZC65JSLcKUAo5kRLl/xmO1/naMoIY5qtV5O94htV0xtHCId5oGsX
cScgch/4D16FinDTSEpijRDqwEYmqVf967lRxuONERQ9fLI+Aait8mPWnQsQdYJd
BqFUuW4c7se491nfdHGbPFyZYvF0Tz6KJeC6FWjnID0qPof1kaMNfbii6rjZpehW
vUXBNL6E/lL9+0eYEBQgFpZdLf8mhFbeksVMPr79d0YLB6veLR0uy4UCii13xs7b
qLXLjXnu2ISZRAkPtsQJNzpNPafzCI2Gl/8i0cxu8u4a68r3jAwQQOoip8B+Mw4o
By8nkkuCLam/Kv8sdyekH3Pc9RmFI8ImFReVxvVwpC0=
`protect END_PROTECTED
