`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gsd30w2N8Uue4PktERlYBymx8sJuPr30o9MWfuxK95yTcm2JJxe+wHfmy/nzv008
W8WrjHd9DMzEGfkFc590C0fVmoh0+nw1sUosTmPT0Kdx/vu7AUqp3AUogBCsmrNj
bIt34XX4igMCjwsdwRoX/6tz5rcE4ZQtmPctp7Uj0UDr/TIhW/u/GTjl2YSSwhrU
qC8t+7aY5YjmOpU1i2MIzB+B6qzK+mS/8WTEK/w3iL+twmC0ikWT5aTXdHG388y8
PyRJkaaH+HSBjBSlOhqLzKguoQDkzCleJgya8aT+UHjlXDz02nQjEJg5TKhhj8V5
mfZHH3zc6bCjb9Xgd7XQV96P+zQsei3nD83OxLyC7EjyQEj9a5S5lpel/jAxMQl0
xZAyb5lDPqKQQas0r0J3YwqA5YsA3C+yU3H6nCHtNbZQSBUqRV238ipRIq+1JOW8
kyhVxVzku1W9ST8886ODlSdrcD0KWcubTnZmRe1q1Y7Y0SmwcXFjvfRLHsUeQYC2
kYDgyYukBzsWr/ZTIqszrfemvo8S9SCmAzyWjhVYyX4=
`protect END_PROTECTED
