`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GiDOYDN8K1Ma8vxFOm4UGXrJ5uFbHOGYKOWtHZQqq+JUoQV4GOxIaUb58qoQzA3d
MGrVts5BT3J1/GHpgdf40NpOMCNi4HilADDFIuKruBtcY2ZxCxjlLwaEzaz9TioR
+9g6nXwoaOxdXr8tke4q8EaYhWVUmxCo6w6k/Q2XGhP75pVjJYQXNVrhkjSoverk
RDeXj0cw1H5DWAxlr1WC4HFhhWXoCb/z2wdVKdYPEkzJHksUhMj4rBItllmTrMPh
jxAUd1yYI8sL9VTcy49+EQb8TSMzRk1uvqsfvhIclUg3HZ7mapEBmfkcha+V72QE
6d88SIcJg22BSR+TaJvQeTDn1KyXveKbkBh1AjmWqwrysmZ8K4WwFqvlHt8cNTh4
Qss4ze3MUNCBHDAzowhy7RUEeUuxdddLK8O0JiJ2Kj8=
`protect END_PROTECTED
