`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iSfxfiaL0u7cr0rZW4/bxLRp67LCM8qrAx03vLp0nSaRUUv/ZnI/EuWTGeLquOK3
WGBc4MQwfLxWTEdbV1JdSqEoavOMOff1LWJUT4tx0CT1bEHo5SXCBLN1Q9qV4Z8E
p5z/b84thEC4+8BfqLdB2ZkVAIxHfLe5clfE4jaNbxf0p9RA3Rhw3QRQOl/hG+gs
BoN+4dRNevpjBtBSOP6g2EfPboXyPLvDqB79JqqZo8LrFWnpbrX3FRMR0AJMFetH
CAbfhYWbcJhGsXXOwHWIp18xM6UDMIzpw0SffIaDC1Wlz2klcSPDv1FlXY0QlvHx
vEnoYvnazwJWspwEHbymK7LGOnFt25RhANS1tq+G4zhiNa8PrZZIBIKSl2tmO4ZJ
PDHsj75hrnsYBDykLTgpWCO/TE2LnribhTNGUoumUKNGdVkQmzQthFIK3d5X1AR2
EJ/HqoaU93xLhOgJfO2AYTr8iNdr4yHa1rbVY9vi3/0LuiDWNBU0gcx/vZBGFyuf
eZfrAcv+QW8MSLJ6Wgmy456lbWU2Sw3Nuyhj1GgkMwhLPGZNDwkoecVsQ71FN7vt
7uW/gg8djeRw8y9J75Evs6SsTq1hH9LgWbwGnMLbCd5btUjAzONLBJDHfRKNgOo4
`protect END_PROTECTED
