`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B2fVJJLiD5oQuP+txrVZAMeFSamhIN1vdFs8w98n1VhZgsw+BlIKZlStx9jT53tf
oPwx0QJwRSKWc5DLf/9BzCKJA1uzAfnRvlgbMjHS/vdg7XAANpLa/9sqwMhE8g8y
QK42gHivKQeNxLFIJEO6QuWSXIBzsN1SmmmR0LjBMLMuO+p28CvsHMgLQRcNeQoI
5tsy7wdpSKM1JN1AT6bTWpISkIvqQkkW00ZhG+3U3LbOQdOboSdIC0lSYlHW/6pc
jpdaEPwgO+zy7oB2KzIGDzUw1Bht7URWYJ1rFVbRlsUtbUbayLsQ6xENXc5pTjBh
RXT3KTcMJudTbYH5i2MzKeeweEEA4fOx3IJVUCRZIo0PzTPONE4ScxfTVCb/xCrE
UCsLl0YF8Vn96lqnSo0uIw==
`protect END_PROTECTED
