`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zloUG25v5Kf+kChs7G29NHUcSz9g2UwAI+1kMmyWxCfmFF1PXCLSuJDTn7rsLZd/
96sKFKWSpsksezs3Bn5m9TZbASljtBdBkpD1s/D/IlI6R/VK/jSu4uQ5VWdmHLOw
G+R9WP9MP8PKb27wih9qRO6Ke9z6MdVN+MnokV0u2ZR7GxtBJZZwc1GTUUXB+94P
peBDJHEK3e0yBdYxPtISNqdQYIP2b7y422wwNOvRzEyJGJnucdK6U1wppgfK3f73
KlvITqqoRvDDvNdZFLgrsS2CiPr0sb7QvY8ggjnT3QJ56O+J09DxyJgePXT84LJp
jCLWkp7mjXs8TE1gObWpuJNEU0GtWKUIQ7BdB9bUefAfy1zM/lQ8Q3Py4NJcH15g
T5x/ZSDWvJ/Tpq2mLrH3wYNaZiBzWRWagGr6DixTt7FdAyyhPBEHsNZaGRMdjZRQ
TmuPcDitEuf3m2OlOuTuG6QPuf1yu8XHQ6JYNriHSeHVSR/Tmht9000pOyVCg5So
cuMCJX/iLsQPHki65ed3P5WE5VIl3fqsx+6fUKXqfNo=
`protect END_PROTECTED
