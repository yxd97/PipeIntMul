`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/usp1gOjZycghc/pVnYUEKlgAM9VjO7ddizg2ztyCdduQrJWZUVkOZyIMjdVXvl
cNN31UvyLasnAR5+Lk0I2YKJls0V4CAbmHDG8jUUxi39OQxGAj0FffZl0bDy4pvW
T3gvN3DSJ5yd/+fqDL2iMwJe6+7MmzPfmY2zgNLvUuGVtEShOzi4GcCHI9TetlWv
uyAnukjsOUked2pD015sOysIKV3lFApQdEFD/hUQbElLF03+lfHbjWk5phqXBcwA
LJ1tfQS0Fgx61WJqgGyKbckHt4FLpHQN6WxE4yndwcA=
`protect END_PROTECTED
