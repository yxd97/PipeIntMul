`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z51ZKyHgztclZVwXkswBGdZK413aW37C/RJEUIul7O3uT6tf2XSCCciCb4K4pEWF
zTy8oIlnwsMMyYg9k2q0U5ArwvFKhtljaDKqpp77tHFNOQ5PEebu0aEBR3Kir4w4
EynNKd7Ck7QBPL0hn4jEeWR2GbF15/rMeRGKc9acJHbvNXjC7WvnhejxEqsJ/xdd
lX6GjjiNadjfIcMh3rVxX6QjKui+kuo84JuUnM1tk4Nft8pIoTUApx+KSgrC3XR2
rG+Ta60EH5DmGkBgzwr6nOhYNTRcnutdfWt7YCWK9qA=
`protect END_PROTECTED
