`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Z/owtejl8Od/aBLvGOV9EtmTZRzdDdwRw2N39JIoxgJjPQD+9Rxo+m2y19axhYB
oKL16CLeq527csQdlvHkLolpL12UHPPzqC7hM4kMdh2c4lL0r4yL6jXDTwJFidBI
Wa9n7Pj2Qjcpy+GbmPe7IprglGHSoDpd1EyfEtYA9rpmehIDf02XZbKkJr7JuXeo
SxHgoVbIckko/Y7RFl7glrnLLGLUHjtHgrzdFL62WsA6ZJit5E7NlecLdp1IAm1V
gWa9QqtoaJ8NfvYRZddCz6H6PkMRyB5YU7PbtpWDPj7JYS9bbksQICX3FPB7KCch
QmiEW2GByLhhS5Vn3N2m4SaRcAhpFifQOUz4iZ6pNC+4bWTTzBKJ0X7yBRr3SwoT
mZh3Gk9+0EhZbCSoi6MbVCjt+oXf6D6NpC3KonW0/RMMzJQxe1JQ2vY+FQzY+7XO
hH3xxhOTNgjOvfV18MQ+WgSlD/xRfj1Nyn5Ol2VOzNtoWKed33WuAGzs7DL13qXF
EmzTE5EM6HrLTRDFmFsQdls46KCFJ333Lp+2fOMFhm0=
`protect END_PROTECTED
