`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B63OYZftWc9PO1to0FEG/ikGhuvyVVtZls61ZjILpnTW6dcPrG84NVno0Sd8HUZT
ERgoH872jUx6XYDeQaUF3oGF7HHCmoVr0zuDUtYiE+VHDEgRWSebE4Bnlh+NDinG
+nC3V13xrWs3Cu+TbdlBqLEbXp9Y7llGTtsbdXI8iNGT72weRMeMo5GOBFngogpI
JydnNNB3zA4IexWZC6dtBQ==
`protect END_PROTECTED
