`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A3BZpX2zce6WSIrCgZRJRH2lvAVOnGz5YSV2VFnV6s0+X6sH++tJLtuNOl+9EdC7
xfzuBFkp7Wa4L4dEDd2m+02Ka70LLDUr/029BwsVPgx7/YLHY3a635fmFej1VnCs
1pn/BdU9k0oerLiKneAwX7YnK63lxQ1TcCpIGs210+4VCU5D1xKtWN0yEAzmpywO
0WDZgJ+UT5SoomAeW1pzfQYDLX+EvaLPXgWnkcwYwm9fDLopsP2/UouNXs1zcgof
PJ9FaHQKOcO1Dd59h4JI//7MlRfv2PqYwTthV32gkxVeSaudQX5MOEWOqU9LWN85
Fo0aXN9e6uM7PqbxxzG2iQ==
`protect END_PROTECTED
