`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aycXc8uKq17eSzpI0D6twxYcVrgmqC6GUzOnbZjKBN7Aw7Yhdg8vB081W8rsL9XQ
yUjNXDu+ddCXjHDJ5wshQcPvhNE+AF4AWrPV2Ky0eMPpMrOmaYd9A4qO5jiVlMsG
AgOYCKzgys7Ne9JWRJh9ezvoXmzhMzmRX7QjFuBL00ROkP33fpBRCUsdUnobqsaE
t6uumvmYE8v0tjU24rc2bssX6qP82BMzYobtg9+E1jwlnz857Xc+Mq+Dl6NTI6FM
WU8Sv2DbeLqGvwDC0HA6kG86++TEVgtptpSnWeerKJJcZ8OqcO1WNi18Mu6BEe40
7+Ta+qknCQt9JU14ec5EeCjhe1LJXUD/97ZzZ9CW1A6eoe2+Mk7TLRXoLCdIiZci
r8I72SiRszDvjmWD+/jWrFRl2J7j3Xk47jBeiV2U9GAA0zS3ZOFsGhPFFCNIG7OF
ykfynRn5MUJ36uOgxmQRqctkhrDMAwCFifqnxTuj8LA=
`protect END_PROTECTED
