`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WrJ2T6Z7PcMkfw0n9V6Gw79bDiRUBB9LzCJbN5/qMlGaYfyQhGriykuJGMe2TkcF
l+rOoqC0j87WMJ2/RXCoS90pJltgo6Esvc2QaO0WvQZBjstfu5tUCIOwegFK/zHD
7CaleG+LmXV00tG+LTVJJLC8Yrj2dcgPORO3gksAAZS1di1ATnx95GdYrg/CYVzG
4LOY/5xNAS7AShLBwfMDd3Na1ueHDsR3+QRmI8/czMTfNKfdggZF7M5iZ6SkTuY8
HCn4hUS2D6cegx2MNQ2c6CxW5k15sRuf5Cjx9XF9iSZ4Yh7nA7ozm8eWOF3n4Nx6
ydM4jGBCjSRlVH4XT1TflhMS8I4l4h46sSZqEWlzNikUauwS2Kuta76kissigLWg
VX/skpTfUOIFN5ueGLz6qW74+hmqggVJ/4UCg8UjTPtT4eY4q5UZwf5iieFKNn/I
5vHAj5bez0m150BEQgFc67zjHOLxHxT/lfevFigAd1QER3Hrwjf9DBU9gHGbCUrW
vWyE2Svcabu6gsY8jVwQ4hG9y/ZXykRHDqVkyhiP23KTecIgQRlT3kuL7DKz5xja
joKp3qs2rqwFOYJuVKkiPF2y+jc3nzooGxi8kwDUSebx2ObH5vOJXTXnVHkQbPT/
jmnCS/Lj/Mhh6OTtbcQ9nDcfLfWuZOJQiNPVWsNBJjzarahSNfeov99r5tvZLYhs
upJujr2LW7ZHzQ2x0Vqr+TQNW6cVpWC5J++ugkbqtfIU/udSr4XXqMqJn1mq4Ody
YvUYgJpVyz72Agyc02H49GJu7AB3cjg8R7m54bpxIusRHk5HjzILhbX8AiBXxYmT
jjnvMBlNHaXl3XE8gqrCD3VbvO+8d0ETWsBukamolKTdtIv3Z9ok5xZ36pEnf4qZ
UO5YYT5p2hmm/FQ1GF/OyWJ7YP66rwhdhkNYv09RTlj28zcscYTSVkGM198ztt/y
BZdhdIjiPb1vhgBsRHK0f7pJkAfrXURJX7m9oATRIxmfrmN56uzYNNAWRREotOMG
LxI5SjEUumA6BM1rQoMH/PB/adiLA+ScJxSxl4S5X26nXQ0zQb0dDNfnHjjQpjjK
hoqWqJZO3dBIEGya4sTFi/Ai6rX/BQj1Zi5Up4QKxyLKMJCQf58tOj1cwSZbEDn+
dj4kUZnWrC5IPpvN8bZiYFBw+UT8OL+uU8GMUAVv3FO/V1CgvRNfc0ADCcFmqCsv
fWDkAF5JgkHi8TMxsNBrEzWxDxl/UgwlTOjKLy8wtJaW9BIjocV37FULB8wfnevo
VMxkSZD+ltH6Jm70nnQiQ4hP3dsd6e5quOIe6pYi4FsTcPSiyw2fTJBf/uaX/1o2
rtrOHWDiTIHW3FZryJ1u37RnvsJdlZfqCJCflDDVIMHUFi3ue9TqOwHHw3lVJwZK
cf5wYOvYhgvIJA64NEYsdny1OnlL0YMojTKqh9c6m363CBOSKQNdZdaXexRHvHKV
rZHg05/sOWCLjypkYNU4L0P+I9JxkTzJUHXJsWQPcMUmkZ7b63+rV0EJjUPIuMEW
eBg3F0kH6uFTybLa1S13X97KgUfgFgtxDfbxkxr2dyOXcsHnf+k7Z9s5akKSuMRB
1SIJEN1BnhOZHx2QAWAoVb8kHXFHWCnVWtfitgesa5z05L/wjbOmnnN4lvLFjI4K
CsVKw9DnPVp1uDgoWhvMPg7VpY3oQD7JAe7AHWNOpJ9QPjwKK9tsudp6ZX/+AFOe
zqLuy5uXCR85FYG+CCzZD1xbEipGkREBjTmU7Ravg00CKMoXi0o6EQknJRwFIVwE
qtBMPRSRAd2uY3FI49uWJnqtqGZ2fDJKd6FIKO7/kyFfpikQXOAjOxA8TD1KaaCA
7/jnYSxYIVPVgYYW5nAHKB+VPVtHLa3kitaM7PadWvw=
`protect END_PROTECTED
