`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zV63u1yFo3a5kX8uIsdl1PG67O9cNCj+l0K76Q0b1QyasF+JxleszR1rVmoX7I/N
7ES0pk7Gq2+S3aCYG+xDi+x290BSOJ49geavM1cLQibtkrNLwHI+3ezvMBsALJuq
/Xfv7ulwJaP3DHvxBI5no8KI4rHIyup4yF+QElEhqGyNaevdN6DaLkNM6iRYdDGw
6N41EHIokHFhUuzJnVbGdYFaNGgnIYP06D9H0L7NKGcgMstrYFZc4QpV8rl7nVkL
lFwjG8VwPi6mlNUAM43iiru2qT8R1NCFpGeXTbpDLRNpnnVTo7CbaVyVkuB6rCTH
WWO2RHQLz0uOLE1dUq1tBmoJQhh+RAItGZ/KxcXG495gnk5iQ4MZKxAU7E9dzUw3
Q9Et5fhLgajXHPnumsflvdLrWyCuoxFiDbMaSsaqPgNoAve01YlxnBEzacw9m0bL
xvGN8gsIyBzkspDoxYeJCSwDMhb3gf2EeCeUeP83nbpllK1twCDbRKhf5AzL0eqL
jaEhEr87xZ+/2UjRodm/07NFJkQGUX7l+xFQjnuxbAduE5tC/cByHBMBUfOiFxKL
xayjiBMYhH4Xb4D+4RuTfrTd7ngIB0XHf6PBb1hFyl7KS5gU5P/M4UF3ILcjL40R
KQknF4ocXisnO9Gb2vBhiAaOecTKIsCtpNvX4JJZhZRwDDExGP5IcmjI5zubZj2J
a6Nh725qDeya7RTCvriIF05+58t+rGkGHrgeZMzE6awNyu3By4sj14hhejzxDvLg
V4PWRYm4DjE0BuCcyhh0C0eMKE7K0pkcqQZFtShsuYApALBE8VUbxRLkzS2BjcSb
bQJEx6ckA1D5pEfAm2I8W2am2+wO0YQoXzzDnbLNpNO+HIhonVYWtXVOgm0/rl/C
RT3RUam0syNdjkU3iX8Bon2opMw+Zy99QvDgrTDVhZh6lGc1PpGriylPeWzZ7Ia2
+ZdQZQEDODpme64qHhHDEQ3a2JXZBE0ta1wVSOikFtLZzOniYOXBubfyr+jnVKon
hD/SRQiUeANIQ/aXdbFRyoakzWc7aUO/hlDeT6bmOeNK9k+mU0ugHlQjg3GpVnt0
D4UajRGk85XjhnZAmuW1rglI5BrbHSmXF3AZPcWFxCyEtxG0dMtR166JxyvwF6A3
mKhhAwuUBYwWHKOeqdporVJ3xSjhjbTdPq6e9vFJsxABrXGKhb+HOeDbrwd7ZrDA
n7As3Qn3qm6JJR4zDhiBoIyC/NsVh1RteMDFXfhYE3B/ulB62EI+o1Po27hFioke
R/R0w2+iQe/NTfE5jZmddsWWBqb9N3ScxJqtvaykOZ1ijczdmxa+caigpUZTOv6i
OJjVCXWW+Hcx3Dl4q9nKXc8cMkRUTgqIeyI5FM+kL6h0YGBQWqfYrMtn0wTEML5x
tSg0DSvFnc7wa9YktTONYWWgqJBkGdA9q9GbJFI+EPMcQuOwxc0anik0L7WcS3hi
scwRnj/jcSKplHfuwz4WYagT9rX+NnW8Mxnyx6utLwkx/VUO3vUfuLzwfnasRFd0
tHGL2DkoKjVv5y41ykAY/xTwbKRaI87AH3nRTkXO7gUIAEgtgI6/9YJprudmasv/
AVRuz/Uf2aDd6E2PKRf/0vlm3LDFYH1A66dsvkh0GSIa24cTzN1Ej2YvppfiNtKo
R/h7MeJOkbWAAZBZEqy+9MRX5XUpfFDGXn3oPd1jnw0w+HXLZ8ErUq4lcRY60fra
wWpoCSg+SwBMKYy9jILa+Npu61qJFOkcMQduzuJy4TG2xlZmG8OdOkTYmUkQDBCC
RHcTEU3o4bMnQE6T4nuXqJZXzGDFB6KrrptbRB3m4NsjPCB5GYdye1yLgArcmG5q
zwWkpVANaodxp0V3iDZ8tmgIkU6pi9X67Q27G5p8XTMugyQFtmChmpTW5bbgLltn
1r8DrTfuQe2FaRG51FyyhePCgG8myD2a4cf93vRG4b2ZNPZ1rk+vwtZshVXtapwd
imygN8BTUSdhfSyFE4sivOKKi9HoztBexgIG41anHqloCZyTYdDaUR2tHxeDb7sl
mthQPa5qZ28/VfYf+Oig47WXRjyXNDgCG7pWMcSGSsUB0PTYre030lBj1V6f6kTT
0r+oj4iouD2jEAmGr+OlJ24C+AyL0LCdp5BHxZ2KQysqCkvXzODDyPtjoYgZML5o
1G3+C8bg9oThmyQ6/2/RGPCHXKgarL99S6x9ShQJrXlsR8k3T22+NfiFfu/UNhbb
/VUCFo5gLbP+PXlIXfKmCvWje1ZosbEiIzRmFHtFP4W/oA+ZcJ4UEPeje2M3VQNx
ODlbPUja0oWIUWftzAQJCaUdS4gfTSWJTGxpQANQLrwDdttEQk54lKGX9qsJD7yX
D5ICL4yyyhoPk03VSlz+4ktiCwK+Ss3YPkXHzMApbj47mf0pE6NwanFtMyPIJjH6
qoNYzuKCp/3VNe9B6JRiUW/+ovay6D4Mzdf5p0kPEUb5wzuD1EmFEX1G3thhHngI
KZSl/sTp6oLCOPqh3duqSTSApNAL5zRn0ZErUKYqMitfvKFDDTkqXf8vglLe+m3H
LX5MY9vaZfjtqKo80yet0OYy6N4BUbm5JYyCFbbaBLNx+e65BEE25y7tr5z5Xxs/
`protect END_PROTECTED
