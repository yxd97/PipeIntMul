`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNOWDDpvLN7FTpKNDhjF7p0uudqTn4oSH2dL9MY4aZfyXjwnRv6VO0dxGsBFZCEg
tnRQ6iCP+G4bQ2bhlgAtxtYHzyv+QYB0JtzgGL4cbANHzXmihcvcSjt5fZpg23k6
e+n8/W44/8akZRmzIP5ypWXE9FA2ANi521iQPv0Xe60C2+zOzuUXZyPrMq/0Vwda
TUB48R+mD3TqxycZjA2vK6fwKNwg+NrQsF0GpLoXn4N0SslMvXrZAZ8FTF3VKgEO
Aj0E6Y3VBPTBLWyDGRtH/NH6ntUWrhAoJKhXc/BIsjsJupdOkoo6X2V+qlCE6+MB
NNU8wgqw0b8Gw+mlbVtSl/4lNCywXc1ur/RGqWoAsPFyoeuhU1jK8YKRP86yDf0C
`protect END_PROTECTED
