`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQ3isChDt0noTiuauQmZu2EiL2yetBjOxu/Rexw98Exsln5PIlxD2YTrpyPTq2kL
V5+N1CVJFD6Sdzb/5gvVK+qn1R6JizYd+VHjNbxNHVhHm00A64gII+m71IRfkkzm
TpeXkm+EPumPwJ/JK8sBXaWZp6tWuCoalQHAdRlSa/1O0CbAK9ERm/VFEVxQPtYD
X7B3UhBhn2erHasfHLHFQu/iqxqV7NbKBJuQvuK243MF/cz0CBv9iEOIPH8H1A6J
WIkXmvT3KL+wz+fX1TcIwom56EEwMfGQGJLDIpV+8cH0NoVE/wBl3HmyFvYVIC98
J1LPvMXbpci37hEdWKilWhf5s7nZz5UavCEOIlfcbGtH0UG/PqBBtAeuZR2NJ8Xs
LAahMxQcLvKE0uMPZCo2MM1McyD2R5F6kgU5LHCfFUDmQcxx0DfgPBkEutaUBOJO
5DIXykuOBBLZDchOMhVXk4QdM6noxicYJH8KZUu0ddGfDJJ41ox/dzkVTXFLHw6g
6WdDDwEOw2PK+7OA6nLF9MYCFDlvtxuwh+zFleQbnhMuoN3INauJbjh00iv1+Zg/
muxxL+HHNZcgRpWLqKNMQx3huvSgKJM/+Jpc37+sdVyFltdrl7qMp+sLfdUwSz+S
6Tng6ZXBm8yE1LCTTPmykOJPc/0t1OC77YMfywEcJgA=
`protect END_PROTECTED
