`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbW+tN1I6+m3cK8BnFlbLQqsspfsYIaY8f/geY+sjeR8Qogv8Ao21ZJIB/l4y0G4
BBM53LjR255CbuLigtyipZe++5gA6HkVK47CklZwiM9fjiwXy9Be69j5WlOH68zp
dEWwIYeDXNDB8iz1SCCbXRmSj3nE/8m7JJcv5Z0jGi8S2uiSZg0FXBfjcvoeEB8G
5HmofiWYMUrm0XMyuUEEDsOCsIVpbIsaaN8qpqQ90U9PA0MMrk9DzAkmSFcTKnp9
FAZsKswS38Cnwo8oiDJU90oXvZRpBrP8JROZX+jAiCbJap4EuKcOBglfLhcFIviV
d8b7cebdO7wBrCEOF8QGFwtLLI42F3J9bbxuZDu0+pxcq53UJeup+qw+oJyHuONV
gqvkh3zgy2OAi3XRvuJ1XopvneCsyYFhrId7ZnXqRBMlp5UeqJjFYwDhgFG0Hgrk
S9wWFornlW+d9i2qTyNqzejLwzGdge9kM+aU7pRvIfGI2tJRsWGimvKPK6WUuZ+o
4qL8PauzdigeVyxC5EEpJfUBrn5n67e9EJTxpOMHSnc60TpRw/+4ZTkVC3thbjG0
UcsVwrKuP/AiflZFw3hXLqH2Dtew88p6neAFREuzWUWHiBipSSxP4HmY+neNGwq5
Hfp1VWAdDwQC8no0gMox+QmO4wwhYJuHBTMUvtaybgAs5YImu2w8l0PUgoSo7eiY
ULyZ8O9g2xVjCS77mRtnlwbeogxUiE24Vka+czXAxWz7PXTa7SfhqwbfmmW1mpbD
F14l/v0AuNDAyHgSd37Dg2lSTmbrAmno/BDr8Y5mckMMd4Xa8WIr+xwF8BA1JPiP
M33EWyRSkAsSgZTKe2xYI46fS2zpwJjbyj1fF45Yujc3TYsEiCh+nThNpgVNHR+t
6SRTqVLNqbWdID9PWQDqib772ZswGzYUuoTHbzuFw9vUJaMfjF8rC5iDXpzwZSil
qhc2DN1a0hXPk+Bp5Ekz1h2f4AGnsQq9Pk7fP/fMUxDckM9dOHCEXqT3inx4LUHm
paUpKDA4a2WzF/AaLtuL38R+nlTKRUsqhkfVEXKCAZxAUaMwYqKr524u/xZ4Jx3z
f3crDUui4hYrchCacaAmS5jEFscI5tEiL6lntBeFGBvy7bzp1k2bI3RzDBR8MzLQ
DdoQIaaiQ66i49RZOoZeZ7I1tEDtV0NL1jVVssT759BHIM09dgzbHQtj4h+s1UK+
asM8GXaT6zSGD/53T0ObxiJOrGKAY+ftxEHeI/RduuFAjvomMsFm9RAH6l9/7AL2
czZmEM8mfrbFrlbHYMkTi8L1qB1L9MUIqB5bbCigMqA1FZ+LuEPEn0jyjNFVMdJq
VC6z0zLNiCn+9htyiwOBBg4znAzG6lhJLC0b3ydXdCS1J/t6LPoTJypHjzHB06cN
EBd56Gd3d8GXQ2BezuBMocgX85gM7eX8UfOfn72Cj5kC9v+e/2DQbBYDDJEpF8D2
k9NKndB+68dpx/w33Rr/3gF9NXcjSs2kB+2fwfW7+en2xfG082BdsXFGf1ThC8B8
j95OOiXihYBoZxskbzUrWJ9qHd71IiiJoSnNicZj874VryoEQOsUkh78hsWO6FQu
kvFrr5rRl8sbM5PSsF9NbB1QaBS51NNtpmYzCe98enFNpZJc8MEvSg393PoAqI0F
C8f9eemIuzoIfofV5q2ZkRRL3ZNqFNmX+GrYc7PXgqng14PQuQZOBW6zMe/hHYtC
3DCGo8VcfxSylq4ZkQ0F0HImvyLtYsFvj9zoNEvKxY/WGrmQIUaLphU1DYlQlq3r
JcBM9BZ6hCZhNLeggaYcNW3iD9nvmsuiF4d59InPhwAvAdVQY68rGNV36QJyPtDs
ETry66biJntEdTvNV3jJLjkdzdRw9rh5wrlChQ6C1Tb2VJlfjMVFmnrLk+QJ+NPl
DxmtSWLe4k+ShbaWPUYmw8deMq7yfhbD2JwzFRbUFzDFvDElS9v4sCbfQaZbiwAh
5XDk9Oi1ASUB1FhAJAulVwM9vOLAy4FVH0pA8wIp96m1Si7ZYvf+c5BXR5V6JQ3Q
QIL53afg5Q5b15B3xrpbgcxsfBydwrMLdanatgpztJkbv1OygVBFdH32Cm8LyVRr
jw9EFnCt3JJVQfRP7G17ktP643RT54K3WREkcPQo8W+z053JSliB2PkmTO0BM8pQ
N0IXZDErAPtfiuEAjxgbyg8nXpS/pPG7oGAslnRZH98maUi2TBt9TAGhI7gt5Yr+
qocN5dNJbv+p6+dYS6Wrda5cudZD7YJccitp9+9afzg=
`protect END_PROTECTED
