`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pa/7nCY8ZlbrlfczH0BySReJiy+eoIP0eQxi8ZaK6Yv9n0mFAbOTjsQyl7RrpV7V
qF7glWlF/QrhLVaMswv5aaSsJ+HYrJExm7fzZmdhcz5k5yWsdJm4+5rXgzbd1Ct+
IRMselQdIhPtmkrDR4es1LVJX8A66zFRAPrcsASSgefrs5bcGlcVg2I2sRJ/pwN1
9+UZVlkvC9en4XSVx+/jMOnIO7AYqLjVckL3JY/NFIutY4L1loYjMySKv+N/glX2
LwNpuapXQwgbyHtW+pEd77O5xdirlJtRjyP+BZvehlFrQ+kCo0sv0kFbLggbnudv
EE8wTO2bKP0WbBh+QKiAxA==
`protect END_PROTECTED
