`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/z9mt5ose4jQxwPPTWoi7gLpFp1nhw/w90wTRDKXsO3poEKG1TjtNQuFTtwiSYsx
o8SRVWwTwjq1glZDfSDyLq9xwQbTmBP5tn1aZx48TDmIBRiMK2Q3zxYI/TsFMHIn
vgU2OtcMRjr+40ntZih6L+mMbF7w44beuuwTl8mU22EemOJAtKypFRpmUQAvZYBi
/T/t9X31KkOhXlEb9mQ8gUlgJm0itt2dl6/0LJSffMeFJ/CL5Y9tl66Pw+cEFha4
Nxj26BA2ky2vkFih1sMlGH/z26p2PXpscW75EufzP32iejicnMndvWy4OwhcomI4
JR0zjCxXANK4oUUkdAYl4innLOSSsleqMdmfCpO2jCrgd2giYaAa1H6w4X5a3HRs
+IpIdrYCpG1KR0KdL4rTi2+NDpVkoDqIe6Z3B3IDdb9rbf6CyFbe7qc5RgmD3jhz
YVZJc/YXg2pxWAOBnhpg5HoTwc2t8l1oQhUe8GmqfVIXKP8yIXudwGEIvVm+felI
vypqMiSVpzjEapuQ5adv5NZBItzOcMPjbf582+HZiGuH5mNU4YsGo5I9oqBzGgDI
Qqw+zpz3dUE15od0tydXFcJ/KdLxp1Apfns+TFlvKedo9VifqJE/JA9Gb5Nae1tJ
hoSgazbR25qiWEf3/cNTRoTrRHno0qBrwkaqZK+2QTVaqJQt9dSacTWilsm/pDP8
rZOws5RO4HSIFumzJUG0lfoi9+/E/4hycLLXUWGiAeIsiGMmkn17/C4gcyg56KWU
`protect END_PROTECTED
