`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1pT0yBV0PQbevuAGzpiuaPElHXgVSkaNvdix6RYbk7j0NzlX/JuvUEBpvje+8lH
sAJA/RNslNWCB0g1QwAOoCVYTOVUOK9WMhRCWPddJJL28r63owzSlXy6lq1pxENZ
0NELNBIa4WO+XjGk88s0u98XpGNSDGk6dFlfJxAX3EMqhSCbTeOX8J1gOYVlBQ2H
YTECWNEYxpx0t09uj4x0FsJzn9nHzpdvYw4cZFIwvVx4tfql/ZTfo9LCTzAh7tM2
7xQuf6PAOGnNHa3ZTXy3IYkz8zDffpEw5aBSzbYdf5WDjI453mHbuOxkbLKZrX7M
1dOiPx7UffBVjLxOwmeyHOUyu1hbxBfLvvfPbPG4ijk7NxVjT2VI4oo7CgGjwlNO
`protect END_PROTECTED
