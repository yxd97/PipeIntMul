`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eq5umUO1n16xQuGruAZX24mFm6pgfQMA5xLWwsppn0MFbLEIdDuzHiDEkx/FkLep
0JtUUy35zBPETHdfNjoX0l2s4UqmAQCT92+QPgAR5cFkUU6akYUKnXKGnmGfpc6K
nI7FeKCKCczmigH5UQvetIjtXEpDdId7Eric7dCZiaJX3Cia7px2553myqVKyASo
zAmIPPe2wAoFRw1x+1cC2B12WifJsEASRTh4xIW2IK/mBFUwB71Mmzd5v43ruLSV
0Ci+PQ6QAD6oNkGLNQrR5/9jpCaJLLTVEGpt/dZNxGw5cfxXJg7dKHUG2ELBmZq7
oGBJwMVf4nGXU8opGxH2ByG3MYa8uERjJ3DCunRfDvwRSCZ2l2gDVBzKoBlkEIxO
3iYoYubbdgR5cmizZiSrCugFM+KKoliRx9uirDNT2CZL0zqEnPIfADICBwSZkC8S
CfaDbKPovSZhouM948pQ4/kLdlDWs05KOk9O0wEirt4mEX7O3Q1T7HxtR8GPLjyQ
EV0SVuyobVqRZeoJlNDxCzWNqh5BWW8Yywooy37tvxgIN1xTpASmyIYGuJnCZgGD
e9en4MzuQy1lo9k4rqBy/XufhTAIFBfkzlDxBJsAO2aqIH2egC2IGiN+UHOgwMnH
ArZ3iHGYQ3Qd7nkkGi6audUSeBLRigCWy8wcwS1XEpSFozrH/IIp96BVAQOP6xRS
SPvdNQOuGi9b9wjW/63+00SwcwX0jZGnXW7v07GQZPyz/2bTR+PXu1BwYETfB3u+
mvgnuj2L7YR3NmnTufx3Kvkhmd+ikZgBbgDaQ+qcn6hbm5Ifi7tHRtz58nx+y7vg
U7tVm6SfmKZFFd1J32Umr2FWfmUNkr+y4lXETzuUuVkMrhJgmgbAZ84VgjcJ2AuQ
d45yfRNfqpHzpQiytRIdEHchKaXj9IEZDi03zk3mJqPuHUVt78cwji2QNI+a9S8/
3SWjeCYbvJly6AaCMXOzozTqVgC37B2DClxphiyVMkqZ31IkaEX/0GR81PsvcG/Z
Ny9gGwRWP/KjNL4VqsFX5cCLKiYK2Mjopuse5Q0g5DE3x5tJJZxRfcJxPfVKzqRN
m58CVqLK58QSdBOsUHIjmzYuJG6ixKADOz3W1qNm+tjB55qswJosx6DIs4tUcw48
mdczAyH19TD0rRWd1kKxC39IGX9Q/2BsKQhyw5xJKivQ/gs+6spTEj/niX+RoqQ3
90SVQ3GbgzeywydF2Oh1YfbskL7S+WRVnr+0aLUbwuMesZaWyzqEUxE4Skg11dC+
3H5q/7N3AEzLaYd0jOe6dGFkYucBlVQtHyx1Iq3PPsnPZ7a1Deucpi7Eo7Bu97d6
t90hJfGUlbyNNnUUnrhpccnUySN5t9w2Aop6lHR2Z5EqKleKX6RMnfxyaOP3vzZl
UXLsU+I96Zh7ocp1WHziVdwb3sAsr6DRH2kblCiZjIskMVa+yb4aIk/14SAPOdAZ
29OfhnuYM+DKMwFd2mLsaqycsnL9bfdOYE/nKaIEg3yo3RbiAouVqemesac/jlD/
b80aGtHr2GYari1bYuA/wXdHNhh5jT+xheF1FOx6T3fusJYSM2KsTG23yObyXKF4
pRice0SKZVgjotHa9zwFAN1uxTVo3uoPtp68xsbqt4oRcXK5rVKhIzCfUQvs919s
sZIxE5PbsMCbAYq1GS9e+nNO0uPtZVZ+Zs5lNgdxgx7pfN9kcorKmTPFhhbwvN38
9RrZLGiUd95mU3yNIxh3k7vwnrVXBbeL+QWK6VIjkeJEgKPoaeMvLkdmNLJUq9Si
ZehpbQZ6jt3mMbubdQzVpmaMkcAvpxs5lV547IckUpD8IKKI8+C1hXslRKePmahE
syGHa22Q7KUC9sPICg4xHgxtxFjrVjASzgL+AYa0+bP6CKAKL7QKXH5N8iDbYwRB
Sn8/TJuzvTwmtB7x7lwrWCQrTNce4ff21iZIN9Eqvr7cXLjzfFJPWxK43Oc+Uasu
57IOJSu/LB+XsIs89AOjRinUdONbamf2nV7IDAFuYBS+QlNUm5dwX8SHkTRb8iyN
vBP3ZMIE8xyIKYby1CXOuhE3XdtdoUiqxq4eM4UwSHbqG+ycQLCklb1C3Calbaye
eqXvsIJGUoEHs04CqTYrT6KD83MyIUcM3+VSMHk+ch6StqJxGGvAoa0rwFbT8eaS
daOHNlQfJFPTdh0Bh3+9dNCD1eUnuruhkrKmzflnPb9av3WW67qNH5Jzhhn5n+bt
2NCUolZ3sZ6r6f/GLQR+z+hVtndC/cwEYvbwmWrsjaEH6q2IJa4Bdw8ls9IucWhC
bXO9sBK3az7e2W2VBFjTnRvNuRW0b5QP6IcMt0s85HnhCKJg0EhSGQ2pVLRRGgVV
Z5d2Wd4bDI4FD68PlMgoKnKKkGoe/+RtXZvUakXN/EQ9w2Owxsfx0W5AqhZpCmC/
vxof4tL2iXAhhzcaBvn0c6WMxHJK5TKOsWbDSduVBPdFX6wHDi4zEETpxK6c+1TH
UkEX2Eq4f5Uq9S7L4h6xf4TvbVE1jBQC1pxd7/VNocI4QCxS+Gd/HNKLFlshPvfm
35NTiGMlguSQiqEMhXidvjjC4SgglL1+JXYhE2hvvTp1DzoYI9krDhS2ixHZ3KmQ
7+eh0dZXHeGTpQyvy7V3tvP0cZwPC6C3Yqe+U7bVuZhBzEPPAFZcKT+hArdVSYxP
BAKXEXlzBe3Czw08HiiJ3HzY8OZ5IEJx3m+0+RuZEag=
`protect END_PROTECTED
