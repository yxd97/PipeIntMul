`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bo+6EP5BBXx0OfrCo+0nHKJyEkJ412zPGTT12qM+kjEW4DTmhLoNE1hPtsW4/1AC
F3W+0I/AMM0YBCFaKw/cKzBBJW5HBsq9HegFrtr+yJjM8th6RaUPrAcC9wGKc3c1
c2s2FItb/CVXOojk8DS0UMbUkEf0zccPmsXL3pn822oz5pxycO8tROc1JNYlt7Ne
pSqdr8iUeyngjZbaHFxjHooYzSRGrnyGd3z6nhj4vSiNbyI6QxgiFLr1uQXFMLPs
/6W5CgZKIQ77mFQYfD3Brk499oNGRVZGb4hIEelf3PHwfmDTdYkcX3oe+Qj1Q3Qr
3jlWa4wk76afYIJ0A96mp+agTfUHL1WUHydBjTqyS3diZSmSFiHhcDwFotBYAS0y
Ryb4WJ8JRNteJWE/2l25brRFz53dwJSUz6qVmq/Iujh/Ljcm+ESvyX2Ar5+MJief
i0eL3Qpmh7MeNIVpkRv8c76R7AtaGSGnfW3bHbL1N4kDMKoe8sHeGaG5SvO4uvWQ
q9scbIh3tZHH2CYStAEjPNuEE+0WQX1NEgGg5VxIPIiv/ukXSgy8sUDCsXuLHVBd
L9nWH9QJvsnM63lpkgLBCKS9uy05JAQffyRX+W0YA/Y=
`protect END_PROTECTED
