`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ByH3RHcqy3h2w4EqBJYbr0B5Y10hV2y/919vTxrNEqGDmajCM/QUgtuN7xZZRkVT
lKDGdsjrFU1Pmgxv3cTzlrxLcks9SZynSqmj4eRGfvSPZvwoDP4cGWyJN0akJae+
yQ81iHirf4ov3ssrHXDapEI1ivhP/W9pcU3zPSDUCPlPUgs16+mh5Dfgb2IlvtF+
WioALsrrS07bLe4NPybp5DUA8r2Z9l+eRHEDkIuDXn8oar1R8/jayXree62xtbCn
t3JjtZcdl/1OHiIeKz+/h8KV9IzfaJRdT1tSBHyxPeveCjohKajz2IoYH8P0X8oA
IZfuzYxH1v5W8K4dp4N+vQetcM/FYNZOs50XG6UDlyQ=
`protect END_PROTECTED
