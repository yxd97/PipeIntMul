`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
677tQ9fAlpqqJzcwFC8yRCwATqdsusbT4EokyZTK8O5+F0fx1TgGPcWkMbuC/lH2
UY5ZWGl+sSVyflXPKlmNLm4gvqO0FRBn8cIgvgfA1lDq2A5UFJe2x6GyMLdQ/ttF
Z61ajBk5eLVK20D3OvL5+jpKw8dFHb1CIlWp3wqcM8vud7f3+7WEiS+f5LtzVgbP
QzkgWyUh5YkIz2/xIq2L9ld6HoGrkNM3fzJbKBtIMsCFnVTK3mkzNnPSNc9Cg02e
+afmBxIs+nCU72BLZ1du3gLgCtrJ/D07u6XEcxPuSPVgTl/BSAUum6osLiuUV61+
aUEcDoxsAQkM0uDfLxNQlGe0SUYcwYwe/HimK1mR1GdJUp4ZhE0PYBDoCOamOjwv
87QcO5rLpSbOoT/EVHPyj4XI3F5QSjYyHZ6NM859G418upVD8b8190A8dtbwa0wo
e1GgT0v/RsFJRgndywnmpfqbZ3UjdOjyJDzPxGN0DEgso3RdTkVDWxcQlmxmo0xu
`protect END_PROTECTED
