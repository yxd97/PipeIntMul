`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dbghz5tfyfFDuIY8WsHuSyJdbY61V9gnhz66YMQFW9Lhe0YnYXHpb5P0JBbXVJ84
sT8XjSZnDsxDMl6Y6JK+UzOe7qFLt8nn7S5cprMLExpJu5YO/5fpdCl6EBca9tt+
AwwFWF1ZRpHHHS9L5wZBGxXzqs39VR+CtGLRRj7eocX1ZlURMWpUSYYwvjypdoIE
Juym7ZxbCuJclzUnZZwKvSxVb2grjeKSbCZ4qeDg6DRWFSlqaKAro6Rqaihh8DSm
HVBT7k0cZ+7zxZ9yEZCrOw2tFDEkXckBqP0Dzzuo4ORxg4MdF9QowFycO2rSFSLr
XeszPJg77EuU3qaQM7ZYQA==
`protect END_PROTECTED
