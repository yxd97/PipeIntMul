`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n2PnQVFNQeygZWOWbfQTJrZXOgoI5L88wiUl0ybya69ypcZ7OLQYWIC8vFys7ZeW
nZODKo1CpD91awvYuAWYaZ/o/6SpDHOpbmNIK2Q2WB762IF5wIrO8H/3RP9Mlbrr
C0dOZOiOiF4qanSnnpDNHn6CYbx/B/5/qpbZqDCavH003hJMos018Dh++0cHj3I8
tYMu750uVzQhdtX4jlxzIWxjdemtNTPDGOBrboazqOItrHugCUeRbzoNHClEXMXV
`protect END_PROTECTED
