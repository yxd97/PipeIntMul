`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nm94RlQzbHvP5kuzHtcUlos0c2o1dZWO0tnLvewWu/jKvRRVGcqMETO4HDQuKnFR
Y0XifJEkjWHfOyDEKgFX8l3FFkrjJqqw2zLUSB4tLZxi9F870UmK5M9V9yxExdga
caumnuhh3xj+wBsNYdvsXS44t43qHe2EwLC1E1n0JK2XMm/GWtZ4FwBgt8i9XOwc
cE3PCrQA0ZofYb0tuKbgNgVTTRGxv6WiZzDbPdPJ9KbEUYWa4xKtId6TDouWo8/n
BvrcbD7PdfuOvLXUsabVHvdaCUtHaDqnwNBAmRV2qOhlkDD/RuIpNCoV2uNVu7S/
eN4qxniaDzlfOusAvCsdvPylJm6zTUdbIqp4FtalZu99LsU3hWDvIG6yiFNJLYIb
d2rr7e5mDSE4lPrddzl7rU0DJCXiCKY4ama/Gh7M3Xs6hJ894rzJ/mbZPmsWvPU7
cRRxPffIqF0IyTaAGt5/yd81WwJz5SrsdK9LMGCI3gwA0ZcatXtxrY/JOChElicU
SupzI85K2OBLAy6JDHZzDx+6o8X4vib9A7wMCB3AeMk6YCwKpEXe56v4FpAUOkJw
Fneldohp88+IL8tfiEl/xRiEGC3OTPKDpk6AZYZivOnNjpgNP/bQByy67e1Hzvbc
b57A2jk1TMm2O4SvFY9gy27l7+5nyvixmQH/FOdr6JfaNgJ7j53bQdOhPrPzjusV
zK4IuzqqknI9g482wHo6j8RwO2Qu9/Cs/jlzjxsnjxBf6749D4Vrx/4GtcSyJet5
BQ7DPY9qQ4/DvsNVRz8SWBIoix4S4LAmzqM4SeDd1sSuzFP8Kzq0DxxI71d7r3mD
IMoymi/ECGPWoEodIeIGyiPqOwXcSiqOBlC5pGjIiw50Qt0OkAU8EDVgE55gzG5/
`protect END_PROTECTED
