`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OsbvN4MoHsRw3EHdVlBtgIxlYufmtv6NzKU8stUIKxFYLKLVI6PLir01UDOVEvyY
vu0gHFwPaB0JZnyk7KCLgeExoQWqAEDiwzW8rxgXRwK9WDcBCVge2X4C1m2fNbJg
u+znYGqJ3BI7ocYyk+lVaBQpl3j4YVhV+9vF+YAB0HDwcqRUmft+WRWdipgRrfUP
HY+8bC/msNFAnwLvqMk1Z3cY0gegrdtKC+OrjhNuU8NWWZ+82w1tLV3klogueUBX
HmYo4SlHkIi3bO6rKlnefXBN2cwtyBfM2RVYicJEr4IXSuCxEYLb0lEVv49HPlHm
fE52vInrFApvU6npdbbhMTD0XZGPL6ldUvzh/3E8Y/uXTSbR54Nlg6knaezxrIuF
1jZLzNxQqfoqHiBNMvMYtDw8OqlELFNGPqbZdNZGgY7ybQ4amGqids8SGzjrjyZ7
9V/hB73l2JQE/NHRUw0LL22lE/zQNJ3Z7N0+8W/zyz2hMe5cpHArbfbzIPbQR23H
Hwl4AZQtCoXESTZBR7lJ1zAAqmsbdOCc4Nm0HDVXk9eWqNFoKAUMunVsVAcnqVUL
5t3iDaix6mID5odG4+jPQ7WwSyInVRmDl/3zshs19klhMmqhbOm4DfM0HPxGRaEQ
kRoVmYS3xF8EY7rCZ3f1so6SXLixDpPJb99kiAc6fWit0qLMQr5AjTp16LGhvVdL
T+PeeAGPm/jBJyKd50h+pU+kFZgk3A0gttR92bk+uF9R9Ojh3WwLdH/SHHJaSJxV
ZN0//LXbOSFmFk8cpv1pwfigRnOj+H4n2igqMyYnYfwrBik2yQ6/uVBE00eVZpIR
zVxzIvzbYTZXtiTC9EdYVPFRs0OHzZJl538wwe80KAFaK3u96dq9nfDAFesDsBlY
ZQJJWMZAFlmhX5qQJ0TBuVL0KE2S5pfYc5WXJN0Nrsi1RKb+mPaRZRTpT5xsRbPV
`protect END_PROTECTED
