`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GuGN+ORla8FOdgViKdn5Gn+HmNYud1ZNRnrW5MssnDdCwF3bo1X1iayyrfhZN4w/
m3k12cxvaosUkdRucsCo2+35C9hWY3+fgjNqIYdOmprOibGFxxaei2rCLwOikbxD
85vALLvVVgokKYYKxrg/jkRo/d/P5Ihlco255w+xvVkStX0TtG++hjTqIZur0Dv3
2YlcQo/repCnhV85frvFf3W3gb5SXBtUsyKttUvRxYh1mxWMl3yDTPdQjOooBSFs
wsV4mgs1Y/Iwjau+InPlKqo7bbbzD1fy+0dSjH1UyzB2oIqlMRjs6crd9NRczOPm
uWD0lyfgtb97+3CaWoQXKibmjy/n6YohQq41HvFHGU9XjnGLp4tYIkBeBLMb7AGH
+EPoKHnI8jySBWqQvjPPb95Wx0DWHcTw6wvWA5kypDi74JW7iJ+7lgn0//SV0WZe
+ZkyAPHUfM00LRgtc4irIfhMnjOMCh9WGk4axBfQPygcd8ox7r3qaBAaSxAPfFjX
I6JOfkWZ8ByfoB9nHkcZZH4A2XnADpgGIVHo26dSOElr44R+FiAE0SXtteezQNPG
EylA+J93bCo/8Df7jEukz5JS3QX4S07maEbnLWBxcNk1RlCBz80/xI44N8HLsASb
ACjnWYE1kMpwnkncdMVFQIP2BrTHrquI0Mj42VrU+vCgOnCoc6hafxJ9N9mdkeUc
7daajv4Po+TYzz5oViqXpeTlOLaVroWt+ZjmUvC05GxVZL2xkueKDoNo6CjQwZlK
1BWHgANRRCz9xM54jtuRwjiY23MBsTUfguvnHgRh9zbNXT7yWNE1vgc7SYtRhBFb
zb/50Ff4Zo2itwT7AsDYE/I7cDX259OySffsz3ccsTxDv30Cb2jM/WdUyKqUhGwa
gDsdeKo2YgTRpFkrtGKQ7thZfWWu6iole7clj2f7zqCqquTjFz8SCrYe2qLZkbQM
dp2022kXevkDqB/nPQKB8fWLsD6sxlwieKY9S/wkcwc=
`protect END_PROTECTED
