`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nZgRX67OA9aupmZfaSnyzCTVMNfWNcgr7Ei9GCTVMq9NvYTjX4UX1fBnYMRjwwLS
de6he4+sOCHNSOgX1KOcfk9FqvlL/t1qmMuM2YQhOtyCZVvPGEGXHLAKMZpfYKuu
1jGeG3EAKhmT//Xe4CkCOsT/UnNRI70DFEVxStfuIbH8SM7n7SdY07Jv+yjMKpyi
Jl0xz/absFPYmdkAQBpyzj6t4VzX88OXMBtW2FgPj1JK7po5R+ly+jJ0xd1djLEY
ym1GJQUFRjK3Jbj7TG2PfZGwOapkkukwlkirhFHUNC7LBlekjVZ36UYRKovOR77G
dfPASFeqgBZi+486lrRxydORcXTeWqa6Egah0Z4m5k2s/0JH+a3DCoI+AOtHzccI
q+IGqVg41bo4D8+OZZu7kHoOgsFg8GLMnmfo3R1l45YYS/IQd8Hw+sjIEiJQgIOv
`protect END_PROTECTED
