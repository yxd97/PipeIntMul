`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcZeRzTpj7GDLHX3rCaE8puJbY2oe8K61nJy5xZfi4V7G0TlWPZhvJN0GDwpvg4F
sDhi7thVQUm91HYLy71M0FvZy1QO/auN1lBso7Mni+kSmIC+roGw83adIhbdJatO
dt2uEEOTLVCqs+suH8aZcmwpRb5mU7JCzDsQmZiGbwUdR2CredQ51SF3PYa1ZVPX
0mss41F0XezP5OxtD/70tKsUO8gNDtrqrko6YfcXMSFmS9Aj9xx9Lt66GMBwdIZm
az9DjjHlt3aARNd/NpNXnlZAqmPSayAF9zkoQR9STVOW2Za/5m1bszy/9X0PyO9q
cRdBeYGgiZkxu8cDoUIIbg7uTI0MlfT5Q70n13ksswqNjwSwMl4Zw6tdLkm/OjO4
us8HgT2hN4fVYycrX4xRdkRN5D77328q828CYqjPKCa45+shU8KhDCLPtae25qXH
`protect END_PROTECTED
