`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EB50oNyjjx2vyqAnOuiwLpKeP9fKXckJ75I4dwCzKL90YiokWw+LpyKQIJgAtF9C
ruOgdl17PopG0k5flYMzj+uFieAdLYSBqszyL3+Q7psJPggX4D4HZf18r5ST17RG
8/yfHWe/4mGuogsbXfWTUosMAL5jhqE3BANKRxYFNUmDNpvDXuHmRZ8QkWXMFHea
c+N1q0UeUrbgbowIZL26M4YAdUZKDldBsN6XlvDRvyAgHHhKD248iXA/HqVLe6a4
IX0qeNM1TlV2eKydegoSaoS3Q56yaD/oqpsj4lXUqU1TJpV4C31Ci1D4/ImbqddL
FeQ6631uStjZv0aX+FiEN+/q65A9h82y1o+gFq4mQFCLGM+YwDw4RAJHy3BXBHh5
eJ8lOiVLRos6Y4tGYV4cKAyaxxhb2LVvGHvzr7DntbUy3PpqImLyRM5QAi3TC3iJ
rLZDvg5BaSmK1v4yeKoSfjzKbmB3AihST4QSeMb02TIbGPZN7KgTSTklmJSjZycn
gUVhDMlzakZ+xby00YDD4U4i7VYEiquwTR+FWiK8wTgr5i4ShnYjodQDAfPqn8YU
1SjWmmEgeALHgWxKqv0p7LXNcOQRrEQ/4xZ3asIruN+ivaKUx8Jjds/Ooije3sa7
jenyHBZ0bN9llH6TlPzjduFBZOmXDWOXdShtM9wRwHmp0UGj/I+gTqWFmBOKRFnk
C9fY2g4XxDTHAzFwIobOR8nxC7c2RDjqscqfcpLj/NyIektAhrWqQ2tQnbCWZRiE
AV/Hx482gRSNALm83vt/wLRAQIMLUji2fBInhwh97Qv90PQ4yLQygPAo52iVvMqv
tm7VJ4isw36EJyrdHMKQdvjNu0SvDCuz3Tg7mMEviXoGKoC+HG9ivqeQSBva80w9
PT4KA2MrCBq/heVgV3ZZgbbNYLZUfic8M+Bo+4h66bO8sm3PiDwnst66VJFbWXG4
htm2x14FtCTV7n4iFnfqtrpS0T+GDn6BPzjVcRlqXw7Utn4v14v/F5itrcSsbQXG
w+c4x9KrXpWhdfxwJi6yFV2JDqZU7Dw2xAZq2MvwV8Y0bBtaw8fX7Yv19eepwgr2
M3jjOv8O+dik+nxvlQ0wne99ZF1JGiIV3qEOJuYoYnh11hsOuuExEmVgOYCKnq+Z
y+xy5w7VUvuJUncYvQMbQQzlaLbBXq56oh9evdJDj/+alnAsSn9Efs78M+ZEaTh+
YFyaXZ7ZuAh5pTPH/IrlZEbfMNCzjZ94p8L/hdX7X7uC3UBR9Vp+BF17IthCiGd+
4fH9LfXwBVK3t06JQqbLM9T2i9mIMGQlnWwd5PWyFBhGhgy6+6yNDmtHBjg1uD+X
ILwsq+aQ2chQVtLBgP80i1COlVpxnrRuRsLykO/FFQSHIKigNhkQE+bi5iZnib7f
MLO/vnYnfkFDldwggwjYvN0xE949R2UDqBjKuqKmEQCbVu95snPomH86yDikjHxD
gj/rHp6/jg6GgFKPoa9MZwqupkhLdw/gawF/qQQHPIsoY2ijujhsDUIZwSnD1wBw
aQwgXiOjzW2leVvRayV/zGC6E/QkDeK9rD1Zo/KlC6VT60/7LX4oENaTgroowUZE
dDdtRqxuwGFLSS3Oi/uJsyHm3gSvx+Umod6bt3xc75aXkh21ucViNhWjkPgW3fdu
bPiGx8uwGoUTmop+3DtyYpBXCVBZOVDoK74H4rMMictk8abYVxbCW/4nmqCWJU3+
I9y3XqGvu4pqaffDfEH1lZLEy23Z5CinJ8hj0SBPxYhea9ODEFE0U+tVZ0k0iYDj
YcQNBx6HM8z1TcQ9ONGyHnpxTdipnTj235v1JynVMl0PBxFKpaapT1iu/3ziHcLx
nBXJJnZJdpQpiGoiggPtG4s7y0HvMb5gF6jnijYV+RAT5HekNe7k1YplmxJTczRc
g36gPYgnrscTK423SsUg/+/kVeetDmgpFnmy+J+CFt0m/UluM4tCAg8dmpaRWALp
trQhVH5yDsKvRGfb1QUpz0jrD/pu8fStleOl7T/czaUEUNPm2SxxIvm2Cda1BKHt
qAwfeBqQHMfKiJxmzAmeYydagUbILBT4td4JBgDXK5iSH2YCgXTQPAc3hFO2ujiy
zFWCFIvl1HhCa1VGmo/0VT9jjz1f3stQawtO+Ozqo7xIer+tNpR9JnJIXlozjLa4
0iWCvi8fbMgTQApKT5TKPqZEE2a7iXWgf0hAU15kUqzlkufO/2HYsLtC9Eb7TtKr
NkRjmvwltmVZdOsIUzqWdFBYxjFJU1jwjtrUUcU6yg/1RBgcT70/Czh9cUyYu5M2
A0GgVMqjJcmA0iFbXcPLOA==
`protect END_PROTECTED
