`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oN3qTIvHksPtRvBDm7oOHXMDyAJ/LLV8vcUJD+oOsxjn//xuoFTbTmZoMQWvn/Rc
p2toks1Ug75Ev3/UNp0VgI5L5lRSnv/jRdT4i+2pYUzeFlh06/pUR2ERQT3300qC
XO+7Nxmxf98Yb4ERIgAHk5AGptEAjhMFCe2wvhPqGwdY2IainB34DvD0GDf7n7TW
74fCm6AsHoM2n8z04g/UH8R3KfnIHQS8giiYz8nePLbQR4wtMBEd1WhH1qwOwg2Y
BqMkqumg2jMQYJQkGU/KCtIGoTwsK3LD6E0MTev8U/FHc55hWTYTbJayCs2vf8p8
UsYAHgN30TsMcJSAqLXE7pByDQR7kPOc6zXkBKXNtz340uD59gYVKeN7JS3mvsN0
fXnl8M1dIE3BShAI9I2GNN5O0HXyBMPWa4ENXgmb4nN/p8AKXIPxCLv21eR8mnUe
+LPFyqbJL/a7Ar/iaRMQo8pLK8O2ulKVXjEGFzlqMo8aMBTQMuvaS1XXpXE2f4pn
2ab9pId+wso9qR0WxEOWOdz6xC/Ig19kES58lex3NNdz/LkdjooRp3s3tCOLKKHM
XAyLNe2SypdZWhiollSIHxCKQ+69j4syZms4GFnxOfWljgQUWRO1joTZHmAoEikI
T0Cgl+jp8kHQXhPZGNsxtemL3bOPAGVjRefp9ndcKhbmsXO19wWIlp9u+PFiJAEI
hB+BN8fUpluLAuLOAcbET0RsQ1YDtlUW1fU1w7TyjSeQa/mt6Ku+uw1NKhZzv+Xm
umISFqvHfgOvPlSV++7xHujjFXrxBkaOltRiQ+izVIUhN0s8/GhJ9Noz8q/gTrIT
v7qTK8GHUrbwX48EkOjHgjJxgDZv6QxHswtgYhbBrqqLgBJAd6eV4ju80VbopdTh
wQsH2RKhHZUxs6YmuD2S48Yixa2Bcya5m+jmtavTzXvuBf2DH3fn76ifXvsxJqDo
Bku9zamef6RlWp1oBcp01t45Rq4a+jccHeD6JILgJwFwf9E/TLBH9wT9ottXFyh+
rTVl8UvSvROGwRihn/6qeOOz8YmTrllTytCDOElOCEE+SPzpJWQWqGZurGTrv+Ws
t+195bXTI4Xc9bsuYsG/Xh4jqwZSacom4PPL3ci2bcXp7iVXsrnqPHAuHHjgIN01
k4uGYevJENk9r+gvxdFvh7ZeXE+PNQk2CvWqUFjQxxNJHN2DXnlupkOnJIxbfLLy
2yIkRMghOr/MoZsZaSwXEr7r8TB/xE0VQAI5bBkyxApqlrv1a3vuUJ5J2r+x53bU
5348uMxWc470nRF5qzoKScTExt32+QPMA1Gp3ajr6LX/i4DKSm3GBkhWunaQ3Np1
euNlu0XMcN2n2HPITLZuTxut3u1wWNvZNu6GxP+XAzQRvLB9ZFBdVRA4PiW/HKCG
3OzBvgLqyyDZoe7fat0lHCDblDmLscdoC0TGknkiOfgJuqKz+BxAacH6MN8ijpf9
Qzs+wZR4ndcJGlVeuxv3ny7kxJJTVIdQXQnCdMGUnvt5it5O2eYbmUN5mvPeR5Cn
IfePP4G3ARgwnXApsMEFJKw1uXY/TIlDBukBXNScj34NXYGMqTT4HNJDmGa6haWW
JElYqhnlcU8wDEXOSDoLGcgqPOr2FVmUsH7GceQzEFU=
`protect END_PROTECTED
