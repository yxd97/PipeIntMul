`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ngpxjGDloDEdr6kZEr5yFP7IeiDwInM18gfp3XQ5rewHI4d2Gg47Fe0cp1LQxG/l
Kh3JnZ8RrsXXgca3Ve/vaiP55YD8VJinNf+uWAtktHDuD5T2/gJhnxaV0yLQ3S6q
B01d6MT/rKvLG+0TqdPxlVfrRcJoDCmZZrd60x9Srg9N0dskryDapvKuWQM62rH7
pFbXAPeCXrWIr/s2ds+/uJGX0f562FpLWiHPXufFAwtHKs2IamZ/0N1ncORJeaPo
Le29ghAfHRmYetSLngVUvrFZM1QIPWZdbFciilSdsgupi1efMUD7cGabsfCm4NCx
4n1lL3wNbVta6I/3Y2vqWQ8RqUTO0TuGdTpT+taU5Cb7UB1HWG39w2R8F4LC3ssh
XkFGjPZ90N/3RUa006YgVkXUQRWu47QiSyzP15+UsTtWbEc/JrmI45Y3aobpPuIU
XXX5d4gGkZgHRXPflya+KBMrBG0kiwRNqjmxvOeCjuE=
`protect END_PROTECTED
