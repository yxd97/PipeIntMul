`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1xhIq6qQUDSk2P0JvmE/3mFah3qL0Oaboy/dwOmRzItqvDXX/oKLMm/UXNnIBvs
C1O342fV8ruon5jzt0nQY2TbfNWnavxzAk2HUw8KrN3CV0ZYpPCnxNdWnJw3fI+s
qlut5e4bQo781p9Owyx14e6T0y9k+wNUpme1S9i5r13R6iBG4JSZ6HHK9YAKKg/2
OyQ3eGzUkE/LmdLEiyJ8xBu6t1sH2lvLiAKuIpICtS/hrwbqfMpymXLEDVsZB7lM
5ALFAaGR9MtVM7GKTBf9ZlfsNW2zIUjGZtRb5WE2Ooc3RlHvGdZ45BNIDVP28iWA
rZ5dqV4j8O7yBD8UTYMNTa6Oq/aaPEcBJo+82ifbZjR0+pCid2bej9GlgndKV5TF
SouIbM8zoD9MStnKGcRlOmT0D3J4QyzMmTVva5j/1jk=
`protect END_PROTECTED
