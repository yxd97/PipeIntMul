`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNxj5AmGpcT4YnX83gRQWbS6/l/TnjN+2coAMdzFebA3VS34s0l/T5bsTorNHBRd
MMsgTGQz1/nCPpOlF3noi7Tos1HF/fNczWqdOmQ73zoASWQ3s9xSWDE4LxdCJT39
e8UQHbA2tT81PM+5NH+5Xq8OtpLT46NPdhBsbDp8bw05mU2VM0fNMRMiPfYEA9bb
h8KwbBgc5n1W35JuUPt+Nk75TxH8aTMabMeRtc23Jaq8HJWWQJUztZqjlcT/QjGi
OKGE5erzlAo3bdyBz5K9fs1vYjAX0bAcC2LSNTvAGWt4pv7UAeXk9iMLdcYZ/Rzc
HtvCOTZXZC2eEE5Gj18jEo9HCUPrYKCUFNGJLzO8BufhB5K9nvfa1VuJH2t9rlte
V1iE1wE79l2lHOuJU1zELYg3GDotlVD6P0UE6D6rC+7WsKt3LircFBQ9hryIosyP
xYEFlDpNfxy0bhr9FPxgO2vkwvg7B57cO8H1n88Ngy/GAhzGwg1MJ1i90jsD30Af
9p9FreRxcBZwLmNNjpJz7ZE0Ga+diFl7UFj9lYwddknbxQxZkQMsLpnzchBYHPzs
m3qOMFXmIYAx6lAgVllCiWvCQhyr7ndY29ZLE9xhyxe8xbZkRpiWO6QzySOzHyJh
mk81qWb1OGelaI04gbC0N9qEhd/5NHewZFvRnVyiBDdYW19rAqQu2Og2UDUJ+s8u
tA3x8qmEeKO+Fhs0PpyGL3NLh1bG+im+N88OvR6mKiMtNDUQKqh7CcqhkL2KRdgD
sW74JOXYS2A927kUuOzSFDOclOHjPB5fINyPjEjQ5LT50d3xcIZ9lD+IwUREQBxX
32caFNDq75hJTW79qY3vFT//XcrdXjgxuu2BMVCXdzP3qiEPqWHzlKZWWZT73a6x
xFCkSYbJDQULw4fU52VTWyjwL473HvuoWCIWTUYGGsb5KyYGo0I/x9UYBTfvoiJV
cMM80e2wpLMQmrpesipzye6wXJesw0ZagLDn9qB1UJ84NR20hfp8GcS+D6stxqJn
9VnnR3+8hlpDfgy6R8QJv7CoxpexedB3gJEyxWue1xcuRQT/v1DksrXRNfCzj+c4
wy7IDncNWz2kb4+BFMfRiPM0EG3sqg1uBs2Jsd11E1eDgHlKJYWmcbEtBqSeRfgM
ULkDuXDczSRdEwpuSqQUXc0xkkKHjv30/C9KVUfUe36UN6AEO2Ro26YA4S+Ofch3
QlWVIxtJQZeFEH0xsgMOJ15LWi5j+Fm55LLIleELFiGG5SUMXQIsHJlsIPcaGX9c
y6gdnP9hVqYBuBlzhKfAq5sB1tfSWJ7JJGBtJ/FRR5gasgv2ahjJi3qEkznego+n
fy/+xkGeBlNkEfP9UQsb5A==
`protect END_PROTECTED
