`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yblGSlPJbgFyy6CeAAAj0/Vj0YvjBISenFSfdIHv4F8/kx2fZNtg9v1ZI8YwXHY4
zKHHSkUcqmwS7tJVQKA2CFFpTtQGHbhmavVS0/CIqEHYOaCpV+2qgLsxgym6Rb5O
6G7yjNEtkshVaUwp8004TYMNyl2aJUC7g6/vdqL29GgzYxoFUcPMrtaQbpoz3Itr
sSgnH35/oPJGCV3Bv3ND2YxAI/YvxyuxoLcHJHO+ll4r+EJm4hZMooyh4Ulp10Gi
j0sjo9OUrZDerFkqB47lJhjv/6qMT4PftXbywhDUna6dajBnxnMQ5aQ1fkidY8Gx
jYgM1o25n/ZVRVyL+uG6rfZ5W2X4/1IMwxGZzLgV6SEfA7J4xVRM2IVIi/OJvMFp
JVf/NBC/eKyTOomxxrMSzngG0JdrtXm5yYELlXc4zaSINin4yTWaG1W65rh0P8ZB
EpX+0JWjom9F7TVEJod5LjMR42zz/EV6iJffw/T7QHJqzDRAxzP2dz1T/8FPif2u
9LV99za5b8clY3q3GoFeqpuHmr5CPa8KSU7ThqjVdxu8t9lMCeF4XOlAnctq1QOF
g8N6TmipRHVmbeHCcRh4Y2SaRQUoNp6Z6A2kRcU56BpWG4v6zmuLpPvkxwfotXcz
SVd/RaxddjDSYiEkJNsoQnjvWz4MntiWqqHJGJuHaN8WY8XaaCncYHNuNrmHRu9B
sIhhWUsPERcK25ct9KnGxQ==
`protect END_PROTECTED
