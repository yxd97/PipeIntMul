`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+GcQF5Us4ih76S4h1+lULWC7QeXqV+Itwx0FeyhxejtPBN/PPRAYX6pPBhn5W8r
BD83wIR2sHWLGlR6SfHfzDtw4xdrBQNUrBNoydvx7WwtV+oWBM/O4EwF92qqyzz3
vE3OussNfX5atHyN0/8DJPZYbXbpkpUMqOR/dlhxSYoCCtP9OG+ntqDT0p1bqp4z
i7QhK9iY4y4cjylFD1BFXOvB3qGd4YhtFD4zaJZHWwkyy4hJZUbAGPWiAP0AVsgp
6avkMv+KG8OI6WnaRKogsGfEAO57gSHsmYBW3168+WIcRYKvac8rwp6xNtWIfZlm
y7SwJWxUXMM7Z6qjPBiTTQ==
`protect END_PROTECTED
