`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6uIPsMiFCV1h7p9gMsIxb9Ii/9Rhue46qnQHuaWihMYfupIczetPJpbyle6/Tm4
3yS322uAffCMWtWk7MSmFnFP8bN4Y9Rx/Pu4vf9QQN2ZBNfptjbIMF7BHW1/LEK5
Q2KLe7WGZhhWRw5sFqYgmKDqj3cPFJZ5zlq2bSirJus19Abi97vCJxrGBD8+9pAo
KBOuseHb7U2wdUzut9PyTU+xPs8OcbPXblJnuZQPLf/T8mcxtS6wW9wcrYkdU1pz
PrvnDMzOP7dV+/rCAOz6OhYwsSBws52O/m8eQlOaOSTyWfJIyMeWs1xyqoti3/Xt
3x55T8/A4zEVzFhbTDstKNeE9Q+gx1VBDCqBYKc1coSQqkhnZ+boQVC0K1amPotH
INMY1CNHz6tH9C7gB1pOannlTKDaSMpIbWuL9Cus6EEOllEXbQkMB1VLNZYXAWS2
yd9mf3IpiHltiW0Y8n1PhUPlF085eMQKXPwxSU3r3fi9RqzCsJSlUEGAjn3i0JvW
`protect END_PROTECTED
