`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zc/jAYBrey0aMG1F2slVPDp2Iv4VHi6YijM5MlDmdi5Lv5hhuUrk4fozDw/xsfW2
OGCJo/NHMV2JFCm9HopoYrirchqH/IMax2aZeUtqvNn4nwfb2ZxocUHDMJPC3mor
ZQciXZOV6kbMfkfK1A4v0EYg9S9q/uTlv5okeM+cvzPkS75LeMGr4Hy5vYIIGe5I
EZLo8UHGYsQdSVHrrV5LwoPnlLGJfWnWaNKGCZC+I7YSWozoabnupg3dLd3P0xzQ
T8LlnsjU/QbNBJ9Vn/LaYw==
`protect END_PROTECTED
