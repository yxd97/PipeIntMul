`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oEPXnpIgWN84eH+02uoxYldvuPZ/iGy0sE2jPZVfEvTl9DqZuLk0JHNj156huiW4
lNddq+tHp2G+LIVb8tnbew7DuywB+KnokEoET39Fryn/7WbvvIUJdc3Q4K6MzFVm
NamUfJO6+ognSwoDy8N1aWCR43fS/hamr8b62QdNwo+0HY4ztF8n9iBjGdaXRKNA
aVpTEV/Mx+eppMWU08+B3qA8vlgIXB33bh5ZF+NlRUBXNY+SJhbmCnsJR6UEM46Q
VmZ31v/98nJT/2sxQV0YT18lTmnz8rhu2s7i2wH8bBhAn04bHiB+pgEviOzlKhn3
BtO+FHGeijj/awCZxEI/sctqck9GJosxAirMRvH4gAJrRvbx64QZ6QBcRszWeY2/
IF4LUd49o/B0n3nqlhmIpX84Sb3AJNHKt6V0V7xYbHf7a0UYjF4KeHH6KxsaIjnI
Ol02B7XxncFxuKw2qnxAUw0UFBK4oUzpzNLUwrfHMSM5PYkO0kwdBocq1wvq8HJm
LjhmGxYrozTrf/9D+Zp3mFGDhjPvRao7zm6WNYucFGU3ygARx9AnFozY4xTQ51nw
ox2hVlG8KREgX8b5AC8j7nyF4KS8QzYHNxTlZqZIRhX2W/OPaIbT+1+a+1ZUfaZh
G2ZdSJE62F9tdtj5TQoHeQH52zdOgzrFtu7LZNaFeTjB9xdmbplE2OoGUqNtt0PT
G1MZME9Ot1DDZ5nSwcp9pVKZ584weoHLjDB3Bd0EokLh2AxhjjAqnYtBio9U/59u
RoltIqaOs4AbrVtl0E3vSjszx+PhzJyyMPcwazxV+7V9iW1Q5BOMuho5J6ZDJ3tq
sSBA+C8HzBuJz15PMABdrqP92CTJALMmqdL14NpEG99K41pTfF3K0NGONKU2d4HR
7X2c2iw4ulU2VtGNcnYhySo7YnN8fuoSjNmITdQk5yXeYohlRiY+VQFd9H9WzzQH
c/SmtCOremAE7XIUsdQ7sxOPOYxrWMisrzwQrm7rbjdzpo0sWV+aJ/cKIScc0x/4
J4FPOzG/Eesfl979IynId2AzC6GRQI3iMNU4ggat+wgDayl6T99tCYivsx6Fy208
vxSO4V+1jUjgWkiXzCf58eV7jwNJJyz8Od8uwkvSooDLGMC8ETKFd5+J11587+cf
Rgq4J9maEO15su1PL61IxA==
`protect END_PROTECTED
