`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5UwqnQL1ruIn67ei/w8HH4AUo70aJCeuNMs6FuUzKX9SCaoNaPB6Kb5LSDejTdAx
SKkdn33SnuTQ1Kwoug1sRBb/6vOB8QugEc4axZXjOxv3pExz2rfZStA7IjOTMSvG
+SdvI8bOjHlUZeoBxBwR9IJozzSMDmogkcQIm7/tjsUa/zRfj4rOeQdzvfOqmcCb
Kev5zspEh62i5m4EhmEzEqkZrQL1wkKakHwEV1Jb8mXPoHFmIzRQ6YYU1sMZMVGD
9TOry+ZJd6xLzXqjqZNanYUIkSIRoY3Aqtzg8cb8UgOPs9YWXld92hQtA7tKozU1
sv/vi5QUTsX/ot1GhcNmaeNelq6Ms0Gj9LYACvzaO1KjKeXct76+/JAcDsGj7BEi
4sVzvEFJ3NpzXunqQbxzGVFaJ/UD1z4RdFunzck6xgv0EhOOAp4y9ygvLKSUApMV
Q6dkCk9LKaI9TidcpGBjPhA46q6wgIsBPEi72g7/S5KLoLU+DP9yxOzhobCgvX6n
VeFCvhy9U7T5BuYOVxJlSZeJcnuXHij1Qat2BrVR1kFb73+x281jtgQPGVjGdyNd
WQuKRUsN8akWYLWfht3hhu4LTu3u47BTJ7ej7xD9W6qjG7Zkrin5fnVb7uAD4vyI
kRFkmz4YfBURhC07QUurYcyYst8AAXa4yNUZJi+n6ef9WHOIcKLh/NoTU/4ZhUOC
BOYVbt125dDtZydPFkm/r+WsMtanEDDOxoBxiwAiHnowNsoHbH5mspcv6c59KNUs
Ou4AMHNHQPyf+DPPSOfVHZy9BtTrdWSCoDRR0wwvA/Ze486n0Me1w8al9MohcY5X
n9GNSYmFATopb5RlrA2KepjzAt7wrP1Gq1wITyo5OxH9SmnWrBnK+VFSxtcHV/qd
Pj6UnEnzWl5sCRxqM+PvkdhXeVlcOA4pWX0z6sLE3zFpQHe5Uxnt8pgvNkJMNhNd
`protect END_PROTECTED
