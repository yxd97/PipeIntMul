`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIZuRM+kZl1r7tygAJ/lMpuno/WtR3gHKQtCRhjo/lBG1XYKXZdbvREB+PURHNXm
NaeEo1Mkfj6tBkUUoGJBcrv9TitT1hyysCs1vz61UNtr/JcLtBi93Y7UTHX6VY/5
I0qJMduJCqRmrRdSfpNccdYFu1cVBrQmdmVhoc+l7BpVwwHT8ZpBhAKg3ShkxKsi
TPaVI3NPvqsT4VO/iQTN3S0JzeA4mUnub8u5b5OxdIZY6op2EkLQ0SRtjfk/qxbv
hRbDwsQo/O0eT/6A7Mi5h5Ck1nAmbnF++CjVYJDm5d2o9Le4Q9ShVc8zW++TMrHp
`protect END_PROTECTED
