`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l9i4V2TbIGhtu7+LraUCgknr7ujHgtZpr/ZX3B7OoHWGeX8ATRHvWuUdHS0BfjPs
X0JYLSUOEdjmjXvO8azKwlscCM8WwZvV8UQwoQNHqPNJsxwcKQIaSorjme4LAcJJ
Nps02Mkgc3ArYYUTsJrBZH+fktc6MOxtF7fhZhscko+M/YZd9ZscOjK1RsCj1aFl
bKICyCooRwCP9JFuYImUs0ktvf6vLZT14h+EFt9xZOAEtqA6aNAJgBJLeDwHxMbW
WzOJvD4ilalkBWw3M9WElynHrfzi5tX1bx3OIoUiXL9PNxfzJGrJDr7HRtEn5YZt
UdCFALMsv7s0vWbeWvwcoT1wCplkE+XCNIuGfN5dN7cqTLo6vDlw9FcV+OmW9snX
axf5ijhrjU82D384+DceVfvdA5O9/F7PgpGM8ixW8fx3Sz0Ej3MUQGtMPZT1ISgx
U1i2B1oM9bprIHBGOtTNQSHSOhrKpGLEhj9rgzyy2wVKVJOza+2VzfD6xvaSNiN/
`protect END_PROTECTED
