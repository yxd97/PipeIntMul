`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUWrlvSQaJX7bhOYKkI9rvbNqULWctDAxOqs7cqR4mO8Dn7rydcw5mc1m9WOVwxK
TLWS0yKOihe0WxYYnLNMMrI0+oMnfyCjGU7loZqHkEDRfBgebVx6Ee1orzIJiXmy
3al2eHz0Fk1MpceVIjjk7w3IT+PXORUoxZKobin/qAGbR6Y/377UETBPUti48f+i
IaeMLYY9saJts5ifG2HdOt8logspzGIANEe6KZH+kGzJHGzlI4Ik4uBxanLypzDF
6bCbhysi0Nj0pguUhtQbW2xcGAS78p0WUvf+0V0DnxSscb1+hxQhUqZYYYnG/tZg
ngiFFe2+G/c+2nJL5/ZRJ2WoPw8yFjbZAvD7FdJzfvs00NWopkbQsVOAm0sQOqZm
nUTXs5jiaf92eo4rDvGOQy0UNU/fB/UPh+H5BS/6T9zg6wJRGGfuuP039Q3ieRzc
rXZNkrTMziBrbsumPLWhq9zUIG+jq9ibb5zjtXEPJNL5DCIRCbmtCPcEwCvWKJTU
j7hlhOOZGWjdrsF9aNgO1pdMtV0n8XHTH71oNw+8ohqLKqd6gg3Ln5nDDJALI3Cu
aXTFO9gJQHPpYgU/6+Exw8LuRj5jgEYKA74niKQEStHuRCSlWGljq/IF1gEyZwJW
dmQafFi1O7XM0u+IMa4/SEynVntU4JZ7VM8YRjD7Oj4IDXQs/S4MeOlld1UZWkla
ElWsKZCpMBzFq6LjhgyhBGct8rAmK951R/Zp8/Mw96qMnc7ZYR826L1ZVKoNILtb
AVfw9hmcIfG0x65j1QZLJyo9hBhpIOCRn5Cz6mVTUfr2sq2INFNCIJotN/00GRCJ
lVAkzZ49526HfqAOq5TF6hqSUwszwioMeXWQvdVEF6IOR50d4RZh7zv97EenYDC6
upojLIyIhdakt5t08F2cW9lzev0Nz7/yImGk7bTEn+Vrd29Cqi/zQJY7b0k8mBpx
qkD/LhlQ5RugOgOlUoAWhX5IdEPrT5EBh+5U0UYtX5w1RsQwpk0htDEA0wQ0ERjs
zu7+cd1BGmqis/LXyBgYsU7+4EnKhOfKv/EQrmNtfnsJQLNmIpRs6pji+LyXh7OP
RZFEiNK0AtWO+5Q2yxrgPbCbeeDnAj5DYLlcY+KnMr6pmIvWFvwlr+bYgCa7S1Gt
C4eIBP8oPPjbUcGeBZ14aNCwl1uoEfHzAkIEC3qr3B9vrUXabZA6P54Tb+dk2Lnb
twoqzI+djbj9Gbq5QWJqFnjABaQlOBcMed3nrpEXcWAwTsHHDA2ArIBSEDmYizgI
jtmBozFLmW3XipfHiItWBp0EMxYbcKY8gv4VqD23S/xUx+nqz82jFXQ7sKUE0A5f
/OGE7SCwp2Go8pNVL3g4fdyD43fgkE+JjfxpSAvBjuQHZiqUVXZeKPH073YT5Icm
CRBZesHw3i+x8Hs2OTmw1afh3udBt2AVOA+Hi7Eln8XBsFvz1FhqkxXVVIr3u/2o
rqb4gjTkNUp2inE8TV+GxB8+JUiEf7MQsVOBsKLkmFrt0nbjfVhdtqWbdLHyO1mo
I6tYJ7xBRGMCE0tKEdfu3LqZonKiktv8b40H+7k/7BOkBaTyMMg5mrNYA1WIdGMF
A3PpG2oeE359BcfdroCb1mT/G3SpYALov2jeATAyNb/vCS4uGPKjhjgJgFUrRUGm
Iuewvk4hmz7MA9AQGQqitP6hFWVIe0ajuex+N48JGdb3mzHi3J15GH6ei/lemq7M
CPu2brXEkzCRRjSehR/giNoywtTrjw3yax87mKSIOmqVDczGPL6JNFkrnynu4JT9
E7AVhjaKRthr0KE3eVHY5JfNY9pcob0nk7AQq4XsgdhUDpYZpOxnkYQXFvBIcS7Z
vpP/eVzswzFtR+tjGs9IprXxWesGu4jHwxzXGcN/nOpnxBnY51NrkS+yyEWy0nXv
euG8Lls81IPuJL8caEYtk6sKw4XC6pNf08Bgd9dOZX+1gUL4++iam7OH+eY4r0AN
RsjL11IwQVuMXZ7rIaTEFf8KRqbdfKy6jnyrE+39XGd4LxSe6EQJGz3viVdbTBMx
E8OrEfyV2bTldOZeg5/1ZFqifTKCRXai/md/Q1IIWbiFP0a1jXicEkOsCJWE1qPR
`protect END_PROTECTED
