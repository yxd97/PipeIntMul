`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+I0sPHrvaish6AS/LsARJXXLRl9VM/HDhSSUgdWb2QwUWtn6/igGyxEL8vxatpfL
XuhHqulIpueUJl8zMCTShNYzBoKuGQTDTL7lR5UDrWU3uu6XSTxrqwTKG3Xews7C
78mSoLeF+xP2uRTpaByoXUGYwbfYqcjVSzNxcpasJVAJRT1d+p7BmLactNxznRNV
G6qvdTFBA9DD+ODRr+MX5boMmUflGhsRxVtkgS44+fr3KPKvcIe3gl7DOVZru8TC
CBtf0pUfW1dSh9MDv7SbOaKzfya4lJQifn1MHfYlbgOMAqRL9DWIt5mQFngVp6qx
PpMBORpb59oIVtbkSoJwoHS49+z70zOf/3X0Xek8Kh0Uoqdz9NckAd/KRmi22DPa
yCilM545wTmkn4VyqGU6DL6p57adDSjVQhHXxLQVDMw0g94UgcTDXK1cvMikzvQF
1+t9RDErGrcBmXgsKgwJbE6PoBAtqDcC0b28dPWIowEQHY3/4cM9VxVEuy+gtjLc
kVAGY4Zi1Js7sIN+Bb4ghDvoafi7+7FdInGfYZVTB66kc5bt3q05AqvsFsmgVRLw
64Oi1QQgXpNWDlQHsP3FaAjuTco1C+YJDa6ptTFxyXYidprpc12YpgorJlFj4pNf
VVqvw4RC1soMZHHzAgKU9hctIyHLCj32qOOBYxuPtsxo/X0kPOIIP3hsTE1p2yhF
E3svOlaoNRO1VZ8L2g5lX3WtA4kYMDe/9VpXJc/iSDItiJ+xsnRk7FEZbHSlwHby
dZMa2eEqrlNcqKPrxV7+gYMOd/YuWZECRThkMGmDnKpuMMxAa5h2+cGlJ6K865Xs
q6JgZhVe1ZmCMprgsVf5fU77sVkjlwSWz/29HdYlc7tg/iikwOo4prwm4tYpA7Eq
aZBpjg1jgYxne9epW/mt7XUcDVSk3mija1XuVQBwj4u29KKJChz+Sp/o3k3IFX6B
+Hi0qZKF1me//w3az2Vfc3/GU3fam4qguHunqWMkmcXUbOYVQwMPT5yZkCfPZ+HE
FYstyQiSSTpV07IDHC5gTN+vaxbpfKY0DK3uBtd/uad0sypRSgnQCagmbEYG7lD2
oDpQNjNlBnVqV6sXN2HIo00ge/IoGhFhLuxeK04tyeO2MNnMSq23bKiDEAUSGpU5
mrTNwkN8v/XFQBJviHd1IV8AMV/kRJkIE12yQyLNXn2/nZu/dgCqmVzPn+at+r83
W0HPNd0OE0FDBTtPuz+qau9dVR7H6AteqZez8oMuP1Tb64hBfumEOJoy7BuPk1CR
`protect END_PROTECTED
