`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7fyNBAe5IKbafx/fdOQ0/Z8nuvunv9hk4IMzRLdZ5sBFe1qsZU0MffD4ZOsUacH
znVu3q1t9HxaUODEb614onkEeQ1omq++oU8Yr1/b4tfyZudaZ40gh3keCD44qmsM
RNFNEdvlK4MpIerPn8G6KG3KOnHYAzU1yl+o6yRzDxAdx8mTcyfk8YG0NzUNZdXn
GleKV8j33ifIN2lVkQiMvCdMSSyIZLrFH48S197wgV18eNenHiwkR1GzUnwghhfK
AcWtdw4wCYs+2fKmia+9bnKcq+Pb/IZi9aGGZx8quW/6oQnMvniiPXP0+2aHaQb7
BlaI54FdLOrxb0Gy1qTtUVmQGcyGq3xsYBe+ZsziAloY05TL87xkKxqSZMHxasRw
E3mJbmsNjy+a0Fi8lwCRYXCYE4IE4EBMavgN8e+yJY8=
`protect END_PROTECTED
