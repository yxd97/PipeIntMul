`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ytVRMwb+gv1ZzOVvqYb8M+n+kzn1B6DU3fp1fpyb0VMhzHhJBG2V9oXYWfLPvVJD
PC6x+xZ99lp3yHixnUcTkDmSMckA3aiXTI6B86K6/Ll2MFxx364YEdwN+jC2ysta
OAFmBDflETfj38TRrJCsuccpro7ebhgI/KHhj1pTKkAj6I6QSSHe37hszAtbWfk1
1n5nB3Gd+Humal68T8J7xQtZDVYeVrZkXEzSqsQAqLasVIX5wXy+jyG4txDc5OFw
OZfP3pwKFyB2L2cuQjdGdZ/KoMsPvhtdD4YLOlxihXRcUjFF8B2yH5whY6KQJiqg
LfWlu2+A2lwl2bykHQiimQyxu2HEwzC8pSEs6KchvT910J2ILHzrWXwr2enXmkJl
9aB6sEsxplFxBmtFDM2P03uPAcHOfHecx1PpdhYPcDnyCtaSUV3ovZ7cGFZoIcc+
iRZPkQBfAqTn+u8EAjFXNXYqHL3vSE5iw8cbrLSQMT8tYRKagbJO+v/M8xM8Ki0M
2p/pODnMqMH+dJj7Vw//cNSuLm9ExCxNTj3I2/RQmiFvsLb1Mkef72VpKAYwV7Ka
Y4jdK/J0rK8DSMFrHcLrsquhR6dimASA354YPX2ULgo6onk9HHOPQJ2NfVQsM4b1
2KKYuIxmT/RUXSAzzcr2TA==
`protect END_PROTECTED
