`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RG2BeHciiIIuSkmIv/V+NcSVH7DNrENTsI0XqFMParg3Ux4zixBUAu5L0yOJyONA
qZEGCquZlfysNtD0xSXWUeuhTF2WdDPTT8wRNCW/6KJWACU8gniK0J8gTMbPmbXk
r80VNsItfkiyNdCSDLjhco3L9i6Y88fhi99pZBirKKBTBCl84pQ0fhxXdWTJ/bHh
XPNWZOd2BguaCu2P1bPWIADbmUfVSjcz2UB5Cz9VboWlBzDua6E5mjOqTQYVI9r/
JeizmomdEuYavHdujAXp9jkSoOuf/GXSwozRMMmLBnVxxaC2332FI7RmpaBT/prF
tqchXusMt5mWDFX4rUdOugfqyi7eF1cG7QnUj9l41w8MLsp757qlnNmO0wLd6c97
MZJ86r9ll8+jLXGjnIIiO5tJ6SQoXw+blpmOx66m9FdzFqjUmb+a2gw37WwT3DZb
q3+HVJ3rL3jiOyFWrdpxs0iFEOUxDXd/ZeUXdgoAN0pwYQhzrXTTYFzKhYmJxP5i
fCjw1xTEFk4K9MdDfRa4vacniiZojYjlq0zpqlgATeVJOx2WNYe9K7ya/cxfJWIP
IeW1720ll4ynB6Oa4po9cuQTEnyEClPdWdjJ/1e73K2j0djkGA2QaIy/VEQW1MnE
SYFLSStiZfCFcrkzkDw/6oyet0PetBA5EqVpN9xGOAGh4Q0R39s7ljYx4n6bXuYO
NmJ9VN2t5PJwt2biZ+rZ2hNqJ84H53yGCaAAVtVOvi5M5xPNgk5uFJTT9ufaQU+C
zb8Vd+IC/vF8/lkt+AVYsG6JbAnxX21eFyst6bzSxnSZZrqDsw8ECrF9qsuQ//yj
MGBJAIyt4r22l4TIq97ibJtI1w5CebjOMcP55zxCe0Tx4/mVsyC1uXeOxtHNnvAX
e0N+wMODWEg7gHfrJTc5q8odoni4FrkMxCZnqUOvboDN/eeWG4qTYPh1PPtRJGf/
/FHsImxgxWmFBp6FaqyYIQ8kYh1007g6RzMHx3N4SRwt/ai8fD3OylBxY6qUp/Nj
+AL5l+w07rT093TNaBnQvGn1Y4CrogKf4ohrigZmAaRPWylcTyLAZndTBQ9PEyug
YdUB7l+ASPhtVCpYZzwb0u8N2Iv5HSqP6QqHFqnpgcz3WKgD+GSeAvgdNJABLAGl
gWbIdq0uvUClh9yugJ0/cXq8xiL/IqQ4yDLBYIJfgC6ZuP8kissU+Gostabjjr6T
SR5azZeNi3S39cpICIGRRd0Sp06MehUTNgWI9TI/sS6G/nBkbYJlvDkcm7vIfv3P
BVjm+xrYb8soaaPfz45xCZZetdqBT23emBANWkFrnTVLOKzQ3TrNoiTY7Vp9rYrx
FFMfE5hOs4cn2KzbolGNtcB2nvK3S5x70mxVhvY2m0aHhvAl/bEFzOFwfWlHVP2O
yzAeEnIfeTXcGGZ8lWk8r+7jCq1fKzB5G+JRAW7yfqVvWH27PF+C1enNhIqV8hnS
LWGVhR66tGS5P8zlAmETM/TjdKfONPDJiRHLAMhDtImnoW0ZNfSqf9Y3lkcVPgKu
IpIqd7zFgd42Gvx7priDNfcrXrywWoTpF5SZS+xebvAuRxDHfkp1J741zn4iTR47
TeY5fiXQ6+H44smUGwkYWpNwSuFBcuUOC8EgHPNukl4iDbbhFMW2V1rU41pcEuZG
8F+BlJab9DrPHafWl6T1lJ1X43ZZwEy5UTlw30iM8r9VX16dWGMzPwphUadh9Rpo
tHaJflkc+FRckFpVN6F4rXeDeeMkLLrrC8n3O4/z0Pu3CL8bksX7ziJIB3ZOWFGG
9qbjOBKO/138BX0gRbu0+mkG/g0O/aiQmRB6rmhpuCNVBouaLC+3JydmMHpI6mBD
+SRfFZsIWYAvMYQyH2yGwdnxPyHg/L2GgqlUncfCkM1W2DLou/numF5ptAP+55hd
c28CgL47nZDql9qQQF+PJnz68+gaphTMAonAGo8frkJAG0n3dvjoM7pEd4Oz4m6J
IqpEEvMokw5t8ylYxyKK2q9wqvnrDGpvwj83vKmiW4p3W9cUEgzh+KkneOzrC1U1
eein78kSA8XWdCDR0QFu5HDfY+s6c09xDslsnkIVhxqzs5fp+mqlRtoUW8bHxcmO
HLVpSQzjCc+o4TpBuaiKFAxo2FcGhn3G49Y4LLHEIdr/3UJlcC6jgM27MgXUzDyO
4ZV4Rotdv367c6t+Xa9Mqb1YiFXkojdsPhNLWqpGi4nhTV0pCfy/p8QOzpqLvqiW
t3lcoq4bUq/DsqWVkyVE4v2DZ48CLZh0iAQvDGUL4a9PNxNVJooEmUBEHlbGB7+s
P6ixjJqoSie7hcA4CEjRl28Vy7amZxrf5WDBTvPjGzWHgcbKsOXwWwIiwKAkCOPj
yulGBFpnJJdQxHoMZroswHSZ3VObumQZ9fmhZgbD+wji13HvIP46VAsqLH39ywCu
ZPgSPz1DjEc6A3CLOxGrOHrwa5ZMi3+HFsHjrm+TUuZoKHSVXczKEV6yEesDdpPZ
z6SpKhct1hOhb2Db+np3oKYQJkUFLjPyLSTADH1H+lo2jUcKxr2+H0/+HUDWHF7J
eooyoxH6njAxkF3s8Rs5/HM6XTkPKGjmUoPvH4lpA0IqhG21iMRmTqZSOKbtk4KN
8fkUJydYMONvtudFUrjRRHh6wrLs8Atl0kkdYCSXdrnkSMQ1Q4c9BSp8KUqCIzhi
98vUCYnC7lnxST7k95oLTGiKrk+5lbXsKS1yx/J+TQzeU2D7x7RD8b22ox8PlN8x
fge9m+5qlrr1kTSpw1SNOdBAdmiulUGziLTUuv7uOOR6JAXFFJnIZ6nv6v9ZdmPZ
`protect END_PROTECTED
