`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5uYZN2nce19KbZNBsZ7q8NBBaP3lQulyELXNjDP3vb1ZNiSX7Z9UbcXhc163b3p
aCvde14MrlKAZ0bytFKwljPr8AUDYIDFJ9kbigsiqfpHyB+0X3zAH8iJ0bf4tMiD
aaj6iQF8UXvFqtZkoAGhLTneflodNycjwpxqnaf4v4RZZqvUMY8awqX+0OEIZB0q
GbO2//PLpmu9SojQ4JU22/ppJz91awBU7kqP9iwwu+NLX6/lm1i9Ih7RSfAzCSZp
Bh9g2sxazsZQUKdLDQMC+EIEC+mE/4wU+tSHTcrxDNw8sxehkhxnVwvQmckLMzpZ
2t5sLTMPgzDFijIBUNqGf4CPJYBHzGarL03Kw/CIqyfqp6+QDYkvUqlhF7jUmJKV
ziZLA/AcRZrwfWjusPVlcEk35lQdV/2xjhGf6RKEhdV5EUq++NLr9m96YUJfJGT/
OhZpY/gpCLj9HXuj1SLLg42g1yGQbjGkU41Qcs04VH/hI/U7BegIxrURGk/HjYMH
FhXRbvfjDnca6tgl55lOLK7b6CsP838tLL+usU+kY8cpPwz+x3252epF+Uhpbj/c
NyPRfGBZDKjhvMwr6NZEWeQaHxZ9SyKRy6H1Gs+FdHzUraMl5JQPdWxcWGaCFtZd
LFtkT0KRzaqOGAvRXwRz5QMWTLF407RNHfpKOCDu09nKpetx0gi0eXzWIFOW7FjJ
BWG+6/MOvr3zIVsgzYsrJoyYmLxEzHlgjuMJiEAQiylCyDFGI3J0C1A8JN3z1KgA
Q7Xd4dqDI4Ian8JGJBxSujw4aYDnhMsqdTTKhmlZTjd78ZvU5J4frpATjfREXWp+
94g0AZIuKi9BAldHVsbN4SSJD0r+GFDCO+GQKGN5rEBo0o45AxrqRGfyXpV7skQw
MdPeaUu8mX+OD05rxNzdxuOiN8lJNn0vkeNrIBl3xqcof0PmgIqMQbZ4yhSpDMLy
yzi89UPJyDM2KHJ6c+me1BSa4fBueEJS8IteAv7Mt7sDY+bwISmPjKk5NOY9Shx6
jkjPAgmWXoYYm9Xj4ArBPQ0lfQCYx8jjqWdaVmqYA5JWYdfG0GMMCcpAoGzjDQf/
igdlOK8UOysajOVoFVe/6V2Z3C/7dUo4MKu5BKwRfefxYaUw9nwM+SQ2OZPLy+XK
/InbZLEu+5EshTcsFtv00A==
`protect END_PROTECTED
