`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iY8beDSZeOwv4aDzbc9AKEym+Ha5rhpgYNpFI5LfYC3agZzQbqis8ceNL7VXtqDb
CaVKb1qSNFL2joAxqpdy1+2qZ55L4pbPKgIZrozSlLcjMUlGoqy4Q1mLMHFpnSQS
lkv0vq67jzYUZKhUS9hiMOjh0Zc0DMAuyRw57XCjqgGSw7HRW0gp+U0wBfyJ+OeB
vnimIQsV+494aznDuR6uD1cS/FKZn2MnJfBXCfeUYZojCYZwpULt9o1jSNzlBS3G
jG5dATRoL/QpJ9CQyFfnvVGcj3eswb1G89LUFN2MMmQ=
`protect END_PROTECTED
