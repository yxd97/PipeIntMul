`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qE64744To+00ygpO1FwiHVHfV8XEtgf4FVx06NK82PJTgseMtB3p3zi62L/kZeb
oaaRgRikduFPi2nqYSIQeeUo9yiczzs701e3nrX1I9JM+ReRZYe/B2Hl+I4kaQpY
Ks2pBdWUn7oltaySfLiMts87jZJHfZSfE2rR//KOYPtbH0ZUthDU/sLmOnrQUNrl
SOkev90DKgsi+68+YSpS3sEpU65+peJ/Ij5FKhgYV5E98SFPxiZGaCNm5LcVfMoN
DAFaZbFgPnUBf0A1ZEDHDelV7Ng8iqwmPhl9dVrjCR9oRPLZH9idarypXFWx3Iv7
MiYKdh6wNmGNrIvk3MJEKpom8/WNguRht+CQhGjCN1B0IIWQ7OqO9c8crZV9wwqF
ZvB0VeKk3kfaugkhqwriBxqweK3KUxlzweGyQamyHoLHU9zn9x6w9TRKHv8y7asg
0qMCeLlDnCLJqZJ0mPnq62jij/MDV9EcmBAjXixjAiSsnHzUPWZnZY5+ieBK65g0
fOUkBd4lqL6Mmf2MC7T9LTZDMGXaCDT6JJ32rYMtP3OpIl3lXya3jKRGYLZJctzx
JKaQ815mHQy8cAfI9aBRdo8eu4kb0lCSjoNiNhCYvjyD02LERzmKvOu45XuuNspc
vJhh/DtERBOgLsepKK0P/v9tXtGg3U6KLTp1Hs0WvwwmEXyJ8l0KupgQbRYDc/4s
IMmrftjsw2DakgE7t8IyppF84wh4PDnF2nD6xMXcP/Hj6wSrPTzHypD30pM5If+h
TTh0bylNCxQK/RtkYs7ZmUEEULY6mbXA1SsYqESuTQGy/o78GI5rSg1IpAxtqaPh
nBJRLYiIYqecOjaW6OBKB/qD3Gn1Sq533V+BZY50BQjuO7H2RRKJAFvvm+iTnKd5
zeBBooDf203LdClY5CaQD6jg2hoU1dnvgqRmfRqynRqL12jTMk1dCf6hd2/FR9Qd
3O3da+KhUpj/EN7ojKBY2ZUitv8PocZbuLaOGx9iGPmzgQrMij7qx4pwG032voxA
Tn7p66paj9ssn3tIQSH1pFE1gx4US1GA33ir2ZLcKBXrgre6bpjO4cigh3VnCWT0
8+KrdXOrJk5q+8oX/6x2jgQMAKbTsq8CZ3ieYxxXg3KFiDIech6mBNrBuv+EalgS
hCAGSjHI5yttWM3sElPCGe7ho1dnd1lG19hRVkN/AyrKFEk+hBPUAvDeNF2UTS9O
cEGcXZE1ltX6YLjN4s5FfeKTbayDp0TgEXwyb8db+/fKyZO4v16Iw/Go3eXPM1Xp
7jHKjR7arGPNhl0PQ9OiZKj5/OZUxyNJ0CUJLGizEUS2phnqtEc2NcZoTFjmHjkx
8hefF2xS68XC7JnE276YBbJ+Ia4R74RfeQ8yH5DaSLh6ZBiF0g95hn6bPT9BNIUJ
qW9+GisFsa9S34uz/tENDtXJlDiRTmwIV1E4KphENGFrnA7mdZh5XxQA2X8F8GGE
fIBqdEc19eRJqHv+5aYYJbp/xA0IBTn6uU3q3pqnjIL0xNqLEyvbxHLtgabjrgPM
l4zBXG2ICy3UAM/WcJLVN9Eo4Y4gP0QhXaFBWhJ5eO7hl4RJGeicaIPH1IEUyugM
QPkkd76KTBcLM5Td9bShXRA8FRfb64uR7nrACp2QTfQQhmAmqyptws8CCcGIY+fp
o+S8DtmlNEZatU1RkeQb6IzbGbJNQEeokGtbCnJ6xZKKmFXZC0uJQVgjOeClZ4bW
Icu19xPF2JcDa0MD8gvntw2+IYakFbd94A2iLOvkaiPTtYm4vz6HqEJ457vfvzyt
WPUZi07RBAcRkTmC/87fNj8PdkGzq0oFmLg2TXSMOhbddU4n3nBp91LVmChuse59
TMa8vZ0kPFodcWtBfTGwkaNOAxGntHNzQ268pYja0C1JmmFsIGnPxAU/4DQZ0N7/
qUYqmcMYUarJE7tKUqCtQYBLZZMBszrdsQInXHObBUXZPask0eEE2JmrIPQTdBpH
aj6coIPeC0QCxNhOtWfq16JJKHVWwD3Gdjp18azkTlM+F4dtPTPKjwGkol9wfMqD
u7/XJdGnBXGXa6t6l9MuH7tdyDtZJf1GXhNZKbc9FpCyrt2DoQsw1OZVCvxpLK1V
ZtuwZ0x7i9nlsV/Uuq8CXflV2hHIwoiCgK+EHuQP11nf2A9+lZnqXwqoLdpIgxq1
IvuGEKxi+B2EwfcNqY2Qp5ZtcQHnemqgzpZKEwAqhmlh+vV1YZ17fIhAJUodX2/x
4ALB09g7sWV27rUmMLdgwLWmbR2Hb5kqou55gHVOAaMRCdIlL1Cr0IsKuO6mc1jL
xxaFmsqqJ3LMWWCW6CdIxr7/Oy8cREE5eSyJFFezbW0gkxdWX7Hmd/S5VdpyViYA
ZrPiL7fpie9b/H/cMl6smKSMdAP3gQ1XMmjlLlzP77vgkYq+kcHsLg328FV0hf4F
ZAosxx33+8GONNsaMmEogRMYQutBdKsjBRRj6ZdvKyDmeIJRwJBpNOtMfJqgWBHc
ov/1+Ojf/SUSN9kTD8FEdouDiYqw4jl7HUnCax99LpRBU8ZZacYQPdvUyPSJN0G+
t19Zpgs2kGQiWYNIKlFBWKvtpiT+daT6cPpHcc4kIN8WkROo3LpjwcbU0ipNoPP0
gsg0mosw1mjxth7Ipfpt+BCuMQo0v3RTYr8FGwbiZp5qLuGYnBdy1sKjZsz13kCK
BdL9FVlaUB5KJ0uFyoOHZF07cOHEW8qGdqkH8EeRNISQ3GpLPBdjm6I7luORF0U7
jur/ejmUbkeCxtE125+moo6DHE+RqAOJMic5ku5fkd9tHWHH3utoMTEZ5nCasxSt
biAqCqym+QWzRD0RiWaelIjNgGQffyxHDGahWMBA7SjE5uEYkpHyRgDf3qZ+h9yf
e2cxrljuCJoH1L3fUId8qelwHKT6DjjAYAay1mc/LCi1M2CaArhw8GWAwkyZFuWa
cdKZfXCitQ6nERhhaHW7FdJJZvX06mSTrCEqqj6zL+BezSx74mlbHM0JTsvIHBzR
jbBH4MWdARIJ1DD/ty+3ffGejwPeZ/G8BrNqX/A+EztBPOTMZcnNqGx1PPWieU0V
ebkmzgsU6XHXQ3s3rbWa8dgsIIUDr0zRKocPCQ57YymUfWuPVxxBqZAmpu1Yz1eX
iMYvPUdzB/1GrrPrMcRz3fYFCPv8bieiCDS/UavAR5qLnfAgl41scG0akIez5t0z
BtodIIPF1GGosbUb1CT6hDCpv7LVlIb/wXPosq1vLdtWa1ruwcx4sBNH19iDvfuc
n/15LmLhTgNjVklFAzZPkhZ9ItjybRNLhkoLPtOmdHGRh5yDjM9KglA25Bp/R6CU
Y2335HFn31Nj4Wh6i3EY2ah9KfAzHMDG/vX7OqgBAbq6c4vDocHKrW3fWinjQ+Pq
XYp/XFNfMI+JO0UyaZwPg2XH56ijwv1oDfxJXlWve99zy7USMRJNZv7ecYdK83Id
Hs+ee6WHIockZtv/qUMaiuOuEt7Zf6mkrG0jiyjibVh7VVNjxVex8dqK3B/xc9mu
G9b/mPkf+NYnrlxIghvRwjnt3z5sZZkX2lssBH4lZu1P0uX2TTUHfHEXiT10nQPw
gEQZfKYkXJtq2GXtmUlmc5g7t1fuV+hnUH4yU4ESUbg0XgRsx6bAX8UlUAIkwUgI
izjZSNmsk51gV7ohIDG1E+Us7ZNZB4ofWxwzu+IkZYJXcHPGU1ZTGYUd4ABJDaEp
/9XuRJeZxadatz6J8sk1ec6JL0H8elLnimUz5bcuyq3RVkH3c3kKQhCBeXpSXVDU
vt87ETm2htekpXjJRi0vByfIagEz2klwLlIIbwPpFs94mfsOsJ5b4pfN003ZuugJ
Yg4kH7C8SpbJdZNPqTeW74hOqQTcihPqgz3gGYwsMB07XtnibhDLZNkoFsfBXJLe
hJZuE8HpnRP4lEABMT3d/xdpPxzExakeJSPilDofhqnFfiMGbEA4s28k/dglTjBi
lmWWysEPj7XnY+/SDwBlCED6YhGuOM68X+zoGCFkhNrVHyfGjHNVW+fgn1wAKMJQ
kThaUfiXsujmcYuEeQQMtvxHCjTTC/uScqEkcSMyuXHnSbBP82lb8jdHOGuTm6CY
ZVlsusxwZ8cXs4jCRSufl/6mPk9LDPGdBaLgmnFKEvFhAw0wHVHIMryapjj8Zcu4
NXL2u+otGZYuprlywWV1IzEfmg7Qt3KAgKyWnHzGLAx9fGRSvSzB4UoX6FfMnn51
2iCbIWpt8MKEBDV91Nl3cfbmnsTgrhK69UeDjGecxUbHkZUnvY/reEKna5rwA0Kf
qGE2DdUYl0sy+qA9Dasi2lJzEjWUGjqByDIicU4lD9V3lmRt5iB5+PxUSLZFbiUJ
WgT50XZveubgMxjQ9jrUeVorB+BeET56ShAsKdTr7JQ36n/Y48zffhxvucZ2ccgD
3iEKFYeteXGXq1vyzPBfY+Wqk081RRw+z5Agg1d/1drtWRwIopgQneNnqRnfXLMm
4KUdE67yMe4ZmVdl26HmZzZdi+CKFW3I1w5FSOYsscpchgrl0Qn8Y0rFoqzinzNY
k71Qr3lkLwr00/iGumN4v0joLZ74vinl9qJxG8sS7fFTN7L38zTj244BboCR2z6X
W4mhnjlqdPSzhAJsv9gz83WHm06o+OMbwSdMtb8McNpCTRlSsNd4/A0R8aauNYXt
XAQxMV2GTpZ8A3cejir3xjeXrHGPU4taKdcxthq7WuKFR+zV77XDHY4Bpr+ZlnNO
jCVfXqraSzskswx2Lt0HxISR+w1ed87aI36SBW5P3VNj8cRbJhlzh+0CO/wenFpE
wx0SESEVKTuofvRE3dPgGDtYxOnnWMOMsMyyXnqaRiwBObbcNMK+5VLvlsDqq0Fm
XgFf5zbc/LBKro50o9KlBOsXb0igzHlf4Gn8ytcBuLbt+aCNhNixCKkgvC/gj/Ex
nW2p4LNxj/Q9qiyI0FI9nLrTZ5V/8t166/86ms8XY25TwCSBezspvo7xZRSZUrx2
jiv/+FTuhogNRqbPbjh0X9y+eWSb7M/s6TeRI1FG6ek+CfR+qvHd94argy1vuiFq
zt3Qy/SJ/abF5g5vrCG37eAtRmGWLuWwaDRJq6LY4Pq1fSAoi9bvODPwZtS3lazD
3612vEcD3GjfUCOo6G1PHAzJx2R4omeYdPIxHK8K0V+VfxPTnKEJKaZWdF/pykdu
SJuVa1SwvTdOkB2iNZbUc1WuujkaBI1+559wxOj0ryUt1GpYxDQFeKBCn76ImybN
amQbZ2qotUnjk/aOSzw7SpOlN+VHTTfkWchh1n6o2i5HjSKfpdv2Sh9rGpxNsuMj
792pBrQWvPtThcTAXObC1/v24n8SwBI4WopOg7sdAZaVu8iuornMPo7DO6OHeKGc
xNMsG9k8XmQHJ00GPk131PiOuknTKcOWNgEkcmrGfqzzTIyv4Wr3C9y0+h7Aad0n
7i7PUUbYyFqPIBfLLfDxhXiHH5V6cGe7S1LuJkPza/4JVDGOpLDV/uhQa5ZYuU3k
5uaI6hBWJB0LJ5yn8VzC/EmxmIPZnVIM9homU3HetQea6334R6HMiVyCoYrVHNp8
OaW3tXe/5Nzyt61KHMVB5BW5JxKymvskgPnKL2ZRtkpj2J3No4PLy/ojfPqj7/oh
ForNNGZDbtQGA98v2Ozs+IcxU9nqXPxR5H2+TmkpXn1ei+YH8IJO+j4l9yMgwpfh
Y1amDoxpeOgupIC+MN1DlLLwhjCirs+dqfgQWaBi121GWvJYVCzxZbA/pm6Dh7wp
0zSQb5x/gycymFDaZZQwPTNz04aO+BFUKD/G4quc2CiFOC9wwCVYZ7jB9vaHz05p
5BEJCrX5yJ50u9zlXY1V/GXlTXhohoNfZdNeiBkVlPBvT5fwOU+kmHigKPRNKX2O
yaLsGHD6bdR1A4t4U2LrHti586VA3TSeE7P2LEqmdCGA1ePX5EXWv4M+6EOJ12UU
CcaG0MpSQ6VUDJBOCAKtl5HVTPEZGvOD4N5/MbjVvnqmYsWMIGQPmjnl53ocA2pb
ZmFFXsf+8SnHVFiGONdeYfHkr7hjKbbAmOX1P58ScuVnA8B9xmPUGCgZwjFPYAHl
CQq9OQ4jgdzfxplT8UK4ZJ5PvP03ecOs/ABqNt10H/Tj9FPWndosFVPozZAckdiA
YRVCzk/YtPWvFYVYPxubrJKwcg+zGT0dQGOXeN4vxUFdU1pYUlkrnfP4LJQSmiJH
0ojP4PnkKjpP0rCZMw5yZMFLV31kEL6iF1P2vyiwQDuOg1sUxUZgmjPdTlc/SUmE
L4s2MzTB2CtF+PHjvCrqlnPNVaK3Gocj4lhlXNDZeqIELW3GlDjR6ToMJ0WyZIfC
2cIWEWNZwmCtyrhWNu4K12s93FaMmhkGMmOC0FCc+829FDTjKSBfCJVheZa4LBva
ymPLlYZm6b9xPbuRa42pTzj2ZjTwmkN1KadLVUUfeqNZZ/w7KEjI5/pWGZN7FR0c
civu17wl+SVYpoiA3b29rf0AlxAIJmE/CBucQIgZSc//7AtYOa6EdT8CI59W+S3r
1pI/WnW+FHJ+AiWCyK8r0RRhURbEsdqIfJub1Ywn58/YGL7blSzE2XeBG6ZTdtEI
xOutM0DbOvbIy6qssZaZ+AZurtvZD1zp9WYvLJJheDffYeDZIlrvr8zF6bTrEfsA
yAhSjMBeryT8nwytkc1XvRn/Cb/qKNL6LFl+hEqAH8cm50pbEP5zQdvDpArdwU9J
AStpwZVnKy/iTX07k78TtLvlRC5IKawCRL91YRvR85/KsqaPieQZTlr7cll33a6K
tciI6C4QcdD6nlluXknDyKzoWQX7EbjHPx27vNmJxbow9l3GK1O2z1PP0RyCHRRW
mkiK39x6PPcxcVPG8IMste4rnK56Xn4xwyD7R0nZl6HGb5JDrBo32d+ZKvFM3waH
HkoFEy3nWQEtD1PbydZEHvZM3WmHpKoDlJPLUIC1kyDTNlnwXjTpvTmB1TVR2U73
wCFdeI4eZiIqxEzy8+c1e9TLQRbThAIrzV6T0QoCm2kK1kqhB6aEZN44TSMuPe5/
R8IHS/u49opB7FMoKTCMXQdjo1o4kRM86lO5aBVtXrtlWY6La/vqoB+PAI7iKGP7
Xrxff3D5lcrYPCC8DkSW8VDE5KG18WhP+rhWHcZIPAj1kwinC+Nm9r4VA7tVi5F1
oagpjX0RP7EQV4LcSpETWDXHSrxbrVYRLWSZgDOiu+zY4LMbOhm+YWNAYWVxwvhi
8x6oKuI5ERukVc0ZxvfvIaxIkD4IHpr6odt4rZfbqw0MN5S2KX9WNcpIHWIDmTR7
mO02MhUqJ+lbZ06ksacyMYgL53BZ4sWltcuB1La7O2LjqNac8Fsh+hxuSxzr2SdF
fcpJuLTZOAUqJiUVJPHs4oBqx6Mplk5CrOVXwnubHU44KGvvThM8S8zFist8qCPn
J0wNRAmCAvpyFd51+9Bx3gSUGetoEdemjNgKa8whoATTxy2AKYAU//tH0EYDUnex
SciMI0HUsKz+T1UYn3WZzDKw+nKhcffjhjDMH/F2Jxe0tlSzZmf9Hw1BbDBcs1AJ
s0tHW2ulBuMF6j4BM5JrKQwNmJslAL/Rvn2HzAof8QBZ5vbGfWzpwouF1Ti2hMIl
7dCbIvt58pNO/bKAPPITQbJueI4aQFV4oJz0BT0ossQ0s5IR+HDD39Cfmga79B4z
gK6Y0XInMCXuXEr4PiX6FfGoeCxE15EK08ueCz6DgjeTOhjeMo6vtUiTTrJLFsMZ
BlNvh+ihxskG48jJXPf0GeAuhFvh71DdJoUN3ZMkplXeuBnFl0OMq8tjV6P4XCcb
6UeEdhwY1YZRW6MdUY3NHirjnlr1xxIJc0GMNC6/NZhZ0BxMt8a8xc9Kxf5vJszN
Ceclyn+LuHGVjKms/EWMWDxaxxm/4whP9tDjOrZYSw/RGfCSuoue603IprOSO9iC
ReKj6SjnIdds93Wby3pKNeYKGUkGiFnpOKx/jipG5fY9Lo3Vj8DsXGu3+USr4s4y
jcNOEHLqEnuyeoBYFaYg3V2qCp9ED6Hqi8u9x1Ny3GaOgp7E3w7W3dvc2yA7u0sx
o9VhjvsKr5+oJjdN02cpGM4yfMlnEVCrxQbPa+Q4mnsCaK6AEstN9zzRsnlRMiu4
0i96tEmhVpDdr1TRofKF0EUOig1S72xLfwz5DpSSqreUTQsZaP4RbLuxRjwCOmZO
7CqRgRJt5cuNj7mf6QwmzhFx9+uQ10nU18wKIKh/QIPAMdIVtU4O+TQ2+8hbwPKd
xpyWVmfstbb/dRAoUuduLA7Euc6/iGErU6QXQCzPTd38gqhhDjlE827eCP344HCP
Jp7uIvB7nNiBFVhyScp33KikoOzsoCYmaxpl+i9APfPJro5CMlDXbuJ98YYuwfNT
kLgDuO1ufY+51uQYxfJtiRSWTDx0LUx/5IbKXfErc3uWl9+1n2jS4xEWJLNwP5w0
YOp02j6FCDn6BtKjfSuomKL9AjaAldXdtJYnQ7wrlGcTtjTypmuax3SKFXCUrN3a
UPJg+wtr6xNyiZxKL6KA2XGIGwTjxUpL/xtZLJKWoxuW00N3evtaibvvu5pFPXKA
PbU0cX3oBHPxJWfNZ8Hli8vMVXfm5yS6MucsAUOe7ujgKQa4CbcXkphiNXUFoRtn
Pc7gQ0NkYp/6bvAfoL843eLX204rnqYtcLj9s+xsKxUrD0EqFACsNHXkt/dKkETg
V7uyYqT9hfsvG1/6eKt3GcHzB4MwN6StMQ92WeM8TvNpiHsvrmwbzj4DgzMymTyw
IZ0HihhOWIww9CknvEnlxeZ2yqF16aWub5mNpha7UVldfoy9hur0GYPaI+Who1ls
VhRqF+P2JDObGVJjCDWttDUpVVtyN74vJoWhpXjaWFGFqUcx/EiWYrBLWKXGsetK
7DPTAAVxoegMs6kkFE/G1kXE8dadY+BZHMc+avMicpl6yaQAo2vzFkwWyssb9jon
v174tqIftGGiFFYFsxezoGcFkvylvNDEDtgQ4wOGWc9UhHXt5Nz+5vPLksWqnT9m
rB63zKrZtkK31jYXQUHKT1N1TWAzdNbeTx7O2YFgDcEeQQfCXtqQhDy0u1fpynox
Y68oc6SuDxeMzzX5Os1BFCU4Wh4lhin6wbWI7kRRD8JHw6a7tOaGjAlvluDUJlEn
bxu+F3Uw4rrRaTSkVi+P9P79zF6fYuBCqD7z+MiP1Z5TcjPpXdhqLhOekGCbvwQI
6Sz54WjynYh8zV8UAhWdhtl1mhE5Pe8Kw9qt5RfsYT5bedQhew4uIh0uPWBon5dh
xBcD/uZmNC3/vcEER11b+q0ARHQ3znN7wHqxlVe1n5TPw4rdOTEv2owB4KpUTw0e
RBliK2zlrb4HggpAmHz9LHVauBkx+8LXk6YluFP+NDAbI3TANp8mNKY780SEai0L
SlawYJ+2g7nhuniACv8dups8t0BSylRamQ0d77y0UXH+jQCnhNvCkQ3PzX/p64Uk
rzmpQGZdbEBx0ArLcpKSYetfK9RRHJSTntWaLF9S0SKVWTFThXN/oY3n+frVFs4S
pNxve5EzzLg3vY2RQa4sOg==
`protect END_PROTECTED
