`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p/tT7cTy3WHIQcut1+xH3ctTq/grdG2wEQnavcmRgilb/PIaCWnM8etTIBZr7u2E
gB2SaxH0i0dfAoZvZ5DuQJmY3DxJjCk3+EGRxAsH1/NsBfLhqY23GM7W3lcxEwa8
mvmYh0Og/mVNCB2k0zgRutUZga5mBHRGV+67vxq/ExmHIPOlSzNQdugbod90Xgp0
Np7sl+ZYf49RXEAttBxItjKibPCxjRB/+FJDKoPutwJXGddT5Ey90YL4ZlNEKvj/
wNJpYiofROXNWh5l1dk67Xf8fEty5mbOl+YnGBl38Q1qHj8kE0dK//AsNKqzIsBk
LcDNHB2629NB2bYQAZWd5/NnIhS7G6xdcucxdZcJ5LZZKLzzcFFGTUCakXHTJWFt
mxGvab8tC1/uUmHtpo6RhGoEJNTiqySFQX3V7i3k1PL0ZTsRfT9InD0DB4u719SW
Al852t92jKgtQOu0I2yOZoU7x+ka5Lgccz77wMcIwehlC+0N4Y1VmwM5v+ldrDzW
wOitwbde+rQq0IJ6xy1PV4P76bNrFk5M02k88HAgUT76qxX8EsfZVDYOyTqEjdM5
T/JmPNfdNbeLcoVAT3WO6evhkloQyB/UWq75DDXaANN2sApu9pnSmb48E3CZGt7y
uIB8tyf3ytHuIHU4MeS5Vgu7seWnxOE5Sfxbbv8eJqmvAY7hX7+d/eyVCKmfbCFV
AE5z96++AtxKn69gtk//bk0ItV3L04y+9xcyvnSdFzHjWfxAVHtzo+xBVxl0k1/b
Dnpei/dG5xVG4wYQgRjD7/I+YlKF7iFcPKM0oNiEvXE85asj4w725z85ooC/Zekp
V5zVbagwvBn1awr0xNglCe440ruicfqfkR47ArqXZCldD902mr+S7w4cWlrqEyVK
h/hRICnCZC2ciRjrblBRP7MbVNmn3gkn8/iR20FxMFQw+iqIho99kk12a49PgD/T
vMrfeBOCvC86oXaWy4OJbuDFVmyJPtW3I/acbK7WcCkafpwDMnGDbvkAe+6GebCg
`protect END_PROTECTED
