`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T94OEQZbzLKu90/rxLMcDE/NyZHC1uv9CTekBzMtOZnrXvqXsAsFNL02Hv9uDBtb
TE8njYY67Yp8ooFvqNUO+0tkJKD2trKpaqy57HjrfvXa9nO/xD+qhTsUtjh8r3CM
k0fbZ2effpdjrpjK5BZ4KN2fdvyEZTGDt5cVUX7cyOwooa8t205AYlIf5rcrxH7x
qbe1357tBp0x+IuLhPzzqTww0GhgAZIHf4jD+W5rHpKkarpHkP5V5WDOE4AwNPbk
t50lpZ37mq99+YooEfNWYrJ78q7v7yCmLlrJkdqzi42IHUIahhl+93UXRYjHOr9c
xAKar4MZGy2hD98xDuknMo2oCft6dLr3U3KUeh+8y1kriAo/tRI0lP+/y3pfIRTJ
rMOgenudIzafJ5Pzszh0XAbuBYqHkwMEtEcDTQiW8Ip66F5kCixGF2hAKCkGd7CO
B2AAU6scBKo5ipMWWo78Hdtvvi62r9xPvoiYKAkPmkwkWaE3k56I8i5I9bxf0siq
+4Dw7DWqO3unZvx6PZHoFfD+3k72/cwwgDFe8Xw60jkomPJGL1WfjOp8HkqpFoPt
GdBZkDiFbvqrsuEhWtV11K3EyPk8EoJA3I0nWOykSmf1P5lTNxINGt0U2NaH80K+
g5jqjDewAgBOL9/e54+xrnW7LX1Qlidq9WdDppWFAW7l6h/RCTg/mWKyVvfY3r8m
u6628haB7oYyD+fAxx4PfMEVJz2p1GkUHIw8AF4CY270lfCpOYH65feNKiKa0C9d
xk5FNEWwqFQnItQOIxTPNdXvdpDtQIPK4wwx4LuVyMOyLJZiqRwm3JxsICToN/rS
f8m/dwpQBlnWghHczRWGg2q/LqPCzZiwoaCxFZ9fLm4XYj+cGdw4az+8MkBcFTCT
XAi77J4X8phfj2M8FIZJ/V7NQaRqPj4Ovq5yr69Md46Ir7QfKzowxYgkT2h3vYLi
`protect END_PROTECTED
