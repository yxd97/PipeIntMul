`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiqX8zbKY/s8Q53mk/AKyKGOQKcP7OqmwRDIBvv7sQnesBS0ST4SctAcmt1yRSgN
XwwCseHJLGZP8e6WSMtZXSc3FdA7A4sNevohoEdWow7BOJP1DfSg3kAPPxmosHBJ
BYsjAcsL4lURtao97Xh8LejjTHBBwkPFNXTfauu/WH2CmANZaQM7z0UJerfd1Hyx
TSAZ0tSb0luIaiHBx1O2JFToDhsZ7aiAj8cWlonCrZiTwTvD/GUdr39rchJqhGHZ
B3JvCme8cladiwFplyqmG88BFlBpe7cMoC9CZDib/qdFDULdstrossARbZ3EMIXh
fAOxQZN+96MyfVyr0An7nplmFLAyZHt7v/pJ1k/nR+g7Rs5xNnEmjRn/jp3yiSmS
up3owrNy/1Ts+xxhUBzeyZKy82HYlYpsp46oIB/kDbWqEhdUK/zPqKw6C7bpm1XW
1tXuE2aFpoIwrXooWgs2hj52kZVhpqPFTUE+xKL71HjpL+f+Q03hXhruY5NJs2Zq
+XusKlLZRmMMB8eXmRQQqAFNe1CNLwtYZqP3FCh1uuc1xVrCJb3P00BFtrykEWOU
6wrqD/wtqFtAaYZhRlvbRU62ovs3PvKgX/ShPfjl/ZjQ6S/P2z7kvX3GyeNL4zkS
DegnAIDjhyxd9/BDakqMFsKuvx3CzTMZTtIsUZ2O8NlxgUMzKaSd17/P6qOqJ8UL
L0SgL5NaOTPcxWLz81x/YAr3xJlwEtU+8pQn47pa2Ol+E8YrxyvXh8/dpNmDjVGi
WUxKp42ZaXXOK5G7ZQVlmOynr3Pm0p+cq+soCXxFqMF7/knWTcAZwZ/CUCwlnLcw
eCr6tkoUSx2PBnqdJnB4jo6nTJ+LXhcoKxoP4/AamFb6gbLR8jHoamsse0QV8LBR
nGayKg2gGmNL5vh7FZzH9ftvK7q+CabXKT2OrvKLVon0wXLdOSfpPe0Ei2kk9IOC
MehxF3rkvg0a3T/1IKRZAYK2aGAEShA1gabneAQzJDHHOZ+aq9uN7YLa3Le37+7D
`protect END_PROTECTED
