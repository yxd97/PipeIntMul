`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbCeMD6hdtjNJUV9bJUG4nBnoa4rkVbON0+452Nd2KhZTithRXdYp1d4V4gk3/iT
035bPJKtfGC5sWpBFwbdiwKpGKTmw5EGJuR4zKrvsH1Ze6jOZdwS0C8KeR7KYKcH
KH7rIA8mY9tZdkPpdzMO4x0mVBqT58vzxisNHsUKQYmRHKi2oaerBkMLDD0xGUMq
pFbwjzEzjqhWPjgdSVqxJRHbwZD4OVUUvPvq7obyL/uH0iDAysXVbiECRegpXtWF
OuXkgvqnwQ9UYTRjQT6BINvyP4ct8WUQXDV7DGg5zKb/6nYwVoDR1yV9IUNW00kx
GhdACoEC5zMVCnf2WEgS3Q6Z9qvWVZlVD5wrsLnAr1UurO6x04pujHRNDE/BJ5rh
zYldLU2slMboloYTTYneJw==
`protect END_PROTECTED
