`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
saD2pIuEjDW6J9S/bLUhd2TpuQzeVqdhCmd8/cZRivfcQyEilRBA4YQcrPBkhqPi
8DsudmJxHbm7yn7SaQNpn9y5EkZXAEfkTArFHLoSie39Z/hhjEdkteZjVco1LRvw
HCFYH2/ADQ0eH84t8XUUSCXUl3p2nRy6+D6JbrDXZ+FWcaShw+6zFf6cw+wsn5+a
pLqHa1JheOmyl5jc3T/OfjNh0QeynZDuH3LOtCMQGf47GlRnylgwVfXa7hQQv4Il
4dP4r5Pifzx6kFlHgnl2+BWLHkWdwynCJNHU0dLE5opgN1SGEnQkCUXvyjtRJNP2
1DzTQ6hbBoLaG14AxIy7/jsd7SSlqMU8W/+xZgxAFaC9cq/hItJWqKhb+/qw3CIX
vPWI8eNO7JRx/0MaTN7VMYG1e2OH31E1ArBxsiaHdWi1ZCxOLHIABVRyLUlOCx3s
39GJgdOvxxUTyI7HeTOiRFijUhUCHqZZD1HABh0dnYdfCP+KBC8kl2s/LiEGgckb
qmUo7cybyIHLXgQhG+kkUMi+4dZ8qaOXp5VzDRlR1whEXZKyVrYu9Rg4T9D+t1jm
rg7QLLcSFYSAvrO07qyuuImDXj83GLaPdw53MH3nGa/TjkJPK1vaQJWebJ6iB9YF
+e0CdLVV0xEYVrzmkQl+mBVaqFxPJlBJ3U5i/d5kqv+HGyin3zy0np2rI23ZYoj8
YjpUO2GHJ7tPtRUbeVWYfnllDQFib1qp3+CZ76aCQiMaJ6IB+n5q7ZNU7peG+YyW
5QfVLJ2hJwJei5WsUWH18AR07Jo5V7Vy0GMxc5+tpsszuBs/m0sOARhse5PC/0T/
1Kku48HpG2hF+DUZ+4RiZYrMHn5g4VVUefFFMIqTbiR0CiNZf+XX1+qLnyDoxKcD
CPAohzZav+2fg7VcWh+XzGF5/X38Byh/b960IllibHsOZ50UGOyrIFiiX1EMnFAR
`protect END_PROTECTED
