`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3QyzPuV8QWuBSBZtuI3jtt7C4aNQTsvSz4WT3rcOZED1+fFlbDsKLjTJMfpjqU1n
geJwn0L1sHCs0Pu7HsppoEppQgtnQ3mhebGXQw/2pGmTkdqh8vAe9EI+E4XNgyJo
ay6ATQDFTADP+FBLdsIq1M38W5i5d+efigIngEZfDdGOztQEcysKVjPbaUU2RWhp
lBbyyXZz6PSuYPCaluENrS4sYmPwGsDlf0Zd3bB8Apc8JqAiL295H+szrTvB8ixc
wldIi3VyG14pJsWljxKHxlPsNM68WvtoNnS8hYY3n3pSZY8h9qfAIPB7SrCHLDIV
q3K/mDaUXj6zVshv4a9IcimVLcQxnWotztdwK72S7UdlmHp6pym0/NBmxmB5Jq0L
IDJ2+WaMWYrk0ofIcEa3hQ==
`protect END_PROTECTED
