`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oI2eecashJylaWduR3pTSIJcq7GaQtAWOXyGiYaj/ufl8IuCv1U0WxxMTsVixiKT
o/2lRarq/hfGO17SemfOBlavmNPBsDk9i7tkJyDJCrJ6cOcVmclhhoPH4roGBWhW
GzwVaIPHmxSSl6nXTuPAUPHM4PMgyyzFIox1t6QGGaxtsbZe+FiQQRcDuLAbRTKO
akq8tWVIivGEFfouSxYzlpc7MvixH+vVI7I7ngHoAZnGxU8oA92B1wDzPkMp6AXr
wzqtNw+xuYnDOohqSgp8U/HG5AHN6d2JDKn/cbwF9LtlsjvDDkAV6V+iILWJMiJN
ejOg0S0mPf9O/CeWdp2X1XZJlBpf+EDM3PgXRt6hnxTwJ0RLHP+6Xxkyti6HGYPo
e1MqgINgIeZWEDZYOPQNT2TSre4cS+LiVmPgKbJ6SzXkUgVlOa9vVw81e5s6n0tr
gc3tEENVCJeCnddAmvp1MRTNkpA7gBDW4Cpm77PV9f/9Gu54qG4VuWpRmZIHAk+q
Kp73aC2FpWoqTuY2Mj319e9FuwfTw6ZpPW+6zfRqYgO3zl4w4hjRe7Zmw/1V4UHT
jsvzp09nONrr05td1KISMQ==
`protect END_PROTECTED
