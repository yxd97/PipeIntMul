`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b3VRkM1QAGcfIBOtTwhs4YzxSAMEiQ54fL3/U0IGJ5yb/NVAmx07aVbYT4fMCkux
pv66LHMty2ePIrlJAx5HmeZtMNE/jo5RrJMoaPJqOMVVwEscPhv/fDdneVVEM+av
iEuZ7Mpt+GVpafuIP2seMkgwsiTX0GZIK/ZEbEo6UdQxiGvHFf2SHOvbdCF+TVtT
FsFyHy5xhS5UCfFv2HTUvCrZmMYxqNEsiw8WgucHdOazP2pxPvUuIVPHkGVKT2xJ
wqoqIJ3Tgb+wfJORAxb/R/CTW82owjHQaSaMIm4loqaCgnt0STr7qCfir4WrSDLF
hPyDmxmxrDBLXtmoLY/yaHu+iNqaiBLovqSYvWJN8HvtyvKCeK2z47Lr78IRkuKO
27pfyl7t6P8FQw4R57BgHlAzkSvKOkT0SglWzOtfRolm0/E6t2dkHIJ3Ysveec12
9uZCzWf7yq8G1J/Oqo99o9pguhITStyoBSBaJkzQJoHYHK8cEC8dDrSDLOUGOa9E
rKC4yQ2Wfbs6HgpGv5M0QqeXNIniHV1tJtczgfBw1dVp/Kq1mdZKMB0iv9N66OM5
vUUk7u9zS9iTirejG3540XsZ4DftU5q+nhle8l4hCuCTLoEEvkQ3TonwKGG5LO85
MtzBLQfsKmLvpSS52XdRLjzupamwpEeSxSjWKhzFmQpgrVMwfUQ3WNyitGzSYwX+
9Diuc2gQHlqVkbSX8/qnxQVRX2p8S1PqG8VHSJEobwWFANlG30zXbil8UmlVeaAC
kJRz+aXhFHWXEFZktEhQjbETGZj04X8Zu13aXZK6euzW/FtnI3PV3/LFSRy7vK2n
Qi/Qo2yvHFdEst/kWuhwa2gAXVzC14QYSaY4uzhPlSrNQAnFPponYQEkD+g1lj3k
WppIHvXI1zM745cfF5Lq8jQqkdnMs0a37uf+GQpvX/u+JFkMS4eIYWODkYhV8MOY
0Sz4jJygW/QIJXi46wl98XdJKWAjvbRdaJCAzEq5/m2eLZmaSWcrAFFec5XAM6Qm
TbGj14f1Y5RXs/61OwbmHlTRLXHfFRWo2dNdk+vB1bMMd99WhqxL4HtY/5gpzvPJ
n6fwDrGqSdu4N2H3DP++lBx4mjOGKHCTK2+huI2n6JRa4dHxDxWX0CcuGp3+ccx5
2Ah0dXOGrxE+w8q7OVfba0XvoA1Q93ujtbc6MeVTsA2chIQdfF1F5QgL9qI2C0+H
lazjJJ4Bt6AG/OQNi5i2mseCOxycHo5J+wqVZZcv/lQYE0JULJuvKsFvEV2PPe6L
XVJ7CWb1Zh5IgDSm6c0Mkm0RC0ZFuccIkA5W6U+6ClGgK3IfTqOawy8b7A/7wuk2
6vYca9lND4BwxPh9ar0C4o6NcDaZdMUVXnhMNR/ZworaFj+dixkPVgGEyi/9mcvU
wDGWD55vZpMi7Hd/yvM9HSWGZCY3+Phu/VjVvZm+rZ+fR75Zy4yMxrSVThhOKafV
5POI5nT9FWUo+n+GohQtHJ+USWVQO2OjKLCES6/EtMQFszRDqOimaeZjtLBpCQ+b
NCqd3HlJKAX2U6T41WpvMas/vHtc8gIe3uz/CofFqQEcTbPec8Y4820O4q/Tt3Z3
XaImTWc021v3Ja8QSLQf5to1Np6l/c8UrxYh1gTEKGk5dnkS8fbJrjODmR3VUvxf
1X+eYG2K88vy8xkvIEz6DQY6F0uQOxYPQbOdmnL+EZ13U8g/nLajSSb6rTaErLo2
ImqbYpA9H1lJnIvT37vLNv1ha68YOg1xDVISVETzyvJHXhvQn7ofQihlJmuItj9h
IZ97pfZDV0degd1oXW3zxy+6eMPghItsW2pYVyVC6sTZIGrCsnGt/k1mIIrZ4sjM
BYWi2X7gB7nDzXtGras++ZQtpVWHOl0UCtp2EDQbVtG+WN/CRaxiZ6JcduUgyCot
t4AahMsYRxDpr/r7RSvJvNlf65wAGpG56hbtOET0kmduOXzdwiMhmVEPsYIuo1dM
m0I8x7bErcl4lHoRqNfL21cuX0MFzTsJZWwx5xsA4ghuZJ2YgHPN8Ck7IkRe9MaD
90+3QExXKVN8JexOLcTkF9Ir0M3iuMCOwM6tOY9EOiUh947MArBXdxDEw2SabivR
TLEvYpyOE8bVqCMusWNRlYjw4AEodWNbSkavapbpqle9tA8lVoHTauiaIC18OpjJ
l+BxQ9BgQ7Aw66trx7ZfZ0DHGdZqLPQiMV47+ZuvO89I973ibPiX5aRo2drYqoQw
Nk3dRCfd4e1EfxG8GShQOcqfT0J95kGXpWZqcN9sEmANGr5LQX+4Tt56L3fa2Cje
804qS69vI2iHCd6YEZoGFuLd9WMsaVUDdjs6WJzVNUWOFRuN9v9oVx/upTjoHm6U
0MKT2+ieYS5Utlgfwahp5p24gsBhvEyW2YPqzywv8slnx2ge4XjjArMRxJ/NiI5A
x/Ha82MmUCzi8+cTUyQmJcuxNvp8eQ9bnA2nEsoFsKO65iwkSWWYtAEFsSYUaqeh
wKb6H6OifaukTppoVJL3C7i4B2tZ616xcgwWvMmALSw92pZyOM5Yl2Ny9wYjJQ7v
7fXQVwiWZHv+UnQvVEq3ruO1YJgnOv6JbA0JOC0YJLk1jz2JSRSdcH9PLlyw3Qzg
m5cKUVv6rGGiWnnsqB2fVFV0fzWH83HHIk4exWdnq1tFJqmqEe+UR8YZcqbRpKb+
cKWtCgdshKHX7Q7VtoPC6ooE3zeyxwFQShKugU170NYk6yFkNQ3RJXYIgPUP4nwQ
Wuqojr0FotAafNbQB5VGg7L45nk8Iv2IuP7ydoOsElqPYY49R3LbR0I/WRPoo5ZX
1u3PtUIbqmY0YfmTsrezHSfmLsn6K4RYyLhycTgRdZo=
`protect END_PROTECTED
