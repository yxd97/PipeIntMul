`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNDwGK7aUn3WjC9bCQDRWSeNixePlqgdtJGPAAYRWkx6mBNlCdIWcoTKzOc1Wk8d
on7EEC0sH1hgfGkDzty8tEGieZYTWsExo1wKq9aOUMTO4O90THrUQgTosJD3bV9o
9+1uEbhH6WKIXI1vwP2WFTECpYswhS8bdCtc0Jd+eJpHLKF3sG5/83eMJQFT7xvU
4C+hWqpRLJJeOK+rl0HQ4FC/XFg7mf38/SWnsvBc4g7zq4jBwyjZ+VrlvGYcDFvb
KvflI8AJO6nz5gK19QM+ZNxPMdSXfa5wZoqP3+69h+cIJ8eorUNxJOoVDdVVhR24
nQs8fh1dSW6lFoN0qAHnMJ+TlJMkVxuddVMDGDdnJ2uuw3MM1XRjE8PWtuPlEJeU
HP9/aKMdfXC8TervuRzHL+j0ugke+6j397eGWkiVEPZGHIvDNthdM4yhJ5miCTVT
S3BCsiv5kFdM0P2clKkpdgkm6vAZ/earw5Tu5uVlpT3TP+Oy2e7XN1Xa31Z9JrXI
dsASFWHuEX+eNzAX5Pxpvtvr94UImrgqex5+gIj4PVbySgjZaaAuBTKyyIfBVvkF
CSkLohllmGWSKeDy+nKX7cIkG9FSMRCgwW/sz3OMaaOrE8+jen1q+RkRBC4QmMw8
++Qm7OBGOWj5eRLc/olRR4g21IrLXxMH3K4Dd61o2H7uWZYkjJ/flviJ/CPm3Env
SQYgLQUKEQFNkXG/Qvp3zekomm7/pK9F1iUUG44G0WqvCQk57eTNZc6zLCT/Bc9R
Fa3pecX8o2mYOxSpG48UBsOWpKy9asgfcqcr5OpX95xGKqLQzGjpHSgW3XCzMGJd
x9jSL4q2mrVolk83kkJiCYK9fnNpocB+OD5kKpYKNzhEoPOnJsa5rEE+lMdvowuk
7/yzjByFu/PM3oGPdHF6GF02NsOI8asVZAZF4W+mAUhQmnzlhVzn8zPDDb5jWjUS
RPhMMNUKYTLTtVryggvpopUDEcMRsSb6LxM5wccGZ0hM8vk/0XVdaAdYJFX2ELJE
v4/w6i3rIJet0037tj+l5aWnbymvfAWbMbUS43ptdFeWglIPXDCr0FFGQAOPq2aY
bIomnLj0kLcQWySpnsIImZQ1UIM85q/Xa3zD3+6sjz3M8BzSApHrV4F1DMNJuaiL
flvAdrSjcr6mwUf81nUWv4DshD7stEQM/JsxmCwpxwOMAOddDcy0PLWRwvcv8k6v
9N98f9nurLMOKJhY/13JMSV/STap8MgT3PG7DpE+FyWJTrE8zFXOebrtEs2NC8B6
AS4Zb4/LSHFUFYhGzQO8F0bIhBuEzQktWGbCdCMktnPQ593CeW28ru7e9K4vDSUi
50xpC5Uxh/+uMhjSe068grbgNYjwV+Gkh5hixtCBinRTbZRoFjRaJbig0idN1C4t
TUE0yt7hHh1gtvbtGt3Z812mDVtDM8UQ/Z1bqQHkuRcvA+gMfD/ddtEionwdxe/h
KcZEq+r7gb6fyrO84Xn6tY47Et+dtXW48aPZoXe3kW0fDNoh+8NlBf8mms3u94KU
FHj6OA3lJ5i5U/MDpE9o4QZS1NmlZz2ZPw4Xo5qZSgehbvKwFIEQ5carFR5/N95/
EQ4tbQFsgJmqrmC8vr7vFlk2V7KQZUVDLKrLIOdEvCq8E2cKYhzpyT8zMgL39YZx
if+wlilTfW1322oCw94vChLpW2nFK/342vFR11YwodTlxOAK8mB6mgzvA2sB2h8X
kOsn6J9CAdvMJMjSKi9T6oxXBzsEqlCxq2osdXatI/CSdK4If6GSbC3A0PL3TJsi
HsXTDFKd/LyBWOk96kWnZAEYGJMRy5PGKlONKKg/S0HBq8KGnwBVqvfJzuBx+6ms
bAdUt9HZuQ3OjkQo3AyFyTZrLwpU4ubTFisVmWUYnNDQf9C/IBWPWVqFBQ45/nGM
MC5UVEYBqR5VjyoVddbQC+c4KklaQxs4iiCW1z1pKWrdsw9eY8sSdEUdyG+A9bQf
2MtBGhsRWE9V5kJXApvBZmGZPo0SonwZrbhCxv7UAIWKuztAs/D/X7HQbd1WlUhE
Jj7DJK8SV1aFnCuB6EjvUON9+La48x3T5PHazkFjhbduc3a1HdSET0ls2LfzLhY4
7YooiOezVtWuoMZ4FZZhsh4EeJvVsukcNvYh8u90Xrmqrgqu5LSR+IU5LCjgAd/Q
WegZ6nOG1dGdXd4/2UYL0v7YR+4JSKB3d+IEHep8B4fqe4uWMbFdZEotRMckBUK6
jVowwyym/nwm0lrrkzM3IRIZ6MyAcxOtmxPVcCY17CO5wRUf1AbXQpZsFIZWeods
29J88+0T2r7UsJBfV/YBbq05sxEiIfWnkbvpiBWe91qwIXtZMbr7TUiI6u1jKZcB
gPqQQadtc8RyA+so1NZWsDBGp3fsD55/kgM78rw5qHlAOKbCCX3X4AqelOMW7dL+
ge4rtOy+kKXkwEP3ZwU0Il/H/d3U5/xNPGDC7xDeFKHjjT8+EGHHLIKo3vayQMCJ
ubwp86FXaTL7kcvPtAYy96YpjAhJQZcR2H7grPpbOYBqTThkCTNqsvEQa52zWCJ0
1xmgUZEB1nZWITGrAfIaWpOVMJL1nZMmvNDoehKJrjUh9K/BogNcPfBJ0R2aMFUB
pCQ+tU44qZ9PtLhbzTIx+cdwCQxy7h6stBvoMKhsCiJfsm3aKKdzOQBBMzlN3++a
X1+LDGtcBeKVmORnhGSfrsVhZrbn6Fqdl+9GWZNpPrmAMSSpISQjv0WbzzIjOF0I
q7IiZOCMSflOUmK2zB0rRR+9bDzdSAAhkDmPBLIS8L49GhGggo/BVsNTDQZkulfe
JmEyUvHSjgso9WeHTLLB3EUNjXu0afgkqvcRNqRDTJraccBndXPrgaC4fGlNr2oG
+wWZCDlViqNH4vYdNuh9xc9aSmH3ugo0G3ukMCyQXDw1p9YKM8guSAmECNsGL/15
ZAGi/ZnKT88mrt72QFqRK33rnOXunPx9GnhnfHtd83OrTWtXr0vH7e6JJU49QiLP
+AzNgtfTsfw7T1dtk+5Oz3Sk/IEGJY4hugCSsWXTeEXYu+DEsSpAdwQxzKmIVuS9
OnZPr+ZE9MdL6mA7o9M1Q++mOe984e2Fbo4lwCFNAbOqf8KCpvxAmnMqCXQqUY9q
wmFJpQInzmYfijqfL5EFzv2Pe9dSnuoTkLI9/E4/Qj/Q4pdRd/QzTbugTpyTKn6A
lZKkZfKI7jfEmmnqd5LDjUk6I2YRq2M8STgp7B27l5ocmNSHGdtAjA33re7T5UPx
CH/n2aU3tTa6/mLQmhVCxvmVwU3nNMjY1hKAvtjQ2sjW14OhqgwByX1hvbJwE8CW
qqEAlFxDQmgIJVufLLFYCZwRLyRxmNvLPbr19gUdgskY3e7Zn4YzCawAZj1V5K5W
p5IUMmH9L3fzK9+xuD2xUaGB/EigwVL6b4mt5BsAA6BPcPkOli5c2Ama7daWt8KB
OMVDtVHvE4nB6Uc8fZpKGX0UwbDUSFAeTzCKpUFk4nby1p36Ya9yuG+FezBpaiN3
povweDnfMOmE/jYWXjxuNaEFXOf3E96sjeZqz/v8BdTg5xDa9SARE3pkE8RqwzXh
upZ5JNbCpcSCxjpzh4J40u/ZAEGIjpoEDMC+wFU6zNA4gM7WhtO3Pwb9+cKPvMhV
zOjOuXrArm/fU1nWeUmgTDT5qksbIoVyS+/ueGSY963chL6vUfcXUFKCCoeh87RM
Mq2z2pzFnJ6j++D2E/xOdkNsNyRgd1aE2GTfvBWqdK0icPOhB4NOPFxjBHxcIdPF
XZezIbxyqimLWUAShbXB17+rAU52hOMAOA8ziEXIU4AgmJGqdWjCbBPp99V6UXxw
QGCNpn+sa8qZVJm6M+S051kF6k1t852ScySl+P3g1jY/clFNV6j3FZ1RiyNjPT3S
pa5ulfL5xwop9oFvVJDlR0wy10IWLVhyBYJlYOKP/As/fRkBTE13NoZhJbatyamA
Ywq4ai08Te0L4PlTJbO5o5SCRvtng4OUmHCvP5CjQB943dgmTBzYj4SDuBnqBVXW
u7+xTALz8tJoN5hknTYazdbmtBUUG5xak5IVwm8n+Jqs7ggFfY9X90cc6cmV3N31
iaK5G11WMn+urKq5ClCHizd4UGOVijJIdByADjt5svVMtsx0/vUAxEn7nuPSDp+8
RIE5L53p/B9btGmIA9WdIyGd5SlNTiKFmPpRp0Ly4a1tBA5neKogXu003xLHGM5W
AW6+54GDdlS/KZ5BTV8GXTb6uKgan2RT/WG8t4HgbXNM+yja/t5MwwS81brMItEf
8PXA0Z4qvYnzi2AuWGEz89ORMn8ACJSRGIVo952xktwG17R+ExwfKeZmO2ug+9u/
0Mf9WehP/4yESsxQULpadkS5aFtFtVIl2IJ8c5GMvIX4wBaD+dwO7v+7mZTofQgG
Pm9RwnsVIVWQcGWEa+ornTIo9QNhfyV405I0N79rf7J3C2zDgFZU3ug4bH1ZeBiL
KR6DzJJ9MKsbSm6RdzweTizroKCmo9eF7kg41tW99ooOn5vt3ZoM3URf9K/Hw1I+
qMurw8Wq0LjqPZ4Bv7muHTKloxZ8axIHTRwaKDQlYeo5LBxIsdRrOSLMp/YP0mWr
hfRavvuTJB/zAwbKytPIKz3Pg7h3iUPw2KLJT9+6kFOcESCsbRk+ebRf/s7XAiEr
B8zsq9ly2CmhQMKlDAiElEPUuIDs2TmL9iLD8meVP5q9VSqqcv88h55jmhkvEWwR
KO7etEJFdRAZJ/+Ee7d3o1Leq95N6yqhTOLD62wvNUwYouNEs9vV25I4JEyEtw87
/nIeO8JcaPLwmNz34nbtGhSVcy1AzAhUf6kD5WM9YGS46XD5np/RjcIDkhsJzNfG
eQ9yl8AL9ewmvkMoyPtr8S6l/mkIj2hCgAhwtWqcaRuS/3FxYGD2kUQWWC2ffnnK
t7RDmnctncAoRTmqV4RU114jePwc7oRVdprqG9IitX96kogr3mennBBQNKD+OZJC
XRjjJ2bcLOJtcZ8L2Tph7fbYknaMAe+0VfbLhBFjRCCy/vGP855euVegtHcYANg4
VkcSlvv++9GR5fHcySlJWfLW4opUYOzCoUq2i4Ga8NEcnDbxMF4lRxaE9/SirUR/
J4ZMvrF2L3lNoFwUnW4RpWnkSzdOZUoTRCYY0b5rIDmcUL+T3G1kUwXBe5sLilS3
nuzXlfBeaitm2hmnxuGa2MxOwuJ4S7qsWitHHGtK/UCiQIaU4Eh2/9yflCB/EVRF
5wW8Qn2bhce22V5Yj/D1Fp1vh5uDSNn+GE0QSSFhbkVJytzQET3RAtjXpk3Cgtpl
fTblgjs5LtABOAUcEZMgXB5unasW1dmR0hvWVe5ZJNvxcEmx3AHbGvQ9lIguiWQw
c8NSgIxFR6yxykNlXYgOrRHGcPyDYtE54Z6idQdIBXuLDlUVLicXuYlXQ3XwjoLc
UO1BuzeGm58e1s2PGIqDGdGgc0zqNgnb3MfE/BZWJLwqXTogazkPK72L6ExzQX6h
BxJGyvR/VF7g/SkHgvdMcgFVj43dQhJi6B/ahFFDwT+tpmivZ95B0vrmrF+GUYNV
Ol2ClhxsL5zENXEEIgHmWxUwCZdmc5Yh8aenHhe8OadVIAG9iKP/cjIDrR9QlODD
SKHklsYcRHQPq2gjPtFQ7h+vmCRAtP9Uii1aSdPHOFskGIzBX1PdixsX6sjtlDhp
HSNy/asHiq66dkBIzUTC6hFd6ns5Oru9/RsmMUgnxu7jekGQwhtuA/5Gwgl9gerx
SiXAfC4PUnXSH9JJxYwL8WbBz2n6/FD8jvaQH+bsrT42xOMK/99dw3s5lOQbWP+e
Eyegj2OzM0RYxtMe+MVTwXWHeze3nmccBVZ356ks35TroBldCpHPKo53h5RliTQr
Y4kkogRBm9ye2ZTMmYKE31X2co4z7SMT2Fwz2Jd8St2+pR1C8gCyf9zJjGiyXUP1
vfirjEk1Yb1bru85GFIeBL6FAQO8sWU12in5TeI4Fux2sAzn4Jo9zLUSzarmXLhB
9jE5k+QTsvw45Gl59gxk6ulFLNXfQRv1hiDdhCWTWlFXLKQkRg7bVsUXbefYRfOh
CqHtCIwUoVDJYMkrHWwx+yZrMjrDgYwibaaRz+/VjfsPmgBkydVH3zuvEmZ6h747
hr9ryTzbHZ/z0kF+MgY7J1speOdSroBvMkPE3szFlg44/FAUMxAHj7RxwOsyXnEW
gjp2Yv9gkg5uuFGHHn09zuoZ3NbPXqtZdwNPSMnfLTAQKnSlrUmoqfTNbXJa1vb+
EV8ViU7evRp2eRkxqpybvqRp3b9n3jB2XSUuS32NKOUYf2oxIME+69MDBEaDz5aU
7lqBJpKALYEUBCV29HR8sOAdUEegaguZUqOQ862SqrOqsnbgaArNHaOgJeRwKkM7
FZe+axkZ2+CWaY11UNSgTS88kSYAd7CvYH1R8vXHJZEKo12tTnfV3fqAfJgiZ/Ck
6kHhV2zDx0IEstF49TLCPgjU+fU/PTZCJC4LcVyBOAx/Cig606E7z+QK5Vugo4LN
mXcHCeewKKwg+v/+Ls3uJECFZQvc7CHJajE0KdNqnNH0rPQs7nsnwDDYgRD+87qi
Eb15YSwfsDKIH0DdfvpZRrb7f/sMwvoIxZ5wQtuNl0/ZLNY7AKr/8mPifmCh6sPU
B3hvqiXHGb37fOh+UnQIB54F6E+gOEQgkxU4+vrv5v5wm5qCwNHCwCfaPqIqPHFd
w8Mz/8G0wi1ylw7vEE888HUF8eH9Yf5Snhd4Yef4hHOQKk1xxJZiqYgnhQf4SX0H
DHw9rKsSHdc1kK991zX3E3iRqtDRwkEnaf+LX2k8gKBWqQrF/FKDanv+Jrrb2Ii+
wnVvtTnET8Fk13EodLmRe/c/qak5pcGk6zQVG3P4Xs3gQVkanQdWJSL3snxlXc1o
z0jq/8A95sVNaLsPgKNqS0BuzTRX2px14KMuW0vLr8istl+GJnlLLp80e52R0OJ1
V913cvJnjMQtyVFEcsx3u+KK4DW0PAf9uVVIxmiFrmbJF+GF5ZRH9zNZAh3czFh0
JczZdloAGRMV1TSg9G1/hOCyFUejeuFYSBzs5IMYYz5DIfjK9AHu8NI2Enc0wfJZ
caG6oSA5Lae8zT6lYbbkt32Px4NlzOFNVJphur+v49lLwxIBr3LnqmO39BUqnvWh
jd/oUC50/oLs5RNvHVkBk4lKu1T/l5nT5XkvQnaBqqJUV/SY9u9fpbXLxnjkW3ZB
VwFdJ3LI8u89/arKaJ1Pf4SD+cCurh3eBBqhAw1KbxBzSrbOCX/W/0CrKYOuMKHr
O6GKEv4WweXyQxjJJ1Lfz5AGkxh67Fmmo57f5K8gh9oNTMnsacYxb0MAkpbfErKr
PoVaO4BeRv4mOa0t/UDgBHtryrPGNUm+uY4jQACg28vmq/N4DeymLyOhZBWdke1C
BJ+EFbRM5b2LAVGS7MKpZ28cGAEMj30ePFTUc0FLgZyfhYrTZ4ow81ZVnoLgwIF/
RCNIggnCtpmkzJnmmXkLD/Iqwe6G8GnhnM/wQudh2KutmEUPd/WPeZ9flug0Pw17
b/krd+cJTAhFUpH5Ct1fQW+UQXoynr3iq9wcLNTrISmRM0aVGlsUGwoBeNsETQI2
MIm2Zb2ZWx1ngneaBzU/xbAwF05FUFeSYCf2u2pFVbwv3lD6lfEwYNYSRpEbG5Aj
oaLWNOgsz1kIt7Ro6BPWAIBm92ehEJJ5EPJic2Wf7W1kW4VuaDaS6u8WS4ISvK1+
eMzNebw8e7mFUqj+KWF5gZaTB1UDquFe+nZrMDZvM3Wk1hvjFujcIVU1GyLqNBtx
pEXQ8eiA6sON8nUkrH3OJFMWhCjem7zlBWvDafR4JsCJBN0pO6aCEhXSp6Ni/uoI
uDuGXJoEhtWVImG6fqJAWv1BRTdo5sF7S3UBRWcPQcpBWPMAHNwugccMsH4SaIfc
sfALo19nbmTEKLDlTakLoX0N1+vlBIUMBaaK2GKcNQcNFSYUrUO9UiVwauMJGvdH
V1Y+lKflMNcp+KmnW+SLIoiEGciJ92TCzUy4ShCMKzU2plxLO6o19yNvjvTeAIKR
EPBw193lDd7KiYpYeoMc+56HnxX93ObSJdtzvutm0rRujdQuT9uAdzQPiYgLF1dj
tbO+/f5/dddnKh1gK7bJsHwmWVRsNK+zS1YZUmkKGrN28MGQyx/y/a/+5IPW6/v1
tIKQifIT4smOEueVrnN21VTwedJOODzAkGjFWvSYrIoLIp1vvHnMKjS2w3MQRj7b
wk2bBNRH9Z190bJqECuGcIa9tKmRzGpR5HhVp/dKnDjfs1OSJNDkD6QbE42RlIwM
q1Lgfpl4Ab4PwURFVN+FXy1+zdxeGrw2nw6sW6+7qoR7HJapabxVPKV+EtYRR6rQ
i3l0MhDGXb9NFCbl7qnyiqvki0x9XDrRCAySsICW346HbSWnvBqT2SYrJ7A0oiOL
+wPbN16P0zv+b64dn6UBKhBezpAitpgPZdqFEdwaSEoFKeaxuDnB6ZOv5OokYiaM
`protect END_PROTECTED
