`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjjZ30enWRlgKQR5/8yUyl0bvmdt1nCd3qx7XHoMbaYpzsnITFzUSl5KEN7NDh/1
HKzis3k6D0o+Jq//twgpjzV0sj8TQpkowZdG1Ag0MTJbOVn04BSQl/G2XcvlNH6c
yCPizdHcIdOPNFH5QXQu0i8E95NCrv80PhWaemEeQFDVI+gWFeiP4g0n6HUzNmdX
QtOhioqzXiq5NhtQfMwWSekOmYwm+OJ8XappGfG1rReqfpOA9AZOg/7kjgkTuf7Q
FFQ0EjfSCW2Ot3s964hD/GT3QDq+lWbZgIlp5vEFyzUzSE6D5wP+yi857MbnC55K
l91ohWyjDIVszsIp5c8GnshEvn3TAKC0aFdPLjGXTkV7KKnKUzbtTbrsfeOIeeS/
M8Dx1iqNiw5QYA8DYcCXgoIaHFAaT73Un8DScOJjMHmqFTfbncQ5BS7Jawh6iAJo
cU6s9IqzU1/yvBTBZTxuswpUFMQUEFBrlsWvWY1NENDi1vk6nudT7JR23HUREzXj
hbab6TSsHx2HR5VtAdRM1cmdqaI0jeVXw7wv8gkJV7KSej1IvVawEtTCs8hQvofz
64D7aHfJ0EhTX2DsB1HwG8rdG4fNUiSY9LQLnky9+fZNEOLcNWPluMAlcE4Z+d78
RUm+CCzOH9cbLJebggnGki56/G3SVJ+Ib+ys3e2+Fpz8rPPBkhyTjr4GPhDlO0Pt
5Lqbi7sjTLLHscQFIS42tJV5e39EQBPXfE7l7UmgaNEz7W7EDZv1CRtGbOLgbnVA
d0TN0s7X45pe6MehV2sH1ltwFIGlZxWBdf2L4VaSNr8wD4seo5anc/2IM5lc5xdo
evNi8O3n/hJQTeTVJmJK0y23bj8Qu7ftQ4rWY6xyjhSI3RkDavYkuo2zJOj8AxFb
sHtm+GwimUIm2tpxrxnoG0RWfivJPdRIV3B15E3MzPZ/Wuhm6JNO4kg5GsoN6oDH
N1hueIMYfyXnP+woQCoCCZM4vhMejT/VUneDZy5b9HqZ8omfVKcgpx6koZS4ly3b
mLrPkiYLiKNfd2/tOJDi9RgfwngPYN88bvXXlfU0RIpH13UgdSNfJF/ISXPjuKTO
5sv2SQenHj+F3PrXzvV8oqPNNathsZgvXtVtk8s8jjAz1/eD6A5kbdGaoVezkJpA
XsVZQycU9ciNZ+LDvHL2thNlDGxr4muUPtrOsuBVK9jMwHed/gWezqaLz0dn3ty2
wnXwW+HRSttc58+BXkhMi4gYazzhUnD4mi/g7+09SFWIHU8QEyDQb/TamBzmnfhO
LhAS3t2CoJWkh87UBoVAVoVwBVyVwD/wDTeEa1OtU8vVvvNWRNR24Uul1tDWaYQE
ZxqlyoCGO4+/PKc9grYJpnhn7XrHH/dqjtAJTdxk3SRuRy75FkDFxH5mpMxldc4O
W8ayZywDRhQsvnMsEn4fohMVSOox1k4uyo45p3AL3cBTi5i2axwbTL8MT6RUXpdm
UymEpE3pNXmBwIsHby8S25QtTs89z6u4dzna8UYyYOTAdsVj1APGBaVDLy/p2oQv
QJt9KRrGCi4VhuWV+lfsHsL/B77fh+wwO0oCRF2HeTQkobpGhAE/oQfJsjXk3qZW
8SFSfqQafnO62/7TdQLAk5bL6aFJR78TvhsmXXpMtEPgfbG4ROtNok8navywukj8
fUCpdBli57o4tmFGyDK4UCTsdg+9GUE3CpkE/jx3IHTRkpp0UiswngKMRltaBiMs
0j0dfZnFf14JOreeI8c9bM8cw1toSE6f3B/NdIyHUE9r2pZWK2GIR9Dv2MpsXNLf
n2rauEORyBB0ldfjHVT1f5WWLt2kAlOStGJLyceYFAqygaWvMXsibYcv8hTGgLmD
`protect END_PROTECTED
