`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1HKnl/4HTmlD/WYqwzPmPcL6d1BPmtRJ7kz8zSNpOKGoXAMc1FrFVWddv5fKCiuo
zD/zBfwN8kGZx0O1AgnSNOJODiBZyJXxUjMZlJYgTiKE92u1tUSDh4lJdOO6cfpe
p/9ohImr/W6KZx1VvuvnO71oQqZrj1S1x48yLblVyZioC+PcI6Y4plllHi8byDw7
gE8s+SVmTflcwA7VlIKcY4j4FawJcKNI+Ra+ZozHUzIaWeCMCRo8IKiiM7g94iQ4
v6jmDYNJB0TnzHNV5T/mqi7y29cqg62sAM3btNyqbJs=
`protect END_PROTECTED
