`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AjJlIYQNleF2DXKyg67pXXSrdU7OJyJfGQceSZN8TPpQdoMv1P9y0Bj3JmgjMecE
WgPFyWiL6ORkz1AaCRi5Ls3NG/YLUVIK7WcpVCL8mcw1JObI7Zpi9caN0CmIasYY
KxFf79w149vbT73883gp5MojJv+6riDjkYoaUNQpfCNmlDhrKGAiw0R8G/ciu6j+
AKKVLGSSL2J6KCdIuTkPOMtdItYjE8lrBfCOsvndGcJJdln1t6ovRHX5+/5E0aqI
+YHMuuUqvHWMIhudQ+/nCJIjKpvoC8u6UqJMHIUA6KE1LUuRFXwW4QqBMWz62cHs
KSyko9HbwEL/E9iHaUa66/wGC1htIHLUouhqgScnvlVVZdEzhPw/lVkcV7aN9dRj
kOttM8IBaiiyzQXlcf14SNHPLxW02jrd+qnQumezgXARiCdiPbml+KEn6E5sklAu
s3rBnEwfLZba4F1dM0XEnjpK8L++3mPSgQ7azLXPbnyT4QByhFcrM+gxwWAD3Wt9
zcvlay9oInWBpPUwkD+EChqrvSGUDfkX9O/AOqCEi5ruWSokgciPgFCnXOeeKHKF
h2hCeBdKJP2jmybtE0mtgkAJykpzWqImHjtOVvLqJozZSyXNlnDmVMmJ4EZ6unKk
2Kp7qSXUOALFg8ZPwq72cihyP3SnfOys/Q7e9jsvCxA8R7xaLceYI1Oa7JA3bkAl
2IOIJiBKBDdm7jQ8Bm+jv5vLo850Ky/oPhWqACqJkWYAhH/Pw0Bp8MrKqV3Y4QF9
v6LddGvbjpaXrJWRBm4/3yUaT/+D+gGVnNxWf8zEE8d1djjiPMslboyI3kwR4xUN
ZoIOKM4+PdoXs7xB8fVIaUEGl1JwloQVwdCLO0B/gGEH8Hs/trcFUCuYV0FuVlqx
FSgqqHldYNNcjTTOPtgmMocv8SFanjQbtydAk99n/mboSONK7SK5DNUnBxcY0RRS
sn3BQZn9Y4Rv9w2fIRkeBNOKCMJzGDxDCxKEb1mw7E6lEO3FQO6Dwhk9D9GF8M5+
7IJjf+zOsvBO0biA7S/z8retTTWnmVeXiHjNF6vW9HQ0KPQyMZwi6x0vPirjW3em
dCbTI14mcHYz5uydS1gLBlkz36nwI7h4k41LNamnA6SvQ2whcbLhoiO9ALP3foNi
b2yzg1x9EfBYebkoTyAc0qsDsbdMKSBsyI7LvjCnn0kGyiRBzE3dd/GS3inrHkwR
9XvXk6VRp10z60Uyv0cdTw==
`protect END_PROTECTED
