`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kD8ltU5AnBMdPi1vIrZJ2ImIqzM/VJgp9VVCZoEPDvrxrv0yVTc2Gv8P/PeHr+tB
0P5lG8JisYEdMB7oTi1YxHGd0qwo4jNc+81orYNu8nnpJJVLISgtTKTncuG9lO+Z
Op2rutE9qe3sjnftvgc468Y9tdDFEROnXJDfmhUOdDelKeZLC/yU1tyPywryRgte
Nw+Fph8ibYIRLKjGPNZRJJwadNQt2a7KuPD6b4EX0zVFhPCnCZluVUzZ9l2Y3VLW
7yHbHfZd6it356telRhqmqJrmEV4+SSHEwBprqFiNc8LFaxG/natofPdYxagAdhB
Z8EpKFk/GtMJyspDEsX1d81suehFKzsaoIjyzGGJ1cJ4MulXOJ1F9Xqv160HxzFN
OuMFKLhvTJk2HL92KPtPxMHwQOEqnl/XYNzo9N/9HmtxQg5q4tfWhhhEsBCY0hZb
l1BYWUeIj0djGpvWxBumesVTwpDY0NvHVbTsbI5QT9DAd18ZVsRPTJYpAHw4AKnH
/DqXrE5a0OvdWI3nuIRvEFxnu2dRMXCk880UIc1tq/nGK5E3Lyfmsmm2ccwl4mkj
0JwY0MBMK7npzfzhCizlqOICkBD2qJaW8BCYxFp2uYmeiLoy/KDgRmkzj4Y06kCq
8GO6nM252/MJp8fV15hOF2pA7H2T8DdDuwFbjzkpYxq8Ni+oODIz4390g2XD3He2
kMUdQh7EcnOE3l/rfbo2QTjQUfQw4JIirZ9894VKc3dzVoKBpw8s2GL6tAfdvbxb
TIFftIZqorzfYTdVviW0cCdIcCgot1zeVKFV+n+bq61V8DPA2+iktAi5tQ00YAos
y/IV/nK60qK0YY7lZrHWGsL4SNpzaYPpoCVA/em5QwNpjiNL68D8++3Rp02AOtAi
N6ujBCrv0q4Zjqc4T5HdX6UTOO9Qy3Mxf+68dZDx9f5+9HsHfOuqj+ZLEpamZQTX
m9iK401zOCb9LcetkUTCH59GPV/ccTaiz4jpYCYPdMSsl8ESA3IidT9dYg94e3/D
V68Y5j/HbDDZpcr2pSFaJIMBV8p+AO0bUoJgp2D23aZCqXVbOiR7HE63rREkQJ10
vjJqwReQNAC14N4/J6v4s04uYhp4deVs0zsB/5qu0m3i97bppnKnPpQL0AJ9lxEj
sge76HtsMQU5K6vhob0eelZexMim8XN0lNnJHbc8KW4YJsLtdJ3uq6LiJAvIVEza
OEG97GBGTz72FoTIyyHNbCq+rzNNFfjJNn4GjxW+LVNpwkn8gHSC2nkRqJKV+EHp
Fko8BsnGp7ioL806tWtH5DaMW8Ee7zg8LhfqG4vVpPj+3eYqnSm3boekO71VU6pZ
7l/aEaVMFtghmtI/4vONPi/Wt302rwlUQb69S6nIeo2+1x51tEgcK89kT8VQW5kZ
GJ7l1P7riPoq9Ccr5Ej/7RqCaGIFtFhZqzO9za6vk6kSSiDT4v/MGJ1dzdz8JN97
2qefa8c4oz9elo28Pt2Xemmluq2A9qxAhHFlAoV9QRNmBYrBrnLuzAswssHkKC2r
iqe9a2E1zY47Zb/VqONy6eeDbp0vimmtIk8+wrS6SvyRq8G8opYJomNIpH5hu54y
jwK2VkV7ToJ4A1EqTyL2EE+tO88PnpPpW6OGyoCDTPKDM/9NmGE9e1eglOIivvI7
BcnAzeeHcVVlOg41OYZ7QZll4+7+Vld1YYWTH3BKTRtWBsNHb2gYykYfT4rb/Xvv
V6xgShjct7EOUFp2atSYG3lzqg/IPfIxNMx42xmlZi6HsQGRl52A0rea1Jyh2XWy
lizGIWG4Xr8qRlnW5xkD9z2J5oyeA45QGJYHTpS+ywtb/UmBN5x6/JFPJglVE+aZ
zYOleV9GK1sW4ReOOe7X3HaIFGOUBWErmUyIhWanvZHFFVFGzzgSXucW4FKiud3R
Pff5BfHTB7+YyUvKuZhjHbuemxzNKAvyN436I8IP6rB4m+3NI3gXZfvhZHN8zpyM
/mTP8N/ys+7Js9BS5JteYwTHA/i3QvCbHU5NzRRSjQdNv3Z3RWh18HGO16b/HWiq
CdVErUXd+5OFi8tElSPtVc/arGLT6B1owkBgX0jUiQu5175Rzg6Ideke1pwwncVN
mnCtU9uXr1ZWElnuZrkldlWDnL+xL+QvJSajkWOhk3PlNeG4KLWOHjw2EU/7YyBR
suZAYLK/d+kVReHWi3QthIMWujm2LsXaWBexWVzNESxRfkoZmjguvzJIa4YSw4VB
RexPe/jpGv05AE8AWXY5Sj+6z+Koy0Bv6aBn2CuEyWch1xEB61WLNXXPq1Wby1DI
2vVZshDPTjSJWlkjMEANqB42RyMUrGAjFLRWuOIVW/MJXep5/BmmOh9Hkjw7VhVn
qZJxfHCMhLkJk0BZFWdJxMTHAPN7bDyC5zl8+rsOgaUYotdPJfd0oTsA2YkDEBOI
1zFRROjFI4ADBm+0ql6z/ZYrQ10v8WK3NAabFhGinJmjx+zE8wb2mJK8geMJTFyY
zI/vCVcXRKoTj7iPQkuYHzwji7vga9a4hN6JJOQVKTTJL6qpN9udCAZ9ESy3+VSF
oDOkd8zEKhXQs09iKvlya+Kfq9cuY7zWgmmL57kY+ucT4XQ9zyNpHrBqNILmlh5z
LssHcy2ywwTFle7wMT6tGm/X36rqhaVoyDWBnJV9+Hvfuw3RevVc5xJRRJiSw707
N/bOknS41dkIvPmVwN3bE6WJoLg01WdMIc5D/GgAUdXU9MNZqTIxVV6qHkbOZZUg
LCfJyC48BTnS44Lu2vYv0lI/pCgodfQqpkRowg420VehehHQfwWhilOQygdJgfd0
lB31X1lxhzpjTyrziG79KkyzQn/az0gh1DJM+VDWxlFEdUuv1g3cS7pWJmjMNGww
iL9ok12YCo8N7/1CqevEp6E5rzVH/Ea7yJLszu32kKrn7UKUvf1Oy06gcRcABXV2
Tco5tRmDCkBjswgXYPk2vCBv54uXHqT2oV2UaBHL/2qA+G9MpOjuAnEyJTNryHXp
ARcENhVi2sqw2M3ehoZEdPABLiI4shR8suRs/6Xpc3C8S4/AXsC+n4WuVNr9Y8hX
Aw6wpuXZCloPNS+P2QF2/ESHCHE7VVdDvlAkGz2rRpd8cfvqmqlLf1y05BUVz0AG
iQmrsuaxm3bbOYg36MLVqgqGHDSI0lrjyz/2IZgYUQAyDjsv47h3vmraHBHEGrsY
Tj2gQ/kMrafpTrrAncasb+v2VQBtBzz1hmQ28gVEE8bGlCv6gVbLcD+Gw7CzF7S0
8+GsCo+sWROEP5ckEDtxM9TB/nXII8hR1fGWPWqaoUDpwevPYtZvYdX4K2esXuMa
azdz0SYBNsgK1pVWwoAaPM8Q4tlKmg/CLAA+LGd4fzwwwXfy9pCfPP8GDOTcCdtC
6++6KmBZn07EXzh4KJ8dD5CRj2e05DcrawPV3pQ/JDsyr4x4bnW9QeLGz0igJwgU
k5RxSjlWbbyeTcwHyNaf1qv+QctDmhdsHteZP+ggyVSAvST8Mj5JF8E7a1tquV1r
G6j7QLbGStG+35HvDbe12RCIf/SKVOOmkOG8DEcQOgR6DExRRgMM5NfAb1qcaraF
9ep6B+F43yAGKIBW/NiBqHW21ntlnKxFWTVtnjSWbaxe8Qwdyk7nat9wBwPOL1Rx
VzGFwMcJAOG3mjYVkS/BA4DCoc2uEu+lL7F4THGO3SO0gwrgVqbnSch4q+8EUi0q
MSz+PHuXAgbJ6IU4Mk0A6UehyVfyxmhXVrJAiTf9MXSUHF1C4s+i7uif91FSVwdH
2CY9fQWX0ffborBNQF5i6WDBYURQ0rfLDe+bXY9RgO4d0EdoDeK4CMJF/jF4lXsu
+J48AGAF/zDAP9rX++3UHo/RnpRmlOQL9epTnJQ60cPSfIEZhnKfOskMngIHaJ5n
3nTelgrWRkVC5eiPZBjdgMUreuF2X3AtdVmrUw/NHg5dyeRzghSJQC0mzYGk/Rgb
/Rcl6Wt+HawePZwa1iO1xqegZ/1DajUSlPp/qW845x7Q4jRC7wOn3Ot/4hoQzrW1
JcFPD2/lkA24TUY7pgSgGFdxpp7EX0L91u5tCWKIxrTXEZ5rDZABLTJ6iM7kp+bg
jKQDAZoLVRFAw9X92vYvWINfr2hlEpAst6OQtAKeoLyrrSjkpVkCuuibxYG5u7gO
`protect END_PROTECTED
