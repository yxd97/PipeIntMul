library verilog;
use verilog.vl_types.all;
entity MULT18X18S is
    port(
        P               : out    vl_logic_vector(35 downto 0);
        A               : in     vl_logic_vector(17 downto 0);
        B               : in     vl_logic_vector(17 downto 0);
        C               : in     vl_logic;
        CE              : in     vl_logic;
        R               : in     vl_logic
    );
end MULT18X18S;
