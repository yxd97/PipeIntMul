`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aqer9gQVDd4C19PKtgZ8ldz1+X8S3Z1pcXeDiqpTz/ffcndaV5QSS++mmHDdqk61
1prtDsviHP+uAPu26n9uETVxyOUEgV09Yq68ZZuW8f82xyRzpr4ClyGm4+j1WjI0
U/ZUSYppPXpJUgTiL9vQ3bT0W12Xq2ovbS5qf0Pub6k0+wNYiCI1Cni4XNXA7gAS
uugckVN59xr63CCRHygdJtG6T4hwIUmoRfWEh5rG7ZJWRnzuClsYHZucs35R9+z+
Bv2tPer27k3wLQNRNipv5+mfKzyPgxTqKFVOLndu5no=
`protect END_PROTECTED
