`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nHP6B9tvmMynumbNU+bRi0nDpArfzjLsZD4x5B/vU4CT89EqH0rEpqACtsHYBafc
lqNJZlSm0ZN0szvhQZocRGoHXYeN32ORq9+dqING5IxCKhwvSlmcguEMR+ZMmoAd
zQHCFdqu7gnr7uqiNEDeQlRRukeECpkKqbP8T3Ym1vJ6mykR6jd7oOsFhbhicIWT
oCFtD8KIzX2wI0NGzCI0X/dR+HLLCDceCKoGWaQajvpRC2khQPGYRH55PvqkXg3R
JTKmVf6CaYDePHC0o8rmQgguC82U+4T+pnZt9klWQuxacI7WdbA1CjOPhaCuZWPX
aER5DqFSjTPvS8XsuyV9PAdz153m/2yGy6sNdUAtvRIYeKdRnsNnf0I/ZBxzq1mT
HpbrqQWt/5K4wRVta6wmMiELfWv1gXyBgbbRh0H/E9WNetcGHLx3R5i2FIbDXjtL
Ql7bhmwNv6HalReOpVqQkaz3gDBz0WU+Qss36xDfW6/4M6gZ+kRH48Wv1/p83Tnh
bmbZxtjROG4sbW41Y+YEog679qXNII0Var6+nVdsDxyTQf5MfFoOcek3bnbyV4iW
RrE2AL0Ss9fBsRS8LjS7F6novIkUKgJoQVhKA3Hj02PwYoyLhNZZ+n7/FjkijMSg
`protect END_PROTECTED
