`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HuTN204BgZJ9hCZRt2FfekMsbTxALvHhzFQOk3tuDvB0FaNWcQ+6U/LCayPVjsf1
LPdyYdXsyvY7azl98fjAza3ojenMSdzmEa02ByR4Cj5ynfawnyWYSPSI3+RSqyaG
ugBmB0M7XRSdf4OSQizSrv416n2Quv+DYqlIa3TmQt5dWvoap1bfitG8Nvz6lwd5
nL0JaO0l/deApVFJjWAI91bVgdKPlTWVL9Sug2iVRd6AistBXX2MmWdghMjWXAjI
xbegxBGR9BDpgDt1vYMq50e7guxUSK8e80LroAERvqe9dojnaIsVvTNT/pb91r5o
v+o70qvcjSpm7x1bDu9mrEGaCjkdUjZJCs5LNXWsVYoc5r0Gi+XC5iPH92S/I/on
spGul+P2pHF/1+mO1D6BYXD7xU0QXQtdkX+1RVKct1UAl9vuHYdNQGYcoysPwM0F
`protect END_PROTECTED
