`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BWPPcQq7Cxyfr1Kyh12FLqHXGhxC/VN2vRvWz5gPGK0pZl9ie0esHp6jtEYZv1IR
ZuJraHuy6eYa2e6pan2YdGoYfRgNLg9HHNFMbzb41O4LyuMdEfK1ZtZStNVHW0Cg
capig+imCvC4eaYucU4Ad5X09CF1/vcZy9C3R/t4z0iWL2bfEEsEgFr6dMXCY18b
450s68g48wBAnL9+3kykPHj2EfcpNtl0SaHM+2se7i+uHdRB5zI/TbqHlZhG135/
DsvviBNcb+EpyA3TEzTF295rS11QOsE01brbPOGGBACdOm12g5oAPVyI/WX/lRUg
zmmq5qRMdNjQAjLY9gCZcJ/XZrKdDGxbmzOx0whErj03KR5x2iwPK2p+mZvSZdhF
eGzMTn846hLAJng+/OgzIomns2lZhrsAiDD+BiFyThQBfHLxJ/EbEvEmYtrJSg/F
e2XL8dMXyvopZwJTtmEgXHS03X78rlw/gL1dsJxHcTO3Np5hodWDN36VW8/o/Mvh
D57velXqqLpJ7esRSHJpJ7OpMlpoZQEOYIT6oLYE6iOVzt70VQQROisQ0ELQgCeR
B3+Q6CTRtd+XW7Up8E8D5gTj3Mnh+kr5cYXGdzR4ByzMqXK1i2nJd3TrQ8jj5lIl
Z9dxJ48vEiWzN1DScu/JSVXm7LLJVwzEwAOMNFSlRwJoHJCv9Kt6bWUR89CQ4p4+
ERQZ8XLGzPKbrISZOPAe95akdzeWaUv9Y9Xx2Pt70dUAMy+xG6bZqJ7dffvgALNV
yih2EYzzrv1dKcql0RFhGD63oOxGtafrM2SLtp68uDVK11AD5gw870LVBD6+rSVN
P8WdUU2gOKDNSh0fZjChhP3mS9GOkSTspTR1HBOg/FZfOiVqAmWvo2aHksdMd7Wa
72sw9MLWROm6KZVc5DWP5/9HTmbLYtCHPQ5Q9djKBOURi+HTzEweKYf2XYVeMfBd
qd8nix65vnpAQNoPf1eQGcmcpGtjpogEXrcfhdwJ3W0FAoKHeiMg90EbVEmft1PF
a2H42cBhAbzU/tHJ8VlvylNnEtMLGsoQYtxAD1TxiYVT5nNT4ux0YwkSGG1dpWgf
FP4DHQz/99h7ipBchuKkVMVKQY20Ah3BLd98jcRTe/biYETNf2z5tSN1ePjgk/Lh
mQS2/n0TRs+dYg7jL+sWJ2U8oa31nyrlowOIHTxNOG7AjEWs75zBpvOVrgIihczQ
eF3GTwZCcS6kIHFJVRLREY778+B5Tre4zgETn6NsOEzlHpHCBQalz9lY77KLXBem
Nt70XRM0nj9GlDnsPVBrM+NFTB+nMr60absrkOJVDy5ZZoQ3HDFhEAHSNFzmILUX
B5OdP4Zhg3SYGzrtCi0CYM4awd2pRufKQU3040OmeblejPHHfDwSUYSPSfV+tkZT
u+tLeKrdjotnFyVlOsXh+bxO01O9KhWAnMDtA5Cyc3N32Hnd/7iRB/HmSHl7UpOs
NpOpx/v7Yy5B/M12iyc8xxEKqGLcF62FQQBcUeeM4VNULpUbK8YdEhKG9uZUL0Xa
jlJrzXqRH0Ne1y7ACe3gZQ==
`protect END_PROTECTED
