`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQ07yZHOGy6An8NA/LmLr81UDgXxZqL+s7pnTtLdhihQVrRVJv4pJADzh80vc4nO
XChj9EjqCoXQOW5cudXL7k3d8ARuVWQMNFXf1WF/8uIFDE2aKkFh67gyJbRYebVS
GhyByMn9Vfd4FY7hJWYIaH34QKXjBS+sdyZKRQSHNatqGBlTGvPHmhfsV84rcssa
08EEjm6gtmK8BzWVgyJBhV34py5Mz6rkfbvmg+134trpyT0vhnLEwvVvNKkE2Otq
U2yFrJl0p2T2IpPd0qEdjr1ZPiq8qod7erO2QCJmTN/V6WOoMvhB0R4e0KRBquci
m97b2TyfdVde1f0xj0rIaaJz3T24qWCggvHj1xEAOvkFClRz/niLkZ7KpckPTG+B
owUicqF3JEKweKMkHSAPG+jrX6sIqm4shGKYIcgCKLI=
`protect END_PROTECTED
