`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bi/oaaGnXGwyV19MlkBhfg5q+MQv3SYduQBolt1hXXzwDQ+4AhwiXMLjRSEppw9o
bW+Hk9tW/GpFoJtYThGpjORHQJ9IAWOfefozzLETIUvMtcOOi/5CY0Gt1DwxvluE
YRcj896oNM2TZAX8FDPoRtUDJneidTfG+GwaU9VKoBMSSiVH1kRvJDrsFEoxYGuk
E1E1+/mZ4it1rLw+sSk4rd0T46TeG4HSsv62D8y0J6GO1zlktERsrfSsxx2rFGht
NUjXzBVLkjkmXyZ3h4j3zrG0cm0sjcVeiqrwBJBUz65bmiykJHY4+mm50F82Uhb6
mUjF8Jf3d6BN/X7r6o5BqyHsnjzi4NAUutzjenmDcbRRLODiMbz+U+T82xApACBT
hMO8JIit40chj0ZnGGEorQ==
`protect END_PROTECTED
