`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fto21HvWjqGE2IDYBBKnjMyMC5Rs2WUzUhKVA+36ip4hDRG0cRhb2xo0Qo1lDEHo
2bCAeGGR7XaGzb4CYGGUVgB26vLD1vkGIOuLp9eOapixDWF15YmGAHsRrgAWyhiL
IDDmPRLpgPN1uFPrT8OhSz4aqsMSSje/+rej2n4g4e4wZL118xiPN2oW/0r3sPui
TBy54qx9up2Yay7h2ra/MqpXhOZzP56KSQ+XJgKmMdoBDjDsEnqPMGv6CJXPlROX
zC0yK5Xt3He88+VRpVWIqtV/ydH9yWcfqSVMeHRKZsOmC4NgYTGvyDtXHoTZN9dO
nKSD/+JTCs5RLL26HUChxi6Fw4K7uhDRf6Ch4Z2LBUCtZRAWfsRQcv2GRsKnEWpW
SPDaHS4fAIJfYEcTZawnCfokJmE14ecPYZRBncMflHk=
`protect END_PROTECTED
