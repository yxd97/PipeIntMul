`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t9sTcxS8jGhhaGBI8eRXL4FdJ2NrpJhuKXbdzpXy88bKw/39LMOUOLdTyWcs/6pQ
brhhnXVcPAtbXuMCWU9IUwwLUi2LFy1WUw5S1IAl0h+cmDHuP5HcJo8esfvKdiyd
mW8qRW7IPT7g8pRO1IwpCA6W0+D2lANZ7BoGAvH9O/xwrEdEQVjoWgzvSzPQoep8
z+EHFJnt0sdae9c51odKA858meQV/koolzdCD84b38R7nf9hcFrQDSiybHLi2c+i
W4WNfYwm26JRD94D+dinIIQ5xIlbQ99+cfdmhEBgV/J5wjbmxNvM2nwFih5hcacZ
MhOIT2qnGq+gHNjEXcco8gcJKVwiMjhlQrsx66Y5c4UyaugB79SLBnId2pkLo5Nu
rfnYTC4TcxkDZF7AD38iv1dd0f56pXFaiY8tf2twUbmrN/qaiBygCC1f0YUxKk46
`protect END_PROTECTED
