`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6dW43dFZB8THEyP8Y1j3Ig7hcyOlzX65cGmIHfU/W7b4fx7cpDKPsMfQta0fvE/8
FhPbcXBsE+c3HbKODoc6HWMmLe9hCHiOPmUy+0yr9jAhRb2rzk65A4qFxB8y17WU
yo5mf+a0ExPt/D/+yrZgboUXvNa40BYti+ogHnvEUeoxFY9Sm9oY8wjXBaw75+LF
/j8UdgUXA1EPUIxb5D7IXlSbt7KT3tg0FWyyUA/3YwR+2CBCd5m2xs/WsH0DXuqk
yJ67Wrab/XtjWyVs67YJwb0o5GCOMil3Ofq+tS9FHRjaxPMbIVvbPrYmQo7jtKdr
IYDr0HW0lYVZCPq6gtvaFPj7Qtr3WTFp6/izQQwy7RePcfBvJ/inRdJrKggf8d3C
AWXPh7Uw97BP2BMzUg7dZsON3Futo1C5OCagNGgYfHoTguqtxGH317L6tO64hrY7
eLSrQE+tHqyG5s68zCB/K3iOWu3MIWiZ0d2QxzVGmEiMekX/c6+m0xNQOvbjjWJY
WxBplMbvtT08wrPy9tntItkJGlrD4Dn/tShkjvekPhPUEiogaxH0jgjb638wwRV3
eY1SuxRKZGoYHiBAtQc7IA==
`protect END_PROTECTED
