`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8evVscDc+wxe/LW9U2RsT2L/ULja5wkaaFbkkPyHZif8O5uhGhUeQ9VWcL2aBvYV
URQEpQy/P5x18h89KJuwwPoS1gQ3Uu7St41dHYMHEUq3tp5wANJ1QOP7IizG7wLa
+RUo6bZwcRs73vCEuNkYceJbbXEyxFTSehw31OyJT1K84wVowVsnXV+7fAXX73Hq
TntFUHNoGkrSy4ihwHvlLLzgFrFuNUD+FFKzPlROhRP2ZGtbt6Y2xBOV+0RmR5wD
2j21Q9jbKV3jSb1Fi6TaGVv/78eyedIoSe1GAcgCih88wkD5x+VxBLbYltIDCXNJ
8VhZONJ5dwhecVNsdBr+lNm/3Fba4+kXz1QkH742mfooqFFT6TW/Cz2TLmLQ8dyq
qmYAXQYKhtUNwEqiV0a+XwwTpVHzd0tsci+stZCYad9TNJiUbvlBsVOvuUn1w4ug
E2dQzEnuHtSFcf3qeHYfYXjuYv29OJ2JU0vb3Q0Hrz1mGJ35OfUEvp1Xxu935JjM
GLY/YtIoXrOY4scnesV4i8xQRtrZF2lyK8+fB1msGMUFdO9L89wjL6RoN3AzI9Xn
T+G4NU0alZL8r6w8EbE9jJzr5QF5WizxTR5VJED+gEBv5N88ua6rFSj34PjBkbR+
GDnFXC/HReFtqd2Ftq6rBA==
`protect END_PROTECTED
