`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOH9cbk52zU58eAP3vpqaRTVckDQEE9SffOhJDWJzFLDQ/Jc0mjPnWEeCQaSprJr
vNThWhvM4s9gTeDFB14DcDPVMh55ouTXOAFPrg+yOjnwBmbJLuwT1fxm+610ic6A
wsvacggn9ufzV+m93SKj6kMSTD9xvSvMmIPYEMubdwr8Bo+1joItBqrDNABtYemG
2XrAW9UT2FNoQd9kaH9yxjtJkA/+JJ1h4nfAxfKuiuoSAUWJtZqHTgXDBaO49Yc1
UQ1UCX74y7zq5lYEhoLRrCv1B8IlbH+GFM01Jxh2qsZhc3z5SQRXOtJQydoaCV6U
hO6qwkMLbe1EpPst1G1Ed51uOJXUADha873GUjggi5ZSCn4A5ekVFpKj6ESiyBKZ
K33DIwfUrKdBMIIYYn4yO92bULz4ciL3Ktz6KhsgFXKcQlLgoXpW/W1c4IzmUa6y
`protect END_PROTECTED
