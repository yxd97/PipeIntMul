`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcKQrRL50SaUeVPqk8u8L0KYhrUqtYT9SUnKMPk0weZrP58vIbNIISYiQlcBQz/d
TSM7yk1N6LgRLPaz5JS64O3KDgcEQT5k6wEdVcgjiranxs+BVmEvt/o9rgbxqu+7
7ZNLx3VIQb6kQMR/EDtJp0XY9IBFB+HyUfqyWAeMSIeMvFvq4vmYSRMB+FjKRT4e
7A7FKo+e+PKJ2Ky/z2oxk6n1kJhHsLQyh0x4eWllyrCqPXCAFkaGy9QTFLYW/W0F
fWy5jbIJBmJGNkzOsJjaPB04rEfLsK3D9Vz+dhAHxYudkiKJ+50DfZJmvlVHmWx3
DaCP/rMedBkyQQcwyFWKLu5qV6TBdeQXw4T07O8hsb3MWzUf4tIoz5h+bOlTF0dw
VpE2Kj9ulxE4cynHWloXlNKy3sXcg7mF20IFd2gm0ZaLhMbfuWRXYv0qRdoIQkx/
WYWAVs0xByS/jl4DgEAwqfxsJsuj5Y2hLQbO3VgKF/aTEfu0ClgIfUKpLGpIZ+so
`protect END_PROTECTED
