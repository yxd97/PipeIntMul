`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGFaY5WZnm8JMubT0QE4kZeDOAiEoBXPwkpGHtDxgGjyHjUqj0MA2MtimUcDITvv
dP0YebPK0OYH/NMHnWFZg3s7IYQAPOaTiNvmYQK6aCOCB8piRSCk80FQHg25GD6I
nFHJHTQiiJXk+iUFiNWwN/aIKI69J9Eo5U7ahZdZLa7k7kaF6pGTc/+faYp267vp
NwQD3mxNRoNcA4PCcH30QhfYp6bEtaOBuKDGF4mWHZYpdfNP+H1mG3jX2Ix8qRf1
Lnp+R5WXoiv8G8DtNh6zamkY3kX02osi2MdiwSToPF+RWXbwILDFWUR94AAkTIjW
Gg0DFIVLUSz7d+9znE2Grs9WHKAobwXTzf1vVhTdCXOZWMO6YTRN2Q93OFVYl3Cy
WYJaYu3GvrANu9QwQkthQN1DOSuh92oz4wOnkjH5VC3pkJInGEFDAE4tHZVWgrwr
4wHjo602t8G/E90cFAEC1YT7sEenyXU2O2AtIPeExVwH9yFJjX04kcpXavKwpnVw
0Zc7gOtz8JmMCmB44aKn0z8AV0+HLq5NoJv4bkoGjIODS1uK6061FUYBlwFulShT
xCPWTUr8jN+vCNeJP7vG93F7h1lydO+9ve61tojfMZq1+BQvk8Y8vQEIbRQRHyIU
nNTDNeHHqZpp+pjSYOTULsdW2jCllR5UnLGBhyFFI459AwzEo+GvEqGP1c0jpf4p
PaoIo5j/Wt7kT9MhIy7a6gL8qqA0CMe4rODB6LnLlN3fD+tENZ1cP4RJcRGk0nTa
QmApQhwQOZagTAZhmod//w1NyIoAq6hTiVgVPrWAZKMDYlQe2JbQFtBk0Zm9qtni
amdqPWlQOG+vQY5aYrplSGICMRRUOdT2reW0KUoAczyQgw0NzgIwRj/wXaQ70SjR
sXVCLhVclr0WHwtQeytQLZLz3ZttlWFfbXCqGulxDuIcMQCMfqwasUd5CXH9iAuQ
`protect END_PROTECTED
