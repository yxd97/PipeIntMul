`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Lw50pYjHbTp/GBtxqtKQZ6nhGEBgrn0zfdpKAedxeApJn82T72wh7uq6veX5T0f
+PHsdzPDZJciiE4ChL60EP2BOQHx/WAyvDnm7QAR/7KiGaSGS5eq6z0+R0Lql6gW
7rcpvQJaGwF+RkV9zPyDpHQUXHiExuK82kCqV+KdzPH+O2Dt9TYxYseeF1s7lr/d
j9ZwWKEE3LQi0xiMYYV2z5P5tyma1623TzfPNM5l2SYkEdT/IIldqkSuTsSJqC+b
VPKx7Zt9OUXKPEIRAgiUEgcvt5LgtVuBlGIi2ToN8jMoU4VbFozq0Huib1T815Wt
h+vU3XjmxLk6qWk8dMnwpyGdEEQic7/oLjCqf9AGFury1jaZBRmEAb094W604jZK
WyjNKWj73j8kkNA0bIASvUwji7lNS5YYVWcpqP/Bo4ho3hrazZ6tTHGxEF6dgc6O
zUSIPbZVyCrQDUIG8cZJrGrwqHeNpALk/G5AzkqmqDUU3e44UhqCayZi5r9NNd1g
XVLPToRwsVg2RT14AFn/TUBEDjlsa31K3GiZrvlEaYe9mcMneOhBhnP6EO/oC8CS
18jG4ukU9Z8KprN84eSlfRAU6D5hjJeQPBra4zeATHI8WW8xh0pjsYKZAotMxpYq
g0pGvX5hRJd26XTIvH0B4uFoX0K6RDyS25xMIM+iXm+p4c/Xxs3zwrqIc/sYxrX0
Vu5tajsMxAlq8qu6yciBKUwa5gaP5EhyE9wkcyfOZzxnwEpl1fmL0hcdyaJsPJxy
MzxsYxF5GQntCpdc/POeqGIhdcDwcNFmF+iJgI7oHQKRpI1GzKgj5efD/a02CvHk
QOFBtwvmy0+Fdvdkp5g1Xu+j5f7C+TfDsaXx554rOC+h2+5kafWd9KZuAEaaZM3T
VDRyluHfgtRgyxOCp+4xMHXTiyGRUeOLAxqyFx3Lr2Lf6KuWmiP3QJr8yAlz+W7a
NOegtwga4O9fs+sAAmZ31gaaPZyqCcb3b7u7NUbS9nXGN9C8Gl7hWgk+wEOuMXlK
I6I0r2/ItYdZiKcJy/uTJYx8dSoacUneQUWVidOqhiEHpYoAwue0bp1njbYMcS7y
Ap2wRZq7Mj86w0yq3I3ITQtTCwMGXxWbhJm+sTKQKS26gWNJF4UktSEjLQvVPLXQ
TPhuFNajV7L5qWDE2AFTjo44MfXA2JmjA8MQjO5mP+gwNF3rz1GaqfYGR4H8fbyg
hUBFno/JosPKYCxFD1BmxKNpO8Mcb7d2C2IoXmN0EwRCPRyZXJwgLTI9D+X8wWcF
Ah+ztNNWc2yKDzGvTyL+TFKKs9ZxFgxTb8KO5S2KFqA3mbap4q0p7CFln9bz2ZbU
MlcQN6K3h4OLsXdp2GpkFaHnuVUffRy2RsZdYx9lJ/aJsHxGkYM91jjcQVcGs+Ww
OrfW6ln3lnJtAgtcMU7gc9LaCyEhXf80aVQKZj2QpWkL8ad5EuAC91vtotguVB8l
n0Vlbcx8QsY41yQazaDQrEzkK0XjKDQExSB4zD9Oauk2WmXkkYzlnP17vAbhCYMU
5AOfPczAtPDcSQxJ4zjxVRQJo1Z67eyTzzXgjkReAptTGL9K755vnO8ItwlaNbgm
dezIB8RD0N8EOlp0t/aYhRPSFFtvGKb+xd40D8ZUwhQWh5zy61+6m8cAkoPosn/l
`protect END_PROTECTED
