`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+maVQS+XebXB6fiXH87j/2d2yQ9V06QhHiHOdtyjTLTCTTBSwRRoYULf7dsu3fkf
W6NelDx1L0mm0AN4uawaWCC9o7Kc3juFzO+TuQaDQzeV4CPjiRFTtq6hMj2xNqQ/
pCLqPnUsCvNlXp4XA6VE4XZAqUOZlfNQrcHAdW8h8/CJpd9PGuRk64xyfG+Mj/+a
/3zoq8In+nSovKuJvvRKdIyaKfiHwgBIsKTNXFywI6/VTb+0sN3B6tVXjlqQAUHx
bY43AmcudfmCX3Hu1JnhKV0BhCN+aTgFhlnzk75dqCQ2lNKyFBCOOaA+ICZzgnNJ
k1q1ybKt7s0miBLKEdnZ2xng2m/Hc6ZViEGU1zOtqownCPizPG7LK4IXsGAG5JlS
p21B8nij5FzyPlnzxjCSK2Vyq3qA+f3FbkBRt2mL4JoceEwB9kPzPF4hW1Q5tT3I
SleJ1FWgiz3UGpNsbSWHasABwC+9EW7JdRm8Rc37VUMWTJGoYjvxE2xSJps5IG4A
jYvQvLS/HFH/FaJuhsAK2Cd5ztFcsO5nqCPQ/RBZXyvz5S315Xv7s9D2F+KGeZGm
`protect END_PROTECTED
