`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZfqSN1ekpqrpx852Jdd8ZVeeuq7WH2rxVXp3XNZvncYLu7YMfO5ZqOZLFHKsGkv
HrXGv3mMi6PaCL3+oOcPHUbUlkQ9mIskh7m+gjqPpjmfplaQpG4HSvv24+H3QjSe
AhfS8A4uSVhtRD+tvCm4bQERjWCu/QPbALVz/Coe0vWq6PeyXpVwVSKlMYjGzWDE
jNnL5yJ9kV607WmMpqoLj4SL0/DHUFaI4wBk6yYLCegdNNhUAQtmVTKvPL/eoqfZ
eFljwOToAS4h4avflu7OAK64b2zu86akPMt7JhicagNxLcAwQXEMT4GThpQPgQrj
dF5d5KcBIGaVi2gjCCK2MKfHIePW5zBQtnLQSAfgKBodNew1osbjU2TjcTAswrNL
HtgQ3lutWENm2lXZll5RUHMuwJgUJbnixffM2/Zz144=
`protect END_PROTECTED
