`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XPo9BLK0LDUu+DOODkChajeOH5qkWxYsyDLYLJPfrc8A7WRrIQ5vwphQNbmvIwU2
9Xmvyke2XbYIJFm+YsV8mAZVJh23SuBzM8nNC+UQ/EFDsI1hRA4bKG5TMe+m6xic
TP2qcRhQTKowJ/1W409lpUt4nzJ4xpf72hfji8dg2+vvlAcwtaNp82fuGCP0++UG
uvK+8QiEsGLmmoLYtD57qoi/bzMNQenY0Y/+XlSghPEZUCCSFNrHL4R6UtYOdyUn
m2etSnlVNtJVUX7UTKKFjupLJBlO78dWqPZJndjTr8twwpFS4aQhT1fNbEcKfGml
QMK7kdi/5gG7qQpRossRMdFyB5QOSfDjGee+65ANtfQgc6AafeFu5o3Xv4J3RbZW
9ewXzcbaC8pLxL10NVsqn0vevfQTLjUCwM9BF4X3qar8kCGmZEsRiINtBQxnIUIt
NvG7ZgCnBQMCLWMSpmmPUFXXktLV6D+UktmZWGVOvzkh/4BnGap0B3iIAs+a/vLQ
`protect END_PROTECTED
