`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vuOAfgzpxqgLIgVrPhRXeDK9+Eky6iZYnFe6PjITWJf3mroz3Wmgh7XvX/WfQ3bD
Oaap81/4gqtHuPvqCCaHTT3b0gImF15f3TMMphqO2/EPYqWvEtA5K765pgeM+Gmm
CEoE3URmmoAHH6eY4bkcSVgPb4UKfQACpZ46k+xql6KOCwPCllQntGyIN56kLj4E
gBc6xaF1B2dpaEjIjnvIdxP7kqDKkOiaKepy4Zt+F+8fZq0HGYwlzgezcshXfKcX
rjw6GaX1VNv+OQCHjaYWrDBcCgLFuuYdiiGe2B/+Y4NhpNLJAPbzHot57gSfg7X0
O7dlRHiTTuu6XtLe1DJgZ08tRG6eDdTLFbB1oNItgCzqtFTLe9jpKip4GoO00QQ1
tE3Nnsej2A6GnZ7h2O8dnz6BQiWOpP+YX6div4mLEU6UUpveNWFSkm4ZM55Gbfem
6AAXFGOD29qfKcoK99HrsfGNXgtohcav/gFWtj27QUY=
`protect END_PROTECTED
