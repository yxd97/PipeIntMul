`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1emx8gVG3TLNGqqVrO73qHP2o/Lzo3i/pYEHXC9af/ObhLnDhVcpbmlFxJtDoqf
zDHThOIF+lAII4ik8VsMDRA5NT/slgnnoNaiWZ9XmtFR66I0rAWzIWY3Be7wtGlx
34oI2yOfAfUUben1XMk3c8CD8C3lnsrbMvGZkHNyQOUPJPBzPHIUm2BlcJ0ULtYT
EZH6+Lrq21qLBOLq7c4a7YZ0fCoXSt+Xb0N/fsWIDUTgsRClctUoteEikBMTbUfk
OGfIMnDYigqaENCYAeD8c7dYjO/sVcB6o9fZTXm3lM6uOS7f6JZfr61INTz61Vdr
fMwHPAjqdJDekR8fASiSA/ajmvIYpIM0UBuTNJrQe+MVn2GYu+XkutdnQGedho/e
z738ejvHJocY5DI41PkX/GgHJ6JhZGWDnvaHGVPq17DSF+GgXuhV67DWk4e3UkDE
Ll2auORDTRhLPB/0Dydloj3UuW+bVBRU1ILxK1Kx95dvwFc7sgykwAPDaQJhMEVb
auk9pB3ntQrl1BrqwMOPPNxdXAqQeAcjKhHIYBmJIae73u/YUzuIGrB4h2yWs8xM
S4Ew9hJZvszGTx1jcfFqc1NoV7uNGe8T05h2v01GGYC/Hhc3weLs9s3K8olk+qro
0RpGrMRjYVmqYbZFVY6cl81qtVlGnyixu5UHWNKCs3u4mD0uEA8GR2ACTqDy4LBy
4PXsO/SAvvpmmqYHcSPQmw==
`protect END_PROTECTED
