`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oRA+VwB4WHfCKTLKbC9Aojyt67/apZDhVQCrANUfmXS4CzF7JKneQrG+V/vk7/sR
BxQybDmO8WbHFrHTX2aHladsYsIKbRjkoFRmKeSQbTqI1PgMT6qtAY9NHppzwBg5
UVdjY9dZCeXMtd6/0JVcZb4saRYURqEEsbYJ+05ZdaKLFburoNMqoTNDer6vLxJy
d7GezhPWM6dq0MOLlCzf330ycIx5whkPtzlIuWbr+7PmmkIFskfpnYoUwf9u0zAd
suwAeMGDdWGePJrxxH+S+cryLb2lGJfUEMehtybMZjXiOmBiTrn2Dm+bM3yn4MuM
eB9dkCc5f/KVGbGt8ksLZi7+/RGztZ/BpQl+dFIHUaPc6WQadbAyokRYsy+tWj3l
b2Fw3fUEPBHDK1l/3S2nSRIhZPCjXC2OyisZJZp47IkaDud4wpqZV9vVBiL+Q8ub
87cqMLWVB270BU55hf92ed4+TDI1JDxuGdXYxnVT52Y5mEbPlX2O0/dQbbefyYsZ
TAi1qCGquEIq0c75tA2BtBo0ZrwaS4HwoQn8nPHJcjJz3JdA/LpVb+/itgE3a4Rv
91qMNqYVERrnXnhb/vMpbE851v1EsFIkNrBs7MihW+ANyP2ibCwR+rnUR2zNejyO
E0OeXT49bCBUTKqz6kr0XFhb6PKL5bi9XUOW6o/YpO6DoAC1qqcGNV+lWb/QF+Oj
i7m0D+QJrnrSpamyxdshkq0W3wil0yyY/zpLd/75X4hOl+pkBp6CbEX7tlEjbdOx
kX4y8Tr7nsgl7K14lWDaybahXreyTQasE/W08/0Af6TELpwfW4+46jJTtlVDvwJ1
XdAdqZ4hmbZD2Wn6E/0XBBooFDfkOvRas69FLXdiqZJTz6fY6wgB9BFLzbP0hK4w
0hi9mXQT5o0aZ/+79PsM3HeNoy4GnNY6q5vSloMLF6ty4qey0XM7MGBD0ye669Kz
9aR0mwk2O+bs61LucyRJp7ZmIQJhF5BpXSlPAp9qDAZ8eADkXv/ZITMJc2LxE4Qd
8M229U1me+SayEDEHnQjxFDwfBhAT/3ghAnp4FXBolnJP6dTVxwUvthiGLzbZn+P
FPdgO4jVVWIrg2aTaOFjQZV6wA3OWrE+xAs95pL5dJCk8X9D6F5CWTOmXVXsL9xR
mTfbE5fgKK2t5f73KhQEjVFSHdyWBER2lwGSp9zZSpHxVza/MJXkyIH94sMDy9PM
ETqb7BE6oib5dwtnkf/qsebS8PnKKIet93HKqKHP0BsDKX5DlQMKJOuEdmSSeVj/
ReRGUerc7i2nJ8Ge0yxM1XGFbJpAo3ZN5aNeAZj3qotoZVypQA30PPN/wkw9aU9+
xKELaAArvnDnNR6/L8Fh8p9wUTzTJbQqYsZgEB3icwJNHVcFd4Vr+yBzPQKz8xJ1
cpauAaG50VBzPC6KlMZocsAuEhmwhNysQzgbTq1V1toZYKlO+Qh45c2jklYv8MYe
`protect END_PROTECTED
