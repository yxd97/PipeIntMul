`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZieU9JtgewzwQ1AW69DdHv+IB8MPL2AfpulvfkKTISsXXBFkt0pwZGHOqcEGpWU2
PgNHtKiGyZsywACVLfLwrN4vDVt/QSi7Vkr2/fT3e4+R5/2Bk/WPBG9fQPprk+kL
XBh3bPT7byrBBILG7ymqXbghbc/DAv0b7YOddrPWk4MCbsnQLG7ZfS/ao/YzJ2Tt
ufKZgUGKUh3MhHk9sO5WI+m8tP8D3VogrZaNTtVcQIZioqG01VhTY+afrs+B1YiN
b9RSO/Gdt2/EgJLg1oKRdnNOTYDjbhh8SM/ZM+cIusi95hf7EF48i+qSQkQ2yoMn
4LXAohEHvJm6XgcQPDzGSW+3K/0T+qZg+wk5KlrLt9XVe1PohMfwYzL71SLNynxG
zMkfXdJNH/1n2kBIsaKh+PE3FoahplCXjg8u4F14I8LZu36KLbA7qsg3/UyLL6S6
lgsFLoNgcDkZYcuXEjOFANGK0HJYALuZfCTT/AbYVtvydL5E68hVzklCElZtkMkP
L63qHgQs3MXiL2JoJaW842Lt4uRowiZoB/JMKu/z1qpsD48Ankd3B1tjOYuKNGjb
oT1dnwiYpnpc/WjZQwyCfq/JGKCiy/JRsRyDNnzWSzbzaX69PD2ut+3F/ELLiDm8
svPiFzKLaAnKgyIRyrOpuHYZzyEkdN7P9jtqyic+VwWmpjG+63R721AcMe/gxkVW
tqV8Ni+E4kURBaRm6y819cNM1m1UQJk9vUrXUHFR39P6wWGdPzDF6oQwJjw7E4Iu
6ElHU7vrePpchfJJIJA9Zy3mpSbvAjDksSQvzztHh1AXXpYsXCnLnJ42uaBSU0Jl
NNqfwK8DQC6X7oXXIXOIT/SCxwrsMDdGgH0MVJ/UvI+E2QT1WJQCx/sgNHXpp4mu
BNk9F9Mf/1VBr+Pi9XQ179RVXNZxIUPSDMbflFu+scIOjrI2yu8j9SiOvWtHJOaF
mMrIjlo5Ph8zoIF2VvOlPDnvxfTG3tP7aqTcaKL9j+z5g6G5G1flM3AEHr2t4jn9
KTZFHng4YCrv5yadnb+VwJZH/m1EM2HuF4JaqV5l7Wzj1CD8ew5zxbomluy7NDz1
dlqcRcRDkrAU45SlskdXesxtXcwft5ALczXjnbxul04pcWa5ue3+4rCM1iAYpzHY
1TOLLnX98QIHs+ohF3NbDv73/gj/WU2Qq+Oyqk8hEam8a5hvF6+X1JDmXOoOTU9X
F9zknBkrTs/xoz3/iWTZDJiD6AVFyujGW9qk1YzybcnT2XwrmZAinI2zri1CoiSa
IEGbkdbdHfrE9IdyNIUVLNr/zzFqg8CbbGq9KdNHh8o/r5QHj08VxAEW4hri3Lzv
Z1Op5bpHn6r8YjSWDk+GTTRtqY6UJHMthfg/VECgp1hf2mrIxmQ/rKyMse0heXDs
sTfW0OTZF/yWz1OMbojhA2/Kb2JWCODJCCJTsKZyw7zc69YGqSjvt6+MOmmmLFSk
eTKX8UdNYuAabG5TeaW3M2n6NBEK+HJERhTiCHdOhmztAWMdShRJyfawQtriWtkY
m9nQQF90elHH7jJ/U0KguFOJ/NXxA0XRb/aQEHJ7z36z8UsfetkZqoC0lzCw83rk
5DXNO8Q5GUb6Efb3GvcJpZ0U/wZ2i2UXf9p1eV3ri2TqWQ8e/XfZuINO/iY0BCj6
PIFZuqO4clwjd5qnH9/FJb9rjJCEYy0ewJzFleNKBGn4fE8DYsuCoO7dq1ARvA3D
yCFgMMXq9i1WHomJ7wqRPpMs263qJt95BhybYeOiFGzUwHCD5dwNsnJkiMiXv0c0
MdWPGLU91NhSEg1uAqvM/rXY96NtqAUhNv8GeB+xGtMqA4BrjUt2Z5o2vbSpDXFX
7jr3XHs1hIxqTCcZuj+uYiABjatmIxciDscUy7/T/ID42e6GXLUk3UW/qfFkiuBc
vZIufuPle2lg4FTzdWHEqeYdbJmrhxMYts9Mjk88b37uuzomNu1Djqvo2a2zwBAl
gvnSualHTTNvwPXoSCS+vrSky20jQx2rJ9SxGfpo0hZDkm6CsypuVbIpo99fh39D
0lXyDDkTWOSO9uAKyF4oLJ6rImvs+xc4NualdSDKaDMnkhvZpZ0X2h9YZYYM2TZs
2uEwC8jV6o/v4NnJ6gAHKr0Z8xxAXJjgrkZNrP7HBa56dubI/sAm8gYjtS8Z+t5N
AJhUIWZraeSoNyXOv3xF22Mb8DMxvigRnskvGbAoZX0jqAP8Ky3mL3jTQC2G1QTL
HW7QRISNxVBF+afOeUlibm1oQ+lrdI3cBUw83FBJ300oRG44oAwm1EPi8V+h+g3i
8RRJg2VK3TkupU+NPjx4bfLVyi2OAdHqZIwAb0Qkmo+DRIhpR62jpKXpMcdRZaKx
TSNgMQ5Q0L2eTBoSqslxMDFy7+YY0Cp7r2Qvwi2k30heefe8kfg2uvoH5V0X5wfF
e7iO6vszoQ3j+i6o8nIMNQz4MXmsoNrydIbKuwPRu7DIvBhNYZcxm8KcQAy7IwEB
2LGKMWYnjb56zNrUtLpQ9JeHrUhxTWfut+EYWMd6orcDfDjsR76b3ayvTRMxCe+g
KFjOz/jNuXqIKdpLHL6+ifxANk5G2rk1LKEqYaF52rCRTNfSKfMkr1NpRi0mwv8L
fIJzk2vodd1oXsMi2h1/NlRKd9Sjp1ODzdg4yMVx5kzMmFBkNIUcyliELNGyShiw
tCoqy9aCIe062bygC07BpHbKw+ULydwgQJ04W37j3JIFkol5Vk3g0GDJ5DR1l1a/
Wt64v6Bd+CNWt1MuLWvJHNRgRmVDjF0oMKKwPWOBA7DeoCU5EZlSY8eLZYqEKaQB
RP/wZ+zOlK4MCS/PY2rOpUPqTmGDYW5MuCz8rvWsJbFGODr8L3wbA8JseVKj5zn0
EpQKDjDV/SkJznqrRMTbIiKSr9t6C6ISq78V/TvAX0AXsd29D3b36NVCvuA1aNjf
8pMoMbXPPIhjeM3EtQrG/lsNQma9udk2A/m1ERl7dT+G0G/pNrv/G1/0uRtuSvFv
qvMFPsSMTb3faIVgd/NMY+UgnBngMQU/R4pZhY+APH3D4vFFVEkeO7J5hUd/7RbW
3jy+hlBHTpt+COtKHDHWJIYtMBNPOxEm0acVtqsFmiA1kQHEDmOy64J80y4KYyp5
edPqLMMEUNZXAm73qdi70LIuXZIoEiRYpw/pS26LP7NDQOnhafKfR7EZlaeaTIaL
65MOU7tPMwl36FOiiIzocDpmRMV0qCsdqaFLODjUs6fvFtTCC24oh0hg1nUnGVLo
r2ZLPb/Gh9xb9dxKDu9NwoU5C6EWoQiP91yU0/E1pYNOuWoaygYsS1bpfhYmeJPL
RDtNJ1KS5QqcZ73IeSUhCdzOvRa+R89XAwMLNQ+0h2p+VwJYL+UIAxl+QEiy3sdH
aGNKYKLGPUMZ/FJSNyJi+OdYOpamAAuHePnTwOF9dk1DBuyQ3FlA4YzqkWQySOqg
gqZSRCMRT/ogS/nCIE9+1DM+ma/5NAOC2+zNbnsC7m++W1maXuQS7D5Pu7NN9lVK
073OTsKz6pPmVMzv20eri2EC919Jv+B3+mjvE8keYBCFXEB2ZGoeT6CSSaIq8asG
3O25ZBkNVMs/LOa8k06f2rDJaU3aakf/DimdjghMJUbAPLdecnE/gVhLcaiLQIYp
3g5FbNeFCCqKrMEVYI9vDhM7jb8id7j7UKeFOfymFCrR1JHL/daPnzLDKNthLb0Z
4vL4Om02Xt6o9cZsJrT/PSwY4BPCNrwb0YcjXC4Pac0wk2VbeMqPCdZPBS3HaVRz
UI+NSnfpErlEinBmBTR24mx90rsSLrVqVeaZlLH8u4bWWN+1PpQVXgO9AksZ+swF
kmXmmF5+COXqYfWRMlazU4PWn/GoNUVe5VTSlnqjm0NWcSY2SR8UDh3+wF1mI7z4
jSXeEEHjkJgEVbQwilVFqlmyLZ2ueRuDpN2xQXLxGamPs8ze8CH3mclVh8FmE249
vcloqWLNA6PgPj8Ud4/g3ANvkQHzsX/zo7/CIJHGYWYSxc+b5JzMm+9psFYym9xX
HR4XiWljrHss+mH5txsWC/Px6pq7Um84rLL2fRRnuCGQP5wJeo33WYKWoDMzpn+a
k02V6aJgbHL1aFhGaHgYJcKl2sAM7jA310UPm6S3SSIyvZYJ6wj7+aVjod+EIOE2
pHqLRjfqwiNkLsi2jMos1vLGJiFiH3MdEV1lsuYTgq7L4G7Ai46v+EDWhbPRLSSL
AKGXIkIBGbX/EZmKS6wkBu1NW/7PDEBETorv3yCmk3rjT9V/3mOe5k4G/C+59YaC
ok5ibMP5xXUpdHABH1a+CZ045hlguU7RvfQB8NFksFv6h73lZqufo9EPMb5QM5Um
um0srLycKcf/o3INCjxTaHz7Tb+gq6W3S3kZzAmu1ITLIJXUR8DkPTS0Mt2mSXt+
KqpEON493N/Z/PdEDDHf6XShJ2TQ0rTG0DNFYjnKf3FAjT0V4Z2x18qDt2iWcQAM
069HOPZ72UA2Pmpzyu0kbGi/QOCHLA7B4ZTUyFyuR9oGIuFa2B4L3g+Jv2EpzO3V
vet4upnbp25vPeMVFWY4WetsfvIOMNYpQc1bR/+dxUTvai4GIuBuK5sVJTxA4AdR
+Myl6fn6iUykK9qO1/KGJVAywCDGbBnIhzo3Mon51ICQVRji93vyGk/evGhOSRMt
UjXRqdR1LlO246Y4V/NEwkD3Sd0b2s/WYKMcZYmz1PkDv/7KB2khC/VpNKB7FGPX
m1OiyCV5Fw2EqXaoQIlcVdrigH7GpmBEpTzizrLsT2/ogp0Y7Zg1JnU9vfweY3gO
SbL65ETuxQIWjm4X5zLX4yKTHvrvTXZ/p24jaXHyY8kYi3ZMirCQAleQNlJE/avj
Iao3mK88BCyUrJojo6GBt8fd14UDfSMDMSgOf6M6yAYnwIKBcDheDdiPlwcV/sun
IRCy65irm3L9vNS4a+KmXib2Kn83E0jMkYj0pnebJL/YxyY+tHyK+q7xpqeAloxJ
aQ2SGk+ted/fn0v8M9hrQDLxksPxDO/afXE7H0aAEeuthKVPuBJsFP809D3cs/KF
+XH97eIZWBFzsPJ9oanPKXJzBLnx1z73BBCJKQjzj2v+Ook1blEEB9LepMkouoNK
StGx+ZUcEwmrWYboe3V+XjIa34MulIzeuq78eXsSIFiH2fOmd9RG8Yr5r6P7CaXE
4EUPpWV9QvXcMb92ZpQUkTyOaIrgHAA53+fK+9iZrh3evgxfFmUZdGVz3q6IKrEb
EEu51B6eYhqwGBaXv9cG2FfSnXgXAbujtCtTy2arMpLUwbN5oiFtIPxPiPuqeOqx
J436r5N8mwk77vg0C+DBdtu733IyK4ZhXgCbj4hMl2KL8cp8nsMEu/9i7/OP6cMA
rWqTNduX3wYqbdP6vAcZYtGZ3eld9sdmvzsmDfueUdBZ8TCblESSdZaAVNDLDVIb
A3U0pZdvCKMjNOiSc5Gx+KVADu24LhL9bgD6UHLk7DdKrq9OK5wRQXEsY1xeguEk
7AMfxoaPnUMS1/M9wmOFujFHs6BPNi65OrVBwGFNUmFE+AIJRIC2eJjYBARLYUfj
9QtxE/PWRt+HE+1pEHRqJOqbkARrHeOM3vN9TugiInBsHKaacjsdpfsFCLxeipB/
8ONIzuR9RROXALgd3iC7KYyoXVIq+VfKTpPT0USqtAxoM/3VV9Z/emVQBTFKxehT
UZGcIf/cN7iKRQWUscRP5XtYj5Sp7ALsY8UG/Tg8d+8HdAp91v9bMJSHCrpJT7MT
lgbFRa3fGi5Uo0gEhSBpZw4oO+i3TrKzR7XzU5GSlG4A6DU3vX+bItkGVvVLzBK7
Uz3NgOsvo3eDjQW22SxAWwOcsUYVSc4TSP72NAxIzIbYTn21rkFIjZqsuHuzETxW
iSe1Ogbwd1hMFPa8Pq/QnlEYFgyhitEbsknpAUhYtT5np3LcUPKc0KkvvwKzXnxm
AmrXxeF3s7NZPWmNRSJH1XDsWHw3ajOVg8nHi5DTiA6R8B2hW08SxpS4Wb2cTM+t
D07nHOheuVRy9Z3Pm/SkTKCj9qUjmkwcUr9U+j/yto2SGEr9OifVRKiJMazMTks8
spsj/8JlcAP6aoUPhvOoVfdJ1GvuuzirZD4d4vuAEkhIkjcPbSPmR4hR+JefeCm7
9qzQZQ3mH4ALTJRQP3GISKdpzWpIo/ANY3a/2owBurkeQESYNZLp4qymh/+3WYZe
JjuyBYQVBo4xOfJgi0DX03/VlBv6r1McENRkHTACVTKQGBmw5dB+Tc2RakHWWaOW
Za6Dc6rhiA8yElW6nGWLqLFCSY+1B18owrGsciQzSJzjyJsnDm9KSQFPFHRlaCKb
qvGstIxyU6MxXmNaUhDZ6n6Iv4a3oqQ2d3FIucjICYRs+JT17T8q4TMg/Lj1kBtw
46Rp0ZqG8dZXYdAuUpRLpDVM3ZHRsFHyoYR/mtHR1vaDMHqX1zDzyyNpIEywq8lG
SrCq8ZH0FoUJKM8jkXy0MHglVbnUVzeZf9HMIxBwG/mL9h60yrIK8Fft9YqGuNCU
jV/5bHU/tVlTUlBSXVPzhNRQdyEMl/bUr9p5t8wX/jDT7k6KFCkgMCAAeeelT2VZ
ytMTlMVYmOCBdDsA2Xv3a0siokNPNWmjmbL40lH/cnk2VC8o9m8G4/6avMe9fYA5
NbC8pTedHRWqV5/YiaWQGywdHYiaF+jhcs9ltUYEDwWwbUc/ggBtCgY4f4WO5qWI
ikG+Ez7sLzUA/yQPdo6DXih5HukyzGKhR8iriLYh1FxXLYIvtyjqoQAqN9e+0fRL
Ej57F6Jmg97knuyLQctocK5Gm9vmTuZmPvRQGWX/DIYfxH61gbsYWodHn3A9jzjz
7U2F4S1cmT+jDz+rlt2JsL9mWxS4rFZBkFB1BryWMUZfsCpEuqJrBQ9iYMUFTqOK
k+EeaDfqEJ7g2T9Qkug0Be/nMeKUApUZXTnEDT8Aw/VnVOvLM1E8Vq3dolTVBbRS
favYWZUONOvBh1RoYjQpjyfsavGqa21WaeSEa40WB1X8GfSa6MqOHW+5nEYDmojc
qVrjsFN3O26Mg566eX8WKS/ztXTvhcTG6vXVz04Zy8xXjvtTxKdUhvRWce8EXsZk
4EdFoq2l6SnARwvcDzNlreGDRXJSQ6lT3xHSR5F/94/f/EMrxlIkgG8PXzvC5x2N
rlo5alKRZV7F+W5gBm2hLALb1nwzZ40GiPGKCn0IEMwQe60Rocub5ncWakZCrjx4
T8CoBtgJ/Cn/S3ZIj2B7iAqujP8BqV5ANm8RBLtnxwPhAZ7Sv8iVrssHA17OT7Nn
FAsTVW1UXLTxwGnVI/HXVg==
`protect END_PROTECTED
