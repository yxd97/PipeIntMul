`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDQmTgANYStzKQetzf6qwZjeuSQhIjWFLYCa8kEkWpTEs/bHpwb//6pf1JqDJatP
03y71bfSHTH0/A79kvtb0YUmVCDbVezIvtAZPhDFw0p3uf8GuaWAn4eh+uix2Ig0
yYipisKYm5GeOGVnVbYd2+9lvgVt3oq434VvQJTzFr5oGe/cHxZ874eiZ2vDhAMT
a2CpyUMdwNcyIe6uizq+Nyozr0qU+RZZ49K1EBG3FdH5E6yx2ZEtA0OT5eLSHlmx
6gkoWogM8aby4Z8EfbT0P9YqyQpwr8gXQYMNkwb1srcHpwL0dItcKuIuo6FdMHdA
`protect END_PROTECTED
