`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ToHxOHCsmEPY49av/QAYlMOkM0Ucah8ETVHU8llv0GlGuCXoMf4IqXql0m5wE4V
DqR4olUncbri7YcahOdGPGnuq8k+Mj9Q4bJewkF3iYoOuhZU3jknqASzwdYTOLTb
HLoIOmCGUC+b4+8GXzsiZAb6i0Ripx+1hRGJPYxTIGdReswF8yCYEZ8aQZDP933d
jPr0RTVYV3ljihkyVELHNQpzoQxvFo0l2/7gY3hOHAnW5DMv9Q4dyDRSpauPlTdn
tv9EFICfu9RtcbNZJT74g3tkN214gt/P9cp0urhjK6kI53wspprJBykBWjMhMxm/
qpmdSsOlcrXB1e2WaCzyR8JweRK9V8FgJbMEJmr74KScgVoHMYk6q2xhKNtA5sjC
nsA9SSS4UxPlCo0pEkv8ty29v7/WEFEsgvTdLDbbr0miveJbUhBLwaCQpbAgTR1T
dbJ2l5bozXpHF0n8XfK5tj00mgseBfazkCH0VH01C7YmMW7BPSALzZgIPvpMDFp7
ht0Bbg25o12MtYX9GBmhrnL6/7GB1zpNpaOpJT4fxFM=
`protect END_PROTECTED
