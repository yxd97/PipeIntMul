`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ItxbFs88ytAr+fqUjlIhxaK3IP6zedBhIPOyNspw7w4kAWQfvvHsqQuRlMQK2o8k
BvgnXAaUgL/6qKbQF/s8YBWZr6UCHd5JUMsZHnmsq96ldlcma9WFUma7dLD8EFcU
Zm31LWNySqGXLEhXg6V7U7AVeJTwPI9XXH/WB8wcVrtbEBgxQiTZ/99tjyIXmg70
SP1LLuV6FlkSnMPYwxchLPB6MOxF+8qohcG7SPzBp1ljf0eLIGYHbMbkmbiP3eRo
rWzl5SpVhKR88mMqn2IKVx0JJK/UG/qwtB29YLgeJPGRYrGcn2lzCLA/fv1WWYIa
/dWsGs5JQCkwkALK6C3XOlU0clGtYlIJnmq/w/2opbI=
`protect END_PROTECTED
