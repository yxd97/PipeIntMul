`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGRXQOQEl0RmHcb7A+7pAhrnk1jd3ILARRsRAtQR6QUdKkc0J3omGOQuLgh+t5oV
pS1iyEh7sByBAtHt4saCq2RWWdODx80ZWPWnLAviE+S8WXNK3JQBXTi7DeJpyif0
7D6SHFqTVcQfluvmZxHi/gtQN1bzeF14EFwfQflwdu2AE5GwFtE1L44Ur954QwjR
79PDgBBy4dBBACWjbiHBR1Ouzkm6HlrLtOmmszusMAiRhpLqnuHmpZZde4cDoMVh
eexRFr+C5TIgWVhJmRvi0Vs0RF26OSw+8i3Kjc0ma4bgzXbJq+XzDlBDvYcQbk+a
NsVHTvECfk3SS6il18wJAEqaqdaQr0RkOdVCuJiF0vuXjek5ascwE0nwdMI1O985
QuZnusK1rQceOxQHRAqcS5367LLX9Xm2kBivwwaBEQSzuaguUEroYLq0JVJzPBbl
rHwc5w1Xlkt7wXJiKZQvj+w8IXtbAyAmPr8XWfUWMiIL+OPSR8MWwF9EilKAvlJE
TN2Ks4mAmsZbe0/cL502y8vRaO5mJ0NHy0vZkZ9CYvZnjbAzm2HonMVSMMDKxK9o
RULcEnzdiMuTfG4F8Y7tXN9s1RTf6+qyXGxv1FigaSAWY/PswAmGIqsY3q6oGSyq
LO1TjL7gN7YSxUqiU17ZF4KMuMyPV1cwFf/LAeLIvw5VCF6doY/yOiEkvs89oqs7
mbhhW6qnV+rCIrL1mmiSBNPv0lvOZ1YP8J1kmeOtKr/LgiWO6Bg4g/jMFhyLGHA1
rd6lEKCU0EBI7ZzZxb3jc+iwlIucKut3WbJi8VWP/1PzJPtuiBigBb9lyIJflqpl
b7GJOchaTlQ2CrOrVUdkM7sHYk451VKfLuPikTyk7Rfo0F8IgN/WAgblWaal/7bM
Houutq2g0QmH5gZfkeCTBIkqVHOguojro9YXt9FYsSUy1FeNM3+gkonqX8v2kqT8
t3vHeQmx/gPXXzE1UrFlnEyrM14dGUVaoks/jSZkv43p8m3UxcuUCuRu7KvdXySI
9eAADS66Iqmr/FNBwUgWreGgZ+E0DBwedGCLgqIHMZ7HwAg99A6yGr1LFiin11Ng
FlkQ++t4lm+Xz/Uvph+62xnkZqBHoNzGgEAPYZaLQOetkIv2oDna6FXbzpkjxKbK
+pSQQy0cgRDTEbp5bWdZaDHdJ7ofER2X7yaA9/9EiXdOCgmb7PmYuTflLAqImpHJ
QHaE6tbXEvUYxTBiZAFk/MRVtWkmKrnmYQy8h3BKmZPvCzd80OZQqRDlDozoNwxi
0LAz3yynN6aaQ20AnoVADd/ZoCDPzDjOVnIzIrbl4g5HlEqBFggx9oJuhiaOg5MJ
TbnEkMvQ7I7FEzzBoxOFQEZb3qNRcirrYJmQsorXn4dpGl9ttGgebo0NayHhJ3++
fnKvwkfspFwPgPtSR0QXoB3bKNGib+KlUJXfBALhd9dIFBRBRCN6WLhL84FWRsEY
0Em+DEYjORwnutMux843hhOt9yfWCeUDQdoa6fBMeWRAoV/BtvH2yRVuEcaMNf1d
tJv3pdumVjLbMgznJa7v0tDw8TnAPYeN8kHxsUSXgcbuUxz2K3qE7GA18nvmA8a4
8fTaUDv3r3mh/389nEmxz1ARYMnObbpm9q1Xd7+6OQ0qXYdEW5pyA7/3usZKi1SJ
VxcfGx1qtJOap1+T6tyxFXNiUCn0pebrLVQKfve2ZmD0vVCvABCSDhJYDhkG8QSC
MoO0QLZr3byvnQxetuh5Eppjzus0pALRmAGYhHSU+ouky+LKBfAQdtoQYkz+rx4/
U3ckf8ki7ZD1i9qoQOVZ5zDGjIjXcAVOglRlST3kEzoy+6e5jtnExaUZO5yS24wV
UxfbQUCNYTSASMQz9qcdLXYiF8NASmz7KtkgZMobXtrv6sajtXIc5bW/qi2rAYh+
egKVCtUYpSymn1epdi+eThy7cFvCQD3yx9KjT+c72Zs3RHwrScIPp1sM7j/nZxU8
gA080EQ1MsJ7tHskMDMBC7SGmgXPMe4WjFfCx2ftEztaDu47kIt6+I/kO20JI1zK
qfVY33x2w/gfv5yCsXOoI4j/duy+V6BRmXS9KBetpm8GWNPrXCxn0kll0TR+up/I
I2yLY4+e5fjc5s6wUgptIvAlsA5IBrUBauVprONEB5/jGMbBXORSDmBJRn2DWKEp
/Yhu81AbSq45a03vvxqzfMwNS5xmBTX0tQiTp5zfjBPb4JB1hUB2Yc46APZuUEmj
HJDVTXs4tspONe6sXOTuXVtZgAG3wsstK1BkEJATmI0qJLPDmnmBGHJmVKMJnaqY
BsoU8SLEohFBoDeo7PJ/uDn/leKC+JgI/722L0O1zOyEJNArDGNaGsdKgEvMGvzl
/TUX/yEejJ/YtnwwbwjohU/lwdU1GOioS92gJjuAvUpAWDlPegfwZ6KPz5NMg7S2
xMkuzDkfdeTTbXtqnKOD3ovaQL5fq8+XdFDX3CQpAr2FAudWWW1Vux/q/EOOYleQ
anmNEaibljQdXsiJV8klINgmwTXoSoxs3DPcmA+7Ma8/wVlIy5TDtkyrAuYPWSN3
+bRq3JQq8ssobMofKNP5s7E03XRB+nr6b1bQI9p2/nGPZXZ5rcm15fXuwk94x9qg
t2JmoAt0Pr3fWGamv6YYIe6EUSQR2zYZODCzE9XimQVJUO+39xJxWzi2QzDHkLfR
HFAhkzXU0ZBtNC/ZYCA08HFSK9s+zMthhu+001n65CW2hAw4jAPAo8i9Y7/BNfxi
hnN7U2IueiE3JrdDCzY9lChSQbVjdavT8K7973CeRYX5FG//lhZvCo7EyMkzew/S
9cIi8msyxxqJEWF1Vx5Kf3M8OT0pnuhqUwKW1J6OxgXVSZvTwD8IEMftyElBmiEb
AIhLsbc685lWT0x3CoUMqQ5kasNrD+YubXDAvUT/6qdMu1Ao5ny8MIEhCJoMajRB
sf5jqBGO267ycP+w0SeXk3GIQ15vjSkam8r06rMGMwRZf5wX1Tkvbpi+snUlhBdG
CTg91XrizixPL2gWObGq3ClG4IYje03yScEyAMv8dy0X356gp51Ai7EzA6lFcrV0
bq8EaO/ATg3VQBZcDe3Iehdpn5oTesMwzpSMO8mBwwYSc440GTdOSJiiDvTlN39u
BHaHJEr35Sk8N4mRmh/XP8nN+02GQJWX2H7t99cZq1cc0UPd9thamUwfWXrFgB0b
/azxE3IynwyZdsbvUVw8A/7bSQ8HN0c9Jl8NxPO0H5URRbDUXhaou5aP3mXMN8Kd
ih1vjGJZbLPgGz0vi1YKoRWmgvb5ZoLjjF8SyLrZAwFD3A+p38UwtfqN/BE7ilNX
0HgTpvknGqKo6+79/h4Wrr8shgPQs3mvt3ztTAxHErkRXNM25S1bhgrGdLjWBpuq
3BuSTMR0f62DWwRrylvTaMYCz9F46uI8/rAD2+jHcmOcr6488xNVUBJCZDCjDPt7
2/15dhEVqqwrG+agOnW3WrD/742ReaG8uMZMYxnANio1DCbvClvzGAK4H5tdY0tO
GB0PFtNvNgf+g+w46C5Eyal2Q2Zs4MSIWWddBfIcWxEMd07WD96eqctP5L/fXc+Q
0KgZ937eIGCfc4c+VUbJ8BFtK5Qtv10WRWOtSbZBEBD8/c7UcP2vz5+EZtTk2OW5
Z50CS/XELU9kb38eSi9sYDxULjrydDkU4D2Bf04tQZi9suQ/b9PsrNwldM8CFO2/
LgydvyUDETBEhkzQjLJQd5e0wBk6Q0dV2CV1JhEKcCzAghM9XCgaKe3jjgvxq7Hy
naiGsHfYzUeXPlXjlQkA1g==
`protect END_PROTECTED
