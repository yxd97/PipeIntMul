`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+FG4gevf48u/OdQus2e0tHKgrfkUMXGBUrujhYmAASLQHfkRg/LD2/R7zY3pEGmf
BS2IUlOW6uViTZgXo12KOfRul/ymEG7yUlOq11B2/ZkV+LbvH6oeamFMLAGuXJlg
so3m+ECA5PEDtMVSLl4eiTBBYNI6fWDpkmw4+JNTkqs4Fk4nkrmFI3/dYB28sWK8
KFuxfJpONdig7hEHc/pQEcRE06Xs1eSJbufti2HPovvEOX9hHvvxrEqZXhiXCjHS
nxk8ECFQ7lkqcuYG9GM1bcdI9+q/VNaFqRDM3N7hI4TZ1c+eMVUAk14jXQYQxadM
k68Z6kEiFhzBDQQhUuoE8r4OU64IaJbBTPIwlRLvNy5zijmPqzC6zL7nj2wa+hTB
MfXZ+cTL2+R9W1cWxMknvNQ+cnx2CPEZ3pzK9OQ/Ml0=
`protect END_PROTECTED
