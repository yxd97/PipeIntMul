`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDQAwmRtSbEI7NWVEbhArJ9X2vbI9GBewnHIotlQA7i1tx4GkeOciR4ALM2ysj/M
UGJi6nXTgRLkLyW6go6QsIajhJb31J8ynH0kKurHvtf8lgFlshKgGVIX38y6QZzA
sRyC7hkJTQ/chJeyu8C6W46A5zWVd7ex/c7MQJo4JrG5gxuKFsvj2qZrCvhn0LCU
zJx/qR2FJFk5s/3+6kmNfL4d5Ui6oyJWfoepqiApJI9oDhJLmpoqGCCMd9MCMeNE
zWW1KedBheZXuBxNZQMU1CRL//A0miExaZHyC5l82rGTSr17RJDVTVWoKB3J3WYP
Ho0vR7tIWoBkfAmhccWA5VOJdI/imWJQ19xnuR/CtFYlX1JsiS0bZdkG2XVu5N1R
XHktCKDIu5inX/g7PcHDyC2V7yvY8nUOBaWph4zbnt66Te2WyT2XvCb1uFBlMeAf
0p8eKpWBRcqPkdZHF4plZQucWIsfWeelT2mh7Eo/w4Lw5s5d7lfynJEJuQoMaLFk
+eDIWjeQsP7qSB2grbwIKw==
`protect END_PROTECTED
