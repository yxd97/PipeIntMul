`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7CcFZM60mzcruaQTUskVR4E0qoNYmtMDFHVZpeZubPXi4wEOnsVZALa7mEV9ycN
TOgZSbqHHkniM+FenTHoWjanvoMIJj+2+++PaGV6WZZi/VVXAiqafqI2RKvTDXD1
K6TxeLeTJejMfqCYF9Gv2s/zTSpA6w/9lO+cBcbDjB7Q4aSkk/RMxyxgQqM9bzfP
4kDT7vTe+hN5pZVqH3HY61cn2arWRVwn4/Tsr2qyvtkjeRl9bASV2ku3qqqhgoPg
K1eSH3gdIkJ+iWCLX2dXyZ60F2/VomaeQIG+c6USzCXltcJW+Rke1vJ5VguOXspv
65uBbK3JK0f4gcaCfjWDAYBe9JgUe5czHFvHl4c2K2RvgMMqPvxqHUojyIt/CgVS
`protect END_PROTECTED
