`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iV5p5JUbLvq0xZ+2qhySsen1l8zNypY7WTFsjN7h4o0lb+Jmgq+F/cf4NHNuh8V6
2fF85r7DUGIzaBXA01MjICPK6N9rcG0gcwA3LbLZx5PddviBKvkgR+40xfBtVlgf
HME8cow+72JfMqfvb8+G2HxmoDM4nnFON1/BbW+iEP26H9vGdxVaT1byeEkMSgUz
Y38p4SCtzB0vhTY8bzzBNPTZKsUObbddvQUk+YFJ5aZxWh/EeNBwsmopw2FwvbRs
k3Nu3hL8pWQ4zq9KJRra1Cx2+InL4NuvRTccKLTvfgDxRIECjSKnNDKn6IWcCB0B
MrJkRHnqiJyZMpWYSS8lUP2dVoVtVLyhpktK4v+1TL/aWxzMKQ+Wpyq1mxJs6+RW
o9wW5OOAaHUpV5ZvqmWV001MmhL8eozbRuhqeJAuVppolPHxM5P/eNRupTQphPn/
u08ZzO09s86GeslkWmfEFI0KhENW0zDOFnGrnEpFBkPc2bq0Cchx/lCRA5JuQLVr
5pfEpMj8SWNKLaTWiGhfohRDko0X+smv1thT+Zdj2XPhGRZstSyRsPo4IsurH+be
ahysAf1Fa5YK3r1HRztk0tMfcYI31alY4lRVylQNhg6opzRFqP1FTMbL3fN1lfV6
`protect END_PROTECTED
