`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SxEuvjjUDr7lXaNPD+f6c/Urk2peT6/Mj/XsF8WJoXQjwNYXomOpbM76zTufvfWy
m7cDoV0gmbsQit5nMnFp2AOaXO2NeG6OMG/tqtx3QWhsciqSzVReufuUxfIRt2C3
DTdYYZfOlg1QIYYd6Pq95wPh960CKg1lih6G/UTBojKiUOOvEhdhUW3aIApTM+pL
GdrDwO3Cwpuy77GqM2uNHRHlxi+uc60PY5XZNZsoZzqj0oq7PCv6M3CqO5kF+Hg2
FX4/nTEQ3thTzbHFxjg+BppROGbUxx4pLcQavnqDnxlnoP0z8Glx4FLTqK7zXJo5
yTVkkAiiJsXItAY0JlF1yggxuA9FUnIz/8kXNdp6a5RLzhnpMPV1wS0POCplA8O9
96hkyVuqy+JLtgYxkSB/VTJ/+Lot1WvKrPFx5VsjBrRPQ9VKPZx1a+Cb5Lyt1YJT
Y0c8zu1fTOIIZjJ2WgwsXsCbTDstFcDSnDHJxmWC7vyyxy0nwmmkxAra75emymRm
Rm8oRsfFDZVmsGXSbonoODfPElgfUdXwjOXdwY3p++Ch4GE7O6BDItutXrnRihCV
v2HocxGmZUp0ZWLpUebj59ePxNT7508fFGIoDevAcxsiR1EdeAoQCItNEZ3s8vuK
TtYndjN5D+I0EXoaOl3kIav2i6SBWEhnXr/SdX5SiAayccKM/VDf2fGaqqJ4HXMD
dMJ83oeR46lN9y8EgHngc/uRHmsFLy5adupIOXaXuBUtzTpbGH0bJM3dgr2rq/ch
ZzXWeUC0FRl6r+iV1Np+rCRVmu5UuNG5F6xdYg1NcTGGHc+ju9lWBhCFXkhlJ/Yg
70qm2eQ3GcOcwLuW2KEZ4D4+iYsRz0yDdUamqZZzLzooOyn4bXKbRiQtCdGeaaWE
Vp5awCbn86Gofd5ZSPwtTbEaZs5CFCD5D77wRcRYNbs=
`protect END_PROTECTED
