`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qhhIEa+Ln0kxEW7IBfkoG5niHZ7DN0joOnv34DveoWfq0ji4n5FGavPbBf0EVgjv
LAIYUA1wsrF6c/8DURLRLJW823oyl6ZRBbq+8hLMXjReRvF0ikk62z6/T2C4/LS8
nHJsQ2GcniHKTmV2D37WdaAgeL+mn7N5rbQbtfAmLebr8oSGF8lvrxbB0f7yGYwA
6OORb60NGe1ta2/rNsYYis1pYQlEgAD9YxgVQUYoALp9+Qm21K2pkjxCG5ro1S1p
`protect END_PROTECTED
