`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSKHoiSvO5LEGe2mz0wlom3v7x1feU2lPk34GvucAGFlUZis+Gt1rRoCQpp85YVc
1CjdExEs+2X1nl+bFU9wuVPjlaIIzq7h+xKaA0hkQhbBt18KqJ3/DNt3JC69QtvQ
TON3G7W4r4W5ooWHXxDZOwPDuBbpQuSi5JgPXr9MDrQG11N1afKho0XlFrIw4FTI
8uR7g2yuh7NVpR32MbL+nelSANtCElEIvoy/ExbwFx6c6kuWosCxi8qLpfJAoz+R
parV3ogpJazc49cd9j9zZcL3jkxOLcaY1FdSNqT4R27+yqyZXpjNtMjmv9E9rAhR
PEZr0DDzBtTVVOsRlVF+kzIZekCmDmyz5UeirNEmTV7063bfoaTh78dfXW29VsHX
ke3O2v9126hWHpolmvAhdNufcH7wQUygwOFy9bMas5Mk5SnkFcn5W1Ic7rYSSMHM
XTUWd0n18TyN27QZBHlTE20WOENUkWEPWaHXqmhcTnM=
`protect END_PROTECTED
