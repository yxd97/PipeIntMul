`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9mqdQEEqf2RLkrwnLKzxJwS6Qzu5TDIYz82G2cPJv/ThIdhRQ+fhR0qE+g18plDG
2HMA8Tgg81hFNbz8skmaEilDGzS7+liQx/qH6aS5ZUs92Sqf0YAvRjiXZu01It9F
Hq4bMOPdjSdHJUAIYH4qC0tlsc0KjnQ6mZeYkuPsUHjlv3XJh4enuT4COFi2CCr3
M1abg9Xl48NQFzEHImdtDn2dYV40i+HYYFtAnJbe85ZZaO25IzLsALEIM/wlLjP1
51fdo1V95HZj/OyOwFniLKcgvF80xa6rELEz0xZk9R4uexdJrJGB6EBSgpNGxs/X
WZ+nNGThuxRgUk429+46MAWIokHASrVHDhGzqhh69DmtHO21/rE8tPsfLRskBbGB
`protect END_PROTECTED
