`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqmhAYUAFN9alZ0ypcNwkz8yhC2KMuD1WlkWj4T30Db+/oRWzsQ2n3HukuM0l7CL
U02vZle9/iSRV+Wog4TKSTtQ4ACpE6yxxcK3XEmwKdJPvI6hG3oXUY0/2BfeEPEE
cKmsIAOrl2AlFujAMlXuRgNGPKMSKb4A4TlfQoYSkXFoPpfhrC0sXewIPuQjiJtS
PGZ0UtwzZGKYN8bGKFpdOap0DmKmpjMkdaKPcqEdPLbPh1k40rZkqjUFvHioA7tX
g8laS/43BdAW1y31Hf+HHwalAPlNYyMPKEnomfgLWkOB4HU++g5swqUGtAXcKg5U
jyqh6JBFR/LN2jkb1Rrs0H8INr8CDw0bT1iEYPAF3zPtIvA+uOGiYq4hj/mwW6pV
+7JedmdtlkDUVOCtUMJNBxV0RZwEdgngelIWfwBxpcI=
`protect END_PROTECTED
