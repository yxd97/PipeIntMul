`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDd57WRNMRaVv7nMv34DMBkuiHksD4ooTPZWPl3S2W0YDLhuZY6GYEjaGZZTF+6s
mRAmLsaNsz2H0iNiG5VdB7xXAoF8wnpdRUBkwANr22gecrTMbbf6XqC1N7HWaaSe
z/A3sefeF9UG1CZlmkkuJ2GiRhCbrQq9YvDY79RtQda/QNaOeeUd6XE9Hgwu3jVG
dW1VfQZXoW4IKWeCUcvmQlNzq4YJhkjwnfcvLrrpH5AQzBy8ovWKclf20/22BS6T
N55CZURPDzNAlFsU6pz+zXR4RyxDmxG7CkZOGnniw5sMnQXNuwUP9U/8uqvSSyWd
`protect END_PROTECTED
