`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9IKDrcvhbvzRDbJqfYBtSJFFOW0eXNoEdx7giq+KVW6Y+pfGpfG8ve9SsLlsxaDs
IYgBIbl2QNVF4zQX3TRfn0pBijOCzUoLhLOgneaJKcRsn0vRfx0e3u83JbW+A10m
hPCLonTRVczuIiXRXNF7TxkkaZWIdps1z3z1LrYpfkGlD75oPA9QExnTIXLC2Yuf
LVGE1d0I4R7SuAw54oQoRJH7BKUpLpWqNUW57vbG54s5qHCiMr60bi+t5aRY8v9j
yyDTF0djvPzTFR7HcLubyZi/8MfKxHu16+Rle5WlxFBaW1FvDN1bSX5VBlUeBgBq
EWraBZGpimJqDBV46ki07C2pV7xeXsQu68hm1290EHI6eWGt36i+munrVvKBloBC
Why31fNiUsV4Ydw8Z0Yav/+MWO9qfcJ++gmjs8/oVmA0u0AJReol4BjGsd1B3dnP
7jykoonNweg8JWCy1HzQylXv60QlDF/56z+trtpB4aAPPfMixcK6WV4Y8K5JMyY0
ylxGMU3zg3860VsB5bMfTIqBNpyCEYuxwy6x8M0mjlS3oguawZ8P/uhUgSlCg3d/
m/0SiiCnpYA2Ejm12ku9HjcxNdubIzcfrgivTETJOUwc3mj8xstn+c0weOeN8EWD
ZZJt06r+kixVlcAnD5cCbWVbmNVprFbDQh6q1E84+97YJsQ2SKL7cm15J8g4Ovt/
fPN/DUH6pRgTvvg7a1OTAeffD2Djd+eob6P1o6+7niwdU5cXrQ7L4D8xGpLQxApY
T7QrQm+kBkwS92ImfcmgBERBGOHiMvEwjJ48jDw14pq0DlWY9vplBlNKancVquN3
zkUhqftyzwLe8phPxbf22Our05TenvEzqnwZNxV5Uefrtmz25/2Ft3PpsAXz0REO
5OQIKjvBhNUaZiGdTO3VGuBnGKa/66nmKl1oV9wllclIajNNhY6PgtSUeWobfyk9
SJWdET2v5PHn0M+FLrNF2KY+FMoKNj+pgcVQNQxp+y/I13iWI7I1JAe/QODCMsc4
Cisu4tFVRQ0D4Jz46SXqfIuJ6/+kiFf9tcmMgvrrTWnVkycnzf53Ipu1Mq/aVHj0
yH7k5bpRcSzsNvOrvTTyDhcmjSLZvQS9ReuOLaoIi/7Q4LDGBnY2tY7Glrqe2wGJ
nRjvTolzDdhQpUyTrcWiw65in984eKq2WBw6L//vnRfUN7onItGajGriHQm1mPQt
8fEhASZpKcT+oaofHGQyxZa3Kw6ppP9TS+/Ikh7gTytPK9dCjMfxGimBRS7fFu4G
EVPMXdZEcV6a2OwMNUWaiMJbo4BKN3ddefDl1Z5PS1aMrS5axp5N2iy3qXbuu1MW
LScbIU1CX8ERGndNSBTLVUeVrW8gfSgt0ddiBnxH1i5K24n6EQ3nKUHzX1AAU7/b
TH5AgUxItjHTWzFHfyPQRqlRagMsKV2c9+bwY273NJT01vaMAocFLb4T7LsZ11oJ
Mys5QToMGuk5Nubmpe19ceyw8Jn9/G4AIjQGIaczBmTG56ku5VEBpzsRhCTudmcS
ycoRdgOUxtPnqoZA5GQ7uBuCmaZ7LUQZAA3SGizMjwmM59ooSzkvQ9BBCFLETYB7
WJoCRzZ8zl5SjPkWwMsvRZIlLvllI9AU/rId3vJQiPa2LIY9XMVtDW9otur6fp2K
kK34G6eL6sO+Ti8WBLXRBokJParZ/xPwTq4kyEYsvmpv/yHAHgd7/2K0yRjr56lQ
uXGF8K62drSEXFtYpc+lMgnzR2YzlN+wGVEiBKNxy0wbY9MCL/Ps+4BxOVrCtMwl
LQUJwvxWg0tvobLoqTuQi9a6ObEjg/7qmVknC0zDVU3qDTctUbTM9SUgcIWrW95a
rXKMWn2QMKmMk5Ukoanj1u0W2d7x17Taw8JgQsLdzYrlcaOXFyXRW564obW/D4nZ
X4d/tAEAhnGy0PoU3ER5wSeGxhGY96z6cMbfElylhAxMWOFkSbeTPxY83s4pnXko
sM9/N7ZEgzvbdO0OeYuEuV1TZNmpuiIsqzTNszSWfwOVAq57XoESqUj/qd1eWWdv
PaNprEGa0nm8xSVG8vqI9Q9uQ/0EEDoHhQRZA5YSbA53dtlj+Ye8gvJXLFxcRaSB
8uRJtlUMUcDxwxMyGK4JL0pIYUcof3pa4i6SFCrVvziqNukthYJ3TmeTNFFOQDcT
kejgwKdXt/8wSZDLNxnpWsLLggm0DwbHr3WocG/5/K+KMTzOZ2IhLLRwGwyVTVdR
lscgW8ACBIy2uCngbJNQpcey9LzXGYe+TutrseIRvY259ecDNe46s4gFviNGehG6
OUqCqssC9pOk5Xr5yBcFtqOVSY1iSyRvDkzDINEVi4SFk7Tuj0JqaRo188GHDHZY
fiP+f3ZdKJntQEI4CSDl8/5aaCBotd7/gcohXvp/8EdrJXA3pGTM0x1kwS/GaGQa
hIsWCLj/hxRJfl690cdqCoeAcXO3AeCkTP+hwE6Zpfpovfj+E56l1v9XWfRyWTq9
Y9kHgh9iaf5fplRHoeijrrWeqbdv5N/Xw4G+iyMnfI1WOJl2QcSr0frf2BN8cULm
HCFIeiiMeLJb5YM/jvKuybFLAFFLGDUmaoyfhiS+ViY8Z+rChjXTsLNuu98BzKFZ
GvCBCbUGsrTOSc2B/EpPxFpPfKchZ9vUVKpeJX9S0O4Bl56vs7Zh1ITz9z3QvIln
xQ5D1FCSdjt7PfBRMqXmxRrgY59eKZGAXNYwsPt5wq+NT1vHeS6AVBPeEc8yxXtM
E5nclWNyaSlSs4ES8M/8CASbY9tMrmkvH/TdqsBqJRLPpovmlqgXp3BCTDp2hPbx
96uY44Pm/0Rse+tbl9eRJZ7xVX9XkZiToL2GnudNkZRGCvn75O+bq4bLl+pPc/Xl
fR7C2OdX+09E3/TTyxycTkm+t8hMtZVzly2gPlUCUTQ7mXVtqXfXGdb27AbuVKAi
+tf/Xw4+B8HUaEoBd0QKJC3pIq8R6Lsk9XE0Yye3wT7YUef9yALoMiyJ0HKPoGTm
ylA0OomdVsTwEX/cQDFMsqJpM/H3sarWWPun3r22OFEr1TTIfy8xJsHLzrV85b0M
JjEttwEORnUMAJo1paLMzMeiEtXtnE/dWhe+Xslreft6f/sXrAK7Z8UEF8bIq23a
OnUTTywdDUa0WuWg2JZRYugyYwx7inxfoiZeDBiog1Y/E0zevQu7jBG0zLTnpcRO
O/Ui5/iYV2tyh24ZqbhRgrXGHxPbwl+m2o5RCClMeXnj3p8j2+wVN2MRyX/teZHQ
KmbVxydKLb5mAONAICj73pWLsjNNNhhr98QmIc1+CLBZjx8mSiEjkuwP+l2THZHN
CQboVMUzjRmYSk3kFInKAO3konERu6e1jwWRo2N9JUdodombkFC+Ishgks/2zMlI
doKCva1DG9QmgOPaqOJs32X2dFlpyP/qe27+VVSQ9doQs8QKakwmifR+zLtlPyD6
OicXgSMgk2UDsK50ItmWwtSEiIg5/qjvv6ZOWxztQU6RjG4cZ9kDyVg6O0bfC+gx
6w0rek4ZR58po2Jhc8HVPNFSktJJhZH2B+xvx3uCEI+Bnn6NtwzCLfrUpVCd5JQN
xyqmksVIJhtrA0aY2//px7z3lC9o/r1n4RpfzrTSAie6x20Rt4i21FuA0SXJ3OWx
2ep2CexzOoa9fkEDnW52KLjoWQZ0N5WCtWawAatYJHPSanReOl5EgYG5aqm8hoNd
FftwlkXPAt8okS60BT+RqL8gw3NRfUgBMITcWLLVqEdLnPWoi3CaLtx4ctSSqu86
VfB0TYmi9LctpkV4qekQumygp4gxFE+9ZZbJn4zma9JTGM48QsBEHZL6X4teCVUY
1H8EEH+ZOHmcVIcO6ApDBabwDfykD2SDiZkREles5DZ1Ua34WdjrbWp+PMVH4nHi
VZt3S/M2GYFmEaXRf9nTBkAAdHrx+wdVwosuUHkutX/wHiHOpWrGKgX5qIaNLquI
E8w9GCVu+hapxKGaCEZySCjF8amgo+jIaD3Du1Zlm7f4pw5DEwBpFwT6yRIRwLKu
pOVQkHe48ADQBXq788ugv1396rsQC7+H24loGZ43CaCppKIbRLh9PY0szWGOdpNs
5ovc6+aoY/5lC+GDFWMkL0qElQq7xypWDtWH8RWWRuXBGmKUrDF9Ya1s98uaxvt6
aWkFa5JQR9caQnKxVruv60HppU4WgSFvLJ3nfQTzZ23pEmlog6frPb1t+0m7cjmD
TLqneH44L+KUl82PKnYdp+peKjyDQQyOEPOwUZsDHC6/MCk5OSCP+DnX9QtNcYUp
mt8zyeigOsONLMkMU2HSe7WO3VPHqQD4u1N/h5n+sm9ZAgNyFc+pMR2BjQKnTSmR
RAArgeHSSQ5A+g2Br6vQEfUktZTGP44W3etZnFEXj3LL5/S9R1RDn0mISi9GZZOn
hywnxsOi2PBLU63h2FCqZlg2scNDzQEuylVgh8D/jYK2AhXNZiU25avacE1yZGMl
boytHso5kCnUzh7vsHOFldZTy8iJ8ho5zlOVOxBUoKkc0dQh2lMZotOL0H3gu4SC
4mWLqtBySvBGRgmokTNmfmS5Xkx2edvBpdsPVaq8Ag2JDu6jjDcx+eNR9Hrj10P0
a35KpR2SGBjn+1sFnR/aoR4P1ca7XQDaeMDV0JLl41Z4/n4Eth/b2rOeAmYUCeUA
yvDCm+jNpyCfpQm4lDPExVQtN9Lyvvpe4LpdVECZW97ND8scIBeEPQnOGjZHvP/V
8+ztClkCm0+CZtUfLTHSU6opPEfMzfvdRMDv2K8BlQsAWck8Xv6xRbI9ANTV/hRc
f+SkjHV6V4ULjIXBi9cBgJGjPxNykL1ZAABA9IF5xApkA5SiZwpNd9gTlSw7XuVY
c+L9sfh8HRo7G/iSmQGNa2/jWXzA9Ciu5TCLZddAMhNsJ+msCtORpPf2yyfA+Zla
mQGCwTF51OJXuM18B05ODafXbvHz4Sl4N/e/sDydGeJG8SxLPfjbabiNQVNwiQLi
UIRqXQjzsEbFZai3K6aKWaht5/Lw4QoxMgZvl6Ox3zewmoqSisTHht86RyJA+IoK
kZnWWQ5TsfIXjhe5eib/AiWT8ld9iRMDljzYXeS8aN3nJH6mgPLIT9rrZBZalElm
P6fD1KVcNEaqPPIK06wqb+lIS+L1RsNjv2mUze3gHf0dXCXagy24vvhGB0LzxqLO
gmJ5WmgAD4rexIEwLbjmoA==
`protect END_PROTECTED
