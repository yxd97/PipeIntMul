`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3UOLVbAzbbbRFQFw1zNsUVpeFErTt5QQLOw/JREe9nByTy4MwY6ilbk45AOJmT9
0m9kP7gRdkexzz8mCV2087/QHUxTLmikwXu4bf326uogFEbaKr8qMSKaay0ad2Vv
cg2jUMZDrf4Ff0sAxWC88bB7wKhAxrh/XdnImr2Vl6Yz30QGfSdeQgCSOqraAyAA
12yIqawzAO/4g+nJtODJ5pOBpj4PBi5bpB9vG+yV2AnqOe+h51gIpP41TFOH7P2D
uqUasUw50cCXw3LAx+gKJG7hymp6bl2OZ9At/HGp+c02mtx4gNTNBr4fP/vWBTXv
S6fkd5jnne419n5elYFjt2qFQlMql2UNcfYE5d9zBcWBhs7bIyWLjq+OJbtc1yo6
E2KVb2TXwtxFx0HXnAnpQ9Yk0NkhFapYt91fjVrFlGh6cHTETo6aWENwNcaWaw+e
x0sjhJSzT9lClPH9ajKYvuxwp7WqF27VK1rzv+XYf9ogaK8Ii067DITtvxsPH9xm
lyBu2+Vzaa3OLThdLrB+aDFv/yiCzkEDRnZQoeYrjnnl+n9G9NJityxbB0M8HO9h
tSMzQo8BMToi+lO1lYmPxEMf5rroEghiCVkrL6SyhJ7MUcHiZU2BPMePtE9L9+56
HZcwUTQHypgCrlCai+5wlAr/zUe2WQyRpT/ypxAdqws7CEMOhlgbrO1Fi1vNb7Y2
M2QZXHiZVUZQqQEuABVI6cqzdvIA20RT26cqKAe727llHP43WHjwugsJ3tHPUEMF
QkST/akkaL2qmXEVYpQpF1tKN2dcyIkXHC+YGfmylrQwX+GwAWqRP0oAQXR4naz+
v/o8j6lbD2oJ6xyDiXQeczArDspirqpUnDOV0VUy8FkMTXw64rTU4g+EeZCaO3+V
B86GbSVMPzx07+F6dSvT1KRdvemTnyjGzonhKed68ybGcWw4kPQBhZXTrSd42zLA
nRmjSH1yrLqStVbQk8CjSgCMU0i3OfZmHdXkUjYdlLFg+sKPJxCSHOYPt4zdi/km
6IFAj9SMLEOysslJ82NRv22IhJQjqmMRu2yGYq8Sf5lIBZMFywJnOgw5AG7dSsRu
/LdZklxxosl0LHozWMpZPHV0oS/yPMyb3FMFQsCw0HfCB+fbbsKi3xI5S22SH1Kn
JZVbtzdBpIwnSeYWAJGmX0gK0rC6TkFrHOJGvDg7sANCkOrQzs5sdYpHB36ZAUrz
QO9ikq6ocJt2SNPE1CHM2+isWkYXlVcHNw74XFOy2sQRF5YBNZuxvFC/t2opO96B
wrIKBn4hfRDgQkUPLpdQgm92ac4wwbrLcQGtq6wg/vC7q7N8e+1qeAKou7FZpQkj
VG79Lf8GD649r45+MwCwqbrEwXB3p+1rzMh5T+/V1qMS29Se56twIsc22+qZ8pwM
fxs9W+lEA9W8v1m2L4DRAxrfqCyrLUm7pwsno3WvPzbbcq8mIFeSTtGVVCiIPCfV
UPpSJS0hZWZRwkF5DaXQa4d4mvT+Jf3V+QByi642A8GNtgYTkGLB7XoyMyfBuAmB
uJSlhPpO3cYDUXMPV6hMBcLF7Af/EI6GuqIQE2Tdr6czebW2LkEq6cP5XmeAu5WG
K9rTqoEIHfPBR7522qLwsjbDDmOROs2ANs2TbH0pB1bClSAS5F4Fx2X0Nb0tSWNH
7xRU7p7Nkgi0MOO7Pwnp4UhQLzzE3lUDdYEuRvYF5/Q2/iFgH06pq2Ldvp+PAL2X
/cab6MC4/BVHLisl1JEJYDS+fYCjIhjvQtBQNxlFJxj/sqQQ/seZ2Kq2cVOC6GVD
jdu+xjjqlrJOQqY7rdPx6zDzMeoUBkbb1f+xtgbDzeqVxqXdw4hhcGBxTGMO9b3t
ien2uu/Bog6bi4REFwb1t7VOrIlOXjuz76P0xWzJ0ihECB4GqY+OKxBWQ5ovtiOJ
OPDeDTK1GMSNGyzgbo9qu86knmEzghsFyXj+vUbFoEDAUQYIONbYvUjWIE8IkJP0
spcUt8iuqNUBOuxKlAzw6AghEAEZk2mx3DzJtx4Rdn1qtc278yGveLj5V1ULeqpg
p02vz3CAro6kmWAHFVm8DvtyeDUyXy2mmgwhWWJwtWJPdwqQ8lc6MeEX57pUyhr+
39g3MUg6X+bSWlUghvUTBwM4buTdfy5wdwy1BGdJ70CmJm8DdQPBS7WaEZZPpUgx
IRjtlzjm9vuxxlZcelrvNU1T5gMe37eYNQTIsNgERy/eQ5dMECcX8w+c0Z+JGH6H
ZRRJ2DJyVVm4yLppYTPHiQcHIBxA5V4dPuo2uQqKIGW6la+EdYjega0tIZCYP0tl
MVCtF0/jLdTb/lRfOp/F0Wr3PvvFj1OXP9XTnOfH53IOGeXw1Uu4044IsF5mXLCk
55S6K1zho4LD1cqZpXRHj1VhJnDCvbHEho6COwxCpPhu3ZWtN59LpuWYl+SAfqwc
mtTWTV0X1np7KkSTZCeKq0SzhNLMFgcQM3cC8X+bNedQZL3BLsqS+RBUbrb830TE
e3T2XI5EW2ciYHi0axsaEYKZ6PZ2zWQjETGzIXO4I/T7smxBHnrOl3A8kwsjWAg2
WPMreD+3h2dq+Yr/w81BkBdQdJjaaFbSsOsCz8dUDWEJPUaFPP4qgxYtPcq7BGfW
2uuWLSG3rtAAiwoETdNZWWuVyyoGkjF1w8B1TAjxuGqds0VPr14nPN6rs2lK6tSR
4J6KkJ9r7HF3PrxPaCZ99G9DFFWo1SPAhMCp5pBLhQPn++2bp5sbzRiO7koba922
LXDSob36BVHEYU0t04VIXh5ZrOhPgoRu3JKUTSs7oil/I9kU5XIsrDrapI5XDM7P
PujEdUHbEiVJnD1h433gYlEjRKWw7Yy9yFFvGZYmfo64v+1GPZumA11Nx5ByyS1m
2U7RYMxNxCpbly3igzuEX7oYTHclWSVoEqReNVJhpbcTqMKOrmQQf3JyGVgVFbpP
7YNnCbW/7sPagylhHPab06j7gbeXA4dv25JlWw2JVWDONV7T5p2B6xyHA55B6jrI
r6f2owi/nzPgX3mmwvFSB44YguFk0x6kMth+SXl1KRrjlEvSFC7nrwX13Qk+Khhp
4s03mWxABicKeYeHf1yw7sfwVgZLyW+47Kjj6uKaK00XV138d5M/eQqCA5tS4ase
hwXuvWWalKhAdFxO+hUgOdk7IA2P805s0a+tKecMoUztCWu/kRNHT2I3g3BPqEOE
93MMl/Tkm8AMwGm/yhzAGtus70w2Q+rKd0wgxT348ZQdjr12Zsh7IpQsUaAmFP8d
bscSNErkkei+zF/sIHhULc4Ew5ovXGU4vnPdtpsh69Y8uhiedyh3UonNoInAoeK8
g95dRYbpKPRXAbWpEt+4/Bfk5apkJ1r8l3oyAQIs87YLs+Dy93l2UjvBN27dQjZV
mi1rozMyEMaZGEzeTAMGNW5gIQyHuG95K78VH1uu2q2FHLl/8oD/rrjlfxXkZepX
q1teQaKtaksarVi8J5D/6JniMkXnKri3JNjNo/uD7e7LljstQmowGmVqC6h4J++M
pbzgH12gykp9l//rOuccfomccbfhlpqNLlpYY13rUWblyPQo9WS4Xrg5Hm+YY+fS
WJkgVk/9iPY4SOAUqKA2R1G7aoBpd4OcfAzTlxOrvEU7mYkmUAtnvHqwk+RaDPfP
Z88qWWw+McJF99vNznON7k4MwZpfEaAXaqJ+ZCFp6JMu8Qwz5uR2Gu24PTvyk1pK
7CqC1xfiX3qPB9R9JH8AQ16Yh7iRQfe55vHuPtKXSkZLWWuO8Q7ClEDFBeiP1klY
hNC0bW/iUMuTUbqEtpfXE0wvHkTEDB+6NF+xZqPAaQW0n0+7lq9UxwkI/rpZALKy
Yp7wiRdQ4SEivuoZLDOfegTRtm4lSfUFgtb3ekDbae0f9IwKQXUYQFwZ/SDGwYTM
6wflsv7YuA4xTcGaeveU1rxu2iFXEDvojSwZYHA2DJedkd74nwHTU/iJ8tQio+F0
PPVQirx7yBQlleGs56+GMZCf8UuZX3g8IYOHPpHdjHA2cS9OWpk1p2oLXFF/jYpG
qlw7HdlPLJsPOeXVAi83yuchS3XdcmNoKm4Sgg3nrfqi0HpBPwO8NHd6Q+leUqtX
QhHSl8VWNqy0xqHAOb94vfRRD/tML0azEwn19Ily/StBWxj25TnEB9vYxnAXwZ3l
jycdj0ZVnMuHUzm5iMh6VBZ+fAtg36oijPvEGmJVg0qFXLNnDT+i2if8lgAlxpYb
lr6JxfqywZocX9v7ZwIEZKBSxz5ESIlGB6mkk4cXH6n/WbhNPyv+dKEe+SkvYDiq
AP6IyMtE2EnwU7VqbUz1vuqs1VzRNR5G8XxRl2titbmehCEBodIf3X++jY768Uso
ijfaB6ku0UflLyeB+wS7EN1yS1rlqExsk7Vp0I/nlocqkhFUUARbK1GsfTiCTMYP
wxRoNtSGa+kYtsJZXQFVboVecee4w35Vud/UzJgkNyrnDCduCCAIn0h34FYRrL0Z
Hud8sN8lq5zZCyTadkro3Sp49bSpK5vPsx5d2WeMbDEv5LeLHVpS8CG1meEcrWVQ
TPhdBuxM5OeNbSufjo08n/GaTkd72LM3KO5qgXm46+1dwPnYf4O6U6BOoVHblBRh
ZT8FPs7T1vvpQTOJOFUEHnkWrI3oN+WAK3QVFRsK3vQk+qNUPiesO7MIqaEKiNic
Fta92JgF/rnjrZwsWbeO6MBMK2CF2UAhGiSXfflMBJ9q0ZMdvK2hV3+Tr1eaaZZ1
bdV7Jr+8XiDawTWbkgzhbvnIxFA720VSVJPdqHWZLczMYhUCXrJ25MmW6NOeDBfb
SzwAzaHI19NFAXnQFWlYTqhzcGAF9NKPm07j8vCfzLOxF76U7t/ZzSAtZmx6sC17
DhcIlpUuJQQtsKmy5BX+jMD1D+yeRfzqiX3JYBliJvmUuSYZGqoX0SUOBQSCJbEe
uYWQl37jufLKvdFyLGSTd61BHPNormTkUbbzym+eGO6YAV1jlF0bRkBs0F2UtJfI
KFyAKwDFY8R4EyVk3nUv2IyRBZsiZ/1RqsEqYV7yNQmD5jnihgsnwHgFkP7c+dDv
cFXme0ba3PlG65KXAgGKExz1Z35b4RfdIb4S0rlLPl0VZxg4Fxm07YYCSjs02Rx4
yQD30fJfv9ygBL1/UlM1kXvZfB+0G7Ai9493GMg5IuA51y38fpAlouC8QOMb59iC
mxPU8UZNLenAxrQIfnGH/A6QqCT79gRAD54Mji1FHIr6aW9jGyu4Jw+rWTRwsEQC
pnT0XadBR/JkQhbCmGasptjN/2AG0riHU2z4Xy6kjOAesgbtDnv2KgnCaiF9IG4J
T5uVdV1oGfXJox1bJDpnpifNqFU5m2bh3/xmzeinqSMxWST8jCRMUsyYRUZ3oAfx
7+t+GMrq2wFhnHzGj9rophTbgHDNyvUFKeyzkumTMPj8SDj1SgFeVhYoHG0wQAM0
y5lBKmTlQgrMTKUqrnW6MsApZVjlKsAXXmldkVWXjORJ6X437DqkRntD12l57XT5
12An1MoFvXNCXOSSxG0JBcRgq7DDL8a1HLmtBBtDmikqIGkdFDLEFZ1EMhOfN3OU
lbioygpYipW5cby1ebfQoZXNTosR74giEl11kd8IoYlUdWXlIBovhfKTMVMgWd8N
zC7OJDCNXrAjKNoMT40CslYYaH/vqy1yP7+2KR2Yk9RbHLVYkvtANqWz2RerzjmX
JuaUbWx9yhIS3VGP5V3yZNJuNPdzeYCOhGzzYz9xSAy7n2YLQ/KiftZzvzLMAoR3
jXhiDLGKZ8JRDHsz1YuG4o7bwhFGfIU+L/qnfQdNxqP4/TVp9QvHKudGHTGxJMuv
H/3wIcvqPwcmTI7xkRh7B16urXsNH+Vrju8XXBAev7uJPgFT+li5k5UxRCUEw4zM
pouIxNK/Y0lj88tcPEmMzCXl6d0kNwA+renMHGSGcGD5yEWiV/SHf6RGUh5Bqwwk
ReYBA7Q6Ygrx2F5u1jF0sBlvhnQNi5+svxxgZcIarv18SbOhFzZ25vX9ehs9mBXi
SAAAGrV8Ea/VDSnP0dU+EMNZkNZKZNaUxqOG62aYEqcMwAkvcNs64CL4O3ctVDju
fC/hbS/35XPaG2Tq+CWuQQyVsab0We4BvRLZrIFQkO3n53u1YMHquangjY0VAhWR
ds7M2JMcQH0kIk0lXhWTBEEfXB8dUZflR3axTqWyljuW2MzIL86yQ+6z7RFieu9F
dkzkx8jru9n9p/3PZQIQRhmoF2nyVU48XBQFr65RaLM/sDEQt7uQ/2vA0uNdtav1
0bZx3onjUfeq0NSTMldfHWYhgrZhAwMkCg2yUB5Lx1k2pEY0NGwggVE1+EmSgrZ2
obmw8H7k5pTmlKH7KYyIiUcQ5I68HrBJ41FlzJVutpoYeU+mKJ7ZfPA9LIPFFqUm
sMQ/180UUeEAEiBRAWEA6ekxPwTzp00sy5s0tsXUA9Bf6ZfNHVLsCU7yzG7bzbjs
GrBMk8LtnuwbqdcO9tYvDCXCo3+b00WnNeUMiENVT1B/G7vZ9Pn5+MHcloA3iMFz
NX2NhSuvDDtK6Nn+VCpRVl6ezZwz4SRugQqEBwloXrXy06pwm6Nm9w7MF28cKYfg
+9nS48nJKXTS7bPv7xmAebYeXeds2B6Pt/uSt8XxFcIVo+EUiPUX6gtGHncCWJtH
FpunG8OOKlQT1365hou8ORaAOxkV88P99VjTbT8U8bzq69faJj5RR9QR4/9bLoKK
OoU5KtgfnciE5aGcOGsVblurk3aNwgKaKpNDW9UIduGQx8RM1rmX5yYzXuENm6mZ
8y1/vgZ6pcoD47pTqWdsZW9LfSI7vvRIRW5N+XSbsOak+JCcNDhrYye5SJ3GG0tu
0vPwG8x9CZKOiWB3pxSS3Qeff7wo6uyNPQ9KzxWe+hNL5ScI+3ghhgF3ckSWyHtV
05DJTrQc4QXJKLf9T8IDf8rJv5+g9Ewp5Q3X7il9nwPHJlVIRRcxQknCTyG6tzSt
8WRprWevvC2kLIuc0xDf1hAdKca40wERYCgA6THk9BOdbpZBCuGF/O7/DdUhYHUc
tQMnQLFu+rBJFNo5tbDi8iVWPhNHDwuUg5irfxVU8FdtOEqBA6mV4hYeWSadRLJ8
KHt9iY5sbh2yfIz4InLyQ8P0HkWKidkdUWuxck926qG3mLbqFfI0ugJMXdXp3gJs
NelYxO3NubKb9qntJ85LBb+9sWlhZpvTvL3xrA+H6qHtkjc0chLSIu/XsSMshkgc
wOpge+EW1xHjZ0y95KZDoDf9oQILJQKrba5YsE7P+S/FJ7hJPOclVk7u3LonSHLK
K/6iv1SFCCrxvjohizQ+50t6WLpC8KvMlIvmbzJxC8vPB8cT0DweU1u3qcqvMR2D
MuDDbZqWOPz41oDJe3FhCAYVYZAFMrRjNY9ItbUfsmBXXO3uaMk4lpCUadQNLPIT
U2klN85HWbN08opbzCx8W+wRZH/2/gWoQW5jwsNoEsl/g6WvISKQfxH5cYBOM71A
QnkF6Z5VK507x9qI0taeXfDM3GH+OVzcoB1AbVgXaWu3bLPFqZoAaPwwq2BnavdQ
mmIPMe+ERPAPHUXL5c12gXMMT/zVAZ68g6LUDMzrDGYaZl9KHT0qXtn2VG2LMnKp
qOlnZuI1JaiH4jCuZ22ieF0OUtS46+EYjCI5dLpLQu26CEW3vX80pcm0Fuej827L
LQEIgmNUMEVaCpBvNGK59Ga+dxgFaDoFP2mT/O/hxFGL7VweVMU9wDshw32W2vPg
Vrhxjjw5HTx52rZH5TEip0L4zRVN+NKyvbA+eQSyr+Ej718aaOZKaZVM5rwGi0CS
A4J433WVbuP0g7g4TbFcsYF6Z/eEiJEWcLzDPiRhScoxSfG92VCR/ATcDK4nDmik
dlTrG+DWknK2rHMYzB0FXd6o63yGj6CWIlRTS5OK9ctYu9HijfkubGhsSzC2Fw1h
FrI4qfnvkh0fIHACxuZjexuIkZJDAHhiYxFRohyOBqbpNhd23g7LKqTrksKuP6tz
jQMX/Lw+Cwznb/YOFCnXIQOrwHLhTgdZOY7KevSk87sYL9UokbXBoRifhGcUIGqF
LgI4zmUflA1DStbzoVnTgWlWl7nBHfrUgqaSZOkx2C894ujXD0mJY4aS0uOT8xsL
oOpvJC93RlrUTZtxQYqRbfhR+1KxDW7tlmZbkO/Tlz2o8cE3kTr4RIyCCaLb3egg
SAvTTpTFRDUGAODPNiBaDVm8OxXz889LgAh6lBLQuHtt1LMC3uw6vwQiyNjpaosG
SAN2oXlrgt6pBNpw7+y9j11iDzE0pDGHKsCOtz+7BK/tYE155lRbNdfVOyc0zNrZ
NQ+nstGMwzrnZebdam/S0Ah8EOa3TbXl/gao04f8EqzUhlO5NVIu7gFqFf1lK7P6
yQ/EYi1OJPpuR5T3Ka2/+D57ppa84zndr9+88Er21KoowaOCZtO7Eqy0YiKUqoMo
CDs9p6mIJ+GWPdCre+G5N1LEkE0Xqxx7LzdQ9LFB2py+cT2DIUn8qKV43nwTt5MY
HLMCiWy1h7V5WJ/oLjKrVOxUb/2ABvehuTu26UGLLo/jn1Is3YN73yqDWN54CaJG
NolEwTi67cx9oSUdiVodfLQ+jYzhTlDYU96cZfkw/We5D2oQ5h45hhqaMky73K8K
jcljVxXLs7VdqnZDMJ73U2mnvC6zN6WDcoEqBhk4qbqRdEN6/NGEfuZf2LTMeH1+
ddn39coQEL1bRp25e31/f3bHmD+L3efhzyNosdFqhLCPRZ+oMxET/gncnM419U38
4LIeFysbDHn01yA3vv9leYUTGUCt6q2JBUg23uC79FR2kGcOa6jAFxcf3Yj9J3IL
lzd0e5qZsYV3ehnOXSiv5k3VsfzR2TRNFZ6DxC39+I3axN9+HC3q4P+DqMnxxk90
qfNPkJ7t3R+1A6ZDVIcoNsWZgE+U8UKLDTf6An5VYlUZcoy65GQr3Mp2c2MyYC+p
N3ripbWSLcPTt9xK441Q0xuk26VmyldgOVEbl6lEEsIVYNrqyCrbB5zHJqQ8+CZL
WwQqoFjr3dA92k8j2x8PcekkcjuLBKjXYzr0lN//gcJbp0P5Uglh4TNs5+fYwzft
ULZMqMxkGQSrW1QlKfIWBVzV3aIyvXDaFEDOTh40pq5TnuzJF7dVaoCNVpqxEsnd
GRLRiCe4e1dNijK5M7/kbr+076imd0itb0gtNY3M1PQnygIMLVBqJakBeYGrOnXw
tUnPRVP1ZX1vlQMuZ3Ng9lLTjuJuEZW3D2KGYZTJFo9cUU0iAa9ET48VVw3LTNj9
iXP8iitUIt0FcoYLZWEncU2TS1aNYYQxN81Khkl/yCqRdCMxq4Sp8kRNayQ6THsb
NU1zRHMfaL2x8A8CftUpcpXARuf4rXNoXgOLXND2zYa1CMMDIKWorxVcOYKnkl2d
nbqB+ZHnniaGVbKpDmB+sA9TeMv56Ift7Uh+1q3GtYZROdUCb1gcNmbQ+UL/TUGp
alwEL38DPvEZ60qgQ/87goFBNhhE0UmfDlt71t8kb3yrsQmG58n9fopGOAZgj/DU
6RmY5BVQ9UQ61s5O32stUbeX2yH48ZNmkypsPdRzMDdMwOllROWs5sfzDNWVw7uB
posV2N+AjWIT8bzk5MEZakf3HynalycXItHcEo9vnhV1Kcj84odMHWD0OgkQFywN
DqGmKa+Fa60btsV+VZJNyJzaigawPQCitFYd7Qdq2Vje6laJ3JHG16t1TIuEW5Lc
xZuzdetwjVpCx+HVa56d16y/f4m8WRgUzWGHCUrjxbcw/lJ1n39d0sBOuP8HLcsw
hwFbx8nU9gozyw7S2pDpgb+1AiFscqeT8qITp3thwILl6Dh4mmwS5L3vn9nbbugp
fZ9Z1nvqBItknq3o2A5mcRFyz1YdakJac3tQ0GDHCw3LDxFtnXoOfH0RGjVFNT4x
dVgRaCVnyxPKuoCajheDVLpKyNzS6Dz6AwnS0+/8Z9mAk8B0A4DCruLIF3ufbR7Z
56aQ3dlEmvsvoUEB3WBK19yPbaEfJysCDQKjowc4mwaVArGR69eKyFeZzymSCh1X
8/eE65s11NcvpOCm0Rs7l4OXBwuUl9KOFtIk7bbFQ4gMgu6lplI+Mrh00O1cInkZ
/eJT7g2XWfzKQUMYD02SvvNyicGxpbJhxN9LrwUShMdcFA25t/1RYPb7xU8LssxR
CCNtHU3brHDugyDWD8evcStXZUnjCs4r059Q7oEdJ4961rYVxMsrpF4Gjku050KS
aunDPnbd6L2ufirxhUW+q+XrBD4e/ZnX+aIgzE2R3FG9HGtoP36fLzJH0ffmKyWg
vM1B330xyNciQXRr5vmY3StkqaogppH047nz6RMM7N+8kfQRoPdSxt43N+NUaFTr
Xiiwp9ReCdD/OoZxFZlUbEL0Y1H2zo1Znyb6gPo+GiXOsXt8MSHSsYh0OhxTgHzm
/665DjcxPmNdVHIazCbPgNFL36083dmRPyiYR+j7ngnxer0K+TUtQWB+EJfvD9aF
2mOuCgdoFVbYbXh3IRewfMRMRytkGKHQGynsHjB53ITJ8OBN46ZvAAce2HjqkrKl
CzM68SWVzsfWBX8BKPn7D10ERC0qBSuVk6JXaEuQb3oMXtnxKkk4xvW+dSn4lS9u
P2km+i8RUOUFca+t6p2leLVMWJ1OIAC2et1ef9cNOGvyAefD5juIRUVEMqsel7cs
Bi+3UOuJvRqwwUvcC5fTe+QZ6WGr0cLVc36F4xGgI+TUmaU6FlA9iiWfmz/Sp6r7
cPPBL6nFZRAzgnuFX1TAFfB4PH5/Ab180hxgr8HgYZkzhZo+c+6e7Jk0XnMl6aaU
Pq9+kqDKRxba+f6fv96EtLjRgwlD5IFlRdHnHaDZr3BfRZHrEhKLk+k9bGwbdiId
sTWr6oFzyRJBO9uc9Yir6cR5PE3/jChnAAMBoXcHi14VSVAYl0pQ+YUS8PEappIw
Ad5fmPCFZ8SgUWF7+RqyhXtAX7xRUeLyIUu7w8iCsrjmGevgOP+G38XuuWN9P/0d
kYqyOcePVeIj6cb6LhlSvnjZVMOEih/fqXSc26XFJjvsIC6rTXJKS3rDKDfxIuu2
3llAYbqiE8MY/tiwjtSe9apw4AsoFQ0DSHvZzgDR3GJpLjc7Kx319BtqJyQOziE8
j0RBzBimNg/9/zsOTMMkjTkffJr8nh43vD6wCO1w9zhmVPV4DwijxRDz1MIE+/LY
r0nUF+vSqQF/zj0BAO8GPexqz+ExmJp++edvlExQ0pmFu2+O3JgNdg6RafUpgGR6
btiNLmvv+hyMXeHwJITKGHg9mAou1deHoO9i6k5t8aznINPzXlLEqIGtGh9cm3pP
BrnzaoVdfWFb/cSqmeUjvUYhVnWUB04mzTr4eKm5vbZ5NIH2ymrrowDSDDUZf+/O
Z3/S2Lk6pKkczKUYMQeXWlTppc1vtkJpHnvU3yp85xh1G6fiAEYTVpsoNM8sAesW
l4RLQLKx/mDM9PlRqj15tULifExYI7VzNLcJCPKdUgTsecTS7fgJZZBcSJki67fB
o0+C1i47ERs1mgQudVv9C78PVG0vFqB0yjRghYA8DjXXCU8bwNZQrxAJXPnNk65j
7RpcMzi4seCfHWD4nmOlHIJ5JE3UJBKEQ/Fky47gXDcZi2XhjsmAskx01PEey/AJ
LoLzzdCX1yPAqWmpin4Wl0kPwl/cWtbaAi36rfXD/c87jjOG9+7yf7y8jMhwLYw8
PjZFcBCWYDhwY9hVPwne2/B3171x6mQsztYRVLhmGcdf0dsWbAU0GqtpAer9TG7y
RA71ry6jGstc7DxDdgjgCmtAFdR/NEFcy1eeoXt8ImPKi0cmXpTwMOjPdSyff+QH
ncVda0tDH49jlg7luBpUtzQU2oxgnsWWlMLhg9D/KO01l084Pe7e9MYbPUwc7aXb
zo1Zu7MsYp1mzdNEDQ12GBIki7uWgpGnt9zPGWOG20Bzo5+h+XDkfc9hcduF2E8Z
C08K2h0Cy402rCfpaVt94sr+Hofodnaq82raYTL1liWHnLWF92HFbcg9u5c5X3ZJ
iu/kjH5gZOdXowCRhlKx+uYB/xvjSIE80TCBy6SJmG5o5zHiR760eqQpe3GhLTgP
tDMVgSfiU6J4iJM35ssKNDfNqAmeG0vKaY9AB2MnftvFXz/i0yIky2Qf2lQZv/21
GNMWf1FO/Cy/2oa0TjjMI+15AhL6kAnE90ze7yU0UfzueidXr0rnCrs4gekbulpO
z/0wuDOffKU+7viSRMs1q51nktS+Nl6zoPnqZTFsAYx0i+ZK8wf7LNGple/KZ7Rl
3GLlFyD0Mk83AkD2QhUtphD9XR5nbJx62edAJDM/oEYmCjKifvoBk7F1LM3fWPsb
39zXTVGsoa9wu+pZYwkw1NcJ91GYF8jrPqJTk/+ULiExPr/k5ScRNSYfyKD/Jicc
Qfg1nflA8qRNxDqz6dbFOI1DAy8eMw7WipjuJwku6llsujcf5YBp58JXzAoRKMwr
6iI1/4AY05YgJdkG9UXRZjqsLlpq41/1F/jv7q3tYxnanVTarcUyNOCmEIkhrDPa
ZIdN7pjECjlEIT/ihDvmKhqqUp8CYPaJ+/Z5ttAH1EJO7XgkC6+jObsHG+LrXwgP
PUjhPfAhaxAKWOloqjHSC0IZzfzjxuBuxgkzUJsZT1hJxrC2DxS6UoTLILwWziRe
x0CtzaIVXkWc0pXRag/DxFyQOFPpv5p+4qXNB69oZoez0jl9JIaymu3opugqTBDW
dTP2XTPdnfSIQGeYbTd9p+BnRBhcK9L3FExGR5gzDXDe3H6wcWNXisNZ5xKeylye
JaEhn5gUGnCIOBigBmbnGT7XeG/GihF3Jr2p4hgkUZpfY5hT0HLmjHrUot8GVKOP
RzExnN6Hlb9bZjsTuJ4kCyeYk5+IkUpuJps01qGFtiqCn0P/TfBjt8UfYdG+/XiK
58RM3P39HPMqvtDgP6rADoRBWQt9QXsetr9p0EKxrSDXFGEU6BGlmbnoTkgsxak5
TKupno9fP+Ok1Q3j0UKrWzYXxRNTQgvY5zeZfMu8rHbB9/CgHs+WXcxCLGis5mtB
v4lxDmgsxae+py2HSSw1j+nzxsEbovOOly+sPv5rRcapyIpnqGTULpGwxmzzRo1T
gho+t5QiDsDa7elcIBh4szFlmFa9MHemRgkixiKZQuUr03RX4stj7lTE7foinUCn
28IVMRTdOcrGDmCAoBi67Gv3JF8yO9ffWXyOHBMQb4p9MvvJu4tDRy4LC/q6lxK8
asv6PDmouzrXmuJn3qNc9Jl0LgCP8PG2L9bUuxyn+4VwuowsGx3OwzRJrDOkax0+
qb7MEMiWBK6F48KNWP5d+62x+Vcl+X8oWBn3bxJ1ccoW/1Eh7E2LlOrSBzXx7GVs
vCY5S8mkdY6FfNqFl/33ZLxn7lLYkxF6pqkOJHjNCcQsKBmTlTt9d9uenhfxAJZE
s1Yll988Xb+bTivdTP/J09AAzewh0mF9Lu6bsc4WZa8CN0lOvNTRseWS9WN9G3sf
en0hWJQzO4R+U4oUzM8DxC6ViPXQdO6q9U+Slpxw2APLAywsp+CkdfwR5h6jXvcC
FkfPfyEgk++xMn4HVtbp+BUQvuY9hIWJN4ez5gO/jiAUH7nu2buon+UTtXTgMzUJ
fsxVQ3sliHGF+Yg4WGfqDeM5kUZ4vXBSsmpRea829c+fAYm2Im1eXaHlTz/SURgT
6SPpAVeQMY1i4Iq8aRSWFGwnUF/d/heVohp+n+AmEJS/FjWheqi/TmT69B5q0Tof
mLP8B4w1zwJNdoqNFDFRTEc6ZEM1nZPMMsnCo0KK/gjc04MsYVFInJ6kxhlj/ayc
ox6cOWuGbY0mpYYhJf1hQ2itLNWDe2IlFNAI2VDzTt/jM82bOuwVXKFW6xxi8VI7
wKiHR4ffj5F8PNexW8CfxRY9lFfl/WGDVsoYW0omljZqXneO9YEAINwN/2knXZUM
vWCJVVUpJb1YLJiyGEAvF0XA7/5r1bb6HYiZIrfUbn3z+lqRkA9lZKHkno1m0LHa
tl3Anec/uV3J+eFU4x+cWHBay50JFh1b1zyEEKOdMACDcPC+BgMXgyV2Ery1jVez
4uzbKzvOgXaiCRIKBatczeT1qucA2BcuAX501QdYIofrzkbZjpI1jGGKePJNqguh
8giDgab2OSBpfeL+QkHfdzUCaqrVV6tRaf/XujDLaWnKKih/J5ZnwKLN41j50i71
CsN2JTb0rcFwZweNMWAYHK5pDiUdKPcXSyvapDqzKX34jsDwNANVKVE5/gzYZKfz
yZl6YROmaqXw2u9OiVc4GxfovkZ5Eb572SXd2RT+aGkss2eSH4t7FBvLuRrvG2oG
y0SvERbfhY6f6ESatO7zSN8gYvDPnC3vlTPxb5N/bbDKp6PNsY4fDWORqlJcE8HP
AZe0WdC+kpysYakmS30Py9CHXOTmVorZcSPswp82RXkoeefpfHSL8gYApfoRtUZC
oNuxXHpRPqEdYl1RuxM4bZ9D7yzMU3Beg76TXAHEZ/YG1jW1n8LIoPCA0PALVmh+
r0mFdIACo9Dc6O39sHQC/Aj7yiYVDqydtJr/5fu5iik7OGLc+X2GJTe6/JqK7GKG
ePtPlvvckdVfrJHzjXceZDjgYcWXoaEEVZBktcoHzlJJZ4lHcpXngcu1/jcZQK8l
PvyAVg+sLvkVU0q4MBN9B+muaWYYcLH3i8qPe9ar8WC0wU4HpPxlXPGervC8IvPe
qdG5O1cu2i1cBqlJxyl21FDtqHaJgMe7UVtlYUE3lHyBnFog5u56RxSlZWJceuXg
w7r2NPvywjczoEnHoKkdWsaMq+6P7NldlACbF7PsZFKWOtU0R9O4qx+PI9SZyr/w
GWyXxUVnkLDVAFB1nLeQrs3j6MrHjX1Ka4HBeNcIUyJG+sXTvmXpfZJbtmluSo9i
bOrBTC6arSkuvhmLFAbI3mAUWC6kbZK7knP2b1Omm+e/CLhGkBJquQSP+TnFgBfC
nVfZqx3qOb6t3nzXnUsYhVC1TfFC/Z07n6pZcaKXzX/tN4sQFswqYJZ+lodWnkkp
lx3JIdYlHgiTpAMvrVpQRjQekB3gn27YHlx+2H3oXoLwg7OcAlacSdOLiuESlmdf
DYDOVAipYBdIwI4S3s8KTAkBeRRUi+Ek4boPdDEjnz2EFaHvWnISGuoLkYPS7YaU
wKxabVgNR9XLx/qIw7syupttC123lMnhTGiTj2VJ3YkYyyvfbWWBsNb5nrYcl8MI
EOsRLpCrt/QXjy9QFB9tNKYMPoU0qeWAYwXrvtJlCo4LH3+kWbjgPhrNxTv8GR2k
TFIv+eDdvI1k1oaofdZa9qHVVbJImvBeZ4iR+y3g/PGZZp3P20+aBGG04BQ74Q2c
7Bu839hR468hzQyO2VKK/5xF21IvzLT2en0789bpRVndbUBdry1/B75TpMpX9ptK
dK/78p/J0fCp/Ck4Tcm5tozu9mviWra8UuDRyA91+ZI52P7I0rfimSDeurX2p4i1
LddmA4Lg5NW1GnoJOSxTTYIaqNYFq5rYB2ougdOxTqHlhmvYrdWZgvkvMYk8eYnU
z8cQ1QMrmylVib1yzRKkHtGyFeeO42IlVhaCxmVP/0LtZXPx10bIJpVZ9S9Iaa0e
RFY3yfio5yTEcEmU1oUDLyIs+NaAi05uxOrOE+whaOPXz2qs7tZILlDXp3zUQN5f
9cJopN/cBMWXJUlEPXB7OaIpAJeF3NcWgIGkZ0kx559QjYTGBCYzViRD0KIP71co
s8RiS/OyMs8CIhCCwnsyJVV0YgsPZw1tIF/ZIXUDPy/OzZwAeXqzNYfhjnexX0CP
360GwBPSo+dPR1NvzFaxPxLdKDQ3dtZYFeqS06ZcGbZoUux/bJH4ldfCHZHaE1cI
WShRxf/xZnaSZAoXE+l8KHVFYT83hMD7BjC7r/UQthGpJbCBk9lO3TjneAhiWXf8
DflSEnO3sBz6rB4PykdxtgBoeKNECesDfMRWXPDaZQ8TICf243p27tsy+5KGqIr1
xedNV4RZDPvndPsIPRxX7wN9NBSmyUkOYRKUzlcNyu30FDOSn6jI+WB6wkk5GoZ2
jVqlLQYT9yTM4uj2y5khZbOojimNtHmW+pVyC/vNWMC/BI7B96SFrXCiTxmuh+zo
6mz7FaTAoJ7bwJv1/hkYPn8qDMdvqM4EZmcytH5LiQGkj/Ke2OU4aK7zF0MRy8tn
Vts/dUCmipnNpixQHN6JuBBjPIGEVncMjfRpKErVjrcA94eLeyLkbkRFqi03kP8J
KmenANBSRzJni9zb7ATjLURU5AmG/KkvqC2vJDeObGKKPqGQd1X9kPLP1Efe/Vvw
ranpzWrbZU/7Yw2dFqn4ws9qdV7bGzNdgel/93VZehfnct1SMdJwtebLStv5nkQO
teXxYJlqevShIqrHLSx4GX9+W0az8Zj2Luu0+XH4bV5zac70MdingjZKP9tp9a0m
l4gVRTG+eZGpyMKodjgh4mVf0XeyKijgD2OkyJWvpli8M4PIzeLIjZlxi5IPpphh
dAZpjHXSBlRH1RGPtmP5lXzlV9bNW93A/5O7eXNMeshW07WBKX+SugOy7GcfgJN5
gJmLtKjPeked5udRAr4mQ9vCrdQ66CGmJcs3jKiFy3FUCA9Jlxnxaj3AwzZkaeBT
9pEpAFjfl+j/wPr3ZoInuYPfdLKG5ly3iFme11B3hb6LWPs99NSNEHtK9BgxtQT/
m+t9Js2DMuJqG4kXc9SBCwLHkkQAW0zDtlrzcmSHVjDRUFmAKYSY4qqjROXZdMFE
1ciKQ0HTZeKRWxSctzKLExi6J+lZi8q2I3r5EGudfVn6904zrx+cf6TQF2xMxboi
/iDOvD2z94+XPhSuDM5O4dCRPsSfpqmqBfSu3UzH5TK9avXcOIjJDEgstC3nTNjA
UigjPVTuqTKV1Vm35CPMnY9hpGaG/p3vbhTxKJ4FCn6/g851gwFwbi05c1bJp5cs
4qLtn0E0RRBeAbefjYqCV2Dw8wgSu1Vo8NPvuP1gxHGEDzsAoiQQlaQrDvfcF3fR
3nPn5ED9DBdJh4yqi7q5F8n9PCtQf8HuFHkBO46xEkyVjcs+xVtobmUzBDj9mNGG
porKGt1mue4BHtH+KaqkNiqPYCNj898oABWz2Lm8+/RUd5labBqx4HuEjBgldn0B
ONdFXSHnPUSZ0iypIqMjjD9i7uORtAWIuuqEuPUv3G7VTR2THKZ0ul2R/22G/5s6
+XPkwTFOnq41AB2OKYX+oDTZYauK4ISLP2asqZfepmU85iu4LoI+p/Lia9eW1Fb5
Uu49rdYFAleDXr1FyJnudnQWO64lQnhcFMs3l3oO5zDZuV/O1PSyGigdm2Ifi4IC
/kRu7kQP+cgXOYNKEw0tIeDf5yitjWI37499vnFu1oklMV398WSGxZBvZmUeN2FW
42G6ZOgDsRwDG+YSvtLj6LUyiYbf7ZVpISFph9tHWW1IXcpa9P2Txt/jvKuGmEGj
cyDGJk7U9FtxkxXDOzVIp8STe879Mnmq21s7+er6ErDi6XmbuCLCAyxpA+xcgjWW
nKZ+ZeJMel1HqhdHB1T5ysR/NIurJ8pgIFY96TGXLJ7qKs3H/PKfvWhErpjqsKeE
EDKaMdYSmVGxHx+MaK8y9hALrxbwzKKF1k+HhtyuwCtJg3jx3sY9cvKl4QTVtyv/
PCpyaCX6haNTpl1CGKlUbiLe2RVBZmGQHA4xLFpZ/WbkCRCtqHguC2S97jhjkUOV
b2aZ7CMdJqU91k6VR9Plv+3wxUGHqIhm42UxXs0OuJ6vI9TcitEUXcBu9RD6PSAG
VnrFRBgEN72A6ZarzNAciEILUAFpz7amO1vu8CVwXAv6vRI7rBpiH6QpA0z0QKA8
CunS9HaSaFc4+JcZ2dQ6szEdEKwcR9fcM4tkS7EBpn3O6hyRx+10mfO+Ra9NvBs8
EQQEchiO7c4/SJm7/K7RjTSmJBFr1BOT8+0mLUbLM81m0HCpztjIZZzjnSXY7Bjf
3Rv6rayH3DrWc5BnCXqWWBv/a7NPgy+ASau8sedeYyrzhMLw5DiP72zPpNIFhSoR
iT2kLkd1UkR81arv9oBctic1UP1Ecu5JQFfAeHIGuicsOO7ScPCP2W2EANWVZ5Y6
Kge26BzjbrvzTPhp63WMRUKf3DJ5aLrYM7ZD0LtVCaQ4JZ5ujpX4ufDf8BYIgEeF
Jehrbm/ba9OLOz6+3UW0Ch6yNlYAkELFjEPLTz2n9c9FasPlRIBbXVse/JxHDwc/
oywrSP3iIIPzE97unnFYCLPFNlCnLIo3g7Naq38Y+bzXkv9fQNSxPVD8Anr1HHr+
/IPrclBQtlDTOA66W3q4Bjla61ENHO/rj5YX/mXqB3Xh+l1rQ5VuXWE5CsmlUGID
hkYgCOOug5H+fGNc88uy/aRgjogQIpfnzIvDaCE0eNrH2TcBgpUG5yLGk+iaNsV3
wMCcMuI7kU2sHwm+NfZVwsF2UzVZWurpmYCq+tIeTr2i86ihvbyBWo9FcMaHCyoO
tdnubNIVuxDRM17x2Z7jVZTSA8QcoWdZLFRffn9wRtX8j6aUcodsY4/becPHzXKC
teuFdzPIrNR9Ioa5KPn3q2JsfiaQoTRBzDczOrhG28CP5dUsWzQopOB86r2MNSoV
zYJe8x1Ndywr9V7zVRYca4ELMJ/yh9Ala02AB/+CbMrcPWgIR+7LsmytI5cS8MQS
tde0xXzZRF2hCM5scRq3Md5IVKNvkZxToHNDXBK1EPamKry0nqiZjI6z2hiaGBYt
dh+AI8p7Bb2m4J/6V6gwUyMHE1xl/AVdKFP1zrw7KF0U9f1OuP9MhVDXIg3CJuKN
qL9xSZ6/r1IMB+NViOD3lDI67xyQtunlZbV6X2DvT+/0ZI8frUOL+XtDskfk3WWz
PL8ljSrMa5szKFzc0gF8EIDeKGzf/ZAKdJPzmASqNEzsg069PcUhTWlM2BLrwKe7
/hc3xbA9lqTtgI4XIFa29QTzPR42L8W6jKyLrQrDHx4DBe0HqtrOgynV5Ve7WbtN
+p22rnAJHLELnnLOVxpXY3T933gpAdkHIzi2zaKCwpVNbNq63OAy4wCxjeUQ1arN
Z9hHIGr+4A7wsZALUSosGBKrVDPliUjCaF0Ma3sK8xk7NndCGpVfAgV6LioJ0B/r
ovEmz5SFBYgeUBmtZ0aV18YGUbnEhGikipvoAfbMfpP5zMD8LSIQG47tTKxudRrx
PHDeDnJRTIpn2eoHfGWdJKBnvHmxcFul/HOBajMG7GORJujKowr+zsDfda07imYs
2YZMwyJWgj+matqNRwmsjgK9ZmCOL7n0NHRwGAuzkhz9Utl+i7Yob921WwCFPYkP
4d7tBJAdswscm7QGlRqxDJL20d26mNQKKn461o9tciSWd1ZYaKMmk5GaOi0FNzTs
xmE7E0wUK6/Ui6jK/UE3LM3CNUno6hR88S+zudJuZJrPJyf1GH5f6HrnzTZ8PcgD
mVt14X6ZzB7ddi84pBOjmJXo09LI5f9wr06Izhpi4Z5KJpZjjlhgrDve4lprEuJV
DgqF7IlnIaEbUFW45/ghlwxa4mfjNqHVvK5sBQYWo30y2sMCOanMwWxtxX/t1bLn
wd6iGo2K33ULef7IlMhozIuRJPcj5yICiSd8h4iTRqU3aAy/X3n/quLVhAF+y9fB
I1+koWfCsPEe7tiTgtwHs4kkxVuP8lJI+G/JGW6RWSSW4LSLPSVbFSPymL0OfhRC
fw5oO5X6JmBn9mVvejOdaFpw527Qx/hrAhXLDrqOc+owYbX1Es+5zpcAbmrKr5DO
PlWX2x/Rmae/KmC40l9n8LflzdJJJsp28PAuTH/sTxipluiWmfQAF/jcQNZMuBQ3
jVgXUZz6GY/7QBCYxP1nWiQLWHrN1STlmM1rl6kPJKsHVESgK/DxlwGTUceDRMRo
xTCneVI/F8Lv9wlkGOdjTfiWofa6uAyX+9yiKCKn2LtP58urpaM9XlDsjvQe1j1i
9Iv77n2KvD3MXB8sAAfJLxDuH1KclFOPpl+uVLaALtJOZQaGvMg2JCV1Os6fEgdY
uX04mNlDQ2KpiDPeha/Njzi9UIrH8Z6kpQXy4ROJvHPdvM4NKn2hPRH76qhq3VVy
EfJqPtzYHmWgS427K9AwryfuKH/Kmg6DNNvz6SIETR0TjUqguoWpVcTa+IAcn+DA
k3ExKGQUeN9VafnouBZ1UCYfjLiXfb4MGuuS7Jn5rBrKl5tMyKLbEefCGpmSZw11
iLF+OoruRQXPD2D+A+Zo6UPSURgmE1pz53E9+nf3RrKGB7VEFQV4Enw8r7WtC6Ev
L4WlFN5mEV3HV6tkcdZlUH4uiQl3qILFqQzUMJQbjKx+7zDfIHQcET3Eu4CEQQ5v
mSCZvB2fbdL64j5th+iefJIXCirtTi45h1I9n5T1c2w6kmJSdpn//3zub8aCt/pb
seJ30J7uXswIvi7Rnv9Kbxs2kcUbBTYedVW6jZMC0Qs6gjjKfe+OHJsL5aBqAgt9
rizjmMNQdIzE8/e+Y9182znMnaSRgT6plOklXpXaa2MIK9boApcRd0yN91F+LRaP
62yUNfBl973DlIK9cqIk3AA2VIWeP5ZpMvJgCVwA5I5OCjPQiporjbzWMbFy/NM2
ltd4lIgu78QukeeDkZTRM6QQgTMnLJRDDguD3m/+dj2vg9nRnmwT2OSocHZX8n2W
+rPhy2nXICUuPveHRRr7A/3qM1b4Z1NkaXpQf/Fs2IgP+34MSyyvW7V53PZiIh/v
o80bT9tJPL6m7qE27MesOag4Ynux4t/rJoDrrExHCz23c2WZLVxZbjznwU9YB2e9
X7IbvUot2kQbtKKlklnUKDu/j3Q5oEeF21GLIN/dycvSQtWn7AXPVBmzZ20XNfub
NrPJhscktDNd0CVswgG4HWI2pN3fJyicQrYbAwdbuhmaOgcq89W9bCT5FF490AJt
/VrjAsDgAZuj/GG5gMlmNHpydtqHJM09GmIyounZ3yRIqmwItRuKnn/xtsX5IrBg
lnYgyXV23YoNY2GF8xBkfvBFr4FRxfhlzXzuhlKRuWEjkYbxxenvztnkxi+r9s5z
sx5NG3Ip8rzKrkoXOlHxG5ofXYKX5lbayjedmCdG6KCx3gn6xXNSYRRD+2Oay0S8
sI4iN2oU3y8whFtdtjCpatlZpmDJ7AhF6mMj3fpqdSjgIR3R5NGxg4377HXcRK9o
TxY2z9tjIwvN5LrARP6VidTRKoJw9hKSh9dYw0OCRBMigUWD3ipohx9UwOW3/fkC
6g9NJQYQ5F8Q7I38rwyUQpReA/pu12OXElIXbnb3fTh5hJIe0Gj/XNNImCkkXS00
IHyDdLbCkq7olP7ujzZtMKIcrnD+Wx5OWUiMo1azlQV0rZRgC3tOUp917QdWpjnM
1XhI2TALDlCzunrrcD6CUvefBWoOmmkjnW4wOKUDmR309/NjpZ6pLZczbX+34NkD
eGG0dNGhTk+j1nzin7gln7TuShaR8k2F86sS9AikOZPzq8CFAwn0HlZGYncFnCPu
N7/CH65wsghANh5sAvUsE3y8DPX2opJyW3xaC6iAjUwC5j8ZyagiG6467SXm0s/b
i2iTHMuJlPYqKpROhVSwZFImd9rf//bsgdYKUmjIQ8GcD0PxsdZmTmuJEOPh1fW9
vvc2pYGlviCf+rLJTWpIrK5sW21ydYHMi46/j1rwiO1FmV8MJ1z1JyCIEobGJ7RJ
oXzusDib8jpMMuFspIdReD3n23I9SeIw7TDJIBOF3vUNAnsNDe2+0p66CiszcUJC
hspa3E9spkqmOS5o902GqjcMJx7zAE96zEYkWISM1hKBDij8/OtBwyT/RvttpMRf
xiQOakzBqOtPvpPk7LjU8lxBemFUGxZL8tW+PsabVR7cE09/XuRxiO3Ne4szIyme
Y/30BdmeVfm+yAzIaXN6Jtlm4sM0eoYeuRCbTfalzr56yhCdFiCGszUgf/0zMXCB
i/a6/g9npLmOSuvKdjaTjm+842+9G9WpZJF+ADo9gyhT7OtyAJqs9HpBa4/0nGW5
HJFqh+K4S28eV3RDN1MPNd2gPRYjW0ahKLq44bV+l9WwlYnCrTgFkIcKLEhCiQem
c4Y47cQiz0pQd08LkoQmBGct/5bMwgmYonohw7IkR/uYA/PQZMDGCroXg3qTiK3H
+AjLTw4mI9Wv2aLOqLnMDvQODhXyw8Ql16yn2FlRtsjzGo5+d/VcIycXxGRYarz5
ibGnNtGIMAxgWtuNXFlh65AnPbW7+uPip/OKrzumW24pWCHE6io1tk303q8omt2p
A/QHfD6Y3qQGlkATtPk7ttI7RCn/FA9AIp207KPkaxAsBrkLnjC9YjXFe83eXyVY
bzjZ1gbymfW4Bs+ADCH5nXOha5LqVdEo+h+4bW1IRWwKf/2wFEQgUGkexRy8RIPf
lZItVWSKX3gq1JveGNWFgzL9anU7kcnhvvIj+50DX/iFXdAqtoATTluwVsiDLWTY
9Pjsw6G4GHi8TPbhW/x7gh79iS3tHGuYlAT2sNOCuyRAV1NQ4ygScYLAXzAIcNWh
n4+gUl1evA3egVuiZZoDd1Z1T1kCemzd+1aBcPg66OE+9YL93C0VeIDeWfvIRywE
V6oENhB7EY/QNrOYWSLfgbivN21kcO/Ptjox5qz7mbcoyo1nXoZkKT1ttyEuBiBw
L/g+OeSp994AMTDkmQKGpJXwYo2PjuoZ1HiZer7t5LTK1ODnREMpcpIm+KMFJT/j
1Fx0YfGB/uoHpGM0Kqtcn6vBcSRDkTJxpbG2ZbUPkG8NV3nBHVIHXlktrhaY9MV6
/ik3Jptf5KrtsQ3OCM6t1h00KojfqTG4qQsr9Y4PZDnBYQGrUFmdi9sasmVwMZWL
k1n7+HNVd/qWd+Jm/oPjulp8j0DdMxvspU/b6j6dPVbbfsaJWpFcS3bfqy6RuGjW
BwqY4UT26aMRrsf1OrT5pr/atzKThT+QVK0fILWoUBrHx7L3hIghm4hxn0ZvvxAZ
wCAGM1s/NCtYgNR9FSKVinbGB5LFN0IqRyeL7J+2vVCSc/bbQzU2HAkBe3X7qb6+
DiUE4H6Ctfm9jZBGmo/uLp/Tq/Zjy+ElRv7sFGMnd6UbNhiUQTTfxKAvBJKZFIja
2xzMD4PUS4TVM7jUfDhVc7vx13iruEA8eAM3IlNfxC44D4LE56Am2QOBPnco+xTL
bvukA4m1RBUqNmQSQLms9drm2kxGxqtqccfzf0iNRuos+wdLlkuvu99xhDqJrQEo
Iupnu2k1Gq0wA4KXisUWTcEI6N2o6EyvN6yzm5wtYIOGtm4qbrnApyF44v5B56RW
icosMJaZ15uGJaLZW05HXWPnT5TDL+Yg1w84Eobo90YgKNa3FCuah3/IGG+/VblC
/wjzffTy1WD23aIGVCiW3pAjopZTiB2B0GZ0teBGywENhPM40rfsnMs3aFx2jXEA
P7hY4MnnQQ0CUjJSg2qcXX9ZSDxyBF3ZDhlNTXvPB3Ytlta4dEMdrZ/yxzl3rKqt
C79VP3bXdVsic2SdJx6DrBXl1UVPBwi8s9pSoYgzxVW0ifcBOKhlV2r9czab2us+
pcuBmqZJpTiTiGQIO+r17CpCwr7/isqTXBYbgWmnMTVMshG6ZPPKW7bQcHdSEu/y
/CHmkJuqMCsGjxY17kblwCXXkrE6V7VwFnCCSdcir5UnJddmIg+JKnXqhoQUmPTQ
8Cl11d4xfdEKEjBvADcgoM6b3PAJDoSrwQVc1KocrzcF4KMPMzTeXGIeQ3j3EXpV
sfVanUdwo5Wgmhhi5/EcEofHkTpNeBIBfdvvAGvsmHQTGUrgTebMtgqarqCjksJc
phsBKO+TSJQ3/Mnxcf5iwxb6ILNMD9ap7z8nPfgP+RiXEjmQGdsHMkORhdLjCSso
phyRPlYiIWK7uus3JpagDsClke+dr3I/jKnkLdpge9G7Z6jh2xCdgYVXX1r6lJtb
xNti4/HDqA4Q/lGMNNz3OxNEjfDDmFRkDLvbdI2PbySZNwCE1LIlnjtw6pJDRm2O
9Vx+KSlwKlYrKR9j5zBGHZNbGtL84mcedXJmYOuu4Q2kVzf+1ccKCzc8/RN8BYhL
QJBovINk4oOKvgfFW+bsoF0o6mTIJ6ovZssis4jm86ZgPyANvKsVCZaIngZOnnGK
inXezvWDxSNW8ksEqrYVho5N1hYYjFbSwQVJoOzJ2+Poyd1cO3j/TgbG0Dva33m5
Lhpe37GdO0UoK0DszAIymL9q0uQuNuiScEZG6743C/tvLL5lrZPrAH1gvJabqVZf
GyjxpvrAbC8KAMa6FUeDT/bNWfpwIpg2qjcL5nO8eBjg0lBLwRnk8hwPqm7Pu68U
wxoIrdvlqpQReWU67dYyNAyLrhffZhhNu619g9HncBh3netSzgD/A3axTEwyixhq
jWxV3LNrTZnxIRv3MbqAEtzbXcGMVWPAgRwzufcyiy4GgMZymnTtFBCHnmltbP/7
4IPtQrUIXlzYPUistAVH0kw84IXTioPec6M+J4ePjm6ZiZZ+XIPM7up6YQcMiA4s
O3hOJrks0WyHn0HRdkynrPZv08YkmwPzo9uwdYnmpZB+e2LRgavTfbG885Ng61iT
HNB13eR1k5JXFU8sX1w9y020KDeGfSiUmVlhjyRXUq7VKQqtKPO5XhybQRRl1igv
NpXwWz0qpzkD2Y4cR/LiYM2revfACZwUBp/N1uLAeCOhbTenuzKenBbYBRscHRt+
IUxYUaGdWHwCjUVG3x0RFz1/HdFGpYeOL/FPM+b/4gToEF05YGESGZ0icRm27Idv
AYrb6F0lAPFYBmN43rhOoURcmQOMStCKFTKYm9nLG0k8JNWO4ek2zsm4lHL1jtB3
PJPYLkQPY8cAQSQz56p1g7J09op2KL53C3KGw4yO8KG0+goXtyWtJNc2eODxpxFS
j0VPi1gPH4c9Hja1f9Z411Q2XhzPdZ0CaZ6EiZ2hDlI9+jI+FG+uvF3LysTc5RM6
/9HSWiC8dyT/M0JcnHpq0uOrinAilBwbzNHYOvd7rLgdqNi3LAZZNt6uQYn2PZbz
d0QokxaM/JAo9bFp9zHVnvLdmmBSNsegMVaN/s5B2+8Up9lAwbi6FJXwChikNoFU
mwEnZ5fdX4tuwjaPes0UcYVWP77KAFCOBpZd9LLKhwZvKooWY1UBBBPs/xjs2Wys
ygQEGRXZQfmPfPv3quvmJNyt3OTwnwQMrFbcJq8Noziw7NV+PQ7HLt54CDK22iuW
gBiPwk7GvsPmbzV7+R5LPaDwVoBhSIJlT7Q8GE96Go0U1jj6jOxpuWm0RtpmL0Vn
UE4cKkY9A6jxiM6kGv5hffKAHNdX7U8nN9yqdh/GTA2ZOEWpnI4l9yGngMVFiLo/
CbljUg67c94lk/m5P42kLw8D6UaNVf2nDnKplJ0j/1JucZn41mwAAobeRqXHpEsK
p2pjjjG2JK7wo8jkOuM0VZ68jojT6CuuHriFwBni4okhPpUMZdTCrtezY2J4a/nT
NTP1HJSd0BNatr6A+iBN2HD/SLrjgq4zYLb7o3UIlbz/JVrk9epU7+CLfSVY7Uh9
B0OaRbh/CCyQXVNFA1cxLVN71lHgY6rQhOFtaDmlPNmNAC9sg57Y40+GgEFJrrUx
ZDs50B5C5COLuINbv7BysI4ldjYhYPiQa5QuzN76zSUdaiVSLfgnugKILwcB0ivp
jI7VDrJzNULFjJA2ob9dLJIaJQ+Ab+dgWSrPgdfjuM84gu6c27gn3e0BNonAzCpL
gwQiXzIBA8PA4fvVmmIBQb4coRJTJAhkBSKbnKhDNIqq6CljKJc5HZ7oRf0yDmcj
Bc01FRLfEy0+qXDhHoUHpJWOJWZcBhaTpolTUzIaqS8dhvbdSffKrW4Q7sWqk93f
J/0G52a3T16jDCNVJloL2yVuEyiZm1c9mURATaFfIUNMSOyR/P6KIXNGMuopQQ/u
U7dt9ybBLP9kxtGvrvUO8i13b5eX3IbgRLhymOg4S2eTYhR/dIAHOrz5lP61IB6B
R98UmWKjIzOGGsZPjmU6EgF9eVfsNbajjSZYAqHhBLo/6IsdhVlAdjvfD1FZekgW
9btsbomC61KYj9G5Sx1j68wq6WwesSmdO9XE7u+aQJ3JIWJA4yYt67fQyY3d6Uza
Bbd9lF7W2LI52lr0TWbuDyJLhfvN7ZUwazp6NyARWiEJDJXxVEJdhlMXF5SGX/yE
IdMxuCFolla4jIa+FdarKeeJTA9YEcKZ/1sfKb/bC3RjYAKCU/H5OVln40saOY/m
3UbpsMf3LrcPAQU6zfdUoPHa/2Fn1rzmA5V+5JW67BBULY/JfYrBfq7OuTwxt9KY
L4fnn8GGZXFB1oZlgntg1CitvVj0ptCEE8g6TTVXnEaHiuxxMmt3cUOX7/5QjRgx
g/Cs5qpzcQ0KkY69yd4YkZenoEuhIZQdpiGp4ECiL/NNIEKCxWvQeDf2aiYudVEq
dYCisvb3UQLPHZA4B8tnCnn/kZeF1okVI+u0Y9yhE5GHzxFr6aJ8g3QKpVG6IV8l
B3tzbFL/V3AxEVE9gugnA6tjW/YdrG8n1kle9dMyKmqPuQPcycGbpCAZRPFlJK57
+xgYhCxNj5xv6hcUQ4tDiMIVWuzLFODNwpH9gtG80G2GMn+kt05ELIs7uyQ4gaZV
KbM6ypRq0KwRxXtUvBYyeah+O2K0krvXBZ5+PKTbCdPBAiVuv7i//KMhodEbzpQF
PZ8ur8jQxnMBcA2j6PswcLJbEPk1ILE29aeI9CndB2cLdvciVC97j9A8+HvKbnpg
BszqYNwen9eSZQo5GiN180IJtXNM8FB+f9qp/c/MCR/YLzYfk4cRqYS3TPP03sBY
ParuMW1+ErVhnoOz/Krdm0Zkd+EbN5hl1qGQkF0oavumSKLA5PAY7awT5BNCei1s
nEIMyWq34gzt6CbU7hbY4wUs+71pk+JtFq3lTGYBBPWkRP2ldMtAb0q+rmwQJv7i
+4uf6Vkpa5MW9hDhxKUOdGnoQzcWU7lQzpMhlcSZD9w01+h+Oj5oZs1tlHA9l7cz
s9eTSZ6h/b/sC3lwRypzp20rGW6Zciv2eqrhbxsiu7ZWqS0pWJ20wq716yBouY62
cwwb6Olv/fHQh0IKWLQlfwkb9fUoucapnSyFpzXOglL/FXr08gOnt3Gz+8reeUTD
Dru5dzbZ8YdZIe4D/xz4JKn0I7WSS9pjoKPTQeudc8ws3zhAFEENWhWDvh8Vrr3W
ujcDhzFUr9iWEN4QNIdqamiMf+AzHhGgSXW/5e0Zhz5l5n1Bgz18jzHgQbysw12r
kc09n+gucMlngYrI8UN4At7+ivcTzWcDTPdLd8dUnMXnPeMmA5xcuMUG7ALnb+Ez
Fb1O507dhOvTRCS4X/K4rQULnrkpVf9bVVCsOcwbPBMKcOWGrB3Zy/W/k9+WOE1l
DTAM0z3nApXMrVH7TZClbVhV9sn6uDrJ8dGGVk9lJcr9Ru/7YiuVi0Hshq62K99k
HDfvAVXsRXm1oAG/dyY3eeqFT+EJIfe78EzgabUvfc0eokQIIwnBX9CR+AeHXpsY
/2Dx8ILl78TbIOsyldYlWyeL0uBCCzoe4ypBbeNByzaQJ/CLdfFGMEVOPKMvRx1Z
kJ87FSPWIOLmYXZsPkZ7mOf2WlyUu4ggw5VDdd2e59FNUR0ce/yZ4RU0iYmYkc1W
YAmidsNdAzsehsLIHreQT9eXSOG8hwFQkatAbGOLwJp2SV+fQjLFPW1aiwZPkvYq
fAjg4ty2JJbyzvYdltr4X5ILRZqroo6UnLq/ouIrGFqci64OJ4529iQYC9z9/xDw
EnLfSWuemJwBIBxlx3ZV5xYB8fVhPp0ltnWUUweP9C6OWxJtSJa7TbYCMQItde1w
63L+CRK8dlO02H0kiEyMb5jT8G5iRdlZXzD0RKaR1E1sS/gQJ2/iAdKwE46FhGrL
B945wNhfaVIfRFI7umyYNHb+xyAndKV2QjfHBP8CYIUMZgq1Q+vgOoqM5EI1FZl2
kTit40ZLZnhYdffV3ZXWKm7JifKWjkrEWEwjIpoqtNE59nchKeUGjo3EvHxF8lGe
RMoA0t9OLrFR6EVVurg3MbDrxD07w4FGf1097uusrjxUqG6CBlAvVg2g9pavxUFv
4sGyN5Cbpw4f6vDdLJAcAyQNypKNbS+79yyst72fdNxAcLfVJYvPFDu3jt/ZF4zD
Q2nXAkzZLggo0YgOlDFtG9aUiLQAlpvAkmP3Qe8/bAN1Os0Z4CAVzsaQsvGPxP/c
yPVdCQ5sSo/VPcO7O2Z6zp473TQOXNrs7FB1CnhROwsv+n3STjV2C0NB6AHrF0NK
l/hkYoCB8otwbef+ub3glMHckkkhKwU7t//07e9bJosoRVb1+OpgZyTS3jfTo4a0
blA0kIjhBIv0sXLGvFjVYSNJ1Wg+9yrxUJ39uu2QvjruKZb9ZCLC5CJ2UyhuYSdp
SdJb+rtvWhDdKCkrQ3MnVs4S5ufbk3baxpIPZNnZTC62wlAU+lGJQETEnrtHGq2p
j1lYU3iHFoqf71YBXAHOKmy4dbbehQwp7X7RrYNakNNAKHlhrDmHrUDwPJwgRSSY
e3T0v2iDY4+5zTfWLZ9tR0kHleRIRFLgugAI2A6KvhnQngogCNKShd25eWnbyvR8
tbjrjXOtv91qMADrrmR9p0CbvYFCtN9zj9XZioS9g+8X/igeg4V4KeweZypIJe9A
rLVuztDXMC/52tOCRWG9s5v58fLT4o+5wAYE4v3iaBMUNKsxXxlpgpsFMdomYCcC
jRJ0JbTQIIpOe1xRrgnGhcQOYXEhEffo6ve4doZXwH89g/4Y79V7WcTxqG2dBFEd
xhuX+2BWVbUuW8eXdirMkjr6WQUNuJsTJx5XttoG1N7mhmpzFyhfP8O5zTU2jsTi
Gesnp106xRmDN3vLG8IJ2lvs5Zm9WI74GgLgweOxFWWocY/HLPnT6cNl8ObQSkV6
EtwVc4uiB9LuzJtvOkPHvdFjoQtG5Y0Q6LjDBGrNpy5fUBkCy8axqsm4TmXWLHpz
weqZLRRJJKokfvWZ+bB95V1dK+Kn3nTuFETY3/uXZ1R/M3rLBboitQwqDVWV/qE5
jmMNw9X54oVkkLxHkgg00lqG4MzcHPlEDUzeiQhFEmhfaqRU41PRfrfui13H+vb7
wz0txkUHN7rjmyMuPkyQ38LlJ3DAEA3dgaKySVUgxmVWGFAu8Nth86MUFWEnSnjS
cZBizKt9ZMThGK9sjQ3jT1/GBK4uajIWJRM2tohUjg/BvXOCiMgbvQqWo+fdUv19
BIQ3kwqyKfFdPB1ghQgUv8igxJZxOJ8rBFbyJVuQ+wGcvH7uJn/TG3fqnvqh/Deh
e2iPsWdaWGSpCido0qEiDRqoDh8wD3Fq1+96wpll5JvTDndh/Pq8wvDIivhBxoNX
4VrM4fQiBh3AXdKaCnooO/aklVSYIF5VyZSMKmAyN0+7F9+R97l2+Vpq2zHHOVmc
FeEPhlRp/STbmSJlLGtZyqn8NbGlvaiwNrQLPx3lOjnBBFEcmGDYbZ+ZOtl0esND
sbrBoESWfVG4o4j5vFjNP38V4QxnWVFhY/bitTjAj0/n4GaaGCXbqykpCkrw9Iww
GbYI6nG7avJt6KmrpchZpq0aIesGCPdlhuPersLMKzW9NXYSUOLymiCCpVeLP718
7X9DINgGJca8yivCe6DZmxGzoiXW/BU7IhjpDcE1c5ocu7hQoZkYfczK1tYwAIzi
fF+t8SfBzvRwGX4XCgxk22/D5iCEKXk75Moc7LuO8DwrjHn0X6iGVajPPbhoTL8L
6JP5mBqxZeD2J9zt2S4doYAeopiT+l8Mo7AasM5IPDBJ96jHlew6GawyldDbx1rG
ufGIQGT7hpgyIyXrKwIYGhL46oIJyVwgOUknk0gcaJI7m35H5cdVf0OmD66J8ISC
HqZvde1jIAkwmbOBk9KoYKQndfvtpeoTz7TP7FWbNHCFjiv0FCcIqgYrdxgcdDEu
93BumILPPT4beikbeI6fliWzAUwIMVeD5O3pGocJBYBki/DEtCUvp/i4+YhaIPxr
TpAZZm8uFJ6ti6PejiasrJyq5wRKuTQ+8hosiWa5R5WE2w1B1VutmZSryTKCk6zL
X7ypELFk/ch8TFCQBDUv6GiLfn4ZJ4RR1SqkIIh9i5Mlqv2c9//uVapwgnf73Pjt
/LHn3oWGCtfhiQuiFzepMySp3fjsmm2HaBIno+FRXqJD7AwsB4ekAPSD7bXMCJM/
LYnXKaDrJEd3h1xMs6iLasj1qpgpJzh+sDdS9N9Kp8jBeu0y+nmflcM6MPnRfXSO
Z99OYXQEZ4G2QdHbN+uZtFpqDHJLeW2Z/RI6W9lekS4J7D4mzDq44oaSjMblee9t
AZ368DirPvkRC9nT8Y4qvRXVfpDVOatuChcO4zz77iY/FViEhePdGxsBx9tx+Dfv
Cj39xXuNtjdF+WbiERNmA5SymtCtN69n3bg1KwfP9Quhgvvvq/TDHaGqDrmU0y3n
UD6xaZaxAF1AhhAj2yNSLLC2jCYZVPs5y0oHTC0zMHxidPFRS5O9sj1QdbN8Fdbs
rYy3XIo6S8VWMxj5+jNcjTdjrCvHjeo3tDWfyDfLApK9P6BKI+Os0/4F/lifnewU
`protect END_PROTECTED
