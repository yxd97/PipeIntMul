`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4mC4AyfJAsIGLPvz6ZBVoV8Nnpd81AjqDiQut0pPPTMZpOZQWvmqElsILB34OIM
4KwtEgcD2qVDJ5DxDy6IC+uT2otqUoU52wJ86fJOPI2NB8anck29UFxtVxyJo+hE
9DpB0vAr/guOYpO//RuFk/ZK7d/XPFKhUdmsfGttZfencB6JPNcCzlfusK6zkwC5
wubMQ7AVQ/NucVmWbKrQk1Aj5VU15EeuU0R5mqEpGuOl4V131Peq2aq8DnoKbFwi
XixTUJNC4n1KhwnpSE9wK9BrI+Xa1840wF5DnfU/R0b2FyfPwc+FiOJNU1tllTB4
sc1a7Pl/5FBrHQgz+lDndQ==
`protect END_PROTECTED
