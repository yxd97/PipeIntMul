`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GYjlumT/oSDAj8SL2VG5vN8A3u4TUVyJ3rZHhEwbNDd3XPjhr2kokGLFV10ALxk
ARMVAlCeH9P03e3whmyByiOLQJwi9SMIluP9n9s/BHfECBCo5bCiSQVb5wgLUr1A
Ot1KxgatDhHeb4BjJ15gWiXrgFz0nR9tNuhF/Ka39QrjLun+FSXtVwlvKX+gr3Zq
Rg8/+NlFnBZbCtw8LXEPE3pwHQQqFi8tyL5qECYs/t18cHDNbudKxDu3InfgEbNW
LNg+alY6t8iaV3jBVeBvZInfGpADkt+LXLOjIPUc4HyVd9C6oOeXeoBLewIoexLD
7FFcTHbdzkelKxFVw7Y1IaBTlNTL+dOGmezSokpPwtUa+apa0/g51Qsoi/cyYnbX
daDQZTLxftcwpVarMwb9RhE9sCqEkwuu4Xl0fXo/HZnznU8aVP9FgId4okOCfCox
dYY733aiDVrYcL5BxptHEw==
`protect END_PROTECTED
