`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WjXJ3lt2qcfCSS2foNdWfY6GOrTXwRwNHa7OEg/yo7Wtx9DvYpR5WsCdggFMho4M
+kEl4S4Mlx6fMvB6iTsWR2RKFSU7lKJja1asnZVPiA0LeFYlQCcxb9c+ocn2ehD1
qd0fo38a5r5aTLZMJvf6LnmIrqdHaVrKbL5WRapBBGFTQ8hSeQ4126dbAkYXdntL
ViG7PS8ryP/oP01j6nkoXK8o2P6F22hgUKnrGYuBCvrM29sLw40VopceFnSuul6x
xBlX6Je97C/KubkSfKdglhLO2stw5bswsSb62dRniw9+Rnp+YG+fAg8NLw9+bMFd
Z1DDurhYk6SfdUXojzSpIL2kKj8St+ravNRn66FBEyKEmC6s68VsL6tpl7nvKTvn
wbRyeJ3kHXJRoG7uNbguO+hBj2Y9+NuyJqyZQJ5UXpmj9KTIbmcUhNOaxbQbMbLt
5yBgM5lWnO7hgtEMVF+WftrFxReO2R1gUBU22j2BwX0DykGIL8SpVGwKFjrVEyiS
SmZZW1oonmBtGev8TqCS12OTPTChIjR0mimZEJntGQA=
`protect END_PROTECTED
