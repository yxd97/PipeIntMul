`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmiXy2jZHMraAym/q/pwWPKL2Yq/83SR2wEDYgLU4rcTNu2izNz/TZEHZjj8fnGG
taeLCa5Anu9S2sY3NiACBGVpxJUl+5RQ1p2WhjURY8t/Z6/Dx52Ozk/SumrC/KKm
Dch6T03OSlJOxeZeu+FTZpO2a4l/PjuG6/YAe97V0hx5Sf4Vqe0ZK9OLj8PGvBE5
/qP8cirdMtWqGGqvopth3IaPXPTfDzfeEeDKZc4fVDLbXUd6jFPf1Zsw3Sr7StUp
HFYjX9x/2jmY653FXATiUHncgq2x0Mepmi5xeG76wGRgDvJhYpb/bZNby3RYHF1U
5ruImeYdXMehlE7U9oE+kiA3qIqHRlkvlPju4+E6mh0a3v9CXkEzxawZofVDMwAQ
qjyvJpO6WAkWW++G0wU8+mza5tlllk7a0DVNMQBAenU=
`protect END_PROTECTED
