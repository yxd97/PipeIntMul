`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7V9ogZxxIJZNQul6JRBFW4DcLWeKqIp2OomZ/r4J2l65Zu3o4b/eZCX4aps1hg00
2kjZkS9LSCFvVNWVKX6vXlLM4wkGPkAvMlRvpjxd/wW5bLbVlKidub26QYC0WD9O
zoNcFBR570qo5TQ4abPem8qxXEjspv9QBOZGQSOnEbkXk5lPoGH2nPOnX6JJHEce
H94nM9sMNgUjfVLK9WFVcwcZLjNIFqF9RLalyn86MV2rTYFiuvFOEO0bCABGH6Vt
iodMQGnO4XBdf+tH2JhEfLTmHCEmym6iWmuBku4VHHjgQoMgrD0xrFVEBc4oGmM6
XAaz/nolzkmO0yPmBi2sgGfccZrkFuSOPEB408JOikQ=
`protect END_PROTECTED
