`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WQqN/fDEYXt0xrveiAaIHf9ovD/JPl6nLZLGXc+1RvjmEz8ru3w6ldIsuQboAA8a
pQGDgVSo/D9H/VoUmAkcziqB5L+eYLKHSohgzZ4c2Ht5Tlfs3zD9gS/TIwYSHu13
rE6XHc5TawKCo0Edj0MyH7BpuKsUuZ6PWoitGaaFp5DZXZPgOFJFxA9PGOEqMXcW
csIKpriTbJnI5x+byI7K1euDk+odyaSP5JBph6V0+smQ8II76Ne3Pkhz9a2fdbo2
hRulXcpEMKpF/jRFQ1eZnSmpid0PY3ceaanpAvgoUFsZZNG8+3IkjrjsqeYusqtu
NNTogVbyCOUVi9m6Ixn5+RmunXAkYnouUu3FRJZqSZsJluNjvG0Bh2rUKxGVYE24
MCMnDWGYK7jR5lzUOtGVNpPuL2XnYQRZLtv4sp63g3KIHHFx6eacvd70OUA8BiTd
SD+w8bplOzEVMO9eJ1diDXnDa2/hxzdiXf6lOf3lrnrbQ1+p64qnQerI3MZ25yUx
ODwSZlADbw6B1xyl2sQTqhi0HrAVHZygtQWWNBLIStg1jf+A1SyP4BCaqMCax/pL
KOWnEZu/2H02HfayhGvYZk8aAX/ou1Dg+otzShLI2CQjm1GMvT8WO9WmbVME/Gis
FGnJE6Wau9vqI9+qSpfIzIiNPy4rKgzpjp2taVpE6InQB9RtnIUWO/myD4Nm/cVG
kJtmmrtYjnfJlZbDU3mKx6UwiIrVOU/aTMxQcnaiNnBD8YKmvvXnKVbLpUe+IQb1
nkH3DfMBIKYwtzNkSsttaMP4XSDwm+7jBeGatmWKkUm/Pd+4a48jY8L3Q0oi9Jgx
uRcoxpGvR24og+KTgEstNnz1/myU220KnbqlVJHDXXgLMHiweShFd+2A8uMvj4sV
IQz9EdmUa4iH6QzbEocwY0T8usmw3N5EoeW2iLTJrhlSoHQA4wHa57qocFYdYHhA
2x5qnKSXLFtoGQ4igV60ocRvcP15WUBy0IoFF7GyiBg2e3V+yt9FwHqARDh47M3I
uLo/DFKVz8PJKNFG0KxHawiN9CmfHpHjc80CCCsYarn+wrbj6XOC/RgB9tfqpcTK
xpRlOnGpCoBIbVJ5Vw4QDLbrpNa+wDw0BWU5UqMTX5DjzAxXDg/OwkxKbTKl1uSn
lkvMKDNbbrAana3OBDR6hc0adI+mWF1rFOrmtOdgWzLdMGv4vn9SNqwVGnPaIcWo
2Xc8sKkD+7k35Cfr/aqPV1i4cWOKTnG0n87GanLlGRd2GWS4sh7DXq/blSlmMikU
zhMD8mfSYwElR/w2ILugu4/SPuzArF5EWGvY2XFvBD41Ty5Yx17frc53fdlh94o5
DXzacwkA1bUBLZ49bA2sxWyDcOSzwoEkAy5PbvnTy/G2l5wPDNAClWzwUCAM7r0r
+ZO5JpcBhca/AO8j3A9owOuxnSLJyNGA3D8w4MDwJKr9TmYEasHN35w9PXY9p4kh
IQPjW7ksklQ0CwwZAduYmp8X7vnPm05nyUCbVC8QnyR6Nu+q66mUpOgMpkHUIjPx
LrUXpsapnW3eRWJ2aRiTsqiDixTspEYAxSaYei6yP2NiQkcFH7n4hMscH7cF5Iwm
xMsELudKxhgWNydkYKWQ1CZAb0it4jdaCMvF5zgMqJ0D8DP8ecrrAxv+8sWzatnz
LRiT/wJ4MS265lJ873jR+z/t8SCr8KZY3v8ieF8qUEV2HBOoJ+wS/uu8K2cj+cyN
mJfXp1pJ9cJ4TUs4AzpeZ320Iwh/RvrIU7Z0Ceiauz1X8eEtKvV9Og2j11esCxNn
vN6SK+ABpZDAWVKmos6J+4ZMz9A735cuDeNdyCEWcz/YzPqQdUO9Oo8MGUAjK6kJ
qOwetbZmrUA0cBLRwpEh35SOJwbrtdkWwXyQpPFdCr63JXSa8iYQSNEaQqxUJghV
7UkpSEaZ2xZuFvUz5NZeudb3+gDlBrS9ITE0RzK/7/wuJVeDfO5XY8OqqiElWuVa
xfSx3xtIjpccCd/GC92D1g==
`protect END_PROTECTED
