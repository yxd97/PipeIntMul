`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uvKWSHrSq1bvalRVSbJE9HkhfNNmEFSzdNBe80NDukwGltJSqsJ1mwY1ypuuB/RU
iaMwgxICYmoMHBWXpbJuFbyOWu1BIFAOb4cjpXDBm90PP2PACuk4T1SmXn/4lECF
MKh3twEyb+8ZSsli02mZe2GOT7+WI1RedLPaHN7nfO1+rH65n2BIhcx1kPiZOK05
xG4TZNHK9s7HRkMZzQDwDVQ/BtKWuOqj2T0snOD4ZZhTlhT6IGR4glT6AeMml+UW
e1yL6mmjH90gihN2SvKSHJnEzp3we5dYz1LgbZT5M+HS1Pe2B425bLHb/brTIK3E
VZOfOOYRO4hriD7uHnzWsTiT3pHAOtBXf1xVbRzto6hoq6NTx9Yi80YcZieUlE3f
Xv//r/BtZ0S3bk3L18g6w18O+tTJcVmniXABmveNgjPbx/FkkqEQi7qKM0cDAGd+
VUlcG+McvyVXCnDWHQKoibfkr9DmEm65LXaZpgpQJRXRy7eZe15WP/Gjf4kiroEl
ihzvZcNlZpyZwqHj/hLN0Wq+4DdDsoyB5U9vK4cAyyNvbaunRBoCxhgAOPQyWchE
i8RCvIufDaxsu5iM5KjiQMfHQ9LOgQjxz/ETHdO5u0/VWkQiZzpUAdwPPIPltCq6
TxJWiWJmdinDttax/bVVRyWa08WI1Ql29yemuFHHsGierKKQw1+tVBULma6UTSob
GGujfRJx2IAQys0HKG1lAermWGyUCTFIZRYPxW/BIIJzWt+tExyVq/jNzxMeiWGz
b0dvGUUKiv489xFChlljEf53EN86By+8DClC4SCMRy46taUkyLHl1z7ns5tEvu3P
kuB0gEPathfLCqGaDvNHA1NsCGWm3QyAQxhd/omf3dcofwRFTNPzNLZwdgGA+A94
C2IOXvjNmF33yg/uqhGIOrnMiROJJut82vrNitEX0SSItz+tB4vp9VOZbrD5fNht
Ufxtmr8k//e029R1rYVcr+nlz932Rc2vNe3dpqIP/K9owMxxpPW1lDIevy9wSHVs
fTmBU8hUpPwR1UzFj1pAW2iM1/6kMqIYyX+FHgFMOHQoo4e/vsAZqKmqyF+VdSdH
`protect END_PROTECTED
