`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
io+7XogTAbCgcP39sdlTu/F3hybU3vsdOhXbF4t1r5uu/fhlz/RIdbnK+gch3Soq
NozLIStOgMO/+JXlfxQXwp51hzD1r81Ryav8cD4R88LcWMuOeZHtQowKZmp3XDct
5QnxqhYKOAlZgW55yJshAgzWW9b7P9u8/GEfaJug0Czslpj9XWCTD8Y9F/2LocF7
iVWoQL58PqIHyIRzJoZoPUnUGyqa+04Y63OvMXOwPOkimJ10u/zGoMqpbTAaxaWB
h8dZgcSIrbBDP3EcJdrJ6XqRen4Bua0gLAhnPi0qFZPGz/8gkhplk7GmfL0dZvb3
0Kftpa3IkgpsG+RjsCqKBVXnAiWDuzon447rBkY8YCwwBkGqK/gAiQTE8FuHubus
oJsAgzg1RoDRxhhbebFk5w==
`protect END_PROTECTED
