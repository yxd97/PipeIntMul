`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJ50/1cfzVQirbvsg6RxOo0y4Gt2WD4gqt1oI7HIuDQUXqB/bmGWvLhBC66f+kCi
PxJWvBEp7qjHNlVYKr5JuAOlqiH5OCDZvGNff89KazxVvJJaKS7mtcPWaGh+ggpZ
MNwWq6OCN1Z3MOOEN8ky9J2XfCDrdc47XJq8BWOi00L+3NOxaEeQkKYXHJ/swjT2
uf5u9428uHCsKvVgIqU11nmcjoJQzgwfOIhtrJOrH9EOVp8SvPd0qJZH1fHfPTwJ
eJNuNhc4QVC1HNcple64wgwMFYKOtaGTF0qgP59pvIxgjf9YsvEagoEGYIvbz5Wk
Edt8ehqvjAIu7HJv+tT1aHbTws2l5Y3P6LQ57xWYMe00AEc46lf9rVLIX2x3myBC
QUgan3U6Imgir1iTVyzk97ovJnNvFwbP8nwmHSwPfCKPlWBL5OCDAe+almndkORM
AuaSiFNeveajTW5ATyhhFsVR1M3eQOvmiZEypC4MPJ3lCKQRwLPoJwRr640O7eOG
nnd4xaARqVVf00qpF+S3GRvfzScpmyjLU+PHZhEuByKuX9nuK1Ks2J6r5zJyDjn5
jXaZe35qa89qw/bvFf7Yz+krMPUwcIwJ7NnSRDbkNQ9TPPNJ017a4wjWvRU7E9HS
RjOw+4eJKB4rxxeo8qqzrvcF9mCKySXsX4U/88fLI5DB/faWjnaxC8ExiB6ZCi41
0Pdvm332CbqzsBKcc1phBY4FhBslf3DoHQSfNiiFG69W7LI2pS3j+y0olRHyxXgx
gcehqtOdPDkvGWmcTbkDCi1WZAnSlZObBAYel149x5ELqUOCMj3f6HY77fS5Hya0
/ccx0hkLt4YCW2doCKSf26Bow/WjgTuyIWnvqzxklAn3FIAexjsN2Jzwn/KEeGaw
7n8rCgZrefFHQxaI7fMZSS0RX49GxHfOGEwWYx61pzoM8VMyZ/vhdiLv3sKfvulK
QlxhtHzsteiVkJTv3YYnXQlttlC2YJkxtLZupfgOdIJIRvAWY9k/S6wg/mYGUTao
fXjJKSGf1IKYHRzjwZeOK+GibL0LuOi5zEXER8HjOAE/K8041x5s1f/p5kAJD8ye
xgmsp8yy/qH7e08eHnb1mnPpdRMqROzJ/k4/ldIpZlj4Z7GSUMht/lWwI8q3q7sO
DqRp6QQBeiNu2isXxudFymKdid6+ibhK9/lhtMBeslC+63Z3k8GtEpvpsnlraNVp
yyoD62gcSwwmrUGhVKcwb5KSgU/7fJDMI+y13UirF0iR7VyrdtK+XGHrEuRNStJ5
sXqZ/4Bo5DR56sYAOC//u46aCYr5tYEHw8/XycXvdbxQXYiz6I40sKMSnW2AwKTn
Grto/wlHdjpRwpScAZ3rxI3S80WUG5m4TjDYw+Wi2Oh7GFHgpemHD4mL5ADpaqms
0vb6iLpTpJDBuZaQS1OcjlbkEqlFk1ENhMAszVHyYjIanCrlMxc4eY8p1O1kku2L
7nX6FdL75u76eEnUj4l0L3fmyqpABtxK7NLLViB61xf1URhbleg71zHj1QNcVMz6
HTDQJoPQL0Y7fTgan+cBDisbokyR1UqSsS0PjFeZF2vJ+pDr7qrcVDW9tYHsQxqE
xMXQTtKplYgx6tR6ZLBCLnobGBT1PY01Wjx+U5d1RLVV72sFkyCGJwfnKxPavu3h
2COCygO09uYv6Lz3Sd6yKdvxUW2CRiaAFGvNkRvYb/ODgQvVPzD70WM1YmScCtoL
lTfYxQM3sFLP76SJWuJwZzoE4uNWhaYkVsgsHqY6RHKYbmG5jyvaA/ec46gkwqI2
HdrRwdtFeADpcqYnNd2PnQzeCIEhtMonELF548O74LORBarWA3nP1oZ+ZBwieWmn
m5HNw7DoADCTEojPTIxJHgvaBtqvTFecTRh8yvFFJpwmFSD9nn/eIZTdOJ+AiqEM
6Eyq4tyeV4JOUktDoyP4WDRlJG8uvkFTpQr3qN7Xl9nZLmrqnnDMShG3z/4oJMpZ
Dy1s//aR+DQfxfRtvV3RuuGf/UBrt53LSsAfsi4l+JbW9uMpXFIasQi5ViaVVZd9
om0Mzf5ws5IedlGiwOiDpA==
`protect END_PROTECTED
