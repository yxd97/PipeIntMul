`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CrcA4PldfRj5ZTW3y79U9Uerrkuewm5y2/Lvz3FiLzKm+DLYBTz3Lb9Wq6j+S2S
1pfznenfcyTAibeKO/t6VPPlwXj0yD1+ep83fVa/Kb/y45l/PpZxCqWo+Htfei/A
xjaKUvPwF3wK3P5iuIV7LX+gMRTF/slwTmhQVEySAdCGCAUTojs0Tf8NPPM5QSUa
+1IYWwS1BH+5lTxAFjOzei4uwhuQeMgacX0uWbO/OkOowrCBx19TRD7OGwM1xywl
ZL/NN3Gi/rb9bl5t3qmnWZw2x1gPezVdG24WOXwlvVuo5SGHCR/jZSV1QAIJM4U3
/iVUTTb8grDdaTPjSNedvT3OQZoohhhnwC2KP60E3hjruVX7+ahx5HXZNq2qzPqH
pIpHo8MerST7dwjqaQSbITxcxoUAZRKVwOoBGMY9sTbSC5+VISTeUwuTptu8c7ia
TkVouVjSkhoZYvqar7N8YvhOH0nSTboJ1IdupoHa87c=
`protect END_PROTECTED
