`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQAsIx+dRIwKoSWcuf8PRwJSwjp/Gl1JpKBPWuTUp1RIc03bO5ws31jG5SvTpr0d
KUDQbEkUQVZtPI44WOyJSM2g/ly9lm+7ejaQmK6iKZOWOulEkxjUbF1xNn/K2RuJ
eFUlKAFivOrxYOGX/fAFXiASSQWWbu6fFdDmw93NzLah2U6bBcKVUiHPgtjOHEVC
VkvZyidYLD9jfm4tv0jPJ3RjUgc1ALwjMFSiZCzQIUaqebxJMRY6yPCzvxXgTAOq
Omuuk2TiJ/VH9kozxzvajRbdxRHQaP3H1mQjJubOZIC21UPB31TV4PHI6lE7gzHs
k3Mnh9wk9+okGrC6tdxzeyOfrXhFHPFW0FePGX9dkxo3/p74QtSWbzhD5weOLgu8
PZasgObSXCwKdJKttYryW8emT13Fm1PHSQzgOeactw1Cv4dx50njPErmZ5rG8Aif
pRgWVykgOxqWxANc595PKa6cXIIY3JZ7pUmW+xhGGUoUS336cRmGVsmtqjKolZmk
eMvJV8zD8Ps9IibsNCK0Mi8meX61ZBOvS8jm9jdZnchximBNtDlA10SgnI/12P1K
6TbLB+IAKofJ04/DWoOP/Pno06031UoX/1GMH4j2sRZD+z46XRyMSwiTYYd/VM5f
`protect END_PROTECTED
