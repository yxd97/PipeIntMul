`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+j5ZFLGdcUDKCrMTZgyWRRyNao0s/rRr1pZ3welCM+oLxbmEhhfS+vSkIzUwR6N
6hPy0n7qH9ndOkQWYCWiJnmwlgn203eUXxsN7Kaxp36vvBuw2VwHBr2XSSk+ppxj
JegTiquGvg13xxbVIYyfVRjGmGn6LMVA6v/adC8yVi+zf7grzOHVhrzjiBJUmale
Aif/IyQ62t+UodI0wfxekxUfM9GLkQxquk4uImXUGY4SWYdc49BB5mwKjMC2fi3W
thY+2lR1/ZqSTXB/VLsvhp0Iof5uHzGzjzkSLl09bGxOU6JiFSgwVVFqfrmDhUDl
vYYJ/dujL/ifA0sQv/tkoZWUqQIQsTvxeyT0dQ9XLr4Qg5W0/x4FmnA4S8LljEOc
WpKxPO8+umiE0GGTJk2X464zHaWiSPC5r9ZCw4hiBhTfKy/0OEuP1t27Z/mznKTn
Y8lsVtLOW52QTQ0+vIBiSd4C2EjrgW0er4K6FF2tsC1Vyn0CBPjg0QPjTco72q2R
EU9R6VoAcM0WoWjbsZYqiUPkR1tRW/jd2aziwhyIWukpZeUa5u7z2pfcOLnsxcDi
1Vta2kz7CnjfDsL6hucZ2z8xuA1HmZE0tSt+1JejvCQ=
`protect END_PROTECTED
