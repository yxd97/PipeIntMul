`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBNxln1TgnDt8ToOYzpkzsau7KbYNiW6Mm1pXy71hACMeyQJNZLUfjIfvpv8Uc1y
oC5zjz3WeZD0WTE+cE1O2CmJmCJO9cayL8TxGmutj47ucNIZlJ+yf4I7aC1bM1Cp
hQoYMJdf7M/t2L0+bOHp4ZjuO27Nc1fp4/nUU/bxjWzsZnuTxfXBnBVSDBKp5eG0
voPpwV93ISKpBKUu0gEPWFfYWuX5JhqdcMXERidFVPtoPhTvZqFLH1iMZlhqOeYQ
gWDzfP4Lk5gzcuM3TXsXl4LcWzQhDxiZzSWp5t7CGqnBFN6GoHYOm4IhDk7iMHGQ
RTYk8ennnkcFGAa408YegtV1CEfrU4bnw2Z8zBFcLcO785Ox9LHon/+YfAQ31THL
FQOUDZgsOVlXrIypigUsZbbiA0kMsHNNhD8bqRZs5m4=
`protect END_PROTECTED
