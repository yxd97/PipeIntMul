`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMMs+s256IjHh5asoJTX8MJcgMxNmDJ7HIR5IzJZHEKjDlS++Hq+WjMhg/veUCPh
7QSwVJpAcwvondnQ9mxEH0c396ix31hnm0pIKFEiKPQcs/MtTCNcMerpTHCdb6PI
aF8YnUwTGv8N07eMvCzA4W3dZL+v52pHM5yPnil7edm8x28wdVpQ8LNhlbBZeAkL
oTyzloiC3HEw0oQvnMmc3mMu7TbHRsxS6dORR59p5FzdsOz7FTHWq93dNq4D9Ghs
ZEopYvplggSOLCYDQ2OCLadow9Xa4SX+O2ubFqzBQwm6he7CYoiIYSITeyh3JmnW
tTylDXdDq7Np0edlETJ1qXcnwq9NBlW8NZBDt3PSNwjAsV8Au3LuT60A2sE1LLyc
00HhTaxJdzmR3DMrbbCYKl9AZvNtxzbwFc13wHT/WzTmnns+KnoT9GFgZ8xPKavg
vZP4LLI7ICR+QkU39Emf5Tcv3r48XgR3tUw5CzxJ3oLuVJCiZ51aWrmfK+PlXMQq
57LFCbdmarFEbMt5Zr06hmly0LHujd7bmnJ9IWkiLHwmtFMpJ0b104CtqyIZrk9j
8Wj858KdDVdZFEZkjtwP7TtCT511KdoQXR68kwtlSL4=
`protect END_PROTECTED
