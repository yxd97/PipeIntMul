`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFxK66rSdksrocX/V2d155X1a9YtSCjrp0Srgs2mKE+o37oW8r4Cknot6QvZVFHN
ROZxvNhNqYNaKJokS1JC0W3K+I0CdPPZcucFXDCPex/giB7XvuCfNOLt5nMSXbzZ
TzeYEpnLwDFVHIddcbaLfkwHDywmccmMuTID/38nEtWgxCoIOfSmFrasSxbysetK
HRdLySBDwXn7Efb0ef92CrPHjfQkFsS4pNMY6oLxl2w0fxgTvXWmSz0ToAqustK7
/DpxJZTOAYT/3kPfbgJ2Y86iAUF4mT2wUmzf+ZCSDUdau050fNdxh/swq75rwS5d
uaLPWOaJPzDLndra1DY9Z8lNECsUW8N1q8nOXEBlCVYRdV9k8jAT+2xX1nzWA+r0
q50+0naDXRZVvtVocFQzsQ==
`protect END_PROTECTED
