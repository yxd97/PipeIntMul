`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0UCaxnl87bPRle0o/oiSXTTzrJ/whX0gYyUuAdXh8TDtX8RIn2V7M33s44Cq9PP5
GTYsoaHvmpiSYfMo328/ynFeQynRoIMBAr6rNiaum3Q0a8UUIEgHeZ8mnxOlCEiU
nM2IJsQQ2yR/0RY5l0DVyWfoCYEKFQnhvO2XWqEoIzzcYheb2CMVn+U7PZXM0s3A
tq5z8OB8Y4hzr5hfuK/px6EQhkj4y+AO91dnvQOv4OdNo2LZ569DuBxdCqTaqNY8
RGM6HZ10wA4xIPNrY2w0UJOEzQkSEPPWSSI474vj4tihHiy2oJXcJdafik/SaN4E
gZjgLwxwWg4lE+F8uQu4ehJXMiVWoH/QvKgsSrXA+t4jtsldGn95dAwjYuGKuEvo
h6SKaSf+xzHLWKuxY8P6CH/BfrkUPWcxkxRkr0aiDfFpLBe9vxatGq9xJlyjfPFn
y6rXhefY+6T1IrjmSMCFvTBZP5cN394i1BNwAgSaxnPc7GYtRAp2NAx3VOMyfQtH
3ggWMnMucd3Pl+MXDcqtwFlCITc2QrG/s0M0YEFs/Ec1YQbplPG+BYU6BjMxTdNU
`protect END_PROTECTED
