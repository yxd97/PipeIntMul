`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2UtSukbwAqdzTmJ09dN+wmpCmiYo5WJcIcrFWanL4Mli4TGPLBM9CSPwZOwbVii
Jiwx1+ISr/TRwUH5buTSIbqFeDvafSaOgJ5FAfANTHS/Ev0e66t7xjfoiL5tx9XL
Tw1sS53W0FR5pczQ3r5RcNKfHLZyo4QoYit3Qmb6qMvY2fmfRzMKwqBKCT8y3f1W
1AZ7gO96K+xgY2MXagyR4iUZQu3Jda4IPHI1Gj+M6gFexDU5G/NZcHrjM9gpWpl1
cC92aNdgLkwe2CS+k7DZsendqlF1RlOrIGBmWRCp2DU+n4DcJDLNwETv4PZK2Bc3
lvZPUzYzaQKY3FHPVF9eOfTXtV6u4LPcEQ4dFv2kDJqKGlvC0fpO4KH6f1i6guWd
+qS2OJRS0a8ie7niyVVI5nVpEwGFYYdNi2qweSSpSm6d9YnuXLCSc6seCWWJ3nAe
7eFv3Jp72Vj3PM3Nmr3u9glSUw5Z8nmQRFYzuMWwHKtIZ45yN+8cBKCHcfL8PWbP
raH4S+yYWKfYHN+Rm2Nc1bzVjf3S7mzNILR7BvXB1YwjFU/JehZ0i5tNLXRMVlps
NSGcw+FYcSx6DHl/xK7MxzkND2h0LK3IUwdnbWX8V5rIQCp6In7kIbwXSuNVxJIO
i3gwgZddPD0/CqjlPKizMVcgU2gjKtAIx5uDHnoHz3w=
`protect END_PROTECTED
