`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IFczVuNoQMlJMLtF8yGJzEmihGk39Wh5UicTuuMdvWrrp1ZjH1TYkn3xtkQdvCv2
A1QdD3UD0d0go4/utCEuA/XNCBG2LXiIElnI0+ZlsSIn8ep0rLIS5YS5pzNQvYAE
DyKTuF+1Cz/UJXR5HUZ0jhSkzFU9D+JFeLC3Qp0Int6JukWlcof4+WVAe2XE+5TM
nx46pjFPe0HcaRgAWyqWBNHSlPkLG+7H0jOV3PyWScU232rY75CUtVB4qH7/oh/+
hmocVZtMfa7eQQFNPbThVsfViPyLRdoMwRZ05isNwXMNbqGbI1TFogaDG9XfEjMi
`protect END_PROTECTED
