`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNRgnKtLuUHmGF4GteKyFBC8GvfoDgogN37VG/OrGaKNIN4oVGL8jFu9tqjUhTXL
fZ1C6egACHbn3qAqf5F0hYOCHp6aQvsQTNQi8y7LO4OepzTlG7fUKrOd6iH2Ab1K
cPQ7dDCWkjsJjcz/QnIVe+oEuCFd1TgxdZJ4yVA1xRDQmH7CghTz584ADT0Nk8O0
M/n0V6hfYa30X8/YuiuuOrtX1MPHrlLkKM89BtCVm+8KhLDTq8nRuY/mjczoEDZl
UDipnF7H4ie/dTlwBAsuwgbNtKYh41ObhBXsQtGiVaIJvvAYKXO7hQCwsi2QxjDp
Z9cC931m1cB3PB4lxhXjbA==
`protect END_PROTECTED
