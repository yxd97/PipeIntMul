`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xh7Ik7CtzZFowtA85FJ3TdGkmdWLkRhCW16f5M2NjVGrJ9hJPzQwObj6Rh2x3i8A
G213kTnfm/JX5Em9aDQ97gv/MITdGdCf+Xxtjmzuo3aGCL9fJWREMcnFEYn4jMrm
OTe5mOJZ9UY0mRXIQXuO21P+NggGzyGPWRNaXjmyvRN+vSksO3zKhZJ6Wb3YM+R+
31wEAeP81/E7edqEmNY1lvWp+fk+DqNY5utZU7/l75JeuRpD+4F3iNjv8Plvo6G1
PyZc+iBkPUJo8zHuj3l3jl7iDBY5qPaDLZCER+6a+G9qOuDhfX2Pnb3K8PrzTqMp
pBCU6F5FRlI4fuaEysJnvFcrNE+uTrjFTH9pqRGEejdefz5q8OL3ccBkcRKj86Qj
h784EtneTlZmtTHykhn2enuF67HhMykDj6+twW7YuDc=
`protect END_PROTECTED
