`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fk8gFB9RrW1JTjmPpa4UqELRzYYASjV3COOF2OUCCagkmpaxKpK7e4X6hfrXrxqy
pqJN0dtlRZVQzZL3WUoc7NckWtot+pGjgXxfJ1SW21Si3qtdNchEzohfZlXYTW8i
GcZCRTQBa0laecGHE/EMCUdfh2zlOJ4TNTTHoZQnwygGEvApTHV0u4eFRPk9awxr
hm0vzVqqADAY5wDfs62saDw2ZgibRRt2Q1UsfgvnTASp/pHBjt3Zwf+L9ji+LXiW
jPaRTk2fCqgaVZMBr0Ujig==
`protect END_PROTECTED
