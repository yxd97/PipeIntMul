`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aMxOkB7h13dAYIvzBXCZIg99bYS+dKYSsTYqbCmrebc0VoL1T+533Y5Cb18/0Qpg
+BzR2uyEoxOiGwjrVb4HDOMpCa+lSqIw54j2meOFY3Xoq8kKublbh0Ph8uM2vMWg
CclLkfFvAy09Fgbc3VjTwe/7FgmPf4IV5VJMHxUJFHmtwVY3gCa7mqioPHz2wbcC
dNbn7V+yG/6OgcZSmd9Em3EvxItdQMBAWRBjuIWCgUa06H0hAXqj07UcLwCQVl+I
QTMNPXErGAA0saNsrSmwQbRwbAznKoeiRgEF+2/Rs5cqCFsF8cL5+ru++KCaOawz
fIq1eh6/ok7/mz9coO2Z7ebcD1erKnk/TPNZbg160WYHBYtMdpr4qhqmB7pt9eY1
g/649eRR8weWztMXpJJyxzHks7iKlHkK7Fd6iMxc0MLhkzgTM6I6HEGMeLQIOHav
aC3cQjNKm14IL05xVMu8xzjvnyN01LI4EltsRDCrMqs3D/2OtsLI8qOfSRlTeT8E
LglTRzyUCF/Isi1uGoiFSkOOsKvhvalqnIiIFZqaUgjGNujodqvGWSjiKPbBq8iw
EIfA3kPL0xiiFPJhNpvPY3oUhyTQpApV1t7HRYRRbiQ=
`protect END_PROTECTED
