`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/uEIKY+wSjmCjMNsg9sgvE963kuzJ6ef8x0twRLHsVgyhh38GQ9QQTGUPtz6bj2
PZO93uNKV4oqFHtpTeiOlFRXKlQ9B0kt0ZjlrfVS5uI5/QLANy+92sw/T1R6rojV
ZsGPYIo6JUOVqWcgMTAlSYx1PAXahD8pWOktvjMFdJF3qq9sByb//EXXjo4h2a0k
O843TIm6391XPHISXaaN6uW/tNybB6zLYJetaUGkNhqvcouQVkZRRMosmN8PWKKt
aW72BoE30DWmuETP/p7SkhSplgWVX4F/ltBpX0jetbHlKOrJhVQEp6eEMN0abY0u
1WJSXDPEoTUNtLncOQqqFwmXCdSXCk0QrPZVe3YnMLQBAhr8sRTXqbJxUPmzOP2A
n/rA53N9u+9oROC+QQqr9AT70jQ+YKrgzFj4RQfCV61QJz3Q9359KKL9LDPyrcCn
UdQwpX1krP7ffmsisx3SyZecuUP1YW2yyBMVAx++pOIgz6YgfFtfwTr4cfNI8qYB
Mp9dWXkFr66P8aBGwqtpFyu7DYjMLbsSS75kw494ksWpisn2ZLFQchA42Lh7nafQ
FybTRK83rku4zb3Ewojv7CRDJP4rcffS2301fMvPUAW5/tnjqvox9e3U7pI1CftG
Jur9bQcn2ZRHAsg65e0Ms0TGxPVNOpnroU898FKr+KC2BO2T6VpTiaSfnbhOD/yv
CdZnuekt6XmCPK1M6PWZ0ZE2+KyO7l+Dr5i2EeIN/XqaaEqlzs1jXsoXabCGYFrI
88aRG1bLZmx0+/AQrEGvPnejuLQVh/eGYyvDsZ9VZO/HMOD4XOjZPu1MJ77USryn
Kl1/LT+rhw0xAt5fgfNrMzvsiTp1MOi04Pa99Yrv5d1jarIN9OuWtC1EKkbTHjn8
C9MdReApq0EYwFjuBd8LtZySSK1IYIClht5RRUQQuUrjaJzp3Z6QQYwummc9oODH
DoFrPKq8QWStm9kP/9oQYw3A3v/thjnewZ0seQLSaR59IStVmEDrZtve88X4rWqD
FEN0MUzmT2cCGefnz34HTAbCJp5tnrURox/enWs/5T7Zh/i5GSj6Xp3lmxU2OfZM
EsVx0X+yldtkJyKRRc8f7fNyYzMFhL3p523f55E5Npcc4ADKu/hi1vp1icSLfbAO
x3n4130P+4OiGFmlylMEFwI/B2ATb/rttRBYc9Km+VKZ8iDlz7z+RonS3lJyu/S4
/QeiJEDsrJ+Mrfj+b7blof6vuh27qzoYk18HtZx0iHhfWChbUfnKGKQZ7HEIvvs7
O8Yh2+y16JqGG8a6CKbLkFbKeyW7ho+nlVB7JpMLUvnCIqRmYNq6+Xv61Ed4A97W
km/D/l4nBX8A+Ifkz7+YqBOiZsIyWiNytMz4wftpfmNw6fvLGuVSlhBYdcpq/fsu
urqorGlvoMlIN9iKfH5fmQ==
`protect END_PROTECTED
