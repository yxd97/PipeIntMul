`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65IfPo0CjnqbXMOlvD0yWlck1r9FdX7QeBjcmi4kpbNPtWFpERbWect4G/XUBemj
858ZT7WR1gJVysPOl/5M/3Exs+LVI9VsSiXCsSGqzVn6XuZHYA9u95WLzLLAMlVB
9sFquwGEqbk2V/eXIde1GnGwNKAjx7+hpViSDizZZ9zObqsvbsf9b+ceGC/S9f+T
VmKNRdqRreBrb/YF9zWBxYNCm10/0XY8MdjRCNJeiGFAywO1n2S9CFbaiPH8ymgx
GUqEdl3eHsZWovFafSzY9iT4V5/K860a7zqu80JdeiCI8urbzRyYIUNSbH/gBEQQ
sSN/Ag9hZrH+6yLU93hyuAImnu7FlcpqcUW+wVND6eCEnrpD8kaKbFUFcznEXltt
HrpIG/5+NOwdsLYIAd0jqXvWo1aX+ZM3Gk7ZkIegvOyCGOPbkeePLYVOJkNfLBCC
f5WG0fbtwb/my8UID+PrL8SElahivwidWSWHUMcRXdDk8OkwzFQfPVC21h9VFY/v
jNdUTPdd2j/N638chWJPRhf1HopIRq7Ww0Sw2H7wM0ZYHfyIGZlZFX5l9T+Ujngl
JalFtfGQ2si9+UkMamRS6aV+no98zQgmKTfeFdM2ytJCEsWzJCy7yI+NN8sc8Ivv
jYfrpEfCILqWc7h+Y2EnPR4TFygBwf0chE1iLhveFRSJsyCy0RadY7Nhn4CkAq0A
h5tn8IPm6FptF869Zd1FJA==
`protect END_PROTECTED
