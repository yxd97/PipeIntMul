`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zkcZiwFw8Lk9yarONBbXhkBI9swt8xmC4jhVhq8SMtktRPBW8T3EU5z6NjvVouWP
KZOTZ7nkGpC4UoQEb3iLJ9Wf96QuGkNhCbV/4jVhSibBDyuxnkRwUzEWeE4sCEIx
qdhhPNujbVAzsXCytvHYxYeXshWd9c6erFln6MHmsO5kt+m3T1ceyHrJk71ZU/yS
CcGMduBpjt0DzeTfX9yggjM45N5IGtRzJmGC1wmkVbHg79YergBQZ/BDP0dzsK1E
y5oX1dNFAPNry918961gJd20rlIaYvQdFu3A/jPEmLKxygBQhAAMjtznfYyyTEc0
nvaq6zhs2S8npmzO+GhGMfCKKyMoFXREe/mnyeMAYqumHF8arnXdKyJ9BflIf+c/
boeantVEv3wUemsxlZKhoQ==
`protect END_PROTECTED
