`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SqLYtD8Tay0sBhbMsRQx6vEoJuN4jfa496sDPYtfTDaW1+MhIC8Vxe0zO+3j6stk
HVBFK98Zls9Nz+E/e4AGpe4WWX5gJ60E70U2KamS3ofwgHlt6bWWR5Lp0HO3EqiS
qsUTOssofPuSJAUwgjg/J6VTFg1pifIbZBIqhc5dGVqUr/PTf77maSXRaG+pmGnj
Cxy0as5DBMficVHyL3UpFnel6a0hjqkZhIz4UtqeAW8aJSNBdB9zjRjSjpwdr8tl
BnY09pTN7DdSkVpt+JXqacohO2JQpfSYFRY/w5xW+Xb5XXi0OdFT6D6IbGs5Hhei
kGgoT/AYYWaIMaCYJ3xeMT4b8o6NFvalOskyawBrdO+ORg8K8ds3epe3loPjccC1
7n+l5G+aD5dwpZ5cjnYKFw==
`protect END_PROTECTED
