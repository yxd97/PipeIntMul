`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nzL7vCOCqy6GQL1PzAb1pFqn8t5y1CqHg4x1FDjU9LLNKLGNUjt5y4L3rH+a+zWo
t9a2VivgpSYaZBwscb/tv7GTUu7fRxjG3ZArsXDSX8p+gmO9adX+s2vh2wCxz4zr
A9FM2Y+mOWMeLxHjpwG6kCq4HwjbQmUcXSYPEw2IurjYIL8XLSj45j5vtf0mPcKk
XCKhesOMD7/rmCH4GEM2FipBgJTPdqsMhpod6wFaWieAw26GJbFSm4TU96NsMkaJ
uTHFJr5s8JPXqNxrUsu0/04PTaeyRTcQXjvOMk8fW5CpPdRu5Shj7FHjBn3bUsvY
qS/x34eyRKK3fF4XLpIsDHmViqyoiArFqnnZrCPMENu3wYKXXiNZq4NLFGIkVDff
GG9hNbyQ9jiHciiErRTyxCfxYzZ0m0Y0sdP5oBFddzA=
`protect END_PROTECTED
