`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+7cjRIVky4HeTJG9Vlu+7ZvK8+MUjjnum+GzfNTC5peusFcDubexrcKlHByVJUl
QsRnybL2+ZF+xncVRqbqKtdbat5GJMizsuu+JrJAvWrheV86I/16lcTQQJT0besT
V7n16LjNDWAwu/E5LUs6abWgr9RUVxOyAJUpyC2cDbK1ezaO6yOPBY/6TSDlrvma
fZbvKd8Nh9duI2qlnMsu0IlKn2lihT59QO3IAA5Se18y4lmYTxrEQyBm67gJFcLf
BSUVrKyuBOu+mGxl+jQDgtiimGptsZE65MJ1mBge9EiXoh4XY6qvmCsq9NXAV7Mh
`protect END_PROTECTED
