`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLAZpAQslqRpCzanQL/0WvF35+Xi8gk+/F9pzheHUwa44l2f/b59NUx0qrOhUOkw
wPQi3fH5EfXZeglgkhosqsnRVTjg59heXPDtc9uSFELmzBNX/GtQMtRr4DKRNJf/
IVSqAL+5RfXUc1QbgBUfNc3QAlDEye8N+MgtR58+2tyySJWBTgaU99IYnbZ1/khD
dBdWD8iGzQz5x0zMdRV8zFAgoDMosiT7lZewlGhUauIhRu+EvSF3EaNdagf8SuNo
zLadC87Z+Fk3lw4eYx+FBQIAf10lUUVdfn3LxyfYlcLO/LwC8OzGz8SaE1URW67O
AMJ399nr8pIokN0YM9XqU8NjrK8uU71Zp4S5nss28VT7b4893PmOl4wVpb4qABqJ
+G7htZBT6eIgnQHK9F8V3CtbCzOAfyBQNttTsmg2Eb/YV2weAF92yv8a4eyH8lHz
YeFYsoyJdOcRGOfllCRm5ANVBONFghxXqny2hBRUIZ3/KblUaTyYwkUJclhSOD0F
TRiiEMUtxxURtYHjzeYIPrG7vkPRTgqZJ7UE6+J5QSMF22GJSQX+ez2h4yPsoXhS
1keNZPmxCESQqpva4ebdjC+gQpf5pd/0hehvTkcveytcQg7me26n+3E2uX3sPwR0
reRZK96C13/7unJ4Z5fLCXzH/i6TJd3eJNKBiPfBoGlmWMog5F4lkK5u2jE2a1qi
CLRR/DAYzx8nxSe1zsPsjg==
`protect END_PROTECTED
