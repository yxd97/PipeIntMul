`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
huWmL93hD7CoYM6fcQodDst0+NZFEFHM37dWrmAoJQHnEqI8dDx5F9YlhT9Wvq4c
4wWIo5Ey1rYNo2ALvGzR1OIHbG34VUQJCmEZx5eEasiVVgwXNZ3hy1rddw6+tESh
1y6NwU+uGMxHYirTryKRRuE5G1wgi7oQV/QUejaLXsf1doSxoPaIFAHcLvAfoJ7Q
rVSKBUYZtMKe4SF/zdINjsC6vwcv2VECIokT2xazj4f4tVeBCngv6d5z6XtZP5+O
5fOgzWGUgtcYcMrmaattfFnH1/LoRcpuvQi/y8EGlShs5wSZDJX7IlPlQq3oVmx3
5oPM3zsuU5cA9fSRm7X9mYCG0fHSlsBRjqhXuBk2jqI0+cs+EO8RkOxYjfPxmapN
gGLVFmXOXgIUiQoPX3BrrnQY6fF1pYo8bMFHLFUWtay7kntMZsKgKx/9uBxDUj9H
ajGW0pvxz3hkrTOq3HM4eAMm5xsP9NMvEHK2N7MHMk3JdIzycVVA4a8s5MS3QEyR
4H8AmQ1++RHuCznAs9ydcFq9Gk92vucqKR+GYm/gfQEpe9tkocMQSnYdR469fyIP
UIxB+I9UmOIpGaGVMm574eaGUC5kzF2KZefDJhZ4WIdsqU9oluj8G7sdrYb2LQ/b
Iy//9h3ytG5gryL4pddFT2T4WA7DYOtWsMLGFMQtEefo2SJ5txqMKYCywtvx9Rsr
JcZbx5iPBpwX712VE5rHdwzOAigL8/FWNPq9Qdajttz0Mao8N4dG521OfgLyAKPi
4vc9cDUp2jTmkDlo3Iq1NS06h2K52AIhhIqr5e1oBfZwk5iE3VbdApF6eKL5qyaR
1jAtYEJkQB2lkMuMiOj2rcWC3i7HlOeZ9yJIg3Kb/WZPiLKiBzo6okvPHQGXJAFI
FkHV0l2Xr5y9n2pSxD9Ro8Bfn3w1anNvGxwtG1lPQdP45tQm9yPHHaMS7+pv/6o5
TYAF4ilndWnrqerbqNezHlpI3T/M8XYQMRzzy4c0w8a5oN5ARdb5yH4nMrp4F30x
oAxQM+I+gU3xAxXoKhvgALZd5h4dMyXmiojW+9B2xYsBnjOKxUZ1Cy3XgbwQ7+iI
9NFw3bvq7G64OG8szWIJIAj95l0jTbIJG+vc31bfdlrkmgMGLwqFSnCelQFb+2nJ
8oXXSyhwvpVQDGkKpV05KRjzoxPXL++TCP//HO8mnEK7NXBtUzNkJl5T/Zb1OPEJ
61y9QvUQhe8D+sY/okMc7fYtKmZfHkGm24uFHdsE51hKz4y2leEBpww1v4pcA8oX
Me3GqS0w5cJIXVfb2PQ9Ygd6nmDTOot03XmEJZQXDcnVYuqOrRmow1vdsZOl4Nnu
`protect END_PROTECTED
