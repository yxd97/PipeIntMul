`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ye1eU0hXAyl6oz859YZ6nCXhT4heS4gqYuVKNxfUFjTlYHZMNGcxN3uf1avlXKbq
4EU8EydL4j9j2CQ4XANAtDoHvSsIjgMWDtdjYjlF7Q0faeokUGcgLPZmUp/gkv6a
EdoQRNNNGKFFugIIEtNg1DePHDtlTTYRdTHuK66j/gbBrCkiFgLvTF116ORWo5Ew
UZ0teYI23llcciS5cvXNX2DP6TnhDADmRUxuKewzD6GAZ2zSeiRgjt2X+zbOjq3f
l6uMspGXACqLXTEB95xCDT+DWapsj3SurkA8ANVWNujFHuz4A0/1SLd9G+qhq5Z8
2B0zGkUCMIbGZbHA0SXpyoeIUjGpWTY5cPlQJB6s5wta79iAio8BSKB9K0W3DMzA
9/vFiWyPHtwiqSdC0OEVFMZyu6IhL9JzAaBEPcj9sihH3yC7tZGqGkNLMY9+W9Zo
LKErutUgcBLgvU8p8b+HX6uLMOVCaVbFx7bacl4yaoodaw2Np1s5sO5ZaKw0IvoY
bEvXnyTfj9GgGFnTLFK6/0o7LbhGcq+8rs69XLi7izs/LHx1T7w5YlF8ZNOmyQMJ
T1w8iMSq3zLrAwRH3OlavEsjdREwHy28TLF2xVobDoGJbfWEumcszc73jS1BL2MU
vwaFt9abNWQcUi3ioW6pJw==
`protect END_PROTECTED
