`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
owMbO83c879au8AjHEbs4N0LnCw+G6Bzc6o47CjpxnHaST6O+8tdCCOndB2EkYxY
4SHwzTZOKUVFEew702pvsMsiQS32JpSO0fR6pdBjGX1QP3vMRx26K3u6lgwLjQSA
Wxh7HBWGYF7fqTvCShLvQEzpc59CUho96WOLVmUg/W2XD9t4GB2izIErymkj/06a
Zz4jgMJVR/fS+gEz/kgo0kSShrwoMvL600hB6CTga/5kMq+BSRh84v5BLfedbfwO
PuKxH70yc5rO9/S0p8vyfnED1pW01sKbo1VjPBFa9bF+YOHoXmIY96PbcT2OPd5A
xwZxg6FydM+E1VSUobItnjzlNwQtur9AQtekUhArhZ8mDuIJOCTdmkXOtAudkm3+
sjf832TI1dFsxXSoABZj7SjEiAYBx6wIh3+GBs8VqSd/Iwzr5ETQP8+4pmvbRRDN
SA0jkYMAxrxp3ud/4NHo2Gdx7MEhE+4nG75jUg6tfDo2/d0P/IBZl15Fn0tOnaHJ
JyqtqJelA3XIur78i74yugqPUybaqv7kRAP1hstpM2N/Jm6hFxSCIyjYwplIRSwG
IuhTAU1E/tfb2hdIM6O7IZcAJaqxyteTAaOOOY8jhMI2lVKH6FOZR1zPhXhllEg3
ZKuZjSncucCWsd7XtgWBhIWolnPJDCmOh8dtJtix9mvZ1C6yKxBi+XZ3jS8eVjdx
KVYik0/NeGk0axzjXgeuOEms8bDd5pcaNnOJRYdXo1O4qOhDIGriVwAKc1M1NmrA
8I50LTA2McLsM5YY2xJwKzL6EYVaEbO2OhGThD7zsQuJSLvJP4IvV8Q5yCRQfY/f
zrGYJrebQkyy7h+RsXmGGz5qFM00Vl9jkFo3sX5jtL4VZo2gAT/SfyuROs5aUdTH
gui9/kgphyJTt4/Xq5NBizotIDU+m8dn7WzDIcntPsidLdDGJdbrWibE8V6ibgMz
PWyTNI/lgu+X/vqRYgKumfefa2OehktM5GDnFklMzCwSktcEWICfGT6uYk9w8Www
VMFSoBgyuHy4AxpAOPIiIq1dmtFPjxPI7iEBregdaz/7hasiK2N6WTVFMFzZeC3h
0dTJTt/ckfDb5z66U99o4r9cfzinucmyYRqcSfDJhVXEBD3NYmKtquvzpYQAMZ2m
Du/0Lmxr4Rbo+V2vcbXVXiGJB5wh1RCRTfHtdHqxtisWUXbD2yOGe3C+2Vx9LMF2
JnkKwsWXzEF4DTB74ymiGuUWfqlU0L97ova1ZATidf7CaAiJuHzdyrkjAH9NSsPo
LhcOPr8iLS81MeFKypgM0RFHDrAJ7pBEGYw1luYyfLIy4ExJGJWUecKIl0XejbTQ
U8F8m7RT9spDvM+7hHy2U6Cf5GFanDy4+TE3NS3pZgBdACKcdtIpi/Iq5pBAraY1
EFVJ7/pg7RIjpstvEt+JPfCJdRn7YizICR/j/35H4NRTgogPB7knY1UkSgnUucBX
HjhNL5Vetqo45Q0D4auAYFTEUiKAGyHqfD+e8xdKuVY1P25L/1bXbKkvZvJP7Tim
4DR/jiwMvXZJyNfTuSHUEysm8dazhCdltS2OSwjjX15hBaYrl7Bddr22r+8IcUbT
lY7VaKw8H6GuX4/R3cTv7gaVV88A8zPhZ0Dvd0m4lSBNYvMwbI8K9V3RSLMOLRHP
mqAeggdrVa2d+EUWJCjziDKPsiXhQqMAIzk47oL93VU3arie18M279R1kFmsBrV9
Re+c6skoCDcl7YUjnqFAFEDDRfIz2SSskt0eVATpCCZxwLQZAUDRm9TJlUHH9BWL
XRUY0Nv0XaoiiB7eeEXPkXY0bwJMzbFPvSXCO3svo1VAnkuVGXRI/e26CvYCxhT7
guEi+oytx27l1aKciaDk/Z57Dr81dgIzdwH0gbj8nak6tnlzq51SclYcZo5fad1J
9BWc8pabVGVYyQ3nzJrW1IB+YjyIqeM9lXBda8n518B0RVLNqMcR16jvlOP5mQx5
Gel3td6JO3NcPx4XMLeR6g70zYeUmYMLV+JySX7KwSX+CQllshKCNZj6KA5NVKZk
puoR2BtP32QlbOowdrHQKQ1vPp6KQSPU7rhh12S8iUrSEnhvGlHUyuSV/PXdh+tH
JpQWWV/jRi9KGqRV4RZuybrK4a9gwdpQa/7l9ubgX7kt8cWovC7z9Ey1NMCD1PfM
yXS62dVtcd2lndSwBXqCceEXG/gEo1D3KJTg93enmRs9M3oPKpigl3C8ZmhPgX9I
d+ASnDoDCQKyB2MBaCZpuw/QlPwOJWjDpTPGHRv56aMSkkSyuHNB7S57DaXlD8Z6
WWycSKPTaNZMbVEPVvSVlys8ZrZDsgSqWM7/aYIHoOjMuQiBvT6ki3olTjeZwQfA
qDu30iuQNgBXQAH+5IL0ynAjUh+77oTnCUiOZThHkwbrQWECn1Yv9a77hNqow+Lu
LGsBFjsJXbIf4ld/wcujvxiOu3QSJjYEhUM9ozj8/LSs//7qHQ5yeQPgWEb0eNBY
hD7j5DMFVcqGiq2OmEqRyDd3SRWjkbjMKO/vcZ7fIV9oIlUz/wR87YMP2BOBrUce
Xi/xOEoVrsGVN2JTO+lVHb5GYm+8IyYa6IpPdx0nlZEW/GFVGUO57urO8KQMRMTx
eOWi22H1KHs+YMUkhMGsn3+xo+dif9sO1m4KPAxqEg7Mgkm+UY4CWT63k7VBMW5k
aLXrIQ89g1/ZfwDwn+XVn43UdMEDRLZeILs9ytx2nq+tgEEssAgpphqjJCLdoos1
KCmzSdNwGiRpl7lUFMY888XgRoVdHRolLf70AKfSXNpDKXejkogR+PGHumAj1v9M
PlDH/fYQ8MAG4Qy77CIJfZL6vTRl4mlAj1vTWH6s2J38MTuk8qRb3Av8pjFfZxTg
ya+R02IM13k9wVjLDHxop6KQHg8Mn9oRg7bAcZAPvQHtdfDQ9Jy0YYBF8JGeWvby
Ii+K68c8S6vmSE+5LYspHPFUmjrLQSu2RamBZZfcAAoGqJ99uqYcuTNoTOutWrq4
PzP4rlZk6wo8JxgGyDgGK3ng4gQ1F7Iet57uGIBXV6SNULFb4qJM8/VT0KYpl3PX
rhMSPd5x46LnN3If9cD3WdjmIpkW7/eVwcqHFaTD3Q3OnLsqF91lDmzfmHdtaVla
HBCnWA7Aw7XH3VeY5xNbE9b9H1W0VGy/QNQomHcLMPpZmd22ughkBONYLHFzCkhU
HotziQIlHm7BsZLMYPeb78S9pyb/iHKNIj5Po+CK6+tOOhZxeMu5Z4/gAluT3rTP
JzbfDFu5gTJ8TiGm54yVM54l4XNCPUtydefrzug3Vdv39Ra0Ax95970yHqAbjj10
ihPvTD97E312sRotsQe0wK+BqkxmTw/IWvE6qRjgeOc4BblHT6HexSZD/EB2RB7v
dskFo/qUEAWVF1PsaFmHTAys7gH4izaG//buvG/QOQKJLwEK2/htMzZQrCaYcrJl
zOKfWc423zh0lMrPZT8WW8RRAhksulEX3uMUW3Vv12DBQkWBAbnvVmP/sBdW0di6
4W1tpjVGKI5eSWLR6hxGpseUnT2DrY4amK/0i4Up/Li1T05mkCCED3rX7WkEcGYq
X9GwivAZfXQ8WxdZkbBq7qSqPkYE5S6zqZq861VdnZoJCl/Q/npMOyqbWXUPYzxh
C8FvcjpHZywoB7fqKLIM2bYUe5e6v28Utu2ayMwIAGxqq0ZUT/uc09B46dVEvizP
mEMXWUMrEDjSgv5Dvepr+hDhPzeGe7RU6/6cBdASfqBmpzy0BPLOB/rin6Y3dbv8
KmZxN1D5Pki5bXlYpbtn2uKCcDI9Ue1a834cXob/ttA135/4cBUlGZ1T6AOokJFx
Mw2YOI6Lo/raqx8uckg73bZIckiktas8mVJHGhIQAzL0OD8lFDOs4Vej1iVkbZ2M
lduFIry7Gc1VtIanssN5QOSqy3WNZwc+qL9WoRaFuinoiTqoJ+5jYYP505zQBGED
gVQPvtbrwCF+ttCvWrgh6y1xk/wsfNcpEFv10p0+NMdGZc/b/SELJ8XtvFFjD9rx
w9yGLceLILG8clRsfmmqDPcNM+vJ42JkJ++p8QK5br+vq72PScSBrfJUe5Mq/6Bz
/7lm0oOyrQ51FY8Nguef5y03jc0kS1asCEaHJI9qiQczbRXUpyShlHjQgWbhO18O
yuSC2YYLWdqPZMPx1HzOs51Gwtd3dZ3bOsskayGYZxZ1JKz7fMs9A2CrW03BgJqU
QTXWXKyKe3bXDaWmDq9rPv0+lvFVd6Qvk6KHdmbYQ43Nwry4SXLxqtPUpjB2JNeS
Qo53VurwbQL7ZlcteTdMY0KH8HT4+Agp0/CuyUHqjJ7OxElQNSrOZW9/crx8KSvE
wuuegSL9DhN7WZpj4N/j9+cd9Kn1RiK/8pqIfnBDkJd3jC0Overaa7Z9ekLzgPUJ
3p7IFdl0NfJMH8X2aqj9+mWzs0ySzB1b9t2v96JoHPW4iJVV4rNvVDyvaTmzX42p
a1AkQ6M8k5422w8CtAJocR6Piw0xaMstNrVd4/WBcwxF+s2Yg6Fq8xn51qgkr9j1
dpXEisIiBKc6cc2U4vTPXdbuDSVTMd5Ejc1ng2aAoLaOOuoHHxd/sSKp2xD1kqGR
RnzLrTrDnla/H2gzGVImyk8BU6PnPj3pUjwtS3wUDNlpiMtgfcGg8xE7e6LEPB9l
7TcrgXPOX+qBR1NfocvCX100lX17gVZqL9FFT1Q3N9ysXRR19p8o5tjE3lF4ghSh
WYjVQti/Mkl/ZbjtTanKjydIoG3kAs+vvB6VQ6rH8MM+ETDApg5Z8BXD+AXGwoT2
r89wqjTbb0Jj/x1BpY6qjF8erzhIs9F/lrBZeczUX7sTBhwT8chifLDeseaAluAf
j0T9EzHznucnaGzvAweijcVdnpyV7yDYyY06yLGaz0pwvvgTmYYhthLlgFCCG19t
e9vf5ZfheotxNSGwpIbClcVwqmdfW8u1l068FUpiU5liKK4wgs37J8ewAAfZhzF9
g4KijtZDeWCu1BzLJwXgTCFPqguJfpn+FYwgfLHu12HFsC7dK02LvZOLvVVx10sM
jraafTShdwXHFTcT/nzSD/J72sPCsQhzZyIgBFZ0eDVDA+h8zteA6b8Ob+KJf3L7
epbSkoAF5g5waR4obCi4a+0bfm4mW/kRKSZPSYO5NoZdqxRBoozN8BnEhfneeaja
wsnCSpmrRmLn8QBcxN1JO6Z/fOflpXxbmWiS/oGDKkdri+g1TqLP9fVCNtZepA0b
NyVWxHctiox2UDNVdrXJxi9W5do8Ug4XOeUUAS50ng1/azClkDzb+vcJtLG/N68e
f0vrCARKCEQavFlBnnlZxaw73vTA44kN7DhqHYnWVC7uNh9CoZvJrKvR3NKtVAq+
15wFtV3amxAlx4IsCmBqSJJUuOBajKI5+ZnFSAhS2HkiFwqbg161oq+9UhcaZVja
4icX9i+H5w0XbEPs4qjPPefVceHsLlFInp/jiyCS1LqF2m8T48XoCj0hqOtXwqKi
LV2FxSuZsZySTsDxWQJ3yo+a7rC7iGEZ3SvjHpyf6Hk6qe0b5gm3FXu7ClHCL71H
Jbzmv8yRYJlAO5hCC+W7fnVg99QaUGACwyB0yk6x+YcNErRAzznMGzMNDFKi9oWu
wL+iH17crw8gSEq/tIIsnBzYIqfqFs1wwltUjcLIILewdTjIMMfrZqyqkjtoS8Ij
jxITQOH+55xX3LJzvI3npn4o9h6VwvdjHvPfWB+kSa9qHBXuIGlnzavPxPgFWKxL
vez9/HeSwbu1ptLZEAnNDDYI8RghP3Ol/MSEEHqSkQYFHreJL4CJvHgid3lYh687
Ya3Ub4OWtPKhtZRqIwtZu+kcowdbJOuiFkA5qoKTRwsqZV+8AodiRibHRPfjXGfW
2fFa6TpwXDNgagW3SjvkDs/ORYIrFRXNk5HyfvysYOJcv40ayYK6drY7inbAICJH
UXvOzrxVaPdcjNaWByM8YTsNSJcFrSqSSZk4t6oKCP4xhMvEXjDasCbXS06mgfua
/XWI6loZxxbK5xjmKfNWVBEHliAu9he3XE4a9hLL2WtWUJIE27EA/m16wy36WD11
sPWQaXJcwLVRMICVWTZVfQ5d9yc+laSLoHxWs0Q1nC7i7hrvdPmRVJlGXPfi4poP
DWWLU2YpZGtXrzXqGBGXijWwyAXEUmpv4avoxrGhrJf+UcaQ+NFQMwd8mRPycwHa
g7GVvd9fLvqVq5wqPwwdfRiU42u6J957kgmtjBsENhAeLhWkXjJYPoHADR3680eR
/UHn850he1Iguxikc4NFGFrSfIFWO2TCltlCLzWZ2E4EerxDNs6FdfngyhF96Ltw
86kYVvNxAIMF6cDjaCQakYjrs+2Nmd+g85DypjIsOm2s6If9KuXVJA9BMvBbCoaC
LYWHeJfeOn8VQu2lPkYKokPuazEs4Ca0/Q/dPbOp+6ubOnPYkQolaYkySye2OJIo
qwYGX682KjdVUhkgtQwruzxMGbyY3yG2yUzecuf033yMgOm42Su4r/k9SeHs5fa3
JCnZ319Np/LF/tQyL3+7248vc2K3ANYlM8CkgLbNrqU2u/7IfveuwvVwEqLMxyEe
kT1KPXVLE/V9XtTgCiQA0dGL2p0vMqRxqgva3zT4eETsKG7bKDxHXGMTB6od1She
jOf7WiDv2T0C7gU0aYl755jti28X6CrVGPlpF5zkoGpZjT0imqMEJA8FrF1Gq/Uy
qmPZ5bMdZEGbhm5KLfME+8NbnhJFOjyYkA0/3Ij/HBcKR4jeYNOhD/tsTuMuVYl4
87SIjcOKknPu+DSMfIO0eKy8fGiUbVUtJ4iNlNoAjbVqADNSSOXDnbIXlbJWMLbX
al0aqgIrZVw6qa/1A6eHXKw0U22nXM2Ua8Zo4lFA2tsBhtWsvTNx6RbTPJMEIjuk
EFRTfnwJs99ixHikBOJQ7h/evjdMLRam7dAkE7AhS1v1YM07TeheCFwwl9I59OVv
9h+17L8TQ5yQbno+71dkSPJuEWTzxFrWEd4yL/fAronWrazClqmZi9GZOFNjYype
32Yc9CONdfji+F3GvE1JUtX1uo0Sptp0KrDy+7Wg4oTTxpYSsZh8fm5GLyoomUSi
QlMqV7LDO/1lBp3HURpfHxsKY8owP1dfUBAvqo7RYk6yUT9+fL5SLK2vgcKwW545
385bZd18tpS+csjDBW5jzhABeTxLsay+SabyysuY2qYLy/kI61mCL6AoVIkbTqgs
qGZ2RR0ok/fUl/r1LpmHknwnC8lkgZoEfa9LTJwUcOVhPMlGVIdRTu/lybdHC4iK
325szznLDJt5hGFPJE4X56VQzEIl5VdlH5H7q0T3K9n6JCy9VZG1HMbzcjLEvnSF
NlPLwX+rZS43y+5uSeDd/6U8qgKIpcRwzCy2jJIViunOf3blelbW62fIlzCwO4/I
iGaMJfgWbBVGbm6CzT3qSlNrURBbgm3okSfpEbg/LGotb6xi92fb4shH0TTKlJDd
dcY0E6PxEh4ZpZzivUqGSvqGKTJZIsURiYCnPO6u9h4toTSzsMD7dalhLHh+3wBN
MvgGunZ1yrZWI0syXK9f+/gNqp/JG9FmFycKbB5XmAV9wOzyCwy6ip0ane7GNzA/
jh4KAkZztnFFUlNST+N0SMz35z0laRzgTNuUHjhw2AeFndA+Se9TKrkWriKDX5i4
egVz6K8N2qGU5hx9ok3qkFogtZCRN5NLaeNIpfMLI39HQAb/kvADON45J+zmRt31
vnSeQCWbjJZf1kxxPkEwesabNj0PQNszKKT/nnckzl2f55hEl7NV1mHC0M+pDOQS
ZZpotvzHbf5nPABfVjAcbe0ZAK40oI2MtGA6gEkJbxyB5IUZ0mSnhS+piJOz8Ylq
h2JbJqYyPmSNJvyIiMeXcSdBXllAjGUwA73YcxP3tsuAx6mqFo15PJqfBAxu0NOI
NmywO7E/ohhSLeuE1+MEgPtAc2isqcKC/6FF7IUxMwerP8yDqLD5ZUZon3sUu2N8
rb87t/ayizOJzaTWaKYiPle6WGgTRydEX0+9sdvERqEL1euYg0S++Ex2CHFY0IKX
hn3B3DE/NlaHKzwaaBfOyMNz/EEUEU3E3aI9MzBpd7i5pzqizoMurBqrtCop3LRy
t2ot1Spg2+5/65UsJobfRRnshIGiqEJdCZndW7VpTgHI234kvrlLA+kkrgR4w5gC
6Zv0OnIBUkaZ8Xhv+rb68xC0OQsEkmeObfm/EGdOh/2Nmil8tOfgW0B+qQ4BijYe
nT6BnnFe0nylkXLRArewNz4EMkFxDat9H0X6qgXgbhsN9aRl6iumIlJ9QEXUOHC0
qaYi3rAjgCbBBcf/sc5ER75Qp0RqyT+HKAntR6C4P166iVX0Lm5JN9BE5/Mj/tcK
JsDrY6vVZhpsWftYG8L/DDHLDmVJcbw9/UDOR0ttWbSqkTUJjx+vnLm8DK5VNDOG
cldti9ZLPq+TiqesRUapbER+A7CJaBjo/IrtoK9zc8LCIzMc9J+NhrRRgTtrecIR
iwlnZvyx9Gma5DESCI/lvXhtn0K4ujyZ3SzpYJDlS2gnOVs3OQ1SdZC41p2HqioT
AyHqjMp8ipZwFfviJ3Zsl8PaaeLmAiHxX2dbnXZGE9GN8wsPtU51DuLoVvUBvAPE
hphxp2ZuL3itBl707SxJRl6m1FCQejmUt/8ayr3XKNjrM1nBwQLAvhVOdlMHNLzs
IwdA37LHdK9x/igAm4OQYM24S/KJWcZfMqFt0tXM8XZJKc4NVBYE1w7ayYa/mmkS
vhodGOF/3GdIt5XmA1mwE/waN3NUyPeuqGBFuUtft6tY8EzsixvgEF5LV2OvZBup
aHJ/abNK+rpQeEhlJcXG/AZNCn9rAkXHY6ddiYdNKz3DU+BxyyTFqfy1aaH1LlrS
Zsaop67Y1Ho3h7W1myAw9e6JnGzEgh00MllUenatgOQ0Fr8zcV5eSRPIN1gRsB7M
coY8WC9y/j9XXww7rbaJDhW5AVaLiI7deUk6ugu2zxc3+gF9RAO7jFG3J2bnfL0U
+M/1fS1cN/0RCYCwGSgM3jchUTDUqDnmbikVi5pY10gv1ZtkPrQ+NeMIDKhHti7p
An0KdAZE+TUQSIXsiBvAdgONtKGJEfoqfdpwz9IeHji218UaW+9K83Q06gAKZP4T
CcFZkoxTuZ+WX4QAXFesMz0Ib8AqkRk8DFm6eWiHwdVgV4LtN9VBjLzeZGkGVQQy
tZIpoKRV1Qgu8G/XygOwDFYyKlDUX+hg1jQHIHMKFaGdMeXgNQGFKowb1EyPM4mt
z6Fh87fMMfPZmC59DthkoizUZU+iNJa5AzAMbPqmD3A5asugrQsnp/hq0IkR3yRB
UdTzctQ8mfPnE5M77bunYkI3biYHXdHpX8zzOyubXP4/zOizcIM9gwiPdLCR89Dc
H1QR4kX+9MUctGhvjgtE2zdvoLO2Mk1x8/GFY1FMNu1ksQHbRVOQxPC7ZdE0Ee48
QkPF9Wrmgr/2fCKd5cnap1pVhB7Kj1kKo2Bri+pnXtEYuzBI6LSMataXITOQS1fI
wswn971zijrO6Isc1Tp0zsHOloBvzgYgudDoCzeMLsj5H1rqxh8XEhNWPD8SCRHR
b5WLAsVa5Luj/mQPpRmcSvTIDrDS027fCA7EcbiVoggnaFOeQL3C19LuirVSkg4A
jYclBkidlMQbsCIOt9L95ExjKmaxurfjUDE41Qdnd3Wq11NIr0/+iAPClBEkBzak
K7LZ7kyZry/fK4mxP0lvIVtbF+H6wR6hv0keA3CO2qzAfn2djFWGSMA2tLRw3Mfy
DAaM2e7hMlxvFNX/xsBndLbs2qC25nYaZi6FmdIcAk6SaNfrl7kFGLpKq/xVaveU
ouM4XUHD/0nyBIIvlVXWrR5CcdoBdLH7NbbZTToDDKbcQH95XyTr9jl20iGKhRDZ
IRU+Lpy95wyALOUiTI42EGNnSU8IKnJAdUgYGTkxO4eKY1MLtT0HvIgXcw31Lq8J
vEuUTFmcf0FIJbUWReR1wzyJa0Lj9Kh4kLT3A4oYWpQ5I7DJbg97MpkOlkh6CiFj
/c+qtzern/2DyHQRHVJZ6ubzJNIZm2t2FUA0pqtWm3qcpMRDIsuHwTNun01SLoSX
coyGF3+wN+v76uwniRKIiz9ijQTV9cBIjYAqUjLLwFo1K6s/Rntd2GhnJ5Q2NADN
F1qsiMlPJD5FOuOTeKjMrUsCuXYtUWsMgjvr+N8ETWnvac5nOS80HCp1/bD/QDbM
lYSEyauNSW1a96DYZvx+zPLQKXgnqk8qYs7OFS5KIj4udNsgzMjOiLSBcoUBosR+
E+vOeWUqDa8FVE05nFnxhyuEfqIDh4skIj/a2IZpSmDkQsusj5dmwBBwTFNlBbev
efrXgPOLs1gAc1wINTJCBTOoW8oe39aqUVC/NRBlG2ZaG8XtjlqvKPTlVcSzxP4e
MnryyGFcGIYX6bMY6k4OAxaXFb5JDrQOPavUbcClI6Rnq3xnlBDtB2BVi5CX+aY8
L8/CMpdozk3ajMTah9xJ1oLdSdR9svfXzu/heD6VCjMnASQO1jRYp+SRKVqtHwrz
Daup5jRUh1Wt98LolcNFrfhKG8f838g+w493Lu2dN/mttdkyS8MK1ne7ONvYOINp
SNQseuy/zHgiGFWqwKy4S/yqAGSCf9iVfG6zIbWCCNc6j5KI4odaTzoKaBEfyOW8
BtGG2MkK3ep/hjf1xO6Px08FT5adRxqnWybajH/CAlIIL4kV2e/QPuyDf0tE20I7
JPlLE4Az4wGM0ostse0JV7XRSl4nhWec/mLt4b5ug8FYOOgWJbeVmPAjwTXj12ym
yDOviUnEPNxj+7AU40cTetb0c7/YUsxcH7IPe7FmQehWGL9gDYyhYv0LVGRchr65
UBphmwcA05jYa3/3KYNO0vojv/DbtzxCIl1wHvCLFr0YhOKnNCB9oLuoZW98KHSc
vC++2mV569Fytaw9vgWoJp920f36ZCuff7DUFaTN9PsUppENPIkEN5fsXZTve2fy
ce1T+ohEMlJVbMlZxaHJzMJG+jNDxIw05ZB4ZUUJLM7e/kGPUpvtqmJtZwpWWbZL
vFnM3qM6OJThgvtxE/BHm0xrkkayh/4fzIjMjkyc7fhe4PIFExWhI8QeYG4r92uW
U7kEx8aF4sxXr2KvxB0QWq9+3zWXnWjqaN7JcW+5oi5qrUeF0Tcxe7V58lBeo7aX
l4yhQb1OAy4mNi1DsrjixLMycVCY0kN1h3tO5qVHm+bj5hDMDgdGw0fQuF/yO6sh
8vLnzHgmWdDrdW87LTL9LZuqlwR11DbftSy2/dtakxjGKA9VrKqi5Ig12pDY6IPN
QqLV9msFhfiA/lg+RhguBCgVytzGu7QnrMMPRHa0/snqZWJcX59NbF0qzl2LwIq9
T7vfTVpxUHPfQW+C56Nnq5imOfMQ7PZ/0ltbpJR21lIOxJxRU+xxqwe8dXwuGFWi
cD61ja0URzFdkycGnLOQVeKZfBiAglSbRMNhDT6Sf8IZpWGqZ7clSZDAkhlt1OfJ
b1Ut7es8+m26NClRdIhQn2jItTjpR437N/aR7UWNEsMsQae0TapgVW9AqY1upt+N
GQLuhDEVNp5IHAWWw51FIOtQALNKv29///fcni3BOlRC7rqni3vIkeLeQU5MX7Vk
TrDvebR3N0La5Bh1Hw4tWYks7IP8vCG9j9NnV4e7syiQFWYWWu9RlklvRLGdZwhW
QLvLJwcoUPBYOrV3vyKZl5gwqpY5n+cLWQTS8u5xLQ5LgMlyfC6MS/OGlzGwfSMU
iJp4RfNPDGdx6FT/JQsmQJaKPa4M+HDLBLuAim5jq6ufWPiBGsxnFlqg0Cf974BW
Da7nW3bL+RdzZLUSyJCj5RyiIKVY1n85efzf1o9xsnaEFc8hdIimQnTYoc/55l3/
iVR9DiNRDk1F7sCPJy69RFaZCtX/0Qtc086Bx+bRpqEFa6lEwVA04nU5FSM1/eCW
vnkUubcIM2cFN+iOHe0KJC6bKv0Dzm1wyZoFs8I/dSs8FJKeTjCYk1MBFFRtYvH7
C4IgJTR7+hnkXMyyXaEqPebTi4Z+GOm3stuasuBWj+ApAgI75n9Mm+Qi9eCZ9Fvq
PFHR1BLkKnS+l3KFO7YTINmwvVTi0zkL3fGov8QWCKEn5SoBTU+hHqvFJak2fg0I
OqNHZFUH1TI2LU0Ps3F8zZfLeLNXpiuz2iriLFQNS53sEbryV4X6tDz/FeABnKwr
fLHEQZHNljmih6XQzsiZEM6my8wqDSHVjS04G/sDnlCWqHJElALB3ptEuaYk3UEQ
khzStWPqr2bhAk2/mKE4lmm1ZHWz35flucv001YPYeDpSME8yEC6al1j1iPVQfl4
/h46Taedu+bgtr/IfQ2MthwJbs3NIRFqbaJ4cUuZnCxHPs/2to0D3qWCstcpdPr5
DFovXB4VFOPPhEWaHK+mtAGJapRgm/ZKxKOd0GwO+Su6UO/2mQPYuw/Xvn5UvXdq
YsWkMpw2hn22siXbJYhW+DV3os2udyGhGReLZo/nXhFNnov8I48jmbSiHgSbqo6c
cZXRbd4cYuU25nArZnBPHvp7duG5xPyr4hNfCphBICSS4vCKdA2v7vD30/5bznu2
EK6O5DFMXdyFjyCv43OgUN3NsvEhn1vUm2QGgWH96LhTFEpGx2ZvwHkviNzJMDW/
wpP9LU0gLFfoWMSRNqg450x1e4WeVugHJTcP7js0dY4DH/vthMHXppClqIymRZ/0
yTMBa5cVjc2JqtFuVsYyNh0CMMYGRLdDUdQb4phnY9PQzvtLA/i//gTYjdWapoBy
My6JxwViNst1dywP8Az8wTS4pfPBrhyx2ur7e6jX/ECqfMuFdugnjHoJnhhYYtVK
kcYq5rV0+dHl+dyzcJNK9tGgk9kA6mqci2ap6MVrxODpZVdmGhq0W1O4MUR2A146
dXiKjvOi6URycig41LCTJEXSf91p/E+bluSqmFbhvVdgEAA7Jve8L3B55kuCny/c
li4IMHUbR8t9rYxc1dDFOwLWFMzMOR1SrOx++wzAx2UXVD5uG5XhuNisF/hy04bH
rS45OtgEcd4ZU/pFm80WS3AiDrtEq7o6mzOe0BR+Vy4XoTnc75+OrlGz5Gg7y02V
mM+QjuRvzH8txEYDSxUUgvVFFwQ6KKt31sN+Be7S/VqL+/b3a+0MZKk4UKdVEKaG
DIi0EBrNobhG9h87Nmx4tCX+MDhzNUF0lnSa8EFQmrLpUaCLBIklrg0StqFU/qLa
J4i5OsitJD4cdfTWTETh8S5MH7i/QANijq4Hf+9fU9jPIFldbMefbmtWTQmY5P/Y
j/pq5b1aHyO36C6fSC/khazz0Ix4ZOX58G0EFcDzVBI5vJXTpIQBnBiVwDIUpoqb
GsCDG6z3GAk15Jv4+t2eDHlVNyk+BCkz990dqbQ85nwdZWNO0JigKtOha1UtdKiu
kGXIlS2j75lkwRJkkeso/deUVE5/ygS3cqkxF0DlkzNLIjgs8e31YDu8VZXR0v6Q
0YpDPkAZIHxauCizIL4Nv99+YNVq9dTuVz8HSIxzsrvIMZLM4JT5lZeiEvH6b0RA
Lk4cqq3XsAu4WogQ2jqIz2CbM8PBKvt/lLwrvqQW3Yi5p8Tk3a+CUVLgsasmm8WA
2EpFdof4wBNCbYHmblSgtUq00cfksfL3H489sMAbyQJm3DY7dqIbHDZT9mHnUA7n
doDHZeAyxAnMS1UcMhata8IlEezpH8vfO3Mzss1tOT1PUxccEo7LhRsyjS2JsGrL
+QeljAuA+DR7EUHlLLn1Rb0nn+m3GAgC/L1ZFw8+kG6ppiKw6XhFrqlzxnMzYI7r
7EOfM/MBDKVIowjqw3gJMPOwbzWkneUOyyWk1vKZGFDIdfLR3dnURokxmC1VO9g5
ro9efh7ONz1PNgtK8hAuC4Cxur2KJXvOKTLYn7hqj59zt3u4uNqi1y5KeC5fd5m2
PRpbMdeCzvfFqBOLjeqF5KpIMSmP6INARD8NUiWF1InY45ydpAht2OLas05qnPZD
Z+mCFY0Xwmqi/fbscgAtUK0aMk8mWEQ2VQEk5wvFJpoexW6YEfTyiYugtEU0uFs+
5GJ4DkvHu5oFT+KNtI3N5Sd0V5S8pN9MLBuJACCAV74dPw7RlzjfepIYr54ngHBb
rYAUBmk1dmUX96hPWXW4aQk23jnMuucA/CKrvHWQUnYuri99rNWfNIP2EjimXmQ4
cyY1xnCnMp9J5IFLdz45886q4T9A82xiQrOzxLOTUnV9kA/S6z6q6wY4e07VYPiP
WoQyhqC/n13FnDFZnBDLPZWFEJ6ii1EzZAFKg+1Wjq/Hx+92PLV4P6Qgvy1eO+bn
dTg56oZktH14lB3pw/VMmTEWmomPNqG2KUBmlsOB4uOm6dR7la4GonAGktYh6vDU
YHXG4QX5mJWEawOiE06UFLWLlGp6L+3WCIMMhdI8mn0YYvKFFx4DfquBSXeRiUAS
NWjM60fqJR0VgPOSszxARX25LbQouUo5aomIikQotualHlRfXGr1MLcZzsOWDlQ6
Nzg7WmJgnHbNOYqOpndxCyDk2ZFSFUsJY3eQtF3eeHG6cjOya5Td0SB3DOmrFEHz
vrT45/Jl4r5+hGE2+MyZPGHN2baixOj2gxyFxHPQBQbOMA7XUT+wkqoxE/jxLi9e
HW9zYqHqKNt8cPEocxQFjDMpGIM/IOqZfbm/c8y3M7kNX5KvCDkw8UUclgLBaEwc
SQ8asGVXfk9TDoT8Z6vh04I3RqpQINWDTM1vtV4Wx4jK3O1tBe9KzoAGK1h8Q6x5
NFeI7BoxMHfMbqbjQ50gkl/N1szf/WTWF1WzdFOhUVhZEY+k63NPJ0UGEkqddjoX
PZ8qOuSFErv2nh0J84F0NygJBo5JQDz2FwklwzcG1vl6oLrS9q0v99AkWOAvdkWk
05iX1cXtu2Fp45Hl0SuLCfS6c0sDeC8mbTmzgnEKzpitwoPZlNkQDaSRnt4KIGvV
oQzXhzCzkJw/sULaxtHO17qnRywrx8DnUvJK4Qj2chiA0PUGseTR/Y8Bd2z8OfHA
0TOLFWjwcORusqTIXBAzl1MsrNk+OUuZbkPQhMhOumQf/C+GFVspAZevnLx/RxqC
GIh2VvxHWC5oraTQXnUmiVTyYT2VSRabxoYmRyNqMsJoreKhxeLoBJTOMf8HJ2KJ
8OcRd2SZ1BpaSmfYVNYa89Hi0kIz07nM2ZWT8ABOHl4g0kBkova6yHZ0smOCldHn
RiNGLXmjajS4ItHVV+1r81iWUFrZJfWQbAL+gXKAUmXmENZVLr9yX6JO74XlYoQp
x3gQkiUAzplSn06nwfGpeiVyXCXBL1kw2mViDrMnOPsXs+zGQprVBqyFnk0olaUO
tFRDy3vwU/d83IWlyCwHS+7X5vAbx4Rx8ic1YgDAT3+2FNY2+gujdmXuyWrM0mHE
ECaJX8b3idn3Uhr/80V17Se0Llo/NKCl0tBWQBh4ncCRn7Dk0UT8R1dsMPdcJ/YW
Rjw8kwK/PUbm0PX8xbxQux/pApclLCsYh/OHy8eLE+iCniTQePft989Lbbc7dixG
1LR5Uz90G0DOsE8Cu8F3d0plyypKv6Z5B1cizB71E6gulNQs9RnOhpX7vcr6cqxd
myEw6ubKcx0iHD1W2wzs5lZ6cMqlHp8emFcs6n/VPmm3Kfk1pSFyYBrl92s97+T0
7PyzQReYWko3HjEn54NMUMw7NFLzk2V+rlRtxjsK3B+aUfCVOTb+wNosECDziOw/
Euch0s/O+2sg5HCEqMShaMco1Il06ZYIfrQNsJUwTDYKBm/3E+QmcB2YGRzNJCK6
KopF/Q0tEL9ElneSfRZdoOlvP7mSxi6vwuNYRvvaZfU2Umzu1odh4+cKmj4hcWFo
SSzWvMhYl4uW9xI4D50q3/egWsLg3JiA8R7Wnd5gnpRYRE/BtNTv9S40zSIeuk5k
xOI2ln6jfA34x+CD8SOC8Es7SVG8+FfcPCB6zbKBEZ+go7TzlGh0h5wd6W/aXOiH
kt7SNAj1hBxuRFnGpodDP0La1WjnMrLmNJ1vShJqDrWzdAA391Vhfr29XScxk1uP
JcTYP0gKjWdNKvjLSm+F4NHKBg6Kw3O3FJcW/+AxcfhVjQIiFwqi6Y0sN1KqOTjr
G9NRNTWnrNwM/esUufCeZuXFlTUKFmL4nnetzZ/kQ0jQ9KfhvU5hco5EwEarUurW
ZGGrPCFGET0pnvkmnSvlYxeCUlwca1sluhN7w/lUc80gxi1Yj2g+CJUyfSQGpeD1
1W3p6k5gGp5dDaGyt3iKjE8okhEachuKrc7BovlcYb/0uO9Tdt6GX6DrXjewplLB
ix9WGMnxNjWxuVPeCcgAUKF/Czwfx9UBSYDei+A5AVKsTJOO1fAZzROd+3SYqFNV
8QRP+VTG3q++3AvRAySrXXCeWNqAidKSnrMton/9o7EA7LyoXlba2Zu/n6ZwNBON
iKznwiyJ3/GmhkS/xlVh17YQ0xWCvf41TsYlHy1H9NxJKef8lKcFIiBzm1baqq/Y
3iobHxz5n5oNoFhD3YTpUiD4TctRjc/+WuwpTxsFuV4Ve3+WFyMsHDjoj6KMQE+z
TYvr9PuqU3/jdU/mNzRcNa8iRtH6EYQlJlGAQ0Yl6QWwHu8KKenhyE9jXco1bh7+
eHjqpoQsHaN0KaqYV7rtAKoIuzcPnpikOM6wr1DN9fCQ5kRqty5Wnp7nE51e8FTA
OpIWq+bV/7N01xjbmiw9JLD4zy42qDlPo2dNha3PqAP3NffBQ6iFXfS6OhIfrWqu
59Zj9E7SZDmxXhYP+3Af7XCxekLwHeGmDJ4yMHUHGTlRmRtM9FBSl0JmasVZUzwg
lKU7UBgosQiD3sgUQAxBEJfnsCbzNh7FMg2mjST98Zbq0dARPU7/jw9BlQ6u/blE
HpSjvnqLvNVNW1AVQZnyHEzCSU2lQ3B2Fem5TiWmB0H59tffZfbv+N+32m8VZ5ow
F72Lf9JBAubG3RKYP8HDDbGrOvj13BZ1mfZmIAG0scD4u5o6l2qgrTuLALxYtt9C
1PC1kI2LMEb27dVHI17SLtYad7j+dUlgZnqWarKuNeBmRyoqGAFqERapKnRRASX8
bjqVo8IuMU+jmZ2BlO312rucxgVKWBU9LUlY0AfshdlY5a2J+1npOlVa4d+DT7j8
hXtoR7A+x4GnDG3cS3e9Or+KJO2rJAAOr30lHnP2UgloAZwg9/r35VDe+DmLeE9P
Ni/tKyc6y8/36MJMlfUWUkaM+CzpV1awmrpaH5CpRkA5i7lNnr1dSDVL3SVxaUd+
6zEY77iJZpPQqYCh0K12VIbtZHhFUqgErw3RteJKI/cywq1ZEi0lAsqzZEcSbP/e
iu36eCP+3gKUZghxYOg2vvGaK0I+69XbJoZWgujZ8e0UzVkql4hKhEAWAEcXUtJ8
9p6rJozuuoy6xjSfDHipnqPnU9/1gfHP20m63buBimSYajTLeRdtjiswzusVJ/VO
4se1Issy5+Q4NFCU7mTj8+j1SxNkAEW/uxmOHE+uvhjbDhJlu/WvRe0K4NDkQJp3
J2/LxtsfEIH57M/hTBraSq7b9u2qCdtG5jpCGNhDah9t200bIKuHgcBrhxuhTh/m
Wv1+0JUgcuKNH30SVW7EMkEvAcX7YWs47panKvI+8/22X1YjAK4/VlMaemgNvYdR
PjshJI/IMR7WSIj5BG2ClP1hRDt5EU1JJ2vbmHYatff7NmTN/G6lGDQ7ozAJG4Hf
o/ZjCfJ3JJBTW4/LoegPfLJXQF7BsaSXhJHekIgLy5L7lWqU1TvGHpvGw9NPo7dA
+ILE9pMBwhvmLI74URrPOOzh3GckK4IdB4xD46o5NTN3Ryye17eu1O/TK0ra3VLA
c/+X6S5bfVqtnRj0yU/aC7PKUkX8bzZNOHPWBAuPrJ9SokJOKoT3ub/KkCktrr9Y
hfM2opmhhEvO7wDEKCe5ykZOiYKdNXab9dSR3uk9fUAF5V0wldOAY9PRFA9npWXT
8rc9mGGpvvUY2iqCYChbyiwOTk8S2SAvEc7uJVVPwim+QaG42qr+yZuoMaGXkcBp
k9DyDwnv1nu8oM2F0a/6bUb9nHwUDnUP7R2x1VVAUKGiLayPw5KEqX+zaeK29Zg5
YjFBv/mAHO5joTDxFDTctQlztXRnbLzGSeTGpnbGf9P+uhHH8sXuqAcRSPFiHdUa
DRn8Dp4l3zSfGonbOIvIpCG0vIypE0JktLd/1bArIFK4trc/mU9UlrmjsDUgh1Dg
odXCYmj1CaKdh6IAv/W9X0vMa3xNESZsx2v1aKywDklPK4nGfcknNcjoZ/5bvKFh
s5Z/W+xX3SI48gwfX91z2nPOVcztkdiilxVEnQmkxNCxy1vXc4lv06L8kK2PhBN7
+B6iOFtRsqIMi2lJ4XRgjWekB9YPSP5equdt5xHwsdKd0z4Ep1F51mmcCchwOqFh
pUsiA0JzPCfYQUq34+uQ/m0n4M17mFslCJ9N22EkUr8tecFBMqFUyYdvnBsn63Bk
cyeTlW8+pUESnTcqcOZ0MJhRBQcznOJYvsrmzKu+Tl3weIyR9zrV267aKbzLtKR2
yDPEzv/Zl1bG7fNwEC826lsrEOPl8kvW/uOEjYO6ok5ai+vFrJ4DPgRiwkI41Nsz
jUTIbpDAf0U404aFdY1ENTBA6+q1dUgAsW72VGjsVYM7lHy4yStffaPyMhV2luwH
tVW+C43k3YiIR3Fgu+k1K4ngI920j66cILgLwghXVmLQepSKxhSgU0XzFRiAlAZQ
p9SgZ+HSNeS8oFUPU1ytzkWSJTOuJs0WtdPhg7tPzxiYssuYzAFvDhoYbE8kRtgR
1IISs4zJl1IpGO/JDFI4QO0Mol8CYXFPlxEJzSDoFOA1xoPYPpqQMksvaDS/5uwt
zZlxw8/T4WV/Eb6StavacT7GcxHRrwx6Wx/a+dnMjEV5gAaj4JW0iVZ9xaxOuY0d
15k7zSxu7A7vopjIz0m1FWnGx09CFDhLADG6/Nwb6He2uiVctuUFvaAM+Qxc6ifG
N+CNwlXGQ5OQ5cI0p744jLHxxvgKbTM+otlDNEw9qs5AuTOO0Wua0MQn80bJ8rUz
dYGJ26Beof3o+Mymav5W4P/7I7wHjrB5QihWhn5aPelRJxxko8c2LDiscBWfLz5N
R82mBti6itVemKzKgYWS1aD5TFXcwVWefnkjjxPTa1l6y71ubO84J7jXPMuT03mW
wOOGRXxFaybGHyqPGBw0QoCvIC0wjttvi75cdBfKotLY0oSjpjzowayD1SftNtw+
wTNNG4EjRLQUDPGoQny1Z2fnpBSXdyxMIIvl/20h4dxBZCCcC8F2ZKoxQ6pLMXy9
SAV6q+NRFvHFYcr1Pasu3k5REbCjaB2SmuaUnAfYiPsDPopx4F8Ix4ySYPiSwCDX
7+bziWzwGtZqX80Dqw1Kh08Cr/Hj4AUSbIdyYixZZn/YQmtRt6PUwZNOnaobKTHW
wXARyyp9GPO/4lCBUnrKjd418zd1bpPJOVQDFvkLyNrsVyUlItzI6ijilxUHY8ww
50qYOPhQb98takn9aAHpohhfcyZ7c2VpALC2zmH+2AyzpWHsm5q5R96hfqNnoDSR
eI6dsYKUHjlZ/hEB2AcqgtcSX0F4i+EF0X6Wjuv5ZDTuPQJy+9vonCgo9opBKZ9B
xMyJ0g/6A+dHODVBAsSHlelyaqZcUDJttFhmu3BD9Rqh9SEqo5EEmykmmXySSDr/
`protect END_PROTECTED
