`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IirjrW/e2LI7HrAlqKAP+Y9EZSFYsnXRfdpdg6vLw3jJxlVQpc2blaD6uQZ325UN
gOEug6egvbI1mc5kfTMwyg84rEeI405ludOlNeDJ/t+OFjq/BPAd2g2sGq9U7bJV
n+g5cn4zl05s1rqwNsiB0mdBFhZu59ED/JoT04lz0VAjRv9EipGmeANPPahV0d3c
5H+sOMRkgF/srzCJxSXWHVeXxpHZFxBLBQVV4p32aJ3ktr4Xkio6q5iKODEK4rcO
2lAGYVRQJnOw3eKkA6OzHvZIds0QHeqYvzPE0lhkAp4MqJp+t2hwRR9sNTBBUo+y
2i+oH1/ZwTueWJR4SJkeTbPZmA8herSbWiLq+e51Z5xT5SRnRzXb1tz5R63MQ3Je
YwdMQ4hSHcBsIVLm4oVJ/T98V9hdn6Dki2tQmREQOTuhMgF7hToFmrnKsYrjEM50
GklDt7bh8LV40OSLf1KturDcVlExmSgWsZ4w2iLC16iQd5DyQZvXbS53JNOa7Wyq
S8QI+NtT8o17fg98hFukXsFyGYC7K8Xp8LLSO0f0+IyILQSCWEV0gxv9b+a9qcEG
5nUfDbI7GVWS4VqTSBbzUA==
`protect END_PROTECTED
