`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+v7OI/W1uUV7j0MYWHJjkOrltg8JQcldBdtcZ7hTtFWyYLOSNzG8snsflH5cVTDG
4DG9mQJuS6Y2reBiuApYBfgPZW39k9u6PK03HAVU3Djdi9t1Rn5As/+MJcHJN0z6
649arrXKvCYq3gZ7nKfP4k26zi+ZSMfwgOAd4JdUcYNIwQsqaQ7TFrDvAfZyQz6q
nsA18s9ScltEakmJUvuSPAPRRfgtBjB4vezks8XF7das2v5r5onJwmfRaScIw4bg
/jEoudh+mUmtur3RNR34ZSSxNIOJTytYemluIevgVohF97yMPT3RWZlMvRMw4Cwb
tCUGeIWq95ybCINfEGb0yA==
`protect END_PROTECTED
