`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ma3c+Pag62txQTRInGGmzZjh8w9BuP457YMORKUIKMKYMC6iwrK/pxTXwq8vmwnU
tbIgINGC2486lgz6CXjPezUJ0kXL/VlzYZZnspyHudy6hFAO2foCE4fEs/keGOop
ZvuwC3hiTo5NDmo9arWwvY002fa08lVGnqCcZAUeVX/hsnZIKZcZpqbhhphN+L/U
ABzOt0iKW4u2hXwLDdM8h/2lC/X0EcSl8hV9B9DIM/Ix+pdj3jVksR/1hBC97Ajt
64hPjRXsr7tyMAtfYRL35kFWecmJuz7h9+7cVZzV3S933SJ6sshfcVGnEQ76L+MB
tA7pPtcpd5eWnF8tU7Hhj29Ig4EyVJQRE+0RMh8zsBPzhPNYSleU3DyBfDA2Se50
ckRPje+PqieyUhj0+diILdO2bBB+1sCQtf0XU5XzN10=
`protect END_PROTECTED
