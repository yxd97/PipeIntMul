`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s27cx7hd1POWN2m51v5JhWmzQdqeMhs2rrxmKzABAB4kkzmNRsXuEipV2O7LpBMq
dB+3gp3pxqCh27sG4mPfDt7cHDw3n1uRHdcCrgZWx95eAZzk8H6sGL8YvRGEvJKm
0mhdlBpqSFdyJpsyHa6Rpm1mXhWYetPkuMabZZngI55G1Tnmut61ce8f7Oi9R3+E
OFrK3oITvbmgdEc5OIF3ojB9VvjVh6iGGfG09k1m444N3Xt0ZMhv5KVHlsNk8xc+
68fATWhXpMLimjDyC5XGMAWZ2kcqFX3utSg+Z67WgmyDWw7LrmwXaqzn5qTjSM4r
Sfi7t4Mj4TZiVGKN/97i7zzhqQ/+57lgK2oY7n+RCRLaJe9IKI2DfB+n6lOvIQPu
`protect END_PROTECTED
