`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EdDHPiaswcx370Vv9I86ezqNRFO32tqqytWQ/G19kDDasUenwPdjL1yDbBTrLD0T
b+OHETk8pOgpTJWIruZi75H7vnA2sCSOKjWjLbuSa4v+si4dKtc+8sPZyWFrt86V
KscovW5fJS9B5ayk1do4jx7j867kLZlZTs0RlyLTFcIQl6uJ6LAHH8Iq0SyOOvhn
eHxBTHw0/mEJDWLq9lJLzIuk838Del0bm5qHynikPK1QG7vLdzNAX8ppq2zwcK0e
IF2PoxhHQ4H119Cqvbl47lXkhDeTQmvXASMTkfD4UTG8KDy5imsCKabLt5VhDFOz
k5C8HXFx/aWHDgpZFBqyONGwfUNh5MMRE3LV2jhxAk0E7jV0l9GJAAUZe3m3hm6o
/W3wWhE91AHYkwuT5zvitM5T+XO8+4XLZSkI2TJQI4EZskQWH1SwkSTBZv8Y9kbR
`protect END_PROTECTED
