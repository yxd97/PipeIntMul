`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkhzjB10chWVAVhn+OMB8AtgSxay4HR0cH66DG9+P3oxys32/ksTY76gGezGsHbZ
w1OTHH7DMDvJV6HYKFQzQsEwn5WhJEsLsT/BvjHZVpTNh10kN19CSDv+sCQsQ/g5
9QYgqSxwsrHzAk0yUzEBeE7a65NOpVigzj0dTlTldhUbFu5jMk1cR5dTiAOlR1U+
M9iigSZOiYDniDccKUXrWv4YP1o9FNnH0/MZd8PHW54bDqFmzNlSd9KLlc8OEwuY
wbG+OJ+BFKhrjA2MkP+hd+T9/SWeFILwOvIBP0lfMhgfWBwEb7czRcnZBFRubpYr
BuMFlu0Ft1eDIavx3KbcI3LVntcBgMUGu7LNW6VBZqGN2qopL000622u6+la6wpW
X68FoFH3E6w+jm+K2VPFoLNXf2TXdNzjZQFTeer9fBb7tranvZU9Ga26xbX7GErQ
/ACorDKwK/+3MpNzWd7UieYrznMK1I65IDVRgYsCM12IgRgDDJ+8YPv6IGFZtE//
pIXCZrGaCX2+WJRK4ZUScyy1GGgOEpfiBdflP66ugd0jHqHvYy1SJud+WV/gnSMn
Pb2iXuhKLWQPuOFHMi9rgtMZNFO+hz6jHXOS2Cpeya+5TJjAnDXVJf4kyWLw7kFu
2SfRvOTxcuHEjoZDsE2XORGFxe7GOj5bOeOfkZiuJIdzXdjM+gqz69KHildLBUOy
Le71rVFDfxGW6sRmCDdKoJcAB6byThANCxtwt8cjPU87uudcmt9RCmfLqdFBzMPD
VPxksMGV5v2rjYnSyCJNgNgvte7lkk8uWM/nX6vlEmxzTq6jmbSKjIldBhSFc82a
nEXlv7ys/htJDxsJc77N/kK7fHwazq9+2Z2cGzF+e52Ilw1Y2KPoOal5KqmIGbqd
AIEg+WHglZRXudZRjkQ6aOZFPsYvnf8Hl1DxTSrpoIkvGWsozsnHHX3ZMNGZfNTK
CooPOFyh/Bd08de/MQJUJQg1x+gtTv0M2POEEI+J94NJIlS97XoQOngxQcfd/F4R
M7IF5rDtV0pwU6UYqswF6upBpubXutA/HnB4PMQ8OXJo/ppPGuOa6fAOtWjfWA3W
FQ+CvSz13zp9ZwCeomrgiJLBnjGknGnn9aLM5DsA7dpDL4dC/skU5VfBslD0hZZV
tgyGXHgNceG45rR6tDFQi5jXQkigin8OrJL/tXCmO2ZU+h3LlOWQMitiuySIgjG6
SFBo5UM1BMhKWONr6tRVy8fNW8l6AfTEeaJpT5mF6qRmQHFUS6BLbnpxancdRjKl
DlVIRwDl+haL9xR6LLw6kJ1IjzVZUmT2gyjd7r2jJMmvARfn08hmnIu3pU1iDxle
Ptwjb/P3pysF8Jzw6ObVRnYqOz/Mi4Hpv0eia6s6D4xkUroTVO5c2vZ0Cp52x8uw
qJoeZSCqpDf/ScPIvtx5aQ==
`protect END_PROTECTED
