`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ExnhJ0NsGHvU9rApNlqUs4QgZbblxsPagcFjBUbrLvpmeivhwNlhxGBmBLGBbvdO
dfwnh3PPZghp405tSEFo8Y7eZtmfqvv7uiuolcQFH2w9ZUdHdM0IX9oqszzO3iFQ
AVesMVVAqNOsRad4oPftybF3quxJrrAuxD6EGadjD+T5YXUHbQK2+iBQ0weuyOCf
isj5cKIWmOCx1DxjReqoxKWwZ1541KMiRKrgJ5Td62G8PhfJPPchiYTeZqRxLmd1
qnpWo5XYDYxM4Lm+Bmmt1IRNA9KOMdAxnqfRlh9wPnvJleoFpehza75IWkK6SudT
a5nTgVpQ3qjcbojdavqptuZ6R7gr+wNCY1/vLCbksCMeZRv3+fsmvUd/fWAQQnhv
OYmnbDtDSRPeKvngLVYKwFh5VVUEdcFmPrG6Km6Rn/CII1uvM2bPF5LPbwPxax56
u5Ti3NEGWkpMKqf2MORGE52HaMkShh3KyuRxwail5pIfDDk+ynM7zBBe/6SDLyVd
f89D+9M9JY2BBXNJlxtXWPAH/AO6IxKinHYtJ4crt/xTIQTB8Q7yFRNny+r4NB5R
yPtL4MMdayNezIb9kCWvCMUza4agJJdKy1TAxbyvb4LdRy5Nbv0oKVxCutlxkmTL
WDMy8auUNEeWOAtuIahLXl/kRcanvjuLNyAZozl/bPi2ZlTuqGSEcleZu4yTyuZD
61DqvfenhjK9uzGLqOv2q3yV7KFqkHSaEfex4f/QZFWw4xIBvscAOD8dkeYI8adv
eEP/bVjqT/nYQ+sVNjN5K+xYJa0RiISp8TE9l6g0bcvkicBRXRwGJEefNYMRFSyS
AvhKZNfvuFOEjiucUl2dDx3eGZtkXlvthMImiCCsx3ZI/ZwIDzpZMwQtAPkCWJ9+
9EOUFFEP51GW+L6uCH/DIEoZiPZUCAqE9BS2A74SwFU+VvwZBYRciVL16n3aPIeg
BROS5WbjpZzD3ilvWNFbY+LLKqKwpo1WaISvdyE3XLR/ExATxYmvxuHyLhmnXJUb
4HVIpKpB3Dm9arB26ex517/6bGKQjg2cAe1atD1afXiU5qTEHurGCCfJ0VOMJfIj
2bGP+9sjzKEpvzR2OaZHv8Li3nFeft7m8YzV2ex/10dfqk9rZv4RwfJGI1wqNbFZ
WPwsLIaLAVDMf21S4B5EUqg2TL86Woy8fxQR4vqj5yTAnbGjrqyHhpK+m4BO/8GW
NN6ycLrLllE4++bUfgxFYtZZHmZBZcCCNaIqMXNWdU4fTRMeqZ6LRCtSkKNSmKb5
tCbO45gT+8RkSHjfxfRmE4oKrwCRevJOvEaY7TGd6VD+sxa3crsqvri2TUI2ec8A
50rNKD2xW1AjyhOg4YjMG62O7GtER7bnBHqvWI8a0KPSO5QsBFshxtObxCrb3ITk
o/rtavEgXUNFODalZTy+IMHH3r+oR8hARM0ATmoKh3xWPYgmpWGUPPbwIh2NrMUV
qddUb+1ub05Uqb9Bu0aMyZnl32+m20kS/FCmdUIa24Ta0JAUzBAJvPr9ICCr2Fkb
kfyzF8waaElW1fvohMm3SqSq5BRzmL4eWRK0oZLIqDTD6Fh8x298IZyKm8CuXIMG
ylgQbuuQMWoVcTaTFhrSwuWc9nnYpX1rveE8K+u3GINsMikMS96kCvggaTPB3g1n
ILkvjaoBEvQXeaXJjsZ4WqXx4WqbXhlf/PGS0CEgluEJXICvn4+eCInukzv7YtwW
8+0+ph3v17cUjqWSCm8p0SEz4AGY4czjUAKdzZrlcO+12bDadVQPO/Qodz2wd9jN
4cervW+2tFGrLB/T5xl1xUglBIuY0fI31tnZeEA/8x3kyPPL91hGj1H+yspT79pZ
H2B0V9NRYVaPknz4utBrUVOOwYr/ApAKANYtN8cvW1M5IFfa6D5mXQZaLggfjjAs
GIReAvVPUbUa7Onch1GSfcKy+hIdmqD4jQCpNIf3TQk1ssd5ja6od+0k5vcI/fqm
xrTvTfT+KrBqW07T+8t1fjC94Ol8p7DLXIv+omcvqPAloUJj0lZYg6lqxq6klu5G
szWmreuvI/ReF/JLrVBAhVNCDoC0+aHH8URr8wGHY9cgJgr7/jairM+OuJ9kvIrf
C916iKKmWXBO8xYRNOC/tyroyQRKV9LaDNmO5fqS57sTbmLiJv1Tb/qMYMIegAt8
NAI3t24uxx98PlwCL4wTahIEzLaqqTrDCdWrv4iRUJ+wDpQqOcn3e05t6ZUZuujF
aL9VduMmQG5YodnIOnkpZvjRFTrIaUJVU0UgB3JFY7/+V4by2mx7yEdBaeflcGnj
3OYfwnH/qC/HTMF6UyIE2GP02eEi6UAr5rNZGQG8oq6ndcZfC9+I+2Yjh6uhRLo4
Kv6B/YOlLesCvv3Bk4XjIqt08lDa5pgcnGkBx3q8RZZnkQ6PcHJBezGmI/KqjuL8
goIoBtgpyRctWAGBrmALVF0BALKwIGQlKF20rBhXTw0pvdbr1ubVvWeA2YjNapKg
6kzm6yRX9XUyySb69dKXr96BaHAFyXxz54fY5875C8BgH2vOxZx82e6DETeY/eHd
n5OKIPWuIxdo6lkNoLhItcvs/o/WL2f9Qb0KVIcrMuW81ucrpEOSPzd2WbJ0AdLb
6pDxL5lb3XvTcOcwxLGFHVUuITqjKyaiOPsTFw82IMmMAv2lVZimVrpX9kr9W/yE
trgUe4II5HKdBggDKhxQV5HnH/yuqFrTbPeFufAyRNQAHjWCTxHCg2xJNz7Ga2Lx
k6c7V/7Qa9Pn5PGdIrrmTZ56qJoc9EiGEspPRzok09OQxe9HLmQ+nnDxxpNOYO+d
4OSx+Ga2n8IwK6DaicT4BnYH7ribhDsTHArI8sJp8V1YdG09cYqz2RjE4PgYR9WF
G6cmhlVHK3N+SoFBlc/u0taOem22fkaueeIo4ZLN+GJNOhRUc4sw0D+V8Xwg594a
HQfLBkqipbdwN0ZEttDf/8tISRyKShE59eF2CSK/9NtVDJhP9YZRCwQ1hxc+aKVE
BCs8Tu8IUNmB+dqqkBJ6CmjDZrLSFjjOF4oPBVWhlfjhmB86i5+DDUmYE3G1b0Mi
U85SVSVe6aQJeQo5A0DKQuIndH2LuAlcRCLeSC7bZh9DSoTRR1N+RyXDvtxoRJad
ewUMNPCAuJkQuQp1m9m/2RLscQSjKw7z3LK/vCxqU5LbFf2bbLB+Qy6xbipu5oNQ
MBff6jw+Ijvyg6F50vvEiE4rs1zaxnXGMdn+6WqDM9XuYbVH7zSFVClvGiHoacip
/bAO/4j9D3DXhZr/OsyFrpYeiV01+9bmqlSDvcaJInLrB+tTMBVpoTT4C6pvwMte
NWj3q89TxbcZF64UXr+ILCkfxbWW08poJ6aqo5ohAHDowM7uYx0dprB4QPI/uK7I
+y79NP5+V1un/7nmdPhG8X71jk7dutRfWwKPy00J8EKlucSQ7YEOQ8lGRFLPZoI+
TVYqHpW1BlPV2Sh0gPmbPyWBSMNwFb8G4JqsRIgSyX72sRS6UXz+861/A9z9LmxL
6uVk7I7nK5E2QwQ/soDlVAwmAKpMOGn2/VMP3Gogm0JzCdWJ2kioIQg5pTBvmPUJ
iAvu8bGoXOlVtLznTwN6IRABKtv9KrF9c+LeS5Gj/fRjypoT3yVxWKKn4+YAUy/z
j1wSzxHnMmMjQAM+5Ysqoxxnk+kUliw3Fe2Q2wXTeLb+wYMKfQbkW0vpZbsF1zcs
0pRDs8h/H+Aghbsg8yQ68AVZe2CVS6S/suKKG1aexvHxBJrLu9EYV4sbcV8AYi5D
PmmWLvVwv2v4UTnFotaqf4EPKrPlDsLl3ws22Cnm5V/yG3giUrimy+Zd4Ptmhla/
ur9Ryruxune5zC2LuA4svooTeoBW3uE/fxn/uTfOpaEJt77SksI1COSzWFAALmez
cdo9XUjPMjOcZ44fDzcv+ZzwMi72nj5Z4RfeNkqF8DGaxhaYyVNwlO6fRi62iVOX
uhD361tPW2rIrhdeFsYR+MjqB1ymCdIk1ofnBrc4rdMVH9IVfgkkZNO8wYvCblkd
+Fkprc78P4UPGlXTE/C539IWO6alFg3Yc1WodP3GSCqXQsJo1jM6BQUySwn8rcpy
iJPAQ1z9LL0NhlLDGaObzRoHhIPYMxPLJSWHFCztFtzk7hXzJghLk1VWiLnvJwTy
FBuajtG5qFFRn+SpQYFQZ7OwIRbmxYOT1mz+K00woLGpNolCRKF7bN/qdcwWoOfU
PAeBs47sx1KDVCL6q4g7Cy1trkbQq1XnVlOuaWB/bp2mFtBnXTmi6HlscI8z4PRa
/Bh9UZ2GzXZwJObi7ZA9tjuAJotE9hC2QBMyetcmGpirjFvpWa/hpkY1wzNmQYRe
AEo9RQmRIndtTI5HcOmodYugLbwIci7eWb0jH2y1QrDxQv9pWmWJqQBmNqMWe9li
mD61JuNmm4Q3czOuiWQz1q7ZWxkJBG1oVfBQ5Aw2E7yXDzjI/qkgU1u1b6B07RlC
1OIESpoNr+dMGuTNEMjc5fnS/2cUewlDMDvjHTPkmsmUbIEYtvYb07AnR3xDAEtI
DXDBTNBagqpzQ21uFPdAe2oiaIw0PAOuwxNBvfRhn94FwHnsNEcSSr0wQ4Q/EM7t
KKTXrc0sVWzz9M2di5rP5gGrCo3nH8a+5Zj8vFWyvMd+t+Ck+VOtXAY+eUpOXHU1
Fnk2MLXdGJGRNjoV/COf3ht5B+KGx+330H8nRWcQg7OjxGdk2UYQSab5HhW96h8A
d6BcCH+0swyGPDmSbOD7bLTt6BwWDmMPGSXFIgZS+fwceVX9q+Pp8v0+Tf9uh3Rz
NzhaaNCGV4sr8nVc0vbhlsBdRD1gTS5tpwZq1q9cqilWsRhC3a9mlzNYyG73x7Hg
glhY36iyLTOX7zE78SI6HtypCMYiqLy9hovZp+OYg0mUKerKnSZEFp8iHnWbEvX+
GtPpyvk8xKa3XiGfQ8B6cYueGGyuDfku4MF+QflLvjToo+dEMoC8TaffMJ+qyRXU
nyTWyVzpkVm23USf81f7iUyZv1gErR0ErsHvjICg3l/YVE1adb5c3yFcLHuKsHhM
vl+3/4QssvFf3T7KPuhwpB2SwjvGe5IuCu07ZqYbLaxEXmjr+f8JATG847eE4Mxc
D8a52ZvYL5l5lkmF9wF8p5w9TBduXjpDJ6sZZC9cgg57Uae3pLu7El0XFwNCqOCc
p16Y+30xoNDFJvNeto54TIzC9jXZiowhCM/GnBd+9cjv+AQKNNbDtyJ6pbqVtAz/
TTCXLgsDMkmsHE9B7s8OS32Dg/XxNgkn8PlfGNtcWROmPuzwi71rC4ggMG/Oxqzx
MMX3MxPhdfYx3uRFmrByjGY7airhcOlZBVn1yG7uIAAlYHu/SF/2g775FhXKUJnC
/K34RqoEx8va/k/6HgpI25lTOptAZa6nnaVpD6yCcbnn1Ye/P6f2qL2nrELD4RvW
R436TDVi/lyNIIHC8+B3pHpzOmdhe+7wCqdzgScWPPZ+zROLiyPHsRPm8R36ANfD
U4Fdhp0WO2CCXqx5O8e6UuXim0o7D52vz7s9BFYWWE/4jnTCLbtiMUVOgI7VaVSr
g4nsvPpknjIXlNG0Y7+8bDACxPGFZHG98b3XTdI3uE8+en164VupW3rIZ5Wlviwr
kKupe32L/emg186IF30ZvX8MYmUX0Syh3S0gdU83bVE+9y5IsP/XxJBe7LdLJ0bs
9ZJ6GytXf2v56Hm0JcZqesdTBnUkPbXls6Ln8fW1ZB0OBMETGr6DrwNs5lcKo/RQ
j8BqGqWVDxRpYfzh8eWRu54ROmvkGDfpdwOYTOUwOAHWcgAr6Zklt/QmOz0vSU6M
r8TeG2xefXZ4a9rrIu4T85pPswwEPbOI/0jEkS92LDsTZPk9ouZkTHxp14kMMxfZ
lJ8qQC0r+VwFZF9aY0ONnNSuTz6kjKZeS1seKSMGc94KRR1PcGcvH2rvPOtCp3MX
F0F6FNK3sdUsY6HzwATaXgGASGjUB3DKrIqfAm6OxsA0vvaLMb6A42mXDErM+Ilq
RXmXHrAK08mjB5TcCRXL4AvuKtC+fx/CEHPExN3totgucFPqy6929G2mDVf0w3Cd
SQdJGxsfO9yFS+tThxja5hEABcZO96tmsg/wTRlzy0+xVpqIWcC9uYMlacQfguw0
rLrdyRDhhI2S1ShVSi0qp9ttxfxP3staZfUNymifWopdq64lRrIc5DEKN7809RTF
zEZCyiNfCqop2DSHNuWdytM6J8PICXT/KRADfxALTy4VUzh1o3l5LAXvQH3ZT9Oq
kafiuBZE6HjiTO4hqe/q9eHzebovZPtDNtQWxqjg8Apo8jazil8ap7wRWMNKwkGj
73jjVz9lqwM8TIz2uQ52BPLy0jvmpOQHd89auQKmdf9Q65RJJGOrF+3Gc/aJ2MAd
YOb5mh47nXVjpM0UOnn+Pn04H2TypSkfm1Uz4xGZ0/qvk/UekUJui4aIkZafcJbc
1+jg3n7QBdP2XpvT1pljfQQ3mE+PJFNNkLfzqvwWvKOky6jR7DK+dLQgZgHtaVj1
I4J84LQoI4601/huETvBF+n9cZS3RpBUcKgf4A63s5iSBpw/Gamoz6q7cmIc+NkX
DjFMmKsimUm/ui+C2bUCyUa6cpKy+aUvZ42nsCgkUge6G0fYl3u4kPc9RCfdbK6X
uus51jJeZLk/j+RYeyXhh4mAUbqvJDxVcRkQ5fnW3WVCjX5sjm3FQ0oSE4Aw4Hgu
bEabdV9KKXPF0HvYNqHGjp+i/9lOjq9RvKatdKgNud9CMNdJo6cflqAPtX1PoWBi
fG2x+QDa5GMdVZ/+38NKhKZnCheeYn+fA4Hhb+Ik2ijHdAFOSvwEKxfwlIirXh/S
Vzmp+EL7v+YdUWxL34nsi/A4SXCy2/3rvEIZyeaVece/buLXz7Fw1ou8Wy91jB6m
GbAOs6ivWvxkF7IVgaEtQUXU3ucoUtcFpG6eL2xGS25jdI3zvYMpRa0r9HIZISsd
AcoQC7SbJN+n65dr6YS1+AzE/W2NbdxzM/ucBoGxAkV96s4FmxwQKIjEMYIx10Fl
gLd/0/eyfWpEGj+G4gNZKFdOQBplLuRDIPZsOxYm/jZ5SS79iW+BNyHlKegNNH6z
XhFUY3aUxEvFTRBMFEgLHw3b+S4igyR72FAPM92lHMqc1TVrevFLHyHIBl94KTva
efZwST5zLFsxZOLnfW44+8nhiQ/zh30CBPex4c41JCPldF96yQN4MkcUsiUGqgwo
124MArIn6mwbzl/dhoIYdqEdSAps0+2Y/tT1BIXmyRXvVpSma6opXCVcuuHdt9nc
XovWJzHKiZHdyV01cQlyjU407JIcnqHPgd1kB212dtiKKrAZEYfqglSX/g+T4PyF
1Me9rJlZ8ZD1fu9IDapmYPCRD/POvTL5ft4oxe1iSblhqpikKTIQVPFfOEip1Y7r
oR8aA5poUXXQQc2E/7864uNqckqUDjhj6wui5wWopsej4MlYIW1DXOskaypj+22c
rI+Y37+PDRHk/o6c5Yi4Ze8EJ5IcHIsSk4GOqKXwUSjr21yEOzC4+8iWnat0DwD0
rGpB3kYLzjPLidEAwufsQMv6P/e762IJF3y2Qz/h6Y+Jh5RexTyFojJB1Zp/4nAf
HMnR3n7yaYFvHtihO/y3Yo3q9ocvvAu6vIRMi/jOhsv11JOpHpOnARaoL0CccLl6
RH6MsqrfVe6mlKF6Uk2HrQpf6/pG4/Xfc9P+rcpbi05+J4e+NhupCW66+sST06KO
Mgj4YAAcPtir5cxOfpjxXcQTiYdX/vc8PRa7eMAKzN6dv03g7dQo3/VsxcD+UZ7g
owXmmPl9SNTeNUusNZiXk+0f+FZCCbV13J/zCPpDrbwt57B8m1c6ybh4Lpi3eGuQ
mzQFQJ7wLPWs1EfoYPC2VxDIDcUerlbQV0jZK2m8prWjtRemd6Pzux72Fc+mvjEk
HWMti82fQ6IqUETU6AketDgX95tmbVMjT0b026V6q7yd9T6vqbQPbmOQm0tDrasB
hBdAzbRI74jR3TUzRH9j64+HBdwDElnaXQxg2eUNfYnqfkSxvx1lbSFDoYaame+7
1uPtUVvnWtw9JIWDsFPkIyJFhL8cKnf5iPr/xDm9jAhuEvMtiW3O9fLh9Xd2LdFn
rtOCNc97wM/yxZd8acw5oeMpEX24bccS9D61QVla1BSjMiRtIowOwk3WQKpBV9wq
8Mkr4FcS79zjc0w1H4jKyU4IuRjppgIAhK1a4IduqIZrh6uITv1wPqNFOXUWevey
1O62u84H3kiI5NYmfZCkIrUJmcVKlw1WpoRcO5s2RK38UuRPJVqp/G+8jYksXFj1
+YWtTJeykQH50WPCVtDOCvYyTtNJPUekaJVbF+YJSVBKCfJOI9K56SIFuWFYHFhr
WoRF3LDYB9P60SRgLOuyWuCKYd7ylsZ+JFji5WfyiiCkrnt1KwpF5t+y0sa5MIsE
t7ofgHP9mwhurxOw7bcCic1gLLFpi4Ok65XCu9mYnEdbct4GSNei6V9OpeBApxVP
5TCwIixvs+Ri1dKrBBZIgBtkgpdz976BIBh/W29exLjYjfIFVJL4gDGZJf1VA/6k
WYV6/DyQNmPrNFWHhV69EKZ2DqUeJPR8PFCuS4YJG5qNGEu8dWdLjw73XlZJ8WyY
SRsvvOS3UkV03F4ABxszCTYnaEa5V1YrgtCyttaK7BHDGL8mEHF2yun5fRZRWip1
1H8PVCb+wXm1OBhzEPRJ1czKC+lnhQrjJ5Z+JM+ay8h8ExCS13pl2fRnH07/kgB2
Rs5PK2i/KtZ/VILe3kLbdeWbpZVPgoYJSMVvT6svG3POX6pmeYNq16bE6/9i32kC
hDAQnBI+TfJ5r0/MQLQSCal0YJ8zoFo2sRxus7LfzEdAox0UgXvJoVDCPBQyPcmU
zaIe4597OrbXaCg1y2Ioy4ZCxkv26G+7JQhQikPyIOw55aFDbWIYBV30zSshy/VK
DXJHirt9otljnimVQVKhfy6NCgIu0mJL/jatsFcaMKp5/2eBjmgoe/y6Tv4LMFrQ
6sOUzxUzjO5YLU465KggtlT1eKu7p0aeIgBu/uabQ2P2VHzF5WvfNWDr419eq0WY
Zaqf6ce/bFxVnRfsJYJ7du2a2P31+gr3xem3gvpYd8+VzAbVKu1gRdWkbzsSK9+Z
IhgI71wVyjMf66fKcP7UOgEl88e9pz3PfWH+V7FBeF6Ea8BSo1SeS2NzFiU6IRWD
5Xs8ftpzYK26rStg/qjQBPb0tdBFHETqk7IWieNVIHrc6aDeuvSBCuNvkCG6fPsX
OOGY2T0G//X4wHZG57Cu4En2InoqfpbxsIZPsIgTkeRsvzbgFIlwmqzdECTVGKq0
MNagdDnDBvlZ6ck+uH6CKZKYNjpT07oNs6+FxQqyh3lQe456odm20FgfH66HLEl2
9gSSozRB02gz8nTpjS0QZMNwql7qyFCj0P3fnIEQo5ZKp4anjJ4tsa8h+CELkZqy
S6IQ+JapMFP4+VfPhihhgDipxHQe6T4fkJnqbDXUc/KBVSgwPwzJyglNTN1l/RUL
UPNKXyFbVchdlHI4HKVWb24DOavMniyXa2sYQiRssM6W1hG6kAeamO4X+eeiQurd
vtdOwoPiAhOrj84MbohacL8zUqhfR7COh+/ztAcXXXKDG28XyL/Qpxan5rqwU6pZ
Eis7CZL+DCUg7nRgCSvNY3X52WEuZfhaIBT+NhG/z9sZTpE1wQdcrZ4pJX1WPF6A
m7BYfml6PkHSWvfLstrt536frA5fRpd1W1366cjdEAL6ljwa6YbDkFEM6ajzXvXi
XSNEqgofjzfsh7SfRgIhxasr/XzpxgEkcSy8GEdjSbZb3FzFx/E4l44jOnB1vLmS
kwm1N3u1MyeaK7mDD0iL6TJtC+dZLyvthe5aN9P20EmQN5lHjSao4VjZplsxeQzL
hfPjm/GRHvGFeuWROoqCKKb47eAR9J/YEEjkF+jO7VBO9jLmljhfJQY3xA5Vv5QK
eFB6hg5cxyYSjocASQ7DcX+EWo6TMoZIp5CihxL/wsORrC8etMcyUlew7DKua1iH
VOUmgP/3ISw4eHpwk5DWvzEYWzb713r4Ho4HASozAFdiDzb8nVzyHi9hQIXDeZYf
GgDheCAjw1Y6BFICAuPU2w==
`protect END_PROTECTED
