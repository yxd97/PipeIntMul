`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCZfAudsPM22tIU/OPoGFL/kwWbH5/RALe0pP5Px1+3GTuiVeZeJNClt829qiv3J
ByiwND0w5YPpzXgjreX/hSIohHJnZ818COE+5VQUaMOrwDVCPw4G8EKVotOaKev8
SlM5h+O4H0nWM7JnXSSfVAsiUpuxZgFF7e6T6yhSGstLBAeuwOqcNTIGiZLOw4SQ
RTCucH3WqSoOPPQNcupuW8uLfg+CpIuqPmI9b7up2ymbPBuM6KkDei+bABsR6GTj
+8JH3PKKp+C/2rOehQ+xbDkVS50alCNJ7Gp+NZuihiWLGFCCwgdwajI3vESACGTN
yI0zDLIUSuyQ12eNr7+vUH5fItsTTsldIjLoV8STYuYBdhdTecKWrkoKrWZMvX1i
MMytb17D5tOSFqVyOxsUKkq+8OM++oLtgxpXR2PpTOew0KehdqKvVq69woVBN1di
kwTxnNgy68FdVrVZNbYI50rAuohh/X5xLQQF4WE/kgCqxjbu0+Fe8bRJSBIHKLBE
huOOX8m5udUlyZsxIWrXBo1FpCbLcRKcp4J1+Qi1NLPSFBJZ+8UBiUZpbquUnXyJ
AYcIVccGvNpB4fQ3p9mSEPbQP2S7VSWKXxra1U0I8253QmMiFTvL+2iMEmFt+fuT
aW9hq5q4JRxT78tJwkWIuh0XjwiSkfjKtZAng+JlkTAnvpsIb5okhnDzdmq38fjs
LfTRUBGMLw7x7cItijZ1evgy6n3GaG3IZ30kvgBa7i8gCnvcmKS5XlBDR5OTVvac
RLswppYAs923fA7yaJtxeCz98acqAD9yT6lXFgOMrjQ+Slm/GrcaTYyfiVisu1hG
oo3GCgcFKstyTXObt+jvLD63T6c1mAHOFVLjKukFNA8d76g8pDaiGpUhhNy42Ht/
JoKCGNqLzOvUiLBFu3ksShqBRxEyNz80APbZ0MXVQA3w3Y3VAywGYeg9eM+f9yb2
LKztl1UUEVYiJlcC1+kT9qqxOiJAUYiLdnrabwciUUqcTH6t5mqldZYGy+49tRul
WR2kjY0Kk2JljGvD/3V9awFLjneWU5Jbh8Dq9XSViVcBM21Y4soL8F/CrIxHTrUU
L6qFDZRiI7e4tOh9UqwNTntIhNv0pMV+rS/3f+ANXLqopmb6402zQMjkzg+R7dpc
B8BkRAo1tJlQry2x8vUFsfs/ZcdWpevefDfbKYFqW91JUYI0xe0AmEM3zeuNSTqM
rb3/Rn4TZoNxj2xmiseu/w==
`protect END_PROTECTED
