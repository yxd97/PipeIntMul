`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nu6G/JO94/IFwjW9pE1vNI6S7PbYBg+OOamISf6GKHYwkonTa4oMcHWxNkt5H7E8
S0GL7lyqDdpRS7cHIwUru3mmkPsyvAglIW7fgf+LSlAs2GqRBq5fpM4J4hfnaUCb
pY0HpL4cfShvY0xExdifPcrcctmnAraG3i3MmtmULod5Mftw95ePpjrOLnJA2uxq
RbefFXb2RL+M0IZNsQlKWacTTt10Mkea4l7FtBHa3Zqof/25zMKpx6Cr8iHJmeo0
QcbROVtBF7omx+SLunAflQmE+uw4DVTTU9ZOn6AmEyLur4udjnvsDFw5S7qCiz7F
pg1SM443HRl57QYbZFK9Ocl8i+N0FUiHRyZZ95285tlSrkH0cdQHW/u+ZoGL8mkq
6g/hr1JNwFfM89U3XUaNx2aq+IKIdCr1x92mDaDd+DotMMFTucvR3/nKcw0DGf6j
tClubYRcvgLY00KFbxD9Zzzx//Qc99FccxGc8pIxcUZFzsUiy9W7/R/OmJbFyhyY
fcmykcmqZcIWmWoqvj4F5uJMaLEXMgqH8SZB8oflQdbY6tqcKuV29c0pv95t+XkX
6Qx3BpILTMOLn/k7OrgjBMXAOZC5Pdg0s1kUVidp76RH50pr4BwgiMNPzZMLCk3U
hLLkpA1DO7+M3Fzi+7+1FmczzxistFQe0wbvH72ZJVVUxj07UuWOvBzSsefSFAqi
G/Ay0f3zNhyEmReaKJD3tUT9nDZemHj2hsZTmvtOOi9wEtOv+DnS9OHaxriEnmnt
q8w0FGHatNzt7Y1qaRbvuP41iPB5pjQ4pweJasoTxy6aHdtyqkfi8ztuJSELVQcy
HmsECsOHS5KrBrXOHRJ+8r6Q5Xx+7gjvoXH36JGBBqo1o7b1B1KovBaCZInP2yET
LZaHd5/jzOvzS4dQ+1PdsXRpZ9gOYFeF1GIJntPT4HdiSWNIN+veC81Wlv12lcI+
tJomNhk4E9njPNtR7OeQy/zleXAr5s4IE48BOEqPpKjBi/8ahP0V88P1xlctvlCQ
ZWgA0K5gGCxlGVJPpJ3u5QSevjdLn7lr3nbcd3iYCYMg/+e+o51YCHr72zvOPuU+
eclX/olu8YAX1mX8OrG/n9qM4/PBhhrXL/nRLxhUCX5wxtspilvEowzlRy7Vp6bf
rj6zS2y6wGSz2JAXW3QSCNFECGY7uo4Ag9ejUuaBTEXC2m8esSXvpFvikc7D4+oC
uOThsZzvkMZ3GGxxPF/fPHG7Ohzd6h9Epz/fIMS2POFKIz5um7aXBmcrHssQ5FWg
6lMl54rwS7hiffdmRRTOqpODsSbX2sRs9hOUP76H+Pnk5bstbAd7ky8DOOPxDuzZ
RrDNout1P3x1NLluvl9ShVV3XYHBeHnzW2idqmjRBVkvll3bLWn87GyVm0ZRX/IO
SssXVnF3pRD2Gyt+2veNfSk5OEWLdwYIFrzBiwKWedfz9/7nYBCiyf+LnxBsEWVq
pDHOQAYrI7y/r7buWlIHPApod5ncaJWZCnQgTk/CCsebLsybW/OV0uWnXwiU5yQC
n2+5xGssgPySTAn14ad9/8Dnwgi396k1yrCOaoVgMUKWjXoovZ5QFnQ6dNqxn7GK
EzE6UDMD2G68pBXvgLgScd8a61ktvBLV7L2NxdDqU2AvXktewvPc/v9tyR1aKOWo
vUxT66NCvzRsdUWdh2OaA0BeKV80cuNH25WsPhbcgUKz+ncRcKZJmBWd+/XebeeP
QSpslWDLzB5NTCwexKJbjTGyk6aX+B/5PKC285mNpwErRRf2UKRJVUoASPR/VNjB
0w/ViCGMaO4Y+81dViZprOJsz/6cyz6+hgqIAhtQml1YXeMHVa/FEoabUyQVMKns
I4Ut/GghcqL/3wCb1D1immv2DUzF0UbUTI4IRLLorn4H5z8Ux+2zI+z7HYG+CRod
RvXcySjd0OVPABE6XauoIVmYUCNj3kFudwEoikz+5tujAhD4ZSg46hcWJQmTu6Ef
ZjjCk/BTblh5EG+vC8hiWylmJIYEqF5ymM0vxh+eBBqUnXOy8v9sPCUOxfht16UV
nHUCIfy/Ua3De2b2i5hLG7OyJBSiHEiqlY8M5UaAF2nhdKAK9/wNcIrXfTvjEqn5
IwLfw/NC9fLw788KW+ZyUqaVnQXjmiTLk5NaYn0HLBGu6Z9SzOuIR9IdV5foIu+i
LX6ZNorrQbKGe3zrQshMywXI8puwzd39k6hfgcWhTq7eHoVKvMsyq0mHmMaEAijW
U3zFzeMDWEUmXnwePCCXDIE4rbCTAxzQbY93na64Y9FpnXH8mUp/1f4NwHS2LXZS
m98tJtf2hOl2T+BTK2cQEtGA2YCPCpqmjeznf19FYMOp447/hVV4udt2VgXGkGI/
T+ByncBKa2go6OfCmmO0b2GfTCjjhP37VvCwXG7SddcfBTn0Rb7nZizzstBs/0Gc
fPwt/aJxGjMgmTlTGNzFqZp1TdBsFcxw9ULulqufZq6ZDpUasWGnRMrL4GG9NMUI
lxpSe2jvNnoi4CZwpj3JPV4dquOw2slMIdSaZ+US/Q+6Daa7SjFIekWXJxQ8dhel
ilVUqVHYlvqvKG5XtMTyywN6Ah8U66sDX+TNojaldr7sqPXKjB2z2fR4LSLetUrx
ae0Ug36avXRHqZvFx7ajPEP6xHA5slSq19hCPmUP3WxxiP0hxgLKErh4deyJcCoc
VlB/cfhL8THoKhBJhMzxuIeISwyJaIrr+AevbtbcR9t/fWfYVOwTQchAMKiYDbq2
NwLqnv2aX017unwJAio3kqpD2ptLgM2yDxFhIgULAlNhuKe7rz/oewJPw2zE422V
92LJRO9PyMU+7i8E9nwGE3b7OitH0hxnv20AJ71Uw7XulXTF1dAOiTbI2F7jmSne
JYtT/OP325+l95Yy2gyJH11ydtrkUH81I5/CUH+jVEtkVsmRNfaM+LIuxmRyn5LJ
+2Q3UcNUsZQYDrW2EwZ+iHKWv4f4eowiFIUXCHqYwftwngqHnu9nF2BUHLUTz5d+
xvQfkw5Eg3xNH4AoGEAmIgi5f6KpOnO8zfzkO9GSKIXB0wmmsR9JwP3kagZji99k
4chezN7WfFsIvQRa0Gt1FYjzMBvxahokXGRZEs9QMiS+ZR02JMrvMEPUfEXxv4+p
DBSFzJ+RFaOptWCTuofpxI7v+l0BJzApUo8TOs6ntvdWrN5m1WeZOBzEBLThD2HO
zpSSllEEuL34M9mANQxvEOe7UQtLZE7Clclok+PqBV6IStArpP+hpqUzG8jzXcur
jZN8QJO/Wl7sMU2IEia3qFeJT4P9Op/3s54B0YPmjwGa7foVcOTRbuPIUJscXGxI
dDBzHGEZ7Brua41xu9QjVFS/BIlovwJBjU4z0FAy+A1KRep5W31L99TNyaUzyzr4
UKGco6Casj4Psws/Eg/t7NmuFBNJ/x0qjcYKibeRSGMf0bMtX3WLBvmpgbYGj6ra
h99D9qBrKPdFWyCBPF7SiN2nGHc0iavvFgG0nw6mdImOJ78QqW03lLBKNl+WhToj
199husZ3KLvBgY+2rqwHKZ8ixUL4crRySalrjTJf3nTq76K/vtGsZJR1gGnzx5EA
rdd6YfVhrbVaBlwlyUv2xm61H2m0rOs5WFF07Hb3O7iCInRewxnP/RE8aTjuFS4D
qMfxnvIz/0j/kRg1WLPCkeX1mQdjsy6ksUixc1BXVYzxEp7MTbZA5zfJt9sHsCWw
kLOiLokuyav6WDvHf0nWb6/iO5aKbgL9F6Apu8tq0tuirRS+nPmMi+eEP7CPRHis
0B35ENZUBI6Dma7xgRD9TcbGuJSxk3JB1nahk8+U8S7z6P0YIUXtZIkba16rUQQe
s/LnUdSKEqsM8CMSI3ajuNXDZvag6VvVCOzweQY3l2k3taTC4mQKZsgsY1rM5xPz
MguV9132Y2UVQLqGxIYP4FjletpwpELi1qYhE/P/PCyobVZgixMNZtwjiDvJWaWh
XWmvTtYPB78sQf6vJMiP1gH7i3C03+IQ1PO4W+HZtnf4Cbd03Ihm9ea30w+xUxYK
UxY1DZmnaExS+QxC2thtmuz7n3mUOfYMusPFw0c0YXJRKlxKeDT0JIzlaf+gtx1r
H8WM3A5+KBJMucsVlEznr3rQuRlkeO+wN+4tUxX+FMiuGeOdiMnWelJmYLU0MPWe
xPdlxFRrfTk1WtDQ9HEZEuM2YJ7Wf+8zrnab1+UrMxmvCZxz2hjgNPwAknVOXFmC
fQXALg1RtogJv4uYxB2V5DLinrfufkAICv2Nolru+uMqjq95sXDSEWQXbpLkXm4d
2ytvtOHvtqRNB51Q3xHwuDvcB7euAClbfLrPWj9+gh1QPZl2jRSyYWoVUxWmMVM2
S5iZzNFaOiJDlnCrbKgcudqKixBAtDcK7QOPKpauZjOexUbz8NWJ04i4hvfIGLsN
5PtgqidhO85/WL4fDOx+31OXlZBKozRnXo/WSkOmj5ACrFYgoBG5/osnG2OJ8WBW
kGVklQW10KSRNCKyyz8ukGdyH4If4r5IFlhuUhdQ6+s/hKABAiMaw3T+1g77PlLZ
h4AJWu8W6VoRTRtQJ8JAHZ8YjukIcSWKg4lyqr3GxEtTakf+rNre2qfDGQrHryOw
GajO+un41jxLqcw3CnOgVRg9WQ8esuz2Qa4V9w05q2iRBy0ZEBOyMGMbdUVNfrJG
IHEmOpAsjLySOcdbOSmasTObMHz88uJ2nWEhWFk9/vvDNd9qnMNsz+hspVZ8Tgkw
NWsGqnybcBALImFUUZlnwk6ZDisFLxrRdqgpQxYfX1qwW1Qx+gqr4z7muPp9zEZ+
YByAMeeotnZsRsbbw4WOlIJUsEivvTCKLBV4oyDKyNeaVBrDjI/xRhnmJD/3cxDr
pTQCuo9xp+a3VQn3p0gQ4OCHLqSw7A42YyrJE7lCjQYayE7qsX801F1y71TDOXD0
rFRc9lVBHc5lcdBbCrU+NCNk+X9jMBmV+Xq2jbpVeEJ8KiGXQYQxT/L7PcfCjFiq
rtuTKvcv2eSFdtjcE1HhK2zFjWg4U8CTyRFu0SczWhw8l96P79uQeoJscLbJsMsb
Hid+t6m+YBlXojjK6sLE/iwQn79x1r35lVweRh0DCcNzosPHCTH3NCFCTbrsw3Jj
ZF/FQzgkNq2hujWvSTZdjiE/bKTjcHmic0x8Lz6Bln0TBMy4r4S9Z+mQJL/D0jFi
uTdcaFqZ824HSP1wjMhuIkDmBMdJcpdv/DLBixyZFretC5qN8X/oVi40HaAPN4xF
0wXcQPNfXNPxBoFhVK80Q8Aggs0MwY9UsUEzmRJw7Ogn/RH56kPrfqInDAotynRk
2HmX1nZtv+U8CVWP2dhZ055nwMCRCszG9RPubsX/1VzeMyixheT+V9hxKLz2NCdT
BWkqo+rO6OT9FAJ89L+NRPEKFWT+bvsHuEmCndR4VlzVR8YikeQhAdYx5kQJOIm7
lFUNNJh6PcwLgye2pYXU5yNxBoX+TvVRE7/cEA9QJRYbGprs0+k+AhrUFGIO0FX2
/PAwr+KE66GNldB/QQZlu0xXCb87tz2iqJt6PXsqwAMUmeq29lh9rd525tNq4wt3
jiwtTs+J6rFr4duu3rsHA4OENfiO9JBA45wyyiw7NMXGtVT2D2OCFbO8AlHsH+fn
DxgcTd251qT1+ORYy9OYGETT3BgG4x0UiVm/14o7J/EBhi2DvOreomvV8c8PyHSo
7TUdnH8ejQVzNhvoBHGYQyDXwRFqjDcoWmZuYuGsiFY8KE8FYRlcZBVsMSPMsz+r
SxjSM14xN0iEn718t/zssM1xYkzEpGsqVuOQv5tDDlnB3JeyL/UTaYgkAyn57OoK
8f61R/eA3HgFBe4NT6hbxIoTStX2VRG/ptmgvABVl9eNk1o7Pc9OykvDzG2PuUSt
WqwJZBj4hEB+2LRVXYxEYa0obuVw8XVY2IaM5uktD60bMH3Yjr36Ue6OBR7a8Bkz
4ft+k3sGRpEDP0mljGoaPK7AyE+uMo8FlN/YsbM83a2Qb3qwVTbsSrPI+cPPcQUU
rgERYMII1ej4aXrC8/dcNGpEmpTKgl7zqod9w/XeNi9eIPqcwZBjCBLkc8j2KP1n
+3gMeI/QZaG4Lny7a9ipl3Kpg6fEKF9PfUczjpvFa+Nt1auyyHxqNi4suRcyAlNL
zHmq9f/AMytNT9Wkl7TdgpO4DVIvoJMZ3lNhjfeq+bsy8RdUsZtQf510VU/Hkdx6
3rjerMqMzWAUCSONArZBs9Y4FmKn9nlu1MygOHzxSqmiDhLcIedqTE5IdADBHByJ
qIP2FaH/l6gBuLe/fF/xvs2/KbLDNt5xXk8AEULaNLfKZSwgZHnmixVgQJCgfT7U
Fyelm0xiUytzzfxbhEeMhkjRxEDVyNSZJo3DDWathzBbf9jm+HeUAP07SGDIm+30
n1m3YgkkhU87YzRAVaR3Fp4oU9/W0Wf45wQOS3X+HSS4pnt2MLnVAdDVq7nhyC+8
sqtPZRhsojpii+X9VnOxdwkLHCJ5z3mb+hQ4k2P0ww0/UCwIdkbBgrFQpLtL9BXj
tS9e/vYmHe1JHvX22tarvOR8lu3cCmlw3oiCOwIpbPuVprlJz1To2h+P+U8G8etB
7cmasSwu7HYo9WsFPZTXOP4wig3CRp083oCvs2SUWDFrwR85Pn6Q/kJ5spYWLdUV
8uTh56091Jg8Q0wI9Q7SHpnWev9BL1cK2Eb0Jg8pkmouR5JFvxiUDWlxTYznOyFP
+qorNSFWnQeFxyMoBHMneFT3Zx6nXpgzKkphezTkzQ6o2wN1QI7efbK0doGyAhQj
A4Djzc4tgN/RexFlSjovOzAmCUJ6Oa4UFvOuTmfVF0sxBD6iVYJwt1Zc+2OG/CJz
Rdqx8VWtI6lbVjX5su2nCgnAicHqx7aBcFTg/fLewZ9lrVyw4pPAY4dL426KyWce
DgdKSg+h/lY0XBThKrMjK7Jbf3s+smPyW+mOGjOF/MR2g5QTfBtPaWtYhYWD7pSR
yZU2SV/weF6sRyBlVYPpaPemDpqM8UCzxeSsqHhmlfXefMb6txK0BGdtC4xPKxg/
xd223DupDzBGIFWldea8lJHtnPoSIvIALRQudmhLv5J748SJ/fRJ7UvjYMOCkeIb
0WYYRRBUmxY7NX2UF9lQnYVDIbcdKFljepQ/3+45WreeDrHKitRJCI4KEpH1nPis
S91Bfee2X7Dzc+ss2EyQLejyleBjWPbRAIhJDNo+stSWUkuWKW/Vxb9tlRqJWiqy
CrH60ASqoMVWXQ7bsVCbigih1kb+r7Jt4oTHRC8RRK7hJM1ea7dRj5rX3s5ZgAax
a/6ZT0tF7V7ADNtAHTK+Rl9a7l0GmVGLIJJD2oPcwQDver20wQeceVVAFi2QM8NA
7t/4wSzWj9mKCDFyJlpWBAxJxeQfyCoT8NhlEiSAeAr9hbGlMOe+caZBJA0aW5sK
uj/5iwGB/shDvIdUXwIgGoKSQU8hPJkuXNR94QdDHwAmEqv466ZyctWXxywfww2t
`protect END_PROTECTED
