`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zvlNP5K8KMFPFgkyTe1JV7w5XaRLlJhmN4RyKns2+1E8K30g5hYYDSKAy7ISVK1G
kjG0XjRkn3D+wGqbi+JQ0tntK6A4DMeuRb+8v0BlZphYYtg0oAjvYKrWTS4GhDrP
KEKCQtBzqEiiZgcgDxm3u+KLCcqxZxlqbEkL1AEKh18tbDmlQvZIdWExm3w4xnG5
4UfQHwLkNCWfICvTY69gIhwvd2mXOF5ToOBwQsQ2CcNvwEiEoOKZE2VIMavwEBjM
aQqQYvgLB8W73zzAQdshphrjtplwv1Qzucj0d5rzCH+AKDsYwI8/8EnWZRUlB8Pe
pajBdy2YHzayTgxJ45aaDxXMbszJqbF/t3PERy+q55PMebvqe2530TcQVbIGkAwN
`protect END_PROTECTED
