`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bv5euTfxbyGE/WVDD2+TFpgObestxQxXxMV5ITs6IcuzjsuwcrgHH8Q3lHU/1G7V
23UEAGx8H7p+E/1VBg8DNy+TLbZmbKSq4UqKQ7lF+/uBI0nBxHejNOeHlcPbIUe/
P7ct8G2uTxmbZGbUBMuVyVMCkW1+mQczqFB+A0CdgKI92TGtFm8nQIbq9jQUM29l
ia0wqqU0ZdzmUf00v6KkaN3oCEOuBdutb04Y4HruLwUnYOB43khBL9vCimwaKf27
8PIGNWzHI+4NG4yoDNldvMWxECjZ+FQP67YFJSSmoRi62U5AmecuvuG2Wh1pXnbB
/CsYU95CUoEmqoGqLVJxt01ZbSGwG4IyB5m+MMauApYy5xWBxbEaDvXKJ9AW7+70
EzFxQxXhRarBVOu9Z6i9UA==
`protect END_PROTECTED
