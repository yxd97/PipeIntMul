`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/8dyVqBWFyV2IHRRVfYrgua+z8Mcb6KsQDXT/wlLCcLxhKlWxsU0csSrDOxX2Ver
3d+VH3QykbtnIiOSoITkrp+mRlPleRjtO1/K3FGzIXNj4vfYHw0PD/QY5D5uib8y
TyXvdAxS702kZdz/rTu3/4GfyU9OtWng3QeaoU+esQyMJV7xi2KVVKoTgFia5bi2
Rk+cDQ+XQU+vrwJIDw2gST5XaxGyoIGJW3xygdIrihLCS4Kt/XyrXKE3chrPr1kn
26D456vACDemweZidLB/4CsqZ+2nOFbopf2EFzda/YVo73yfmQE6FDmm7Km9ROF6
BC0LuOcFN9oJWGAZGj+DY/zlRhtTe4xh1if0p1VZMFpaaf1ikLS67tG4L7lg4UDz
osLu1oQ4lokcIEjoFR6HbdhZpJ7M/n98m80vE2ffwTwCUAVpc94Ntp2Rp/B1twxA
pgcZjcvBosnNSnxVm32oBGiU2Dyt5SjgdHBCoos9mMKXgUobccSHcp/DN1KJMQND
epVc0ZFxxtHbuaL+Kr0AQJQqZVJ6EQzezvHiN7D2jy41+091u/s3v0xGm/p1JZoT
WhxG/WWYVrZ4fIl9wV3/pgEHWwgGzyGzQiBgjAd2u5hxhY8gz5dB7EsXKpHBZRQQ
Sut74hhYRf0vJQsHTh+2sAypi1JboJ+DYpRw9SxcdC2H5QH4tx/xnV1Bye8d2o2K
zDrrtexpqmrMBBHP+MKtWe6eERBlzwgHNAJ1cmhQ0AROjYpv11KSU3G2q3ki4cfq
7ZuCM84TAGnbeAl1yuJdS8QTBv3G8TZPKrkcayH14eSruuXljFIJ9oaOGTBNH8ss
IjdzIp9mtms1i5ny4wyEwmoGAIelOFult7/UMNW+2gSJkPQ2oHa5FvRtyhFVw1Ny
gqAZFFwGUsNGvrt9Tj+Z12gNmA4YpKcKjUARqltZqKy5BxBgL8if5Oomk+ZUZInE
2uQioo/1pnIApTJ7AIqfjOL1tTDaDJJdk8L8CH0dFex9hkUuwx92N4rG27AX1oNS
rp3FAQKDs7YAyt4lzVCC0N1dk+U9KgbzvuaICKh7kzCnh/3kmpa0q4pm7xwGMHTT
f4DdONfGR13V7N7Z8vuf7KrePRLsWgUibpaYgxcKiZJMoBpuQO4Vv6GW6P5rBXJQ
4Zfrc4ZITrIJFG6dCgqs+4wEkL2lWJJMZHBlLynXXEtYKSYkVXdi9dVxOzqwqS6f
9AyVKyBYuvQwZvd8zlQjQSOcDUrLO0urKgug7J2jEb4MfR1MWU0DfVkTqXa3JZoj
6SMD++ugvOcFHFF0RaL2M/555VRD247cbyvV5sbFBYj9CN5YFURnAMNuuzuAYk/C
9me9d+ajCedBpC82BaaDTwJhYwkOwI2qjh2shDGqIQCtHJomxpxzQCKdiEVYkPqs
/YelLOOp0U+Uq7fiA3eYRIZT7l0U+R0+S6YTEjYHS6+vdSVHfVwAd5HxMLDUIycD
xH8GHfmx5O1WwO9hCY8SqOI2S0QnBRUcP5oRqdg2XDqyZLmfo8g7QLAtxMffNuoi
v+UgVzsMj3bfdab73+BgtdNhO9ZzD8dN/sVkmWZLV8OGDNgXdFyurhFVw+iKrT4c
FY2ycRY1HIWnl8g7m4ozcnPBO1JfdliY1VGHdfVvIJch/oGqG9TXryNWuqxyvcpA
blSfplciIL8bdyV6m2aQe/LEf0x8sG1LeaZjSFHwjBzNzq2rJyLheY247iLZuwj5
RuYgm5jt4NoFzSYYs5P9LRaSU3pmGnhxG6rZOFada23Yg3dPiJY2ynrWq4fO5Ywp
GPkGTcDNwXJGe0467N8DolA2iP2N3CKulGukBrnNMXwlwb13CYtJkMOPrvaZp8Xz
7gPhkqldrZoht+IjTq9fYAxAfj8SVaPGHnFO/WtacYaMM/UYPfm7+INF3nr6KSlF
oElLpbqgjWp7bjtnVE2GQs642WAvfC6zH0VobSTMZMYfRQL5nEV9mHr4BOaOS1h0
McGbB1qtV2qugArzq1sYInahHcrmUQW4jMLnw+WzQDe2RUB3KcOBLTu5ed2vVGKg
IsiQXnWmV6tL89yuBiZ+txAWpBt8E3Pk/G2VB5T+DoCUB52wBa3b0Gmk1v2Htugi
n76v0okh5cvJ1xMBUfTv7hIXEvuvBpFwuO96+5MIMDv0kRs789cnZyFz8NH5l9Yw
DhA55eUJNIDm0Nc8ONYYxAoaLk98sgFr9n7bS18WLNQ=
`protect END_PROTECTED
