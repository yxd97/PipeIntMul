`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1KGWJ9bOHg0Ppqx9Ruf7QUS7Y7LHq8p2ou/8AZ8eRb2KrGQ0smCQ2vgJCUdm7B/Q
08RDFe0m75UwpZl5+VL5gUuAX0ur0bHq+AIt30+/C9tcDtILrXIhkXU5g8Ib/+8m
jiOBTeh8jtL685p1pv4P1gXjnhHddYEsW57kgfcV98fdox09Fk6JFi1Kh/fTvvQL
rxx6z3kA/UJ8xhet8mbvkt3xBnMyMO4nrtO5m3ybmuQtLQ2tdfz2A2kS0Xurg0I/
SsL1QHVY29RovL7LRLHv+JTxV6NO8PXg5A8WlYuoD5a/XTugD/B09jyiSyHr0GFc
rZr1G4qKlEsNmQQ2XwJk+8hFj9AUGLT/nVpyEOd/cRgLDO4mPUDW0BiDmCUqn5i8
XTZAt6zjWDQQO5T1+c54yeUBr0qLFmiXlsf3ckH21NKze8IaJJ/g+DqyGTrB/8OR
`protect END_PROTECTED
