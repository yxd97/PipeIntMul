`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i/SXeG6yHkaXD7zUBHAMy0L6JCogZ17T/umzbb55e/z92DVYXcg5i6RF8OoCzhYn
bH+ebfNeBnc4Yujxgz2eZ9CwGuloFUXmb1plMvZrT9H6689TnOSf+x/DpBBcHif6
BnF0tZQI1lkHj45ZF7kXgtPok52zIEC3y1e3WWQvVvudWQ+sb47TefkOnmNRgw0X
E1OeHZ6ImtJ6amFPHUH46Cr+NjLHAaxj1H8SGpAwk+BcZRIZWZn/HCwL0m876osW
Rxb5wM7IL9OMCHruPC6QCrDfJYc51aehhIgxx4xABzczPSZwx9X51wR/QyjRsoSN
S/rekLVTU/VlVAd6Z5DFvk+eGSolcQz4AvR2VHKiTqp32fpVkVDlIWltOHlOak3f
NsSjjYYYDqevfHn6CxjlvUChMBsKAx8rx2ILhq0DbCYpMFfBVGsijNYzpBAeMZ8s
AzvOAO0mhYygpL8vPcHue3+D4R/ICOcs/o7Ut2bpq91TOjyy4bE4loq4nRxOG4Mw
vNBDY4qDUe0FNCCGOaO1lJzlwSDBg/PNCwK8RN3Fv7Jnkdm/CMelLDhG4J/Zsx4V
`protect END_PROTECTED
