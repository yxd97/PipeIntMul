`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kG7fFL4rtX7fS2CY1L2CxMWLvnChXVdDRABMClMJ+BWxlWIm/3gvy14jJtW6mpuy
s3c83ZhaipCa0PFZRLxSmDgRZv94i46Il/YQ9Sf5ahpYQ47ZJG+dTzSYj2feoaBr
6eLOPMcSIdXUIaE1nRlmU3bv+M/WyImES9CQFsFtQ4pv2crRgYXl58UZEwn40Vji
RUKjpDSqn4gCWdZ5vwnO+dqxDOEccKsVvX6NoGIkhEH70ipiGV/yl6MkRqMsDoBL
iGARlSubg2SRccwK9n8Ol2OMyvg5GbH03K1NOQcbs9VlDcPNYZKBL2OMqGsN2Ovl
LqcD73IkGNKKxZSlt+N/6QPIOK6gfRGFFnhw9zKW2E9kgJcuBQuE2gms5m1n1CXv
u9VqR84XDdI1HRbQV/0e6dFPT5cl3kVYvQVQxk+mo/Q=
`protect END_PROTECTED
