`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wB7a4CFsMj+yQt3GBvLYlXnC4gmYwdP3P9KVX+3rIZPHO0CBKCkr/NsJJQTU7bjd
3OUt+EKBUaXO3kq6CfJm8HxBFzyIWu/m9y/GVbh4vkux5X1CACUhdeqhVL21PFdI
A/Fi6pbee1pDgE0oYnx/flhWO15KNHOQamVsJ1SEaFv6ywXNakXxW2xZesyYa7pP
pYEu42nowLqEOnUN9U5dc0quKU+MmkJyOIRTRFOV25S7G+T2x09HR6XOu38t+Pe+
Xjz2Ly2/gqURX41eN2ztAqH90Me/6hd0E3kPy0s0FMxnKsWh+h9APPbaO+nzXkTF
Mr+r1GXfDIAZtzMvEaMYrQ==
`protect END_PROTECTED
