`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+6AFG6OsK4CTaNQrHzhBuWpI9A6wfL7yl6Vbe8cTcV5MMDZQxdn9FMJ5pCyEfFq
3WsXTReikj1UT8iI9XFtdeTvDNIaX2klq8ufFCvef9TAdPQl4j3fCbM9o+hq7oZZ
2OujBBEtIyUSHise8pIvi2rnVnJmubMCmKdLDR7tfE7e2+57FKZ+R82a9rHnXmPQ
hhAXIUaqHvtSvh7Ks/sd2jyPOZQ0prJzzlteISA3bbrhPhHw7i10p5G27cLpxGkp
Zqey2t+0dByrzllEJjJPm48AqkmpCTEuP7JsQ1uzEb45DxAG4N+EtS+mSjqpP+77
U97tyL9xty7beg2X32+pNEEqiqLoquTFgs8ss1e0pIQRCRE3H3RnnbDe5bMVmNQO
iNcxZ1/aEpIbKP7tcpdOiJDvBdbLr8VQhiboNzSjwfR6dfPdoh94shgCH7oHq16v
WZAPnRH611mMvpFeI+OoT4N/Xd5EXxRPS8xd/lSny5mKLDEyYpB8VS13owQCXsa2
dhkkTDVWfkSdZA9Rei4DD4tn07xGD9O4DrvsqLkaW9cvQyOASog1nJRj8QWZF3J0
8HUn4SrBhNlHxa82rkbBW2SLS3VuWmg74PHt4LZilSEhR2iLxurYOAVrLirTOFT8
OhRhvBP1lV6xI8PG1+acWCNsn87a/wOFPJkT6a2UY8/ik3pzwp6ayBLl0bSbSRBE
6RbHVOqn3gsSdpsT3+nX9pGvKloQ6RxUnuHBf13J74HwR3UsCpQ3ThD+FPJ71Fqs
5dD/aE0OVMgoYLY4d63rofm5Mujvi/tpzzH98/sP31ECqUSyC2ogWa70zFRTKIl4
15CUqA00Y+Rqwkxitq3bve/Q9359tVFnw9SamMauquaRZd4kj02z/1OzJqOBdUP7
SgDW+IVXLIE6ucneo7zzwuPicSYJuckPrc9etKLq76kL93EP4uxe5EwFz/oa0wvc
+LVSOSGiA8xlTe/npFHrIbEXBmD3j2JE0w0E67bm1VEcDIhnXw200IIX8K36Mr3H
`protect END_PROTECTED
