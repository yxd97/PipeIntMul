`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Suzu0WU4xyjQRaFDoC2IoX/SG5NB4HEHglgDkNNcVZuXjWyN850vWMQ2T142bDxR
NqbfwboTs+8qnqidbnH9ERmU/fOFdLgCREwN0XYENEszvKNk4snU9iTIInhcRxCg
Y2f25GpTS7+P56uL3hEN8w74V9ZrU9l9bT1JktxOCG5toyFIpDQVHOwLMH6r/A32
d58UNhS1ygNbObTa1dMekZ3qQQjnpsbuhQwQKPOSar8mISx7z7Y6oBFGYn0XC17O
Pct1t1086xK/nWze+ispLr8A0Ej1RcezdSt+3h91+rO2m9eEzkvU9RA7sV7DKqvs
8EvUEMRjhTdxJmBjcFhF5TCFzTJ4nK2tGvqR1uW9OBSxXWs2QgZr9OaT+TB2vZM/
iyAEANnr9RUjFLud03elNQ==
`protect END_PROTECTED
