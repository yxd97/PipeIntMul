`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BhFwVgPpwq4GRNMWTQCk1utbe7RecqjlOUrSyrUdRLqu4O/Kpq2Og0zd3v3sT2IQ
TE071EZC/amaeWNpzyJPSLk7whjZz1DrMEjUKX9bJnl/DzGlRh0NsikxS1MeId57
uYwTf0XlZsVWBNBkSDs9exkV+5EAt7kDECPEze1hwpKIb0A04cp6kkzFy0Z7/7w4
o9myNQKXout8QmpilL+hExhFbJtl2Z8AciqX8ll48bHfSU0E/Jx3Cfwu9+mdTV4R
wGjFr/uR6T1W5vVwlJNJRRcGjE7rNczGmpK+RjGEg9a5Pymy/eKwdMJfgtfqfdFw
vLQDCsORFHoStiJwulaBTQZIWAabE2pYw1caYSwhTqRegfZ4MqRF6kOwplRBpzSB
twEOOA58UUBpGuvRP4Jw3PSzAJ1b+udssp8e0DsPwen0PLqg0cO8ryN07GwOlDB4
XkvCqREEg5a1RsCAmIAhrHmy+ZA8j4OKQttZNbQ5DTvANerNd2q8lZ7m8zfagBbm
w5HWFeatNyZQZMlQOzgTcPUdG3IMyWI4Qr/AYH4j9y9sNzrXgHoYwRcdXXQ4UPv1
iUg7clniVSW6jZ05daQaJOXsM782PaB07epLMpeyDdLsVeuUHPAlK03Y4OWslv4J
jTX0ygGTBKAko1z6Ymp2LNdcac4YeNPOZrpR0IXHWt0iIN9HdMwRjqSi8GqakIlZ
o8JKlEjlHGOWfKX7XmAuDnjLfCzkB0muLCfFyb6s5fEB+qZ7gOtK3yxgwY6ZV34Z
IDKBnvwrNuGefWNNvlSyiP05hymrSbt5vDFMNzszXPHTMTh88J6pIcC7M17esaaX
3mxsyKgXa6yd5B24y2zBSny7wEmhXxV71ip+xcT97YDtuPGVzC/HxHAG/oPCYwUi
dLjO2uNWrmib3tUQtoIq8nlX8bW7Qtkl7D+VlcUhI4Hgidjgp07VNP/EJMNcY2cC
Ose5rmo6GV76i61+nDF9OLM2C/AJJ/EjS1/mMGSIiohdi55mIo5ZitRnFFKNZHY9
0TQtVkAhGo1D+WsPhkP1v/s12QFV+r51C3bVjXWA46R+aF0FeO/67aD3jQPxw6Xn
F+6aNEMLXPi18S7lpV08KPmVF8RkVOeje1xG4F+DKKhZNEf1g3cMle/134gPwsfC
s0KUm5k8mSyXr8ombx9jcQUr1HOyoU04eL60fm9hLm5VGpfcYZU0y4jna6jSN8s7
A/9mQqdPGo47KfDof+Lmi9WuiBaEn8NVME2gPbNDDWfnB0b9bOxP3fqVoFrW130m
t600aRgtR5CJHmkDOjXhstNM1PQnNcLilDP2JBH4LrKILvG3a02i/hSEVhHEVW/x
GtD/xOthHOfahoR7Ej1PnS8ZWIF2dTAmtnKo03VuRmOrf/1kb3xdBetr4CfWCvb7
9dsMZnaww2b5OLjmJTykGw9VQu+zRcfiZ34626fxyZjyRqFXxhRM20ZQHinjEfXS
y8eSlzKQ107Shcrj/Gkh2REwlfoydjIbsCzTczGaQ7guYdbhgYLGpzCqmKbdp2UR
2jREDh8YleC22MVv1oldS9V80zIZ+DTgunEc+casxU4CuhkIxP9Whs4PXd7pkNx5
QCqINGskp0jeC5dV2XuHcElrkHNgPMa7XhBaI2X7kiu0eZ86HJRH5mWK8U6pRs8J
RFNmoQl24LuEbetlactCaZnT+LSdCy2TTAqHGOJml2ySTZe8aeKjowLEZ1k9l+mk
jKvO9Ete1Fp8LGpptreBZcNhHupuAtrTA6w82lQofzFZVtsOECpLPKHSlRRjjyTY
9TkkJmROmpOXjHQxZLhgC0n6dqWQc+DsJiBXreQARp+w01e1HwSSjcaF/bhloNUV
+lvY6QAKVQ5Z/VMnu5WqeImJa5kcMezOeIUyk8thLuISeEouzLGsfR1NXhfATzXh
I7CXIHuNQ/w6eNf9YaMb/Y/zhnC6eELB9yqhffqOa/l5NXVgmtdWwCP4brhd6nlI
o6359Dm1b0OeOCNxWxK1bNLFUMJiUlDIPcm3JbJlv1gDFetf1XDmx6JF2QB4BQ6g
fLONpAW9OLMOc/YNpqmIIKetmmuOdtQq8lTCBQwOcR/0+DnS9XnC3AQfzGOLhbiv
IWyEQxCfK3fq2I5x5u8qCWvi3AmIWhMswra29ex6YHIk5UzB2iM5Ieol6DYz2gqy
0GPIrt5y2TtHYVQtG4cCyAXOByJbNPo3XzWuqBfvr4n6P+zhy6sfHxhkG8hw5k1y
W7yGsbSE5KDGzVXg4o1iDSFtEqWXKQBCwOhiQ7UrrxbAJ4X6Kbg1c/iwDq2DTxN0
xEG/Yjs7VNrNwmunDQkBgZp7aanKHKNLDnRyjXU8FfFRrIFDNDyD/zDSLPs9K+tQ
+nmzZA/2r1+7jbZPliAlfkA7JEUWFH1ZkF2tKGVm+1aEmKihO0w5JMrDqszsD3p/
40kRUIq3/NBccuXQ1x7l5U5i9d2e5ODcV01uJWXwVuvO6Yg60ecdnDaqk3++E/V7
C8mdw1XBH8uFw1qiNEkF8ejzvQBeRmYkB1p7eUTjdMibCNEBlPvg3R7XTnpIPKj/
J0UM+CJdIribIRVA5IzUfX/G037i3XyipXC3IX9aGQR1nHEkYW6faxdoy9YxchB/
Eku5dNGzVWkrvP+3XlYjs4yi1ZzxDOI7eIjFwUCEF67tztsQTRBgockj7nuT+xkr
oy1vwAIrsSazspVIvfmS8OFsOSGvNfSWlzntwIdVM58StHZhBjaXaNezX/bT/7ys
uLmGykFdBeNQnkk2xtwZf6/z6Kw97WUOCZJrJwo7kuS4mhFN1+zHG3qCIpaSe5yr
BKnUUorT2cZGgbxeiqJvVM8VPIMoNaihGLFOoPhi6oaIM8lGRYBvMeeTEjEWwEAD
gUQLl838Y3pjzGLLsBV5CXH8Byc+mHAOZUiHHrkdOk0FOIYil8LRDAPpGtCCsx9K
FGlx4YzAbc9LJGJ8HYQJcB+s8i8stiSkHkA3+lb31bwPoY4bw079PWqT1v4OtWEV
Wltj6BCZ7Mq3zFl7U7zgOCp+0MY4WmSLh1NTqNTuWCWUJfqfCrbxQUOQxoDg+o2H
1ocwsLqe5FLdxiSPsa8bFAye0EvFEMT2M373s+WZpmdIASP3T0yCmZmiSgfQTnXc
GTslEJGf4krE6CRU0n5TB5jzp1Mq29Yci+xcrNPVZBGxSeijWJXdTZoU3dgWI3lb
jPp7oDWMv2AoBvoClAO1ya3OwJckNRlhSjESK3Cx08npumstYGGx5XzE8Q/p7R+H
bSewUMA7JmaUzjaVWPUurov9oyaFRkG+YrfvYfufjYj0lOpWrSwM0qZ+92CNGYYy
elFTiJcjlPjnFbi8MYWzPcutM72aqzGUDHKoXbWMI2a1AiPZ1xJ4dt4MCI8u3HyA
9+mGRAdifOd+Flq8gTv4IOjQvu/YKl8ORk4D4wHtajlIvdbnL3xtDYaYQwJI/UzJ
zD6aP4mxKhi+lNtPyZtEdpDlz9Fib9KdEiEKfHhz0MODSq3Guvrcfk2sdTsweFLy
xLbq6ACmzsMmxC2EI91dbJCO20kz6+0eiRyFCuY7bbzq0uTjt8so752IA46LUIqe
pposZky4hWivUCIKZ8LOnDPVWc9D9KIMyQ64oTkFWgGiMAOUTziJ0PiwHAnNjYo2
90p75n7GQhiXnpjuSdkczYBoOvmHU0rcsHyJzbrhgIkUxpba8TXbtbZ/tuyWejUd
hYIxwCPET+8YR+XEi2MkBqH0BELEs1x7vlW3MuqGb5GBUjfrKW+DupSbPWLiK9Vi
j6chUG/HSfQUcQZ9Z4uQlKV1K/wTNa6z3RcMajkXwIQ02o7N/JU7C42dN6CX1ABx
JskL6sItVkMK3Q1UyYixrxXd84YvvezyrLQbFtZCXhfGYdxlTknB/XZScv8PQLtk
rnAeGE6wcoq+iptZEgqRzfG0ZaIjRqaHOH7pNYwSb7/NrDgwZiFCf8rKWA37u8M3
MGBO9cjyKwq8aLuF0CXTTYPuJVdEg83JrZElapQsEQ7WfuxJmcUohT7jWsDMb4PC
Zd/Pr3032Tk5iZ6p+LYrWjhWUjP8jVveOXfpkOD+kDTd/xk7NkRCP3nO3l1YuEG0
zmIPc2qtq0VjNzscjGQIaEi2vCSwt68zGIqgwS3yv/lFnUmG+lNhcpPCbrwLuFNy
YOZGWZT0udPvP/xRQAz6b0rZvg7uJj91XpNNoyN1FdE/fl3T2lsVjUb1QsaN2+Fi
stZOcZwjnmyRA94Gc1zwmO6MWg1yQCgHtiHT2wFHcD8urXlCykpBrCUJSyMQVLr6
uurQLcXfR2vhdhZuBrF92KRKf1+trtJ4/4FS4FJ09tKPzhwE2zhsrgSZtDLNexxw
fZto1EgWn+Wc6IRkhcmM6sNgJob/hKZbAg0SzFIAmSVlnM0+d4vnbW/GZJKw/VQt
aF/S7NlFlcPNKGXWBMvVsqFVTPYwjvB2zBh6X1i3FW+2h6dl/2zOfW+Ar65cCxcN
0aYKvNXt3ns9mXjvKfavj4uRk1EWVKi1Qf4rodJFqItD0ujz0cl+6fsGnxZpED0E
8uzQNZhPL0IAervpLammMsgKbKyi7ZMfRx/42x8FGTmH6QQeo5p09apVn3lz+LOy
urM+3lafSi25bQRrZ6fyxp21WSBavVYPrqN/Pamh/dZZC/XPzcT3XaDMrk5oBBkQ
Hmk765FByQ68FVLPyZr2zpIleaqmNNOZOit+ey3x8IBVmIVgf3KVcavX8W1TJ6zI
dnl8Tw1Ymx4ByssvT+ELRIZrEmwe1qDFkZ+3hMOv5rcnA6jW9CTx7oMd0ZItCRjR
xwMxlHpnpg+UrfsGnIV1DMJBhFyesFYmxqzgvEMRa8xKEx3gfZ4MRoSvspW4K4uB
P08TiOGzvwGNGjAKk4hZ/ltrst2/9GgNR2+wNs1knDZuVVx2D0VE83mjFu4nZRmS
cMMR/eWJPF+fEUMno6fEvE0zYZmLaZyx+NfuENpZu/pN5L4ub9lKic7kyljJTnnh
WyRM9MYESukWnGnOgmm3yh+yBS1VRRNqpHxREw0dNw88o926wg0c40z6wmWh3xwq
iuzUv9rJ7FyeMmusFuRXLBtlCGPr24cvLUUKfc60IC9hf6u+CUQZqxAwvMRWQBhP
twq83frSzmqxrMpIqRlNp9WGTCtETyQ2gOxj4GVr2FMKW8j5Un6jYH+oAhZOZnEw
LnY+Bw8pOl5tojlwerZhBWcOYfxdbb/DlkY64KfJZnwvi9vNJdRnI3nepJxQCinQ
D78iUVJImysRW8tJWAjSNH6T83t1EbKqswYtZS7Xj2CEl5b6kc3M+0ApoZSIe9da
FHXRn2c/v5ZvrpA+zzvhZqJ6KoPOHGyBE+33kqDqrwBPQiA8X2E0yks7D9pxqzpy
GnwYq1JCiD4HnQvcDqYrH4FdwcdFUkJWdbRxSuoqjQ6g06OkbtFxWU58AQJzydGd
qtqBFDBbidcrr7/jL7CKBdzn7OCn0M8jyFGPSt2Ko/KgC9tmCGjcoMdYm2L+yzF6
MlazRLRSa7vQEjgtR84Fv8XCcnwqKgLACb5g27kxUozgk7Gzwno1g3wsdf2f5kuE
Kf6t/b15VvUahh53fa1Xc/dikd+ri6crELV8N34cZmhv5qS+VPCqU5QYr1cWtglj
kFj/OnYurLuCyyDiGrCgFTfyuX+3AH72NQ7i6gHUv4l6TTFkwCct8JnwDCxsF7+m
Fuw2LEjDtTr8wXf3HIXuNi7+mrDfbfKH2LjuplYU2IqaqDepiQGgAvy2bH5pv/hi
dQcqMe4ERqn3cQbdR1IUgJ0X1tw9ALm2xDz4VqZnTVQNYW4KLp3VF1k56ke8CpTG
Nw08DA29BhBXhIo2CEs1riNYN2B839OSlao27hpUJTw71A2qvnHbAECXk/Dup9pA
9XdLD6NBNfq9Dh43xy7ld5T4XRhUElssBv3lIDwYE86L4X1HW58eL8TvSlfit3qK
yxGn4RQO14Qm69locrb3nPL/NKwfc4gl371gF9VDguwm+skYZWhdSDko4unJ2o3t
YVgQ98lPmbwqifY6C8w8SP9Muok3ApbXLtQ45Ls4H54hnygvse4fVpx7zYhg6ZUq
iWntspqbW6ISyosMcFpyrycVf4gi0zJlXnRsGeS9iK0LmhfJ3JTJ4p9T9Sjk3RG/
qrZwF4eLWGyP3sDpd43F9iznstuaQRkvlj0oodbrIrNMp70ynECq+xjV0GlegwiZ
TWlkTdSb+Xd8yA9ICvSv996FoYhDS6mQA5yf5X6h92ZtjBXIjSbwLC8Z/mD+LRZW
plUsqeyu3mCrWLzO8EQSAHKhnSZf5Q21GZ+vLFJafMjJRjUQKosjMeUZt8shUoQH
6EuI2f+yRC9mZP8UUMi0pi/gU+o7tpx0XyM+HdRL5jWUsRzzM2ZNfKk0CqcQ/clz
14+NYoxGz0vPvweAFy/4wgrf2HokTpkugg2f7QgCh3TGNoC+7N19IoQcXY6YIpHh
xOljsmWgQATE/Vf+vq+1mHCYe3WPID1TjlnP9o6qwiTB6d44k6czqtmIIR6HEzE9
3RNk1tCXyINPDw9xdWhkKjR9uOqpc6jSkNBOGT/V1+6x2MoVrELNc1NlPORK9dVs
8J7TY3Z5+4QwVNeFqBn7kal6I3fGmEHr0IZZsvhoGdNgg0Wuol92+1x5Ha4GVLap
rgNjSo54caPA9/5zft3zrpxNo9fhd5qLVEeQLcf+DlgArUUc2l7hn9FoQilJVuYy
PITQZT41V2wU4Gc7gfGHIgod4zq/Q6cPrBCOyQpYzpSf6Tm6NNRbX7n8YQvfpBgI
gDSS1hlAeRB8M64I4vIlNeSLn9g38N7MpHfQ9Y1SmSJSY8KJPgCQ8LUuArTiAxUk
mhJFTQ5SPl3/6lneKBIPQOsLfxk8FDJZL3VwQaZL/Tl0hTkaY3tX6KGjq0HmIxhX
PidCXuRz3cEsvQbVdyk+YnYLDmxp1an/3uXMZ4S/0AvngiwYxk2V1GtVw3zZ+o0k
PQ1RF0P21NW+XrPjTN5thU7uaa2wpjmqFRz+LTE2J7HjMTmppLryqkARAf1IXBVy
t2LhoF6RHVm3DvPaw8ZHnSabUXxFZ8knnZ74A0/lT+jMhLJtghk8SlRWkCHoFPqp
751TWZL8V6jNnP1GLlMIsI663ahC1uaFJqOWfEDYfw7ZNiyDqa5GMduxqbxiOQ+E
oohG5JXyGCkpBrlBX6Zfqpzcdqfv3YdSSOQD6NWYxAUKAzfUqRY2zyOFkT6Xw5e+
jBDN4/ixvaz+zkaENlznHd4yjbPsbz+Q1meBqWplXLBFmX8sTjfrB8MJW6eC9iNw
FENraDDYDFmLu9J62yU9g0Cqg4zfHJTb+IGZ9N4OcxB7VhH5GnNxEl0LwUJpwwU9
UknSxa2JSqn44Iq19kUqc6odZ5Kwfa5j+K6BBnjruUXGO6M58YMMw5/kAov8OBAa
U/AHfLCl2/LMvGS/zaSp1cCHbWHHsJVbRTqWq8pps2KnmHfJkjw+Sx6GALxXqjf/
qtL/bzBrxgAqMtl2rnttoVF+yakEFnvGrQ8HZtNiLLzMuZVVDN5Iw7VMwRWXiLWm
`protect END_PROTECTED
