`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSJ2GnfgWqyNDc1mTnnxgXpXpsZLVLRMLKeEdBwlz1mHidqlyqGHjWi0enUEp2qa
KkF473p3Gn6Oz4yL81qZMX+h0t3oIWGSWB8rQE5iuZ3JiI52mmMNREeMvaT/l39h
tjmbA4Tvyy0kc2s3MYk3jdP9kNTsCKdOY2L5JeSJ1FEWJeBuQJr8PGxuOkyTCyl5
XgMOD9FCZW1eSIJUPTSleVvMNs1mjRQgI3jPLC7vmD+HshumpP7wATnoorQyIcPR
fSG0J0olZgPQwt2bvcohyey2v/QJnwssbR+9MmjBTjIMRQSX3zYaUNwb2VY0mlNo
8RU6733wr90YYLSIwfFlX0/kh4sJvhmuRgkGygAtv0/GfLx1RwVhW69EXrNCh2vM
KNxHITqqr10dOXFNokkS3g==
`protect END_PROTECTED
