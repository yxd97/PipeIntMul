`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aCnXPQytbDkt/HuXhkp8JhPUYFihmAF6beE2hmojemzxANiegYNJ7aBlGLjkLEDC
1JONKepJzHLgbig4a7rLeeSWyDV/Picc+ekGxEOxhamLUENr3DcTY+oY6mQuqruR
weJBTEvWhlndLbUupkVgFgrdF1140Fq2LMuNfcI5Z7Z01ii3BciMQUaqfRhKJp2g
gxtLmmvqD/GjlWF+2KkP4zSNHY3EmRKCHTCnOPVkERmJyTbVZ3w208+79jKe5z3/
FLkIi/D6KFWICpxAlo1lhhSIqFShDAk/FSId4E+H2OSgihTP0/uBh7v6jMLW1mY1
0lUFGPNiQbWxf6/p2EboWRty6v5IRtfiRWoSWtKuQQI3U9NT4WCzXS2VnuNY4eYX
ZtQrVNkHwgkkFwv0Icw+2qWPM9NqOP43+bE43S4DGPoQdS2UaUwIJCdl3fvl8qF2
YjEd45nEVZfvJ6c88sXFa8Q5UFgCCK0BBOCYT3T/mwvwP1kWOgdA60aaBlWyga0P
KoZQ+r5pGktdKF3KbDecryuO4s3DF6YsQlWs4Ndps1QH6zu+uQIJPpW3qWjlcsEX
Dlr1oayr7kMqyxbEMQftOqFTNRbnMAWbCIeFuw3N6dF03O9zXba5XdWWKmuxM01l
AH8Qeph53+GnAtNTmX35tfxDYbQZSkheERtfGGB5i0gDI5B6Ar20PSVy5nnr/5o9
`protect END_PROTECTED
