`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kcIAtbh7EXHlPnMFN3OdTK9eQtYzAnoISOrLPY3q2ob8b3cuTvm8uon0YEj9fUt7
KbX9khXCA7YnRPSNgJhfgug2PMgaMkpCoXuC46FPhb6sxe+AdIPiZ++wOqWVMg5W
70E9Pqht+0swDJY8wmp3ljsmV8UDOV71XcIAPIBqg5BMMu0aoanli4VzZeXNN92Q
qf+5nqDnjuOO69ChJeGN0xZ9gZCt0fdyaY7VhDfSUDWJ8MQhtFbzMRPRFEevtipT
Stf7HTkXslCGdJCEYSydpQ==
`protect END_PROTECTED
