`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cdbpjQRgIIS+zgB6duRFBs7+0/urRZv6uk78wFLQcXPpYkoYhzQcnPPpiUoQ6pr1
QE8SeWHrgO0GqUBp3BdBnb4IFmg3KUfAbI3VP3oGTvRTWOL1fkBUCBZSoaGRqU+b
YuwaV2bqZkqeA9Ygt9cE7nmDBTUU9n9E99kxnFbB0MI63cHFlhkDk3FKRosFyZIb
Kdv6AQ6u814fF9sl9yGC14Kex8UtVh/QH/tQ9VdrwfFSrVZWfdoNgJj8ePHnF1x7
aF7TQwC5/6Q1dLO4TjaSC5KmC4l897bCTDTySvJl4RFRgbkx4MiccRlfQ4Gocmhr
gEi6Qu6Zo2qvNCfMlegb6fdsLuT65kwN0vjQ30E6yx81HCaKNAQgl8Of48ZngFMt
ETJH4vUyAp/dscUBMZyPFUDQk6tXpIutHvUsAaOASE8glcpDQk829nX14AdJbIcU
W+v09aGg9gIME3ERSBC73ii42soRuYS4M2IdfZeV1B5/IRR/aCF40OIWFOM3I7hP
`protect END_PROTECTED
