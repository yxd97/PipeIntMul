`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84bV4zunqbYhVgD/nmXyWoXtm/6pM0IACWa+AUrzsqeFumU/jf005pf82Uu5QXjD
yh6CZQxvaSfCEAJZJNhfP8c3xZzMDmqU9NcDwXdq/xW/7X46PYZyQykZOjCtSy0E
PUsQeTXyM98goehoKuIZIQKjIVwOUxBefDZXP0RW0lYIBOaoFTnMupYYxYDt41y/
eLFi1W9wLsXQLNPC5BfK+aQ+Zr/pBmAN+i6Cz0tEsTEV8j+ticTxh0ifUvi4ZpOZ
mpOl8ysLGsQ00T2ffCJGM2w70jSLVbWOAU4WLwe4VRsq7crMj1otDZHF4wd8WjaR
HRvkw6KlUxFQQj4e0v0/T+IWjyJX8X/JsTwo011t/K7yfYriapH8cpixCl0LCjAp
R1Wv736rD3bRD/gUPieu5QMpNboajikDlzDmboTOtZM1mH9XLqaFbNuU8A6tB4hd
pOT/iLALMGRt1E+cDtsM/7vXRLiMXTqzhVw7rotP5lk=
`protect END_PROTECTED
