`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+dhZ9pDZePVmrXYs/xqzEyU5S9Jw/diKnwNG82W6li6ROdcWLSR2ZMNvrhC+oST+
+VmeQs2C6bZS8BRg8XfvgvAgkJ2E7HlGva6h0866QVvb/c13mayQ/e5YgNRh0nqk
Yaz5oEvdoTF73i8QND8Ahh/aXvPnIOhk7nurss+x7/o+HrKLpwJK94mRBFSNcSxC
RpwhOiWFHh0+62CjtSa4mQjLat+kUyqH9GXFwe8Lb8hGaVpxSynvwCvmQnZasCtx
YXuowB/RKwjXKryQdavT5C8OeXMTnuHgrmApTe4R0rXUS/mn3WUUguE/4En4FpSi
hcuR6u96vJK/iFTdtXg/fTqBWVEfE32exMjRCyxal+v0B+VcltLIGBKkWsACs2cL
AFxDwcdhLipl7V0/lassSZx3Khdcv3gJTwGWSgwady32z6/lJzJ++Jf/ScZ9aByI
kEDwPxWz9+kbGYKR6dZPjiZjcWugB35NMRuKhMsyeluifzQeMWhY33WhCxkbv0H4
oRVY151mKdJLB3uYslkojJPFkXyH/QEdExMtGEGODtrS5MTHGUlL7KAuEWsUTdvi
kztYu1jkvOmQBey4Gsg/pikY+wpifS46If63Lts9ZNjObxWIMwVlzpCmFezSJwnx
w1fyjMS3tOV9Lth13HzStw==
`protect END_PROTECTED
