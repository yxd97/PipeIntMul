`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOaFATvG3jO3YwECLeLf9+6ms86n9eYlzcVmIbezHExj4F83hXaVgcyAICQG1bdt
czqGMPzahwV2A18uscPDfhDkNe7JXYy0QWOIdT2yHBAhE6qQbJFNhfOSEASl3cKs
9OREn8Mg5JSEXlidajS0qi879IMzjSXOTYBt3IuiDfggzs0xJqKzaYASu5YoFIAe
VjmVn82QPZ0kBjqKncxSQqdYZSjk03Relxe97+LSEARTeSBpjDIpmdSY3tHxfHTZ
FqlAY/V4vRWxgtfHCPUFgjWJIZ4Z/c03ZJSBam1l8uNQOmHWowQ25t0MhuJYx05u
pTXWodnNjPmQOziOweuwjA==
`protect END_PROTECTED
