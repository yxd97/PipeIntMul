`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XOKJYiHaC+HU9PijDVodxhFUeAVywLmve8TPfry3YP4vs8YOu+WL1TyxxGwYTQHn
4JJ0XZyvzFO5s5P7CTMDmbNE1A1lOTljHnBKQKqGbVc5i0wjK5jE8sxaj4UNXP+t
nBrdLqMo0clgLivnRCQViUOsQrc1uiHbdcw7JAa5DEyzzqyRA/wiBz//vGHdWNhU
nlxsqE/Yqjh8aG1eJihtorNhMMvIehW5fwmYEDMUP8ttGFiL6TiFw6XfCQOBFF6e
BwR1jiSSjtbelvEr+hRYBDL2Oh1zXjg9rukSaJ1sOqb4jNquazNgX+UDMRfI7HS1
VS6WwXsMurB2ar6nuT1ICq5poFayRQl8EHyWDwc+nBQ+Wjx1XuPS4BAH8VuOKhFG
AJ2fp4EPOzhEdgnRjfIf3ZYHQPIrURukuLL03qdQdic=
`protect END_PROTECTED
