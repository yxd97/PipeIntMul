`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nbom9V3cZ5EmYFU76j5UcrQb311+ipTzeoLKHW84OVLWEO09vNpDIDY4+FDM+Uii
+M+k5bNT5oMlDSlOvVmc08kyBTu9i8l9/YocPF6RB1z+H158d223Xp3YqhOCQNQ0
bq+PfaDa7z1cgu0eRaPUwx5afvd62NLSKbJHFBAHpfbnrOY7VIhkb5ESAWbGcA4x
bxCQB9J4iRUQSR+txbGxRXcVRTcEU714B5qVcqI8aztYZVLRSHDbot/aQbf7bZFW
Qc6TDMpy+NlzZ8QLrdOpGERdnT5tu7VDEEAagGas4ckiHzGPje4O/XNfaHaiSq3l
F1CT0M6/6sjNkU3xr4A7eJ+BzDM3nW/CybqMyiIdHlotnN69sDo6+OgUAfg3bK1Q
qeBNTgeuwDZ7uUeorTga3keH3Dzl9XztXLHjEQ+b5kJZ50b5WMZZtIBTrKsS/qcO
`protect END_PROTECTED
