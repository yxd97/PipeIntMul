`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+RNUTPg47nxfuZc5QV6GOvJ04fhW+gni1Ywr1viRdqp0q5rh4nVl/ZMsf4DKDfu
zdbkTm5MztcSOJxCjI1RFehxUgXodR+N5EyLxC2Dt1RHo56kan0MACKNaACaZ8kI
c9XjMgPpXv4N+FlNcBX8eL+wDRsVH13Aeu7V5Y8jmpWtaPBltUYTSoA0Ld+JaGrU
zfqvBf2wy6NS/rwHmEsDJvw4FILkElOcVlfSl5BLcGsIfrVQlZV4S8Ok4dDs238o
CPLKE9jnuNKkOhnLEuwUOz4ytE2R0INS4Q/8alFLnxaJ89zTkugFOvuB5GpbXEHo
ucYb53/xr7WlqaqLx+pVU1orlNpO4AzYFCZGaUpHSow=
`protect END_PROTECTED
