`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+xDLM2S1v6WHbD568ct6r6MrRtzOPJ0tp0NwnObahZqEgw0eZQ0VgjFSuk1E7EV
vZ4J9uta8MgTIdWrtHArWKp5lmdQiiCWKiDxG+Pi6W4kaViP397AOmeEJzYJd2v0
cV8cg9sAEVIHK084rUZkHBEvbaGBlYrZgwIrukfesnKeeTiS0LvH0S+sfrBuh7lU
MIdNrDOmfIqptLN705BICwSe+3LJvnfCu+t3ITPKP9o7E40JKpBFQxAjL1quhUIC
E5YXhXgLuSBBBs0s+vsEqefYpi6e8iLEJGmLMPKl/gYui8tVy/tTII/93bIF+KtD
sdgUgIH2CMA7zvWgaPubCtKzy746slUhrnjPcO7VF9XBW6LeuK8UxwPXEJM/91Hu
08lT+inrRSz8877sENcth85xOujfKNTcy5eVcIoKXH0=
`protect END_PROTECTED
