`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlT/MOR91ffOEYjvAkhsvgr4KJ9Bk2fbPZR1eTQB8VZaT3DWakFq0XLHdDlf44d9
IHlozAd2WR9KqaI2i7Tl8YLXoJjoBjnHbKmGXMx2wuO5F1hLpYLqhfmgPOnUUYtO
5cPq0KrxaQknblKPKGwncIoj5vhjRssVK36QaUZOkHUbSaQvgqjtYFNerjX9xxxt
wcVPuHlqy7Yd1yjsDoC3o6PDuXyablv2siEqx4nmn0RxRLMVC/7wpU8bnMZ1grD7
cCtJYT+mkB918y7PhTPcRMh7BGuhltI+WZhiZPtP6pUFAbRrEKK5vD/o+Y2xqn8C
yMdGTkYaQKTvxjUB0IsC4OtfMpdM6UsC58i0ArbAAIJcfbBVVPe8sZPstF8yBGou
UdgwoIZxutBKEmehqtOJ+Q==
`protect END_PROTECTED
