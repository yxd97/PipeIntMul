`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wc7FleDa6nZKSMquHtoHKKpye1ARv1uxuZ6b5hPyZH168dE9hmRxIaGfS2x5/hGU
ITsA2HLA+i99eINWCUFL0Iq1NLNcFl0ozvCwr2RctFREcxRGulXMajaBJodETX15
jEvpXwyTpimsaR5S0+iFZN1PNMDBL9RiVgfpcL6NE7xyEYE3SCd6TdNqTjdpcTal
Vo7sM2S6JNQXw+g9WRAr94m07TSP5UOKZ4DWRM9anl5Pq3FLMJ8R8XEfY9hW0vpy
KgBbyEUWA9BohBbSjMCrWolmZHuV8tRHmn+EJHK8gThSjDfBFARATdCgWlC3mgQ8
0I9v1/HEdu9fTJUe2XKC37phSwAn6543CmSvALzZQa1UEbOcK7A8xqBvum1fro02
PqHUs+cQUJE/33dh0mfO9efTuVZXHtSfkr1z6E+bseFDXNhCc72k083QiSVZRRN1
XI8F+rlsXlVr/q0Djr8jBlJQXghJczpWUtj81iKqrwmI/CyjcQLicRyTOpNuThj/
Hoi9zjoU86Q1pdyskdC01nZ7i4ZD7wqUeGAEQMAihC1aNjZ4HCGm7inwHTUJQCYp
8E0KgigrrR6XgQGB42C3FxHe0x9VX1qkniYwTzQPHHGCwWZC5ayIPFcG5Uc5z3j7
/th5HdFbrq1/FyesMeJj9r7PwMdR4lgxPt1IcA8194wg0PJYEKawfuyYvMRJXPlQ
0VINh9tpuV+XOIfYHXfkI7/509NSw03HQSoLVPe6pmDraXGfTzpWcsUZAxS6xBYG
Tsz4TUV9vGCD4u9M/d0CNMFoUB8J9cVkrxysRPGOI722GTAF9jYUx+FQP/FNHf6I
Vme0/D5WdBofIwTXXZ3X+8YMQPPw+3SHqgVhFb9bVzCWOtQYPObm7xE9T9llva2t
ypuzfL+8G9ce1jD2k8xRo3xk2KmGReMXb4LgAXgdgKSyPnvCHuucrHpxXP9RW7Oy
VXEHVY9Uw197jNRYj7OzLBpuPdJzCaQ+SxXNDxEgtTMNf+OG4Btw0ZJirPyUyTjE
c9eBhzu58M8n+rIxfjZhSJhmRldVqENwvGa/9EP9vQ2jDJkygQoCFkijmO5lcp5s
PhkQIV5FdihTDNx87Fbw81iMRUNMzGaPRZ1b2dfVx3lxugFBldYN113auTv2Iat9
16wJnxNO6ZgBq7Z049EoZdrg9IWiR9mKdrILVkeWfyvd/PFN27yr7Alf80l3hy1C
4nzcStkmuJRcoYeUkO26XgAdbyqzW5OQXHatvo/6vaqoaRJJWWzcnQQ6q9/+iwo3
`protect END_PROTECTED
