`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZmzWeTvwBccRPiJl6KSiuoQ0m0i/mGO/tiWjEt/JwH5dWnJG5xY49IjpuI2/uArP
LeZz9zeDlXxd/KD8574tVpQetCPqAHpFkmD/kE+GdBSeoHI3si9UgottUfijtho3
iborITtwCosRSlbNfqaLNQoIqgyNrXCcLof3a1vjyyoLslqudiyR+xpHFrrMeIL8
6L5pPiYuNSXn06Eref3gFNErOGv54x26kSuj6rKqNdXp+4oo1ti/0Be/SwgRO31M
v9INVQzm3HMdq/v7dhfOjXNYnkiGbT4lYrQqfG38qpR+sH87AV8/mueDrlFxBVi3
xnXyMo8Q3CTg63JEohUk7/8cj9Yatkuyupd1ze8GcZNqC89lz6zxzwpZMyoUTJj4
RiVXNik/vyBnvKku1lcXaP77LxZkrrmz1OJ5ciGwD1Du6KOvKVFTVPPzRlUrTlRC
lONZKMB2gXUWJJx6o9gsfb0N5GV3jIboReJI129LroPDaKDkLyX2oOl8cGhUB22F
LPc1sw/fyYDyMKVzq4KX8JT8qMOYgl31L6QC2FFjMIAQzMbo5yGu20k1Py5vyG+X
EzP2/xLKhfKTk/0HykPl2Nkb8+vTdQhRn1nQu36oWwy3s7lPv+7iyaP/GSX8kPXV
kjs2NwAUyA2fvMz1PJocHHyneBjSet5IqwUnuODK247TH6CPWvMIjjwewUoHmENS
f+jWekQpR+Yu9RDdMmcM6N3ponWZxoMlSGG9gzIYgf8BneGztzXOkvYTZ5ByCNQq
zLsUFdFRtSn6ZuxofGTmnr/rj7cWOUBUgdl789xFyfJp9wPh3yZi6FdMnHHH7wkZ
3ZUK7FLGqIREsc/w8oErAWiCLwVlP+T6pfxaJTksSqAGx4QV9EMbICbYt2IvhNac
ommjpd171XTYaTvlQMxlyCFiFA9WNobtUyy9VPhz18QyvWSdOz1/b3K2VKE6Gg96
wRuzIvd5p8hvMYgc6BZPDHR23gBtoBAwEIUZrgJsvYBCHiZJoldfyQ4JabsWZKZz
vAXKfigx1wLh5vbkWJGpfmQUXr1Yu5uRiQKEqmDoofIupfPh9+WJj/9Dz/mqLHm7
yDa1ZR6ajq8ZJRWfc42BA/05c74PcM3SEt62q8Qo82ikZ7XWXRzlw6gRcWxaBUFC
tY/M5hSO9H6tVB8BQDwUINgOf0ylpuzNhUvPgacyprGyh8+q21n9IzGf4EW0xvB0
wLQvgytf5k4wbyO94X3/AeR8Txfp51N8Cz87Ak2WoixEZMINzzUsl0XBB9j5Y1S3
Wf19ozSq8d3gfO+C2z4w1t0+uP6Cuvu/NGMGjtcvW0B/r5DAMimKcWb/+xQ+wvG9
y0RcZ6J50+9jOxbeL6IgOJi+UmnY6soIvSxOIXPyQ+TMKp42frwVlJA4eW1u4lre
zDVCUAZL1aSXoTa0zu8lp1RFPGt40+a2ZrLIftL65Y6qI2CfAhswnzLzNXuRbLaB
fViedTZM7L7rRwnoq99GLiBhdAsiLJD9CCw45M/Q8qcByxEE51DMOjDEnwSG9fli
uTdvx+/D57gIEjHbTKmWKzD6naBdky3nb+JhKW5AlcijtU30YfKiwfUdWh6pcBam
rDRBssM3JHOgydMwKBKhFpjj5vRVt4bWi6v43PLbtwdFOfUwTZYwrN8K+MA18Zkp
HaAfS+KA1uQWts9lu+5xN8SHgSyKMCHRD6BztaPz077jiSK14U8j3ejmlbkKYhgg
10P9Lys1vad/oajzQwFPUOcM19UJ4vhrf1HxtfTlqcHSq/aJpXKS7k/SIqZi5UVQ
iWRtfcMk0tdSZ7acHWqAFvgUyrwZL71GH1K2GY5pFdJaeXN7jZoO1/WYI/Z4a5OR
1sdRlVtACTzM4iJzLzVylR8jGDcbx2rhZKkJK67f2O/pxsCYqgleW/wKj4SpRR7O
gBOBVINRa5cR1phpNHzIF2hyZGA/dwXRMizvukIVmG0PcLjvivBpmFNHG1RtmBpc
`protect END_PROTECTED
