`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mRvwza6JLaIHKfO8Yy7MZxNo2TIC4NpZ5O1q4iwZvi51I0OcmGd1Hvg05MZRH1zs
sIzgJ4WG8zaJcs7hpXRNUkQM8tWk5DHmodPNqCwg3R+iN6OXr9SSGYM7KaO21Qjq
fEy1Fava5NCmQrT6bzFaqUXgDuulRs2vlDOVqQjo/EO+coDCfToPEhsCc25pR4z2
wGPyBOm3gupxfayYu3gRQ81GkDqxlBPSvx5uVxpe2sCqJqF3dZ/IhzyChwa+TVqW
3yoSPrXDXHtoVbapWhdw496SDZ7Y6ZvFKKvj4K8agqChEocRMNnwjeOr9G/ML6Jc
X7wYVWjb2OlDI8vOJTZFxzV1x1+vuXSQCA8Q8LQjAKsJ9Z/qlAdc5Q70Cll8O2rn
8LTrdiuYDvg1F6rbvF2KTxeCamRhi3IJWz7Loe2QtJS7ZUbyHw+u3epwaWMnDIir
mOx70wM6WfUT7RBsqSEqy0PDg480TH2w+wuQ401XJEa7DipvktceQlFZoQxMa5uo
ajG1YXAv0C/EMkpld2MQ+AYQCJAfQU3mTuH958rvNwaKxzFPElZUN3M/nE2TeNqB
EFSZQxrSoIEwq0+OigdIrwP0wMgelNVkQ7LbXkCUuMZDk3wMzv+NZZy1zjb6djub
5cLIIeHUNj2U87uXb+dTEbW5l8nmhHmUlw5yeWZkiw05ECdicjb0Vh9gG99MoIqb
tDX5x967NHvUX1/TfiH4c8IujJ4dImxZsTEbwKYA3RZPfIGl4uRMMe1lQbsG/01B
f5mo2F/HdFeroxuX/MqWzaQN75xeZ9hf4QjknnLjNhFmxBM0AjuKLkHwkXTFJzEJ
gmvmkSZ+2bf+AQU3SiV5XRYeep2TKDfTOawebe0r3lIl+MCxRLqKhgBB5Fvt0yiA
J6222c1YnNOJeI32+/urhZaR/OpvqmfBv6oMTnYbj9g6WGWFaFK3mZU81cgQpNg5
/5yWKq4pUZ7u3p/yCMQ2ArzCFGx8AeLg5tVKb6tNJ74LOE4zS0q1smFK4eM3qnwn
LW6eS3fxUudtsWD2pzw3a1Yo1XWDsb/ZR1Ig5b4VvHTq/TKqQTcklZy89CtUyF+D
Ev4IHZSiLIaEUd+dacopQYk+ajL1JblJJiBymaLVhEZU/ugt2UNc/2w32byn+dSV
Az3jUqIa0lt3g/0hkHL2AIqC7ISkEPLwk5H6Zw1PNXfJRVZH5mA/NcebqfDCtQ+k
MY0sMinkLHXNrImW0yVdM9ajHy8O7LC2W6clT1D7TnzY7OXgzQgNHB3AG9gYqXmK
j7iGgxouO5VaDAM7R5SysQnDmEAQtlrVhlXkI81YH91XuWYkJsiyNf632kEN/Fbj
l62vARke8/dpO3IT9N4lr5dDbJCvM2zAvHL6YNOlGFqa6urFfAzxsEDBZ/KZ4tEw
bIpm7M6cUIIZQj+ROnCy46bzLTUg0LzrtRpMVgJVLa6tDeDGDDRTB3KwRdsIgCoo
J1P4rNfl1q9a3VVQejiTBJ+ecoKIiepOupn4R4vxEyEeI4SeplIQK1ZsHmDqWhHH
6Mnp5YpiNl74hor7OeYLAFF6lFwhTN+ydwHeYRpgY96KVCefinrReESJHXaWH6Z3
GmLSPw17DrfzZ4acy/AfYzOrFNawfEj40lAuOfbRB0JN8C5iHABMixM+m2wY04a4
9X2Cdba3A9SiJ0iZhjQhUMO2X4YrZ59U5fxr5Ud80amUxpJg2lcZMwhXM9ndkSp1
koiNSMkhhbmTsMvcwDJ2i58lPI7bauTpGWelfG53+yXb1R9C3g86D673qe3kdz7e
ffRZXz1xaFVr9PbBeUNVuGH7Jlzg4RGkpSdqSf4E5I+ZUWWdkKRz1CSf2yhrH/U8
AGXMiDzq9ndLYQNPfPVpKbU3sz/H50rounqUa40vajQADXmScspvZqwTnUXw1GTU
eb5NHjmsuwTGLiMgdZ6FXxxZ+pSHP0o3mAwDNXnDBLYv6pmfWoZGje3srwBiCR/G
rsCGXWM8W6UnDe6edVAH5OtEVn9FoKnSxlJP6XQufR4zrFFI/zybjV4c13q5oJf3
4EvSbHBnyogkGejUSJgolp8P4gOpcT1KmRfm88ksjo/PBlyWpKmKzTFN3MncYZ9h
tH02ndKaHLaWw2z7aqxsa9IOUVIHIeSefxl0HPVa3fOlrNk2159dqx8t9SaAR3g0
XXOxQrMdngjUgqRNygdv6MBtw8gQARzHq3dF6I27jgRF3dvbMGb+j2MVuUQ8qyBn
JwhVNJv03SN83KuK6vmJP16r87Kka2SLdMms5clM7lEW5OdStmPc+U2XxPRJXzHa
B3ZW02bOjRYbslHTUB721HqRh2CjlDgHCXlbKUSQpyCMfHBojO1/p0S1tx1y4Emz
Ih2ZUb7w43+wxUl9Bnbcq8GCHf9hhp7NB+G3/wWpxQYX2Qsq1mLFKsd6gH47Gzs2
wIO01cbEob32ZI8N9yFC+KtqmE60fZ4wbYa4fU0p8qHzMqmKXZctmjoZgyGM5Gwr
4xR/cSxRB8XZUYDFAhmT7fONiXbL0wm5W0Jr7Xu61su2C94QZOaELXk/4ymjc8HB
pCrlEHaMb5DNyHEs9JS3SY5AhA3WilkcujmZjnOBIr7nV3dFx0nrrhdNRNmsYR6O
jqZd/ZI2doYyWoi8CCf5Z4ZszW9D/J/ihcD8MW6me0OFvs1vZj3/5m8uYWsS0YoJ
vIjyOWjkyC0JXk3/NdvnXp8WWiJ4D6GQwf67uq60tH6/I1cnyqhfhmEnXI3IRL9h
FCApdu1GYsXN1wQjP3cRk06P16KYwI7Yo7Bl9qUx0QKCx99271/01RJLLFlHCs1J
TwrVcCLZklUm+d/SWDzAGyb8wKQ6Mdbv5MAfFKYx+tDLbudtmaLpQZFMMKid0dtw
RYoy2ErgGRUR58RyBduiK8CWIMqmUuvo6WbkW8EmBHm3Hki1d3B2fa0FdoTMJBYQ
cgcLeM76TRqL+Csb0pXbxAkfQoug1DWbwTQ1s3mFEK07AGF3ZMVHWULXASpcLNf+
mFEnwl8FaBGWKl+Ojf+dHeWuXWSzOSvYlvihNMtyU1RqF3tU2PV0W5JE1wkyuGgl
DaEbOxI8hBVb4P0pezWe2HSfgGva6W2j+gowzdrguILCOv6oVvzLEdtdfDJ9agjl
3Av0uCvKRwDpqnSaZKTO5U15fnX/owu57GSoJQ9mCsxMjagOWgeFHAgw93qU/WYg
KckVgbker8XiVXY7hCSAcs546bap5nCpmDY99HysEZLr9z6xqzV3DwMFKamanngl
FnU6j8S9VVZzuvJGaO1jtD6uTb6f+j04oDN6eekis1vWwhnmeScvr+Fee8hvSnIy
PJie6/NCzWq6inykcrPkKyP8rQMvrBc3tUlm7tHJm/YKUIyuc+2kBiUk8spM8KZB
lX8Oe3h4jErmUZWp6+0xFVcjYwLGhaS/6MjIK3XjomF4hiYBTrrPLTeUrChQsdSu
6b8jlNpbP+wtjO7/5L/dJpXKGxTPeaGRAa21ROr6A4Yd4SOJcIjAe8n2CFMchdxn
6+fhvQrnkZ9JYLzaVs5gEYryv0AawQTtMgAO3AJ9Exw7hfnfJoXqiQevdpIddvn3
M+vSLwcmxPsEeeXTEh+zvs+49jEPPWue8ydmVrH4jX59ImYOjIOZOwsf0Am1qCA9
xFXHBhQYolFntogFdJw4fnRwkgzaQzbJqFVhpHvcfX/5JBO6AMBQvqG6U7RjByF8
tkZXdNnCgEYfp6HDApGXQ6WbDQNU5KJhjJd5HDu9qKydZiuR8E9yOkS8tcaDUo6P
TYIgX3DL0v/nQoQYYTTnRQ==
`protect END_PROTECTED
