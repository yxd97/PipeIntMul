`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mqGyaAx5XnABMuVe2lTdPudu2OTefwq2Fu9PM/dNkQo1SnzdRj1I0qL/+jrPDn1L
8okJQQxM9CvF3L2EJs/8ylcK4qsHUAQkxbhW+OmesbkU56Q8Lhb/66k4gragArpl
MzmWF1oIBSJGCO/Bo0HhOFjcrZ4c65TEGg3xcmEsUAyCB7+fG+zBDliglWDZAvmq
Z0m0hOPv3fBIDyCtEMJD+LY2Xv/eHBQT7fEvouia8Qg9rVW+DNq0hUYm92F97ySx
8S3D5gTxuEkok8c5mgZDeuMNvyU2CNQUJ72MI8qfZOGLJlVApJNrDr0NlIsu1IJv
hhknRmx4v6QnnPrga8e9QUHAV5piNtI1BLtyjR3Pdnt1l2MeqqEdQhzXOAP3WjEJ
8HE125UMnthQ8N32oBhHLcw5gRtZpqx4sIMIwyW0Llc2LOR7vo7kMRKCd2nWeE1n
8g7oe7cqinDb+EJe5Sx6W9gFxXatjfZO9eCGdbSjjFQ6Y/MPOLieQvHY2GrEuzeM
MVCh/797dcc5EcJBPXoUO7tlD23QfyD36gMjs4ED60IjD9rLpcl127GsHYhQxKHF
clFXTjJK+tr18RsSacxBlo0RZG4QouYjqtd9Bvgm1hiE7M3f6euPzRQ8XjMuV2m5
HzumSvVkIAT0Zm1zPCg04Q==
`protect END_PROTECTED
