`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qK/p3Tt2vmbQZbq56GmdEaCLHzohVxow1x/50xSBe+bzTst6eb0gNVm9vRCx4pr
+84q6IcftsTEsLeiGt5bqwgpxSHvChOWEsDk/OL4bFT2NkXcfOkTjcoxdY67tlPU
d6ZYLW6WqAxY4L89+ph3KXeVizALzkTNENKdM1yVK2aUMUhc9O1iDEQgoSm7EUyR
TtwTUS6FedAjCvRBAn/rQtk4pUtjP5gKhLKQL8PdpyuLO6yNdrSx6dgPOmBXWUJ9
pG91+weXwyGf5MYMJskuk5u9IkiKSAxyiKUXDFPhT38ge+4uzr9uNTUjIUHUXWHs
47tmEbDnvZMnXjssAmCz1XOiCzarl1Ga4F1tsoVOZnoXhRo+Fh27wYyCn2Bo9SPB
+vjhMrVNLjHAvGFzLLkccIOPS2deK3chhNr88vgOxw1hgDb8Y2gKv1SjMEvFp0kx
`protect END_PROTECTED
