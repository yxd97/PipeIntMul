`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGPDYEDJPBlaJx/08E2bb8znoH5xhsHHHH1ht2RvrJmpn6NGzrdfrJ+HxIU2VGit
Kvd2Iddl5HJao36ODMX0hYPbhuc7e7hIqy7nzOpf/e6k08MMX32jSnizgNgloXku
WD065egAmpnY6z2rLyMF1sCa9fcEAN8YyOFC0Llx3N/v4mtMNMyyClZ3bys0osky
Q8akL+Mfrlqrotpa86aCLLr7tc0lnaOwgSalAYS3/9DC3KVq1o674ISNCjP6njBJ
m/pybt6CxQ9Avbtvjn1P9KPbOHu68W5II/aupnzGurovok9zHgC3PDYbh+OehDqb
+fiBAP5bghkyaXRUl9Q5c2o7hBC/mTljWB6m4RuwKir1qJG+sY3iq+dhKVEaO9J2
54+oxVy++C0chU1BVEYR0PMrN4LX+mNJGLGO22mtOSwSm3y8UtqAFR+mebcWItqd
ZG7HVNuCFNz7/vxeDKjAZRbuC0F7q5uhAJlJPoOICha/eyIaIkmZSmuWQgNnA3Uf
`protect END_PROTECTED
