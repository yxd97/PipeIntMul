`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ja+0m+fuz3sKXl++cDwflGE/wD2Tg6Urp0E0LXj1fa+XfkYmpsLXit6zZ3eT5RTW
bthTtQIk8I1RxpBEw+h+65cvwuS5nWNONHWu1qmaQ0gMrQnKONIVW/IsWXpF7QEy
WD9s3T/wI25eBemhrMwgzlKXpkdGy7QvyJtEk/YIiu9OHIkKDLlB0dj7JrRtrWba
+XwRXi2+9AsenaSiEbcdT3xNa+UX+fG9DE931cTarZyC4uvNyZbHRU7M6E1kdY6J
qlGMcAKLRBWBEY1+rs9HSItt4w+9PbiwNzzYfpNenMFZKI8hITi3ECEPjFmuKNhZ
JfqWewEjEKSoxLshWTh689DWTZGFERpQJt7f7oyxnSm9NB0j+J/Y4qeE+uRSPw4V
e2e5wm/jGGHZf6zq2Kpgiq4bQym5SbsqYnJOykfAT2HUM1cqGuX0A2JvZ1UVzHPK
X8lcle4srOjEtfXSRm7y2q8H/r5YqbQ9gPBMJ50NmsnbYhnQB0176of4UAudrmCm
AWOBViic3lYav+M/48Fr+MbGL3lKR8NNYGEtOzyonwn+zsuV9MD5aicmGlEsYCoV
e6Zrl5a79ndjWCnLFrjYRafiMHEnf1faxzd1hHu362fMeVrjOcmLk5JUcEiHc25E
rWOivRpuBMnxYmzexd+KBfxNCTHAjaoA4ePAW/Vkb8zGCjA2z9M/lnu6oJzl/dul
coseW/FOQ+6JCNTGMOU8wQuhhe1qVW4UicbmgCfJG8FfxfK7Amz6oKimFC3W417L
NKnf3e90VHO0XT7AhVMBNBZU4dK8AOFgd8rAY+FnA8YhyDc6oxuUIh4wAyo8SHD1
ghqS3gcaTz6QAZUSNQ2uHRTYOzpSwQL79IxLT/l3K33/MJCKecNpediQ21c/ScMs
GCFE+CsSKFZDSoBpL17QBcJHpd0COQTemb6MaJI/cR6iHOd5eFYScDRpSJr+fKq3
dBkf8wGgy3G5jwzOThlkOdVVBWu5xn8mAFkzo2Y8zWSNCVPKv15CV5qb5U9/m5ao
jhV4TfSKOvOHVicb4tLpCpN0fhrQ4d+tkzksNJ6c+xGtZitSLpiaqgEUwih2PRdf
M3qsg5Ns1HMm3QByr4dZBusnJB2jKswWs1GYimvxR5/NXdlJoQe5kfPS4nVj4QeK
YfUAE0hzBIbfnfgt5tJVhW7ilxC39jGFRcvZjtwJ/Wj6p+0afAXzU9zPrWMFwS3C
YjYHOoKIs7IP8nn8fWPxyrpOOtZ/cl+0mNb9YTYuUjjjknH4OTo51TCFFvVWf0g7
AYFkp3uOBQYfAqqGq660Z4Q993fjKATKehBKVAQduKKyq5zAknx4AQRVbRQr4CdP
x1KY26Wc8FRrloMtqB0vH4UudIH9U6cMQ9lON5QwS6hMNNEmAcRkzQm9Tqszz1z7
C3vLQdaxAPd4d5PZyOsFktNu0oo5NrpFWncP5sILQGDlJ6tx9IIcLXyX+UzoN+so
5GEJM6H7v/GwEyNcZ+YokEoxspqE4oMrOaoYCE/Z2l94ITzb84uhUPnUvYhWW6Dc
5UoDNVku956Z8ZldPzUZeHQu1eL7Ai28MeefMjkWwNFQm9gQMnwiqwxJORZEuW3k
R45238nAE3XxasKW1i8xMku+eEhWrt39L/SaoHAZxGLKkBUtnhLc/+GD3bQ8d8RG
AdvmxQmHhTRwTMYgkSgcGaKnr9VbqR8/tj8kv8YdcmN6V0xOGaLpk9msr4in3lHd
A7ffmg2rj/6Ock7KgoJw4p72TH+fUU+5mZ9WMQQdsyMIcbkspzB2I6klWsbzePqx
z48e3Go1FGRZ7CvrZUcXTuoLIgvEDlrRC2T82+6ZvQ0JAdfiE/Uf0DIzJ39jGrBT
+y5YFax9s1XUJPbwfN3jp5gfMD+Zd5Z5cw95NSdW8Wm8O5Dewtm5Ssu2f4q8Bk/I
iRUI6qDmN6BhduUq1LlMMUianHVhavAFC51mBrNBujgbStxmbxOCFO8UIlgxqUaj
5XvYxtRq4d6+y8asqoC/SeYch41nlAUkhSi+7oKd98/7SgRXXgfI3E2PKDKwj3qk
J+zPLsK70WCqduU95eet/WO21NejgxIgBv7Ne83Rcten9NLbAV2uKUNcO3/g3CtU
gnfG8YrAoHtv8Nm3Fe0HIIepBEjKZ4fsW9QIjQo3vBflduXFLKutKOOl1Xa9an1P
YN3EfMWrGanDqda4swO69YD09J20SEtOJwQwf9z8al95kmggb/pMZhcCpfSxHfn0
f9M5IQuR+fRkxNt8IMmPAhjKA4MFYVJEG+lL9MeUETA=
`protect END_PROTECTED
