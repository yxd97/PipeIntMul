`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQ+L8jPUNLLnNzWEp4ep6NRfU2e/u9GtAgOmqTAlTUH1cuUbmJVWuk+sTcxRPRhQ
ooAOgy4nkbVLjrtaxVxr30lp3zy+xzXLF6AH+4cOwbxO82niWBKsLDHJJYF/PfM4
n1aeTcQ4P87RMMImEwpq3uh36B71x8CNoRgEahtdsP6IMC52RLgex3++sUz56EKa
KAj8q2wvAQ3Cz3I5z4HrsryI8QFLACBsqS6MiclO6rd8Mgyhk4yO829zXvg9/vDx
kDi0ie0XSISUK4IxQAfDqZuzMiJZ4yfQkNojYauKqNTRK8FLXe4Bu4XUB+a7Ecb4
395I8NDZGPwtkDebiKLn+OPILjWO8edYxpd1pj83HKkG3UwNuBClxtwV6V2/3DHH
cT3E2stPVSJjL7RJlre9D+89b4EzpMzqICXxu3z65FekJCZUn0eSwhCv7jjwhDbY
E/FVk5q+2XXR0mgxd6EPoibRENzOBxNP2ptzfoZ+SdRdnSI9M5gQHP+gMhpS5XbY
HtDiRHY06/E4K1rzzyRr/lwo2eNmgl46BiAaRPJOaEip77+gsvRinuy1LzOXzG6J
DDcb6IFPhE7uHwt+35S3H/QusJoZZmER/NLcirxrUK3yiDW6OqbGsdeKv3ABvnYD
inGLyOTYF7np8RNto8BcChBr8/995eW8I8SoMEx/Z9qUK0IFBOd5GEjXk65efMEn
`protect END_PROTECTED
