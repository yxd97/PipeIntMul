`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubS6p1QVwgXSnDeEtWSHd3OstJgvFAzxpc10sTuucH2rUMKlZjdYmgTuSMop/lQJ
dDRzOxpZtDcJ1RHJEoFFkzjMAnLps6W6jbm1iFTDqJOmKXDbE2epILRa8HSxXQpi
jctfpU60VnTP/4Pzw8ZBz17m1PEZhIBLtDKZHofuw6ktzvx119lkUgyftZ/IKogF
xBaYa3rnPSlraS2EUpwGRLskL5YlDCbZ/xLWPgUrWXEKt4pCWEqw4HpvLbfAuYiJ
wEjmBkaRh8UIJk2KEqs1IDB0Dygq10Fnwp+jxh9AGwT+vZx2rCLrhI1dgCQ8MCht
KAXLS0vXMGHbcuYYwxxSuOilvSZi/4HiFL5VcXAirKPZfK86EViHhIKU1orzq/X5
HZEDRxYhq0czuoAi4I1DzR981ukowJuaBxQKECcGi8exoDnrVwY4Z7XvL8zMTDg5
N6sgwi+n8XJrCmwoKCfvql922wGGAixm//MuP/WaJ5d3F6lruzt60PY3MqVQRpqu
6Ke4dlpFxsroyRwCNLZUwfjNz17wJL0qbnVGJUGHJUfZNPJZh7v6taIZz2Lt+SmD
6/2WLKcYdA6QeYQsAMwl6ko1j96VOvKAoXZ8EsRiUcPJy/MnRLQD1DxW+wCtOErM
s9gfdqgWpxXIoCmHwra5UJsilD/1hjUH9rtvAkV1FcUxj89lTTbPL7Xm39eUY5u1
7Hjp7bByEuGBZdk92PySz2H0sHiY/BDtpreHz4z8rIiArTQH2wR6jCjGmMXOBBS3
OjIaW512whtqB8cYxZg+BOM/IiTk2cHIEJB2QfuASTz+cgCXq06XCmDMPG8eviWU
L7d5L75ELgjaBKPGiZGuu7U9f2G/FAV1v7x4QoSrs4Zf7suFCozaCmMSEfX4BT1g
vk18m5Fj2Gf8IMSoIHtE9Bgc96gXvGJAxisFakfmJ//DjgYBPW/G0y90DTLHph7Z
VQSChwzOKlkSJaMVLUs2gZUSxVbgSD2hxayyIkS9jVico1A1kv+RjqcHC0b4cJM2
nSyTOWNM/t4pCD7kVelTVwcvt3xOTY8bl0iLdUMbcNXNfDB2CSRtaXWexSm6el5e
789ubnUI7JU7jguNFgV+afGgKojd/jdQKwJGYeH4RZN7z/BHBPiShYZGP6o7HQvK
NL2VSvPIC12uTyBL+sG2oVSQGzzNw+UhMRQyN7hrCIyKL91vrtFK4T9fgt8wXQKx
95ZJPOH2o+d7p5uK/20ILE0XxdMx/44+61pn1DDLZpzZQ8mwYREUa6XY0nzeoTwy
9X0lga5uiIUcJB5YN/nEExgA99zjWI2URItHiKeiL/ClTCQQaNtJcr2xpc245t9v
Zz1s2SzitGiYu/+MVlVaHtdX4FubijDDNKZUqS+l7MKFFY2zd73hMqXU0+eBunjy
HUaptg9Z6xCP+RaJTxbwlTrnAvTjRT+qe6WAo80JKWPrtZ313LFzcWM6aDy1iF4Z
P2RhclnKwm//cPXthPigHRjvwL9Ly0PluDjNZEYkE4xmr18xivKXDgceW3Spovfo
gwI1bfYKPAI0t7NAyHn3Ga/WYg52VE8Mq7st/VTCLxRcZk0loDaXT61C7TsfrEhf
4wlifvR0ZnhhAvcl0sAG+H7dTt+Qk18Z52yHKKu/KsBPRV5n8yow4rtg+ax+0IGH
OWNExRxauWxVI8aymbhQXq86YupH/tdKTDC4YJuHCoviHEfuHU5hAAgVhfF4HVol
ARtsI71jcE74Xdf6+bjSChm4HBKXgb8QO4RFd/NXtwLmGTdj23m3zBt2Ikeeg9HM
XeViRT888/xGXL8QZB+XPKPSBkniIPuSC6byaz4smGL5Tjofl709E30krFKEccQr
+I5Zbkq8ecKm8Sx2mYWSuFLX+HtIWyRv8DyZGNlUIZ3uTqreWdBEY1H7SnTbsuky
4oOP0s7a8/30FTapnxG70BE8lvq+/JztgD+X4dJjlwvX2Nk9JBfMiK080v5WKS9V
4bAOV8/8oMOaYVOVlGLjbYXLWbPPUMZRqLEjt9R1p12iJsbMwHq4vEDWVWCoAIWg
l+y+TD+E7up/9QZcIuHse1w+N9HecUNYQ4zIJ1TIr0jRYS44243MUuO4/i20Im0O
qIWWkOrQmfvY/9Z3CpiGF+m2MTchWnIQ6XLYD8rfDr8mlGIvCUeoQp/pcwM7SkYz
2aT2SsI5ex++n6NqFMsem4RngEeWIcEN1aowBN8+o++rfhty/c2eA6L5R6o0Ykej
4QvQ3Ua8vNKJ3tOae+WCJVkJlggEyE3WUhjXjHC77McyI5Jimpjyc5SY/0RTbYbh
xF/vkfs/+qVxi5aKIxuCpTHOQRS4lyTZo2QjN61XNa2rHiKwCm8Gwh4ejpSEDV30
RFIFvwqb1Nbwazrrd2tyYbgNa5DavNwglfI2feHKOB7ceVX5Zo3G/HeecslgLxc8
ONbN8ISb11Y3BEUORAEc53fKHK1xjR8sG+xKV4xojUMTeqs/Ard0IMy2Ff8stD8A
L5P8Y2GsD2haBiIaE4iMbONs4XoZB+3foyAefqyepWjmuKYrQmP4nIITekRNRZWZ
Oi0Sp3cifp6sfwxdu8qtspC1yIR1AVqhqBf+ag+Hw8c830T0y+6AHdjuZhz/LTYq
7D1ZEVZOUrxNqrgavPghXwuT76dMW0z429WkKOZ+ov2+pIS9xbHTQD0iPieTXJOd
0+TkzClzFsb9Ax9mMQ27RV3VcjokxbPEooMepmgo4QwZ6N7ug9dGotqQisqKuFlK
LE2l3ixEM/bYfClp6tVvv2upptJhQ0b8dqCYipT17buUnV4tpdwQggYP9eIE5e9i
9ErvfszlBRrBXngxMJ5Rg5zyPt7o91YB4au633r7f6OdX/dWgvBTAYAWaE4PXMbu
Y2lzw52nRfY4dkF9zhGDVzQmdQIcLTt7c/TWW/+FcegUat6XsC9AnAp3irjSeL4g
dWb1Oi+HTXQ/f46+rIsB0Q90lNNf3JU56A6cIRI/aCyvFoRfcKr8snlXG040FUbY
eRUlUEaiU6mewuLXjW0+tbmTo9U+0YIlJF1T6tafcOwNVI7jQUU/hTj6I3JTDK9v
/fijRyYxVAkGjyCjSrTjcTZDcX2M7cfXLfgTShMtqM1mEf/r15pToQo1HobPIl1Z
TK2W3ASvnctRiyGHSGDeyHgF0DZ/kqMb+Ge5wzZVIRGHZM88DlTp1SUxUjyryjPn
TWUoiKHOqKyUI+fxoYmtdLv4Sz65x0ymKFoV1gYJ7IJNumFBEzdrnwU97KNLW8bh
4e1KRVNmZmgRDm1RG5csgfUUxXJpj30fuAo/6d70eba9jpjS3UNSXR/iNLRf3y+v
wToGUh5OCaZw/u4B3nMTBCkpV6z8+/pg4bBUDHGB1gJERH4MWg17Xg0hXWP6EtPP
DP1iF7DXHjw4evRT/lEKQ+GjwlM/+ij8osYLFevi+G8fhZweZH7mR9IGHQcrd2k8
uSXI6bpPPQM8xmw+/t+bOsyfxVOIN5cg2QJcREJvZwTvZbEL+uTWRgj9OxQwc5jX
DqrHlbz2yDopZiK5JnYTwqXDtvQmGOiZ9/R9qc2a3C3PYBpjLOLF1SL/Xb0z7Mjj
abQfprg4TlWyG1GyQ2x8upCyEUtqEF+jVfNoH/cxY/7P6AswxFofiDltHj4ni1rx
D1mFTxr7YolKbqwjO3ueJXJXjoSqcbip2mdhikwVVZ7oxrX4T6yOdri/dpH+MvPQ
dAihRtrewwFmGPEDDYPpLgh9ReiQ0y4BP/0Wmkk8DfoFQ1KigJ6D5z767lTTEcl5
0GuTT0iX6GZwJS5mQbMs2wssZnWPHavznislT6bz8sYqiWknPSiMlI7isTgmlE4f
V4oIQ/aFGiimEbpgOb/MF3F97P/hw7JL+3+UKfZAC3K4ikkrALzio80vLl/Q211F
zfOQZz453kT0nNRhCAHRjlJvoeh3g8rix6WhULFjtoy8ygm7UONA828J3nHfLNQp
OngWJ6/oSxxcL7uvRvxrED0iRXK+uGJukWDO6wL0nsWCzhdySu7NaZ1/pw+BBfiB
s42Y5BhS3xIuUI1iJrMNYV1Sl4ERdSo5/VTPPlyRuyI2rJY18m+CCCYjVXFdHlGm
uHIczAm8l/sYNMdj8cvbxsOZy4+zC2nfr9HQKEB7YzbKZTKhPpJuX9Trh6LXu2AZ
uimYgfepdEmbuYd1mZqEz4Vc7YZvPdtVJQaZmEz02P/CgrDu08zqik2iz+dJV3Ml
qydYjOY3WIje2gj7ocVrRVLPgFy7XhRl8cpuOi0qXTliDB6TdXJxeYrxlYLdPoMF
uZ8rjsurvT2DHvHyZhO506dBmClf5pkCF5ZpxDxSPm1Qc1GSEPSO7+e+XICZU4aZ
CLZcPwzJM84pQ1QQ7So5XLLWfG1qzkuzrb0VCo3qApCqmziV4IvycQKgbzLf7sua
hGY9oLsPOMvYCd7/7uA2LTAGuj/AEtNJSk0NyRfosjCWXXmIj4nST6tZfe/BtNqS
C7GJhfVEu56DPsqIY/B9Xdt/qtRgdXBqWsP4znnXtjloLkNVjj4zg1nfZtAvYhEG
+VxBtlmO0WpFUHkGs7beFIwoOLlOMzKO3Dx8JC0IdPSsP9m0R+an63eXSC68aYdb
tPChbGdKMdD+XeqZE38rVxs94uZ/9laMCW3vVGy81IucXEW4RgM4kwgaN90UQP1y
z5s5mCQZWdGM6Ys9lV23tEj7dF6V7j76IlZdHBB9/woBLTVRQGrBILUGnXFaSFN2
bm3SyDAwHFdOnoY/QJk/JotD/UNgM52jgBf4Yqb3JTG8D8p97bYo64DX/70ljmuw
Sqlh4p3bJjiqvUtckcJ4omiC98AEH6yyYmKpupABlB9Wj4NGbK15msheNe4VyHDO
/G9LJ3BE0NCPf8hDEBU5fpcIjUpkcI1AljRUgGsr1qpEeTzaKr3l6e2yvSOAsLzp
uEvqSIz27SbkCMj+zZdUCABc0fOcNdXOfSuME6FORh5UDqWPZvbAAavY8Z/K2R2h
VzxPuwuAEUkxKrAYYlk0s37MhR40iH7trLv5DuM4nvacYbyfMV8KZQ7DB2sgySBG
`protect END_PROTECTED
