`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TosLkHcdz6wXUInlpiJmr2hFtJnEvycTI1e1aXRMsYMyDiCA4b9yQ2OLpVnULlhi
bfsTlcUcEHdjGSz+WoEPMUj2HMEqz+5Q67Z1Xk76fNT8uQL5yBrNHsrMIHcKbpUo
kn5xRAXwVWZFtNixseSSl/OgxwEf3VMqE5lRr0CFWh9JxZ1egBgqSTQUP/J+93FM
O8MwCXYGLGMCrjM1Sd2/6ao3Mim/rmKd4ZzTzR1IWkh4NEIXJLHHmgSXYIlfJ8t0
EpFx2F1CGzXrR6pW2RdmXSp+YKE/OjTLFUdk34ORrytnMo8SbCS5UORx72EFvZIE
m8BZM4obARKeCs6ys8GjC1TDVoBJXKBArzQHpo1xuV79C7p4rwmkVKIJHG1T1SYX
UlKrMEONsptxbY4+j+70DI0x0jxxG4dIEsk2USiG1uuz1pg8AAtSiIw4/995SgYj
GuFWr+FkI83BTirfvAbBXMno47d6VuzYjHwPQneHahdOMbmI9KbRjiBsVNkBapjK
ykahsCIvK8/cnV3t6sAZhGIBu+u6vCLpXYo6b1/E4xx211po2Jf7coH5U7xvIOLo
wkbldwA6PASP/t+Y/UB3gFzJtfohTlZKCM70VPOWbEXkzbJwgPYmWkLnafdwQe9S
a141ggEaX0TsSJO6xOcxMPxvpZL3b5owYZutWR20hbX04X0k7cL8ygHnoQRf+xT1
UvTLteDkWMV1/CMY3g9Ml0JxwfXtMSEIxCEMN2Rw1hkifzylBccKp7Go4RCilLlv
LXvF1J+7zQZkiWX/xeKbrHSEqTx1PAHF3REHoKra2owKoAw6Mvhnk+Upvob6rfKT
z2wUQWs/+cu60Lo1i/EQh0Hwhv2RlWfXS+5i8Q2op9Cq3F5F8wJQyYwKFZKUT0P8
yXxtLOJd6mqBaq74snG9xOY3EA1YLJZySxrqPMYc26dGB+DexkhQ37CMz+PEKuhY
2mlOvaaZDdXYu6u5W57h+K5ErX3Ch0IAvqf2MA1X0lHpg3XJAVU2APRQRTQdrI7W
rS3lagQ41OlkpKmkHRgglev7akzd8Hb+Zww1KPTkDZS6UoCwk2F/av4ap9DjYa8m
xxY5cCQ5eRdq6X12YMcHiwyQESO0aeXw22OjflfQb22lrZq9eLTkk8G7yCac95hb
rjyw//2IwP1vAgWH1juBbKX0cY5PeoXY6ihSCfwlSTP1bVlsMf/MMwzh3k/ge3Yn
euLRseL+VnVIB+kBaD/El0aLcLdx3J3M+w/dsaVS0GqETfpyJup1muelQfyM0bcu
qcFbt5jGqt4QlBhObswhPlYgvu7yXxzxZwDYACH/iC08o1gOMYRbrnIWWg2O5bDV
kbX5hu0gZV+/E2W+9bsM+ZVHRq9w5wxS1BU6PErAJnretzKfyYQ5YVmx3dk6Udwu
CCPi7ew1W4s7AnzLhCRsB69+em8hhdOICt6kqzm+IszAbF+i7txl8YmPyIB7W6rH
H6Lj9EgqhcFN6H2piq0KzKD9Wyleq2fKiBOMWqQXn6XjHtHCiT74FDQQE6BdyDE9
IoRvll52eK01zPzultrEYSorYJCrzrOJ566y9X8zoJSeCSrCB41csgyVVIpfqG36
WY6E863Di+VFPVGXEIUKWhZtcJEem/yPRlWnP5Rm6AYnhe8jqaxOWhppsklrPlwc
ZMDlu6v2tTEfTh7HAl84fLWp9pvk1VeqTbqRag8JHkFYTTA69sZHCwgqmymKaPS1
Jn4VibbJ5hI1Gc/YAGKYoqz0sorPbwWpOIPa5Uid3K8B7feBC3R0vmfJrd+5B1oC
0/jJ2q65LrqAmP46HhO+YYXUWVlv3jgOwt+MjUEELO6NKSpSFJOg5z2DHefkbVyG
hCBMyt/vLXGxTufkrPZYXOIWWcDncrejOkCs+yEnIfZn2R1vh/nQanccO0ZBLwe1
dwxJztVounT15vqvW6Q6pciy+p9Equm6J7b+HxOw8u9HBJ3qPL5bTCMEErF9l3cQ
ZRUmE6+5Z5SemA6QPNyrq/99i+z4DUyciAPVZ9vLkVSGrclsLwXhFh6m/N6BEBQg
gG9t0ctBw0ihQFqSFb45WVyshz8nVFpfg5olrnwE9Psiap6SYtgtLn+tX2kQUdlE
1AhycuPA745PMa2ynBCW6m+9N9icLshwkDB5JFkxq6i1vQ8B+fWgPPQcxf6137MH
U0gdcG1TAaw+jfQMlm4GMZbmL2bEfYey8NcpVnW+3u2HyUmp+/HM3Irl/4pV6O8G
/PQlP5IpK7bSQaHv7Is0Qim5SIRLzCCFKgMdgyHsXpL59mWrqa7ufANQ+2gwsTd3
wUx2hb9JIxQY4lgMEi5v8RL5kbmyYYga9PQBhJfJPm7ZL4q734uFS3TdXdVehj54
zGkExPPVVar0McuXmsamB4ll7LUIs+qAQmLPJPWPznDy8MEZp2QHH1hZ0ekzvLgT
rWz0U0Sr7qYQrLiKVdJ6QLDm5yDNhH3dhd1XhwtpDRfiWCYcTLl7FF6GQEfG3qje
ey9aU1D4Hia6INxVgrSqn5vnBNKnQMdpVq9Dl2s4gGmsS9wARXgeOUZD94IPnQ1z
GEDvwXC/c+QFppMPEV5/cYA2SbyxcHCjbKKCVtmloXYchHh19wAw1lM+hu+/kB7k
6QcQGogzm6IBmBEWaFus6it46WAf6EKAq6LTfT0GAO/pVJ/Tc9CmFaiMWcuu7X+K
vvER73VJpVSr57VB9hQrY63cYT1jLD70tNW9qLxCdmbk1EgUDQ/v/AZTvV9+NAh3
qYgo+yyKtwug1HlLVoSyndnenZNcECbggc9S5DT4UCjPfAOHjAFC3SD6PjyZo3oi
V/hxM7iwAp3y669aWxxyBBfBgQYJt1/2hbZBrL86CSXpFwpE8mVksuWt/r7FqWvR
lz+HzMX8SfEgJ2VDOpMpKhO/FsK/gYCrjLFAcXNkfHlH7P6E6inD04j7y/R8dIaN
tvkspANZzL9Fr+Vz2aEKdWF+pnu2Xsw3MiECG3pWgolwIOeSN5jbB5oziO91xLQU
iTppXfCGsdQc4/FavnyL+ZXyDPi0tkUlgVitxzH8scYIXdgHQiFQ/A1RTdl7ICl/
DP0i2MrcX1OqfqYvho6cLS3FBY/QbI4BGhrmPbA0vNnQMiBRBhHNeI71MaUS59YD
CIXnDmcuHwXrId18OdRT6VsogyKSk1PSMbgR6CRonnDuyIxzLaKMm+PxvVY6MFKJ
ey92NbfzMTdbQqsbwm40XoYCXMW2pEtqA9wzaAx8eLVUnPSVHTlvo5hJyUx25yMl
+1GDvsSuwH8G98Gcgzj5JYll/iDripRsaisC2WSNiw/3Kk3aqR4LGt62KGrvZ3Rg
cBEb1LHzWUopG53/gdEx4Gt919nQINEM2FNiZJi0DZCyvnK34ueEX/tZ+k4sfK6e
TXJ0QBKpD7kRF2ooi7CHZcu+V3ptVFAgthw9b9BL1ohbTUxp6LgQg77UeN0ZAKwb
pifcVmD5n0sJYl1diPCDYp+rjPQuJDK6vX4lpyUOW7YFd+agFxvGVh2LvuvY34Wb
76ZRdGbLnuZYDKkil6Na34jvPIf7XV++lGej260/4Rcfl9KpxOCvflIChDtzpjf/
8Nba3VcRvCASFdjwezn6gbcMU4AIUM2q/c0SKhRPrMcJpMqFElbQOfUjAhHQj726
WDQDOhOE4UWe0Vv3ih24l5kfKi/lbVY26pxv8iD3U8YWSeRCDRuWXS7M50Oup6eb
jn0xrbKhAepAwDQKMS6Xq2NssDrt8/9H9AmORR7A9oodAldOS0Mh/zHXNY8iK0Br
InhtT24KPVRZj4xeEWpBXtyumhLH4qUzIb9ZSw34um27eYhcRoVAkLaRpMgVjjqE
D6uvkXeJDHO/00V7A0+KZh6Vhmx0MfHlSmCY+fxYgxmBJONuU+dFjt5ys5iEoBrW
8j874eAx+GVFcw5cq50HmUCyIeeyCZslDw/DQKdzx6YNMTB7F9wxhvmhS4Nj0/YR
p0RkutGisr1HtlDOg3PJELd+0ThdgZOW3JYOM7NEQ0Vwq439w7pMTaxApB8oTNC7
oDKQYTvCQbIIMue2XkKcyzBwUAHxUMD8tdjJcnWatA9LWt69s+Z01/nvEWrka+P+
tf0Uem174UvFhIgoGLrcc6rL6FzX/F8Wuei2OREyazuLrr//ucjrQqQQlsmcE2Xc
RjY3Gd3JzrReEnnylM/sxJTM7A6vkA77dv99XqFGYhGOvTpSyacax0FXUtlFJI3k
gTwVkkSrDdpewqdzgjjmtPLPgImqqI9+V14bUE3wRbJpVtv6QHnt4V71bBqncTf3
HMQOWRJ6kxsH6V0vgQBuhZK2bqvNt/vKGSeC4GJ4sfzEiebGjX7fY553Norsm+qO
HjQw0j3vefKkpNE1h78dYt3t+guQm6kDUMASCeVjHEmZY2X0oW1trrcDXWyEYxP7
JRiBoS0coH/kWJNcpMG5e7R45FGpSQ750r1Q9yMYaZyHnbvl6aRb9poJkKxAPNi/
CHvXaLfhR18tKREWAnlYvbYNwsgCCDEZPJetIv/zaiYLR9t+3sxEhxzQFIh/IwZ9
2zlH5Edlf3VHf/QwTeTTwVOGEdzP6JDc/eUXvKRIahY9PPW4FZybgDokXdCo4Jhc
IJM1dWWtZ/DyrIyixJBqLF+HFgFEWW4mVorqKV8fQMzYVR04+HxPF66imUCAVkfH
7YwR01HSxoAzY+SFBTRhgfnKgFkEC+mEH1RsngTvnFfNqoBXhQQP8pRN/y7LgvJH
Mlx1uG262XmKkiykGEK6q3E21vp+9aPBf2ojB+5jqqnrb8v1qR0FWcWEqkkzpqbr
zz6q9rD2dcVrxPZZkepDskWsSVo21ZjRmhIO1T78M3IwfECo+LwG0gW+cSjgoMMs
QplTqIGVhTRKaP5oPAYi9HWF8Ke0U3Ar7ndDNKmLLwxfmD1OpJT6kTX9nqXnOkN9
AzeLIAjsMBpYG60eEuPnriIuPxTuIHbEQHIljMM02nIyZW59+0lq+D/Ybae7VLGv
Ev+DX6OV4zhqBBj4AINPdsCxGccn5aXDoBEmk80bMw7nMC+y4CFUYVHLhzjY3Mzt
nA8+sE9p82+yHO8aaNfaCBCCHC0a1w9C3I6BNj9mqetvotqWhOb4PJ0idNVfFglZ
adaWKxPVzcV9zUqwzbmoWHMPnIJq7cmtg34n69Gl8QD2yn0Zh8WvZGZ7Drkskhsf
zjIOt+LHNRo24Mw2CxN4kcFR6HnLLphGVWn1fycMACi9i1vcuyc79XRe8HiPuSoE
xjC/cpI+Vlfu0coWJs9Nv/bifAtaOOzImhZlZyj2y2bIuVGSUP+uL6YtYzWqZBG5
E759p26YIDdJsw2jI3c9Nriz7FWtD24vvhTiuYDR3Lxcz1tTWWSimwki7De2Bk82
9cBGZY88ERYBKRO0gvt+edbZghdjPdumZj9QEcn6unXRvmvZjgMpPxmOkjBz0Xi6
bFINj93szasqxd3IwkshGzkSxrM1/SZBv40ZQ8Ee7xOKfqsJM8suoir1q4lxbGem
AsSmPrS8UQUh5ORPm5mlJusN24z3AiECcP4ckIuAOHLIJvMiF4pcRxmD1DE3YLCd
o7OpbZBokaz0+gGStysyZ/W6tKz5Q/zaSf7Rov/4zN7lU8coWsHLu/NzYmm76F3i
/VWxaiusFU7blIjgexmHfE7q+j8xZd2QiWhBLSjMgimRnPknZ9azeEWWMJKucoPq
/Qsb+sh31L27GK59MO6FZAbzf6qGSRcdt9Q6y01mZuXjfD549RoxUUF52CwHTZQj
a4WDbdtFq2Wv6gsj7fTSMLMGbiCkCpvfyEskztY8+ooIYChQ/0ZMXgqJ4blCnW9e
1AXDRyackF56J1p/stXp1R4VPX3wDTp7yJ0A5FZhvxtZX1tP8yyG3hK1U0USywlf
qPOFQUcjIQQbCQWzwMP4lyuMWrmv5zY9jHus+6XEw8SYeME7vcqv9xjNEt7+92gl
GAib3x4N4HMTxd1Zl9V4L9WeR8qC9UHQ0Awdkdd9Ny9lZ+XKjhTmq0QuQaJjuBBB
k9G7Z/lvSc3F/BtW6wggD9MpJ93Mh4wmTlPmCH3RHCmRMEuozHxsurIfxnLw1968
llt480/om0McqJMU2HoyEb0FRtLTymUvn4YPYXE2rb268Q4o2/rs0HeAdqVWfLii
h1QavPicYH1yDCloshqj2fDedyfPoac5dgUlGoD977V3VK7oRtQ+4bBx/tmGTjQA
ZsC5Vo6lPu2K/3JFZhZgdUqogYjGqnvY6qeNlkX+pFxE9vQktxQAizWZlqC9BSIt
geDxPyW3eMnlwqetrg3cXf5cin7fGH5x69evy9s8GptmaGLlxX4+brHlVSLMn3V5
YwWOxKjBwbMjFlMQ2SFZT+EOlRXgHXCNZ4ISt16prNF5heh4Ha7KsGdqdPjbVwBf
8CV6praQdwpax5KUtWG9UdiwCvXdsXdRCPRK1OiBjDnnf61BHN2+R7NoxZuIXH7D
w7CL1hrJo3JXfv7JdrE+sdI/GzM5+mAELIoaYXs1MHi/+p+fNgBt1ZDzDtPUsWbx
VjOf2nkHqdMuBaNYj+LrAbt7qVnqOsNdENHtezisTFCm50yui6Z+NDDzbXMigPbS
YijPhvLjItWnzacsSF/9Oc7f3yHcBXzIKf3EnmH/CGYJ5MS2X3uBKx/Aklbo6bob
6ckF6Foaa2WhyALn9FB9ZQDJmhLfUVCDc6eRsL9zAo1vY/iIOC3fL1f54T1zmqBp
HJS61Vg5eU9oveku/jciXpfknVu2k7C4Vkp34obSgf15rK4aMUZ8g0SsIGfnE3xu
H/C1GLyL8q+iEAKIDkvVFu1aw1MGG4x+gkCiCTPVzPuK+Ga7fEyFzKPMFU72Ezez
i7F18A3cfjFepJUI/KaKP/1EBMN2o/4T5Wv1OuOJPXEviajEwZOoZkQ4L8DhwRFL
KBygTsjC2OHenNGD22lE2L3t3aZGvrEQZBetJAOc+hYvZk+EhzvOh/ncYRNQMCUl
E1GWQjIodU7t+Ld8Q/ZhTYQU2US77ZMDxH8XpsL0pbjYFwk8zIZLpjaqyPtjy0Dq
r9dU+SKB8tQlsqNQ1qhvWCcL0LvzwZnO8WDqhBkQVBmBaXuk/V7Krzuw60oe8Ug2
Gw4piJqHV1zDhctIq6hZb4jLOHcs3QD23OjFTpBIFRvnPvhNC+zSrgupQ7XuZQV7
72491EHWpJoMqLmxy3sTXTqP/soEjNmfZY0FMbIGP0GNc1te31N73N/OF3EQE0Bl
sGnUo/zhckW5BthJj1rC0NTo01I9M+eBx7Uq60I4quOrDh7sHN53oJuCUE3VaI/e
HjrGUVXC/8KsMtlA7w7blnGAVnenP9ap2bP/OpFFKPplhdJM4AXXvqDXEXtp0wdt
+/0BNbWHVRUvSmXwKX1lKEZcwBaF7/eiAQyLl4odr2rML3NlcRprst2FPBAG8iB1
yhpD0JzCqsilgeXwZmwimFwCHr4QhiTkbuyIoH1TnLLikIQBY8/wkJCqX1Yws0H7
Y7DILJa6z7liPrDiyZn/j5rr0hJ3Kw8A9QfDlQKI23rKA3svmdybElK+7xOsYMEn
hcUxwQZscpPBIdukyxxszvXejI8hsGK93cKGnFFCByv4+ekSgGrC3Xi8A4ejxOdY
b95zO35smi2wnwjRaxdfq5sLtWTv06tZ6c/sz35Yl9xYYc4BuBXsN6btRFd/MmNh
seviVLl6N4bngy5lksfjDS6Vv5ushvUuTTc/klUMK4UjWeaq++4mX/NMqnZ5Pcro
yq2Tx5bYJdQBG3MHy8uhXe6yTSQCZEiUQDmCGz7I4dNTyeks8ATaSnDaj7gQa1TE
WxPlPfoHqX2gSj77yGgqUXZGeqaIkCU4x/mSOPPcskmZ5JDDEftLEB8NJNRbNqLc
o1MVVXpJL5GXb8rmbxr+pP+PxArGAOPHyUIvYqmMUp/AOIifbrIONMq5ItNWBWrq
67bomxkOHSAKvC2Fi3YVx2FsajipeQpe3hXnViSl/LtELWXyj9dyAdRzBBmv5HbT
0rXDvVPXkg/fvdGJwzG+gYEDw2ZPmu2fgtxgRlI1l5J2FNyJqq5PT3JLu7/XrEyN
vuo03ABBLpYJDvf2sf4FcV/lzU0WCxLiHLoUr9eJR2fDDw0qEhSPJwzQwDrcDf/t
eab/Z+nYMRNKw/hs5R5FLepJ5h1y12jidvdxWQCIUDn/uBepB2bmDjqg3NgI2HhJ
1nD4iFVk+E42jYZV/L5eV2Wnq2mCVd05y1ksjGomcDaLegei26YCSUn1Ga54P8sY
nNXhjbEBV7DahIm+S237Tr7jU9juCpwH8aCP1IQ/FVjvBkgvnltrr4Azq1yD/55n
/q6tUq8MSRsabY0NSHnI5+/AHEdfPR0CfyT2SQOUnH2ZQnixNZY04jHCVFe1lmLU
tZ/MxN0bp8+ofUZmg3BUIpJjpifQxjB/zow1xgceJRtJk2a4lLy7613qo9duwhG3
gbAG2IKqtO4G0yPfl8NQKdKcrQaKa/We7yDojmbplPogFAqjWn6H9rhGlhOItRFo
5ZVuDtOL1WatnlcbA+MxKz4IjmXWEITC9QOcpiv2O5RahmXtxxZMtZjzmy9dDt8e
c057xdjgs5hMGyIjw5Y6BzIdHoB0mz7UQTcEwXH53PFRYkx5gDoowhjbMMOfnGYM
/o2JBMVGu3/E1B63HgypK8tDsDueRp8yaDe7FFKIRoIiSLDaWfE52oabpacu6t//
uMDKEbBhr13ugGbkmtJoH83Zow9+kXF93MpDc3+vKCfy2NBeyxzZH6XYnOM2+pe/
/91MmT+FWJlIyLQ1JGsSijLi6Vwg0REK+IQGNXOe1+kDKB2UyuHL7M67YCctjCyi
1fet5WKGM2nKI+N5hFTikIvXkkks4Chp/BNcNzrjxnaQe/9eZhLcr6sPI4EZkDAd
ssGuxDjT4kw0kGJWKhRQODt5HnLVQfJk24y5HCaK2aDCXFt5K0j/XwKB8xyINKBK
y8LTGkvECd3dXik5ik+TRhGaLQUUh0yj4wQVzp0CvBPJvwvhGnWEHIpnp1qK1Cpo
MmRIlXRNm372aE0r7S3t/PQgC8ebK6CgC1k5KTU8f5kf1sul3UnX00Frjs5Ve6Dt
yNXYNpBwIfTbUonA25liPIY/QJjhr2e779V9OIGNqqx7C7mQ5MfuvEo2Vo4/LeWj
PgDKmrNC6phNaO1N/M5jU+NSf/66E3yNSVfb26XxendUjJqTIY/DjO/a4J/nFayv
AQNigXinWJf667B74xkKdR6jZ7ZMZqQP9/bGRrgbGRz29UiucFHTjkAZMzOo0M2K
UiSNzAIL9J1BQiMbOq4swFtCiz1n/uU8Rvh1loWU4JPf16OS07tBiZlyiFDbLufx
CWx6pHkq5Qgc4msWPyu7N7XVowjW64SS6WNxW0bFdTXolwOEAU7k9ZUCGJY2zEtk
fSsv657qi15bQuknFrTpNPsHl8S0fDECzA2GWnT6O2OF2jhoA7CWMAH/CqyfBmFt
PveZd8RwpBDaCjshYpi0KyJ2TITG0mKrZM+rUUO+kb42vI/cY6R8N0qvXIw55MyA
5b5HB945bz66W3FEwS/ha8NDTzxOkNDMx/qnN74cB8ZMtbTBXJjKJ8ofJshPn8Ub
zWBt1fLysxxrv7jphDn8vHXLfhrPJZjF3cLAF6oZ4lY6JgHVJHZc9gxfXQj5pUEq
/+UEpu7ObUlZXOgaHs7Lp3ag6FuzpObaCEalH1pYK0uHTS/CldEYdnXOUMrlJTuS
EFD7sR/Cebe0iYMNSOqB7DnSnouCylOTjOfCzCR8I+wEnxaT02rx2/DtuzK45p7f
uKTCDzbKB76bLyCwGgn4ZT+v5ekBk1251U5A1Y3/LrW05y86JSBrJPAE2OwGFXDO
9P9CKmWUTsCQBErI5anH1VxeXuc04Pn58zCiKfHRtVdpnj0bMAztQVq/4ZB8a1ff
wE6XnGVAscMPQUJobpXY4Tpm5CnhGICaxuS8TQgDXw/oy5qJD8buzNYH9zj0b7By
Wd1DIuhxZwRQDZ2rKOYcshIVTJzyR9FwH4dWmHZ7lDwut9O+QMqHWw0FTOwHqvD4
Ct3K2Bs81UzIoikTlpfttEsjAG4O+mOMQawGL1vQY2OXtfFJnRgxqPhbSYCIfjax
9rVN5hO+4uiNCvY4bnn0RnAOs1WRue6NczOhqKzcKaSHxjO9qQMC/cW8VV2uLQxJ
JyKZEf0+kAN5OFRSTQNsao/Pii40zbSn4vOAhEqQ7TFSyAnFwvtRDcc0p58Of8UP
wJGr1wWCvLvx3e92adZGmyW+Wj2Rd3hV5vrvOZrdmOlKDV+ztiikT2rgOg8JVmf+
BysMCGC+NETaau/1PEsA6hPaP3MkMKdy4gHVfMOC66rbNViYO8y6o/wod9ju+n5e
yR1xRbr5aLBPkltGlNEbye1C8hn36sZ2dkiQLA5D84wG7COU98V2oJj344jU5NQl
pO6Jx6yqJjjbdIUc/7f8r2cRJQRYcKZzpoykmpghAEbLWSOSYprt7vfsGfPHP0qu
029az0sRGsnuFGTq6pB82M7J9Rh0A0Assauf/n0iXXqJs8am9H6QP7SdhE7lOKHp
fXDSMo8WDC2w/daKyDf6OH1W69N/lJuBTdBWkUxt0aEddR9tubtZ6DUsnCALvxb5
hVVsQW7lJgKWc2gL7N5gjKMSgTNgYlCopnaQxfZ5ExNSDvKhjJCqAm1IxY8qEVm/
AtCjio13aORkoagJToD7fn6gCcw9bx+DF9ha8DhHBJenJOAeVhpZsCYHRz5/tQlx
J83OZQkUzbOkSnu2jbyCYHHF5lDy9JkdiLq1kGEbXAewdEMzRpE3k4wR4TfdMAda
a/vZSJriWA1ZXxRcAEREusX6NPq4xN6xU3tOO+4jV0uA10bULt3KCg8poCcBf8jW
guDgW2K/2V0SrxI3sVFd9FWeRarajgJdVuI3bWp+ifBtosEJvBcK6AGWBwf4Mbj3
veXDbMI6M4rgJLKz8SXaHmVuRWxpIxMBKrL+HPop33vdGgLFzLyyyYcYAz9Nm26+
x0wD8EPCTe4L8QSShVoVzcXIKRLARUl/jABUbbc8dU9lew3IMLHQylKbShRIkOat
0LRKxUUm+PuCr8BgpZE40Sihh2YL0H06Ka3Sec6YKQIRA0cMsOnf2C4B8oivxVnt
i1Gp9ouXOncLouB7xK9q9/slblvnZ2JMe+CgQm60ZlgCwSeiubjdwCBcJjQYYu+d
J8kMoCZuyNvtYJsiwWs7u6Db2Y65ZkQml9G6YoNgnyUu49O7yoMaiqDh3ma9f+f4
Tiry0IBdUkvVDrTWFCraHVJJPwelqcY/RBgUaDIdAKDwzwwrqT4DbOiG8qW/Kgzc
yE7ET/j5u0rtz5CiimS0IlaNQroc+Y6Clvgc5QyISeU3SzE1lZDKIh1DENtJMaAq
/ueIqxWH6nkoG0AtHNvVldAPj5brIpBJtKAtMnUoYpUdbNSLgKoAY7t4ZqlMYYpz
eJ7kVpJtUv4s1IEIAzH/pQxx9XLhlFSaL+xciQb5LUXUzjrne6umqTwZS4qulWZy
0RQb9Y8pzdvZybYnYeGCXn6TXE5GLGPHqomHaCMamZkw5YzqUR1AGoYiy3gB1mR7
6lwTsCIGfScBEtWswtSut/zmk+Eadly+DydfEjQ/5PCux7Zp1Lt2f+FpURZfL+rY
siM+Dq4Uvp9mcWk6/7y/HSr/qz3qgsFNoZKuDeCnP5m+RJqNNPY5pBJWYKhLY4mR
w4jAibOrBY0uQqCN/PXYVGr2k2qa9yKkP77116x1snPSXopnBON7GuJSbkExG7N1
RGhFZYcluYDNy8mwXqydq16+hsN+/CTzqIjZvbH/NIy5gkgsAg85qTc8cYq5how4
Uk/W/GFsu/L42ATS7kX6meTmibkQhMDm8aWOS9gANV1XVegjtO1N0oH4IPuiURs5
hLdBKvtMu9e3WnAm0vPVpiJMuGoPkuEsMQ5iaYKWX8OipXDBVgLE26q8cEUCC8WJ
HzC5re/MxIxGHk52fUrBgEzho1h4J/pFlTi7J0Wu/7hpPTPjbP2ZckM/9XlcRGWU
XYEE0UMJS6v4KDKTsYr8EZdvuWX6Rb6/2xQiED5E4UQwhg9tUDKDYV2KK8vRjYob
AQKACfZJzXagzqTwsRs3kko/9Od5JpU35qdkbFFqb/RlnxAnPaj9x7J5ocWZPMQT
Yp0NluaaYCeyIyeq9EgAxy2+K+xlmPXpQYm59t85aGRgKViYDCcBION+OwtVJKfh
F6tPwfK+EUefu3YaI/9cmHk3Sd5mUCuSBXhQK8fhOsVGSa+8l3XE9LVSJnXaSE4Z
eyLBz/hc4OCV9lfq3XVdyr0HfAo0pVLtflKMt8dqbMyhvSt8TRp7ZDyTl+X5178z
UVlXkLbdh5iuXbXGH/CyqxC2hv9Icl2uAi/Ql+x8PDq69I7rWC666heErya9RAW6
Eclmvbd/i/BKUCspoe4T+DNxgeeoP9z3h+EO+IK4pYB81w/3OQVsHPfo4iFV59Qr
3Il02AJFASQ3qz+3FmSuEJisWueW9vBLELHDDLVHpK+2+9xDb3mZ5gDOo11PHPBu
03smTMWPI+OiKC9F8WMxq0+F0jq636LiUE5aR7JqDN+/BhYf6kh9vnYB4wxKy6vq
AJRZB/HTSvG/EtbOA50a+gwWDFPAmzvvbsJUMfFOb6dBRKdPkcxDX+vC/jbjd1o/
9gB2a3Jt+7tVOYQAz1ASNjZFcHf/PmAOQhe5iJDftPZO1c84OxAJEuaG+K6NEUDt
XQNIqWorcxbghRoMa3xy5sYBay4bmcvtJV8NUjZZW4za+uCOtU32NYFqh8+PDG7t
nLnEOrW5V+IrY4O97f/qQJ+OYUCfCzcUPHf0Oq141wpJPh9YEU/E+nYlvo/Xy6Fz
HHebwzDTJXNUnunuNuZjc9YfmWBITt4Pe9/64Vcw1fy6uX7EaAG7bvfv+3vf3kKg
99hmaV77vgsZpfESFzmQsueyEZB4PFePL8rWs9XrG/jWzaExl4Fws3q1XMHSP8Py
USNHkaTVTATekXf2IRXBweGUCVT+5X5lyOmJ3WxajhKthXrvPfC2FRPbV2uumOYw
Q0P9InZHZXuIT0aT+H+Wl2pb+zbmLeQqW2lWWRNruZTOjck7AkgsFzleb6OGMAiX
CS5etPU4GbFGb/hraezH9gDC1I+QzNjEx/Fju7e3B8h0sV35lysHI+lwoFozgstm
D1jgt4n8rc6DnEjq38z9Iyjz31oH8gdZUQCmBhh/wBk7GhSHo04RBT9f/5eDtPLY
XAJSQ3Lu2jzTI6GIA9QZmqMZoq8jwWXJVHq+pdNXtFCy8++tVKE0KttuUfLE+suo
UbltIzFSCDMoRgqkeAyO/Qf0iUKMuYWY6LodwdWnDcnhlFKyuRHGNhW2IU/Zj2L6
a1mwi5XATrKbJPZZ3d+kWVEHCE6BheQ7Gx5KGVRxXvIS/HZ8q/nx1DhUtkBk/UDp
rUO+6/9D9RqcWWpA3iM7LzSrfy78NXgccdUkk1PvLpzl55l0Vh5wNrmknoCPQ0B0
xfgDiwxiFowhjodY/IT54T/QQHB1KX6mzcJdLzgxhMau65jGBZN0LjqHrkOE0Fdh
r7BXXNP65XxHZ0qHgtgZ4Jh+XO3mTC47ht2kyptjl+5BA5383U38KVlp/uDgoW8n
lqzEt7c6d/jgyZYEzHt2Y40gSdvoRc8iIJGJkg9Q5ThkeTjwH2HrnCP2gr+IgXrf
KJ0Sab+ADUKOd5nBcQXFf0jMlUqiSn4MbGauDP95QLX8+OisNYdmVbx4DeWQhtnu
GVF3jQochRAkx+eLGw7u5tibsbHsC/7znm6xMqf4dPuJ8hRVbKfeVBqrsMwUep2X
ck2yFOBB4PmXlu7RFFsh+OnDITKUmwGrPBhr/Sjvy8iCIrxeuFIzr/rgYCN0SuQG
t+T4Acjv1vF6xuyb0/iVtv+EZ43AvGHYbTQxM9RIwEIySt8H/row/XCZWAwobHF1
1I81nYqZ1adRUDPbgoUF6YZ6PDiP2jqv6sRIgV87FU9ivE+JDkG00OHxoQaBspZM
C/dC4TauiJ8ufGHL2/YFNwHx4oQLADKA3huUaG0iUJs26ImVU5cra8MXOi6lfOXz
qcZUvi7ve/QIVxFG8YBctDfnJ9HlXf//M2afsL2PY1Us7fQyY709rq6c8PPj+RFt
+2KYoiM/vI0cCDTTfM9UVnxW/Spbtc90z+9ZyZzEorKFwDpQaS6FE5/h7881XUK5
Ia6CgLgGYgXBPOVaWSKbGOWO/B9DnAJrpzoW9zMkjRZ+kKgPq1EMztgR0apZ9XbT
60PGIoxsWqgKbFfLlUjuOIpYDabAZI/iyGIz2IPcFsmWwc2KdRFwDKXK7gcLr5fY
ZvssSpw5HQpB/kQZvvJmwwb114HL6Gey5FKIneUft+spfHKgoafBeWj7WI0qPk+3
yVHvkjiWpVmty8Kg3SpUJuhIJPPCj2Z7TVTAVL320UwR3VtZ3S0nwTMYxhfN30ea
BwpJ5MSiF/GXAeQvK9FFjk8mlO1TeyHnJlI2eGo91I5EFTM85Xd62uHAnXAoY4bo
CvZYTuUSzYbnBXuDTQLZASz1KxWfQKGi3zbY6ktSr8jCJtbkH+ihvUnl7nU629XW
7hRRvtFzgZ+z+8XY43lmjCS/6cHLR8myghM0cpn6/Afa9L34OqwGpjgwifiI7RIl
IED+1dC3RAGDblhWVW4uEEKapOOzUtAKIOcw3T3Vst4U8jsl2TaRIsz1/ITRNPXR
oVjJO/MQUlTX7tW4HwxCEZuRXySGI2lfK+s/rRcOuHsyF/kX9arkfLjDtzBlgM7L
RvdzYfp8E65Gm/Ryww+DVC+fG03PBTBMDWx4+chUalCr5Gxoj+Je8mZwJsZwiYbI
/OJweyuXD+2JivPp8tblQkmX3sViAgbOGBMotAh/M7RbCpGOpata8ZGb5no1r7iV
mViQNGl9yfL30QCbd4cTqbJYlToSMdgDpSyQRU95J+Eiw8TsgDaDvdvq+NxC7C8d
IBi6WbFupINMcheAxbS5iQzqQK1FNcQhlI12SZELBiX3fRFEli7p7bkxHql+EC23
eS0V8jx3l0tdrywxPSP6RBCcQ08ZSg5dHmIP3iIA1SxcJMclP86T+vPsN+8I5Gmx
QsJaRlePKgd+u5ZKMgVXjMF6Rp6PkmvR7Z737niGeHdtnJ8jXnlkBLySjMCJmDB2
aEPRIKSU09b3fBqQc+vYUHquvc3o6z9kaH7jTTJF35DTr8DAiFlYqAVnIXrHcpbl
DyN0fJKA1yIo/AsnLxtddbyMKkAVNL/i5FgDii9nk9CKtca+rOen/oTSW96QIE2O
QehCzDhp6m4rqwQqm3O8XAVqDyfxXlIMyGfeX4ljn8EzhrAlstLz2rhi+AR6nNMx
85f/HsbqJr/x7/7h9bXDwwlp9YlTT8m5hDt6ZUq3kz87fCWBt3j6o+gfV1eRupTA
pxg+ZaAIXTHk4XRdCMm+76oYxfGc+D/EjiVXduMyPdL65NP737OqaaOIGyRFXEqO
wzam+PQ92UyBcRr1ubyVqoSIYOxbGLtWzlIjBO8IFCYL3AB9DV8CQI0TfQ/w8FlH
rZaitq3RbN8MKeb+MxkTbr8xDNmxaQQ7gv9ytzWTYPa17ePuNYl8g3akRC7+EErz
j/DIYfDl2BYVmgw+2iKrQqlgcLL1DIfe0VOzvvm159g0c+OqP22FxZ6SAJ2CN59M
J4vhIWAPqIhT496YQa65iGE5y+nS7qXV2uwDAKUexXwrr4CVVkgMIwLLNa9jRoRm
hq5aWeChri0SeFUhqVZPn4WIruFqvaFljz0X+JmHc2F5iq3AFy8FkfQw02ht4okB
Wj7HjodfbwGWf2jsv8yBPKCRF5kptRae8Bc88W1k74GHCdALeTMvDELJe21iAfUK
5j70Bk3D67BKCbDQgxzTAfog+e/vpKtznYwAsI8F9skWwcionUDuCVvGk87/7y1a
K/bWdTdSbloLb55JbE8J6UWWEHbiR6EeZVsRtqC/djwxXF+JOlaeq73Njx86nixe
Kik/Lc62Kbj7hcbumfxc2DCK/a6pymRprTIOujV5+7osUTFD0LQyj+Qn/X4KAbyz
bktBDtE9qgA2qQNaNVm5kX0kWTZopi08FdGq2V1jViPqXgMsFEDl7XSz4sAciyMq
CHPWRl6ZDi7XmD5djc2elrS8gPOusN5cjqCmTsR2fZeN98thFLUtynGMmFADVvCS
nki1DfQZyrpeQQ/cMvPkcSEs2TGuKsGM6ngb+KpRfJPbCgoH4n8CStW0jEXyu2Bt
E+5ZrvUDNBH/2gyoKSiZPaYnSlcxo/dwHS5XOoFx8VSMhisiPI97lIFUe5M8Glru
Dv6SMeIQOeBJQDmBE2DwwQXdpOPjni+0zc3WaMJCZRkt4VQxaIVfiUdeZfkiMu6h
pEmHSc+U3/0U+JUf9byJWo+Q44zMgLoW77OGt6uRFybcDzvrkuGfbn4yUUUqQTCA
PYSeviFqZpK99DczR3SrQPTsR1MQrtrZfkcFL2cyUxPxTTc4Oq9lqhLY5wKKTagU
QbBXt1t3UrK4Qx9soXEsLUyUDL5F/zp+Vk4g2W4fpNrGAKvx8IfjdRochmmxCH2r
F5f/yZp/hOLlQGj7LFUBdZMlcdmP+Ec+YHf0OpeW0XN0DrsPMAInh7mHAvrmoMw3
WA5TsNjNmCbcZo5cOw7T7SG3x5rseOoTIAD2J0QE44Tc0thnQWQDF33CDmcx7hwZ
WcCQS1bGFJaa+OOYn1HEZqlekLThoTFZVILgvCAwtX1KQLCiEhHyecQkRlYGNs+P
Ijnfn0wY0fs1J85ObKYRioFQGMvagE4bRA0TC+nBWIMrJEM0+XWqmRWpv/w8DdaR
utktAZCiq90+F2u9svx1U0mSv0fMPmdtTA8/+3iNjunKfnL8IPdqg3q9ijkpJO9E
kGAUuE0OOIU2KB0hPrOjxetd7Yte8JX3WOA+dIf6SHfsMUKpJw2Dsf+mNqxfYAcr
G8SANmdx84rFueNMr0G+F+uunwINZrWSuK1BT4izpi4aFO2vfuIQf7t7PovoXC4Z
zktOL/qtM6PJzuQSSj6O2mqwB62ZEjh1m1kgy0gA1FczdwLJWlZP89SVq1tLDAHu
LuQkCXhlf0UH2PNe/j3zw2J1J3HHYSmAQKLA9ZyGfFhHefAdc+y2S55LVtJ0ZiPB
+WAN0xOo2OVEkwvUf305B4jpfIy7lpb7MQ+h9zz/ZwPgpvIJOoJ5CwNxQwawGgsP
FnQ36K5HCARln7AFpyBTuDylhUC++xgSb4OYbbUeMVXU30Tllq/c3+GD9jUkSs3U
o0F/MACvYU5nwiAM5olr29sCiMbRgDau/gPZCTpq3FSDkdI9cggbxFmnFCB+fqIB
8LKPqTSVng5HGVHOfOVHsXDK8YO1aT/I40SGMAoWKLCEPuztFshoX0PvYteHBgmN
OfTdzq2DSVtV+hnJyVxxDV7CX8TXxmfKpbdHpch5CjZ+/iGTM/ftBYT1fP2Qk2vX
+bRg59XswRN9QubTDSxf+Bdv2BmtckV/Klmf37n3vnnoi9FzbZVlAkYeb5LrUl1y
l6UqdMsXfOQyjUOJJofcKRUDPdg7C1USQ0ucsz0lszOUqxQCP19y8sGdWeJ3TJuS
d3c7xjEBBQ0wwFNdEe4UXyBdJMIblN/LPQIYlNCvzT/YJb3NMQ2sSF22xtcx8FGo
z4vuegSUKywEFtBAldHW8WJHeWnwrnkxMQjUv6tJ+agc4cCKi8IG1RV3zoWM9vtZ
U0zrXWQE+dtZtmXcwhNls+dSjR+yzXnIhYduRTNSqOfzEkTy2YGx+Jv3QS357K2T
dJIArHuKzFmjzpLkp2Y7LYQwTg6f0UQ5KDgcuKoX4VTybpy+HlIfM/hOOCvEeCVB
PdZsQHRzgEH8OrEI294hah3gwYlv7haMZz7mMUnwSJP8Ddmj+0z/nOTLbRusTMsw
ZzB69WwAbnfqxAlVHol0mVCx4S/RhzpBCEEQND4IOQyP2YQqcgeSfpPXmuahkdKA
lko7FGVuhk8zzSaBX2SRUMPpFvw53qLuwsW7ebSb2LnFBrPminWAHtX+u1jnPTSo
nMMOHIcveeFQLye0f15Mc2lda5KHi3fd54DiK99tpHHbwwS0NUWD9DyXgs4z5zRP
VtK9apjGWDy1n+VW3A8L6emG7NUKKndTN92l8v0EjLy0QwSEw2wKwkXQZ9TRSZsV
xL+z+Y3F/o+eUXAx8ev2QNcSSJ76PWHFOkkOlSgv+ck+OMYII0MkgQx/GZCQs5Ba
LR+DJ8zRXhxaUvcmuamQ7HyVNawSQVfe/F5wav3cYotPfYVeswK1mfuKXeTy7ZLv
0op5KjXYBHNj3DOcdrZrgpgGhSib6ofq/h2vhe2wFTx7PRuCOvqGL8Rp4mW4rPkt
GVR7hGHhDhF17eq1dtQ1EBM0NqC77DmMb6Pg4Czr+8tZcckHq16LtsnZKv4TQHT8
aVV1mWpo/EuJK8Vq5CnJe+rNaOUBB3WjbkwRdYh7rlP6ODN0xUgEK5JFJdX3m/SF
QcfTZhBjWhBxFBVgfcOLKBwl6HN2KJQAA25F0TfCXG852URrwv1NDaI8pS2yDV/L
47CBGwc82J+i0aBiFHfy6n5fJWemOGkC60/G8bql7qPh+aVyrDzsCmvl4rGDOINa
o327mzn7ZUqVRTSAh34feZjIR8Mtr3KgD4gSfHUCnoiRlVm/t+GqS6wli7H7lNb4
hGDdCcGks3b+DUm/ra36wSBz1AN1tEldcEoG7CNt197/+lKE4FcfpUqhcGskysp4
EbkMA33CdJqM9jAZX0D90MNFdegewdQhbXz8BuHkqb94L9om5ZR5e9MeVx6KpR7X
lma1hNPFM0Vij3eN41pv2m6FTT3hVyKa7vLrpbxaz7UJSVoT53QNCZxvJITN+MTX
Rj+3f7SrOQ+YI5ASMA1l1XvBhHg8YKs/NCw5BVag/YlcDTQ2XtijLh+UHaT5hryg
vJSp4SwDKVTLKBaXV5uNMI38qxmsInV0tmgOUEo/Txi0c694kyOt+Yjn1V7OiJoC
RNIwizDxdUueawkHnmROSVotQsPrw7b4Djwrd1PzKZvTZJk1z50ZMvKPSdcFQbD4
Gkk26LWefccR+I2luab0UCqoL10YvhLk6pFEI8iNFGnTv8wR3ux8MidTEm/BUOUd
u64h6Eq1DJB9SQxJ0WZf5UoyTwj2RrFmjxSudKdq+tikoco3ba7ui3zfd0w9FUl/
Zmi3wAxPkpD52Tflx6sTZOyEuEIkprndulbG5F3W50hMC88xEpE58WfK65qm8O6c
K7L5BONS6jcSU6OtQsm+6l2teW+aFrIoI8KJ5u4haB7iFrXp2ZuYQzowHSp3bQAe
tmA1sm+7EXAd3HQxKJBLOGlMjQZ0DiVqPpxNLy78JCJ+77GhWeYxIdDEZHSwFZiB
eO/rp3sjrOswz9TSEV+nbhC5ivKDtjnjaqyRBxqkXLCTZ6BkC7wbrJmOYYcR9ePM
uC6vKAFwV8Vq5bJh1tMCFYcFMtZrL/fEEAQ8TV8nLOnJvcgjQp8kau7vJ5aFqBcy
k8XIzTxCy7vVhmIjZ+eLZS1HQX/vGNleRjj+EY3vv/E92R7SzXqfCQsUebBq3Qaw
P4CciJUxk8uGMl2FasxUV8Cf/nsVuFljd7s4SnFVHKE0m/5fRMHP3ZJ4efapLgwQ
rIIxbh0Ceg7sHUEYve7qgAP8sluOiIQH+zi78LC1OV71ofBx8wIa5Fvv2ERTzNm5
GBAN9xHp1ERoKIVAnxX1scVDirJcOzWQ9tukShipnrdgoJ6hpDB0pyCZ3mAhyFb2
6QCSm5Gx405QCLmDLs/Y7zMJ+6nYlad1vmM5iJ46aIL2jTWJBFetgVlDVdN2r6It
lCAHsJyHQjJXnCPKv+NS2egRHhMgHc9tbNssTiOC70ED3iL15BZCq2WGcG57/f46
/DvmumS6TKV58muSJhEFWdDZBl7QLg6uPAmkBmcezrgrtTfoIN1SIrnd3rxgy357
Q1nGPDWEsIN8AdHinHygwNLjtlvUhJMhuCrigdCjoec2UsBZebw59ancr4Vky8DL
hH7AkJMWurExhP2hVApB4LMGieGJAdJHhtjXX41WLURdfFwmtza9P1q7+xWu3A2/
duqs9U/Li47rlQLWoLJF+XG2SvVnbeAkwhkyRxM0NkpmDr0ho8l1P8WxqwEsd5er
Zg7EaMcWZ8dD+pihomXT38zf5m18qyFPxHB2Tn+f394V1RsV/h8flEiphZJugF56
CxzgSBldlIIzjMVxrb6Nr8jNy2zCp44K1mFkZl7u3Gycx8algTKg7Y7pjFfdrB14
6R+caB6JNCn5/byoq9LnWo/u7XPRwJmshTdg0ESJNWo8LENTm/StpAudWt/qZJzW
2sCvLf3y5HER7yudmtbARuUph80Z27HmF8+gB5w5zgx9JPQo7pbVE6Wzs6bROSkD
Xwlj4jRri0cDUv6KRhqcdlMb5jFtng2B9NawjnRjj14pl+wEq9tHFrTfduWCXAeg
Rp+J0lbTE1xOynBeeAa8AInTh0Ld8c45t9zwG6bf+KDLT5P+BUw+EB27PitpjyjH
eEnM9MKaE572nOd00jliWSHagBbNTifmqPKuSIM0Flt1Y8zTfSqbTvrWUM8r40TW
qc2Omf51QTVBGgI4PMUd7u6IumPuMeE+W6S6wQlORAYmJxGobcOpeoiB78QLXmeA
I+iBG76IpDTtSAzv4l6TK+vPhCHIdOV8ywm6QutLxwQIWBainSrdhPKe6OYtkp3c
D605f1NZB36KkMjl9NmqiqccQIEFlDQkINpgN6nrAbZCAzi7hv8bAGpmJAXbfNoe
KC0dkLYiPSHzAo6s72d0j5EBIn2Wqd/vFSC05jBoZff/ZCGeWsSwq8zXnEmU2pbX
lMhmAVhAZ28tF2vW6Rah6Dk/nCFaf7wZm0TH7PK8oXVROVF9hFoW+aKGeW4tFW4D
9aRp9h2igj5n8u5s2ueQ4/idmZfET845BmsNHF0hzXshJ4k/82xkCQ8ItnwHuRUr
9dJruR7IKXyrlcMDLj1yiemqJB4S8NKk1ZMR7m9QPQ4YSO4ZuJcnNjhkFdFX2j+9
KCq5xpx8BUrS+r5i3YBN0O3SPvCFeKHVh1ZzMb5KjDmMiK6Ez7Vqc4OY5TVzYG7H
Uit4VVYHTlhG05tXRQ0XnVlJDTbjvO6/W5WeCgsQuHhi45Ik41eFFxGkWYzBXzSg
DMeMCUx5HZgR5js1C5lM477IKOzAOk00X3p/sSvp+XcIIU2YAJYgxxIMiYkyTjji
5BZmiyRL+76qhbSsmmK0hR6wcj06httwZh4NmNzuJwaVNZcMm+DagAyH1dXwTbAd
ExYdmgwOTpTJ1KslmpW2BoOC5XIc9ZlF4Cy+vFR7VzHIf+LMdwylk6NrV9PcjXty
9pc7XYFRN80NxgQ3ly+LEXK9IK/x/TZxiJZOVzuhuIYB7xYs6Gl8ssxdEt9MEb61
6cuRTOgTumTHNnnR7MAq6/TORqKp2ztDtHAvNuAy9byhqlc39PekHvvYrfi7Tehw
5/Dv2P2FvunlOMLXyJenelIFKJz7NYpWL/AIiCXkAVkKKImqQ7lOuYvLpddZqygK
4gT5+jq5oozbOcsb0CYdBMrSHFYJnXAPa9Uqkkh3i67mOJWuKN+qopcuasV7uYCo
QyCbXIxIKwtDGKaiOMWrMJO4b3/d+S68opcrqTspXDPwMPLE9xXW/DoK1hzsPkdZ
CL2kc1L2ON5zUSsBMwwlgkravnd1Odj2joD3MCnTchXBHZQGGVVAkvtT/cmfpenO
bhnT603ZFvaCCbPlK8LA9oVNtQsl1N40OE3AOy2K7g+uVs/kyZIPZygbxUnPhWTS
7V2eNGMJRlaQZSDi2w6FJwZc+NxVxo8Gns9TIZpfqM/UplrExWWk84E1qae5+yO5
osdTa1S3db5Usv7tXxrFaBznu4HbADbel5APlNxYET7e/+VSVBrDRETUqnYAHgYh
UuAKg6uIw0h/Ih68Oe1M0T0dXtTpXovnC7QspvRtJ37kECL+jKVSzgs1xEp5B1U2
0oQ8Rs1mu5lzTmXR7Xj/CfHsqFNB+wNa75Ptyf8Zr2irS8MEN7A7NGbY3iY7VKwG
sfyWrAnl1vpU6IbhUTqG/bZ/E+PsVRygYdu40g99WrDgoWhitwsOLfGeSmM1dgw2
snMOLh27ESvlXpNPRtTLMJfRMZAk4GXOR9dqQ4IIrYfXeKEg3LFtdant8E+Rve8J
qwjMTGYXwdY3fRMoAWWAkeLRF4qNLpJFpTwrV1zRHD3lviquTKO+XqgXkFbXSoVd
ZfbeXolVnVEpdKrtuIZUeesxV9GIGK8gtvWTBBofDVTpDJlz9/b9OTP33FjXjsQh
LZ+mQdrtRBBATi2nxMB6vYOJ4jM8s1i5fj1eer5MdwV60UvqWejkxM5k+gEtG10p
0fGmq0APabxl8NhA9qINuNzBN15qy/ELx7S++6RNEWYX1iIBBf+qAIkOF5zLKHKd
FqZyA+Ib47MFrFTzJ7TTUFhBHisQRsagW8cmeoH2RIuKoBOZA1tuyTc8wEELfAG/
HL3hONxIcZRpM9nT4YkoFRfnsP2k3RA+NdrTrHugOdv77gi1l6yNG9T5Y62+CStX
+ubMz/LSV81BEEECRPlQIY04p0guEAL3iw31SJXVrE9hB9D7tsuCXOBu+1CR4j6g
j4SmUZlTB2MFhJPMxcgQBvpdRDNE2gJpHlNjxHsYbckzk7QX6s8yCEgOtfKdUfEt
K4u8HVdbLwvVfKhtDae6WCndeA1n5V6Zhcwh56J9XUiJafLJK+b/AZCVcyziqONP
jlr1wQuBHjWkalgQz4huxTW6Z8DKZ7c/qI6u08aXlIB8Zyv9GLxuL0uNsGdqfSVx
1FHckfrLOMriCJEf/htTUg1hmneQywwM/2LpAkmy9JBbz1yCJ/esq21NQlxVFLkt
o8cUmtXOe4/5mwV8ZCBYHFStSHxeKgDRUEA9qVfWjPNRsNpd6COOMKcn1JiT8z/P
d9LFyREh1FxzZ7yaJqt4UscEJVV1EqtwrDDe+1GyRGMvehcJlV6yyWJ3XR81QcEB
VWhfKa5gc3xEVMny3KOdzntCvmNgT+mjvuuu8igwnpraD3B6IFO8NgxHjRfQUeGY
tDnbk7rNI+e4rxGEgENH1+4NL1wG5ZaC9JNsAXQaFtiOY26mDs2LP8C9pqRXJksQ
m0C/Nk6tflXp3JsRwc+wkjgboFBbqCgA7szImMN6DobX50HaUo2xbGeBNsd/ljtj
HP9vpzWkT2KHfaLtUD1t8WcR3yZmQT7EV2+hYuAMwjgdzHbtaE9oCj0P6U6tqnB5
ZB68tTFRy4Wg+Xn7ADoz0dqv75VgHn/cu1MdpSl8PcjHEw9/ogGs4oeQFDAN0HdC
kUp8sAl0v/wCH9lUfpEygFSAx6YzUojE86BxHRw6mvW1DK8XyP8b5IF4dHctUxDl
aL8vdyRk8M1JpoNPdZuvXOJIlIbOTIiB3w6UekZ4L/5rxarti2oXRdv5o5EyXjK7
ReYGe+3fumB1HH2QEkWpNxEt0ZdrC/qi9Dr0yvuSXC0IDLL/hBU8G2a5d1pvAzcT
/YWRwWPSJzaPk6EL1fHik0kOmsQQuGivSjcm2oKCaJaxUQ5c8xIR7yFzXZI4rSWz
4oP8j8fWSsYB3XkaPI9V0PwXlXQwdNfbMTB82KtcIoTYto5g/I3swG7ZWSv8Yqpe
f5NVjLkpNXi5IoMiccscSipanXgT8OnARInJ1f8OSuhQicoyjeENPqcSrEFQCSyl
K44iUCEDzu8fkqYnRC1ppcKRJUDtGsgtsRq6HCqdOxt93I2hRfkfWMCHn76lDhGc
9SnkrhM9ICpF8pD2/a2wcBkkxdawT2vjAchiYoE9l6APVIHNFCbddmwuvqkN1ueH
prCtrtdjWOotw9/p4+/F4PSUUW46cQw9O4Gzew6CCLeqhBinm8uGpnb74nHVONf/
fcWYAVmZkVpHwx3bmBUE6/auUtSw7y4aIQz856Z9QbLhyuyfhFQxjqD3qh+VZ6Q6
05Kqsji3ii+tnvR0Mf2comZT2Z0JWlfbvwVGbmInORpEUI8vNVuLb9pbqJtozenp
N/M9TFfcoYpPB6WtcNSKXA15s8whiP7i5n1mI9nmcMlc9fB1kHi8vnVtZWeF+X3h
nPtXI7D0FRkUMGsR0pXf0HxCC9knenXyw3XgzaiRyY610vRR8o9ZuJVvGg9k/CXY
S4OJr1d6YDgepd9HMUANYSHm/6PLlDIcdmD9P7tlr6yX5MG2zEXbiZpRl9eHL2VZ
K5MWEQUL4fuijQNn0rG1XMLx0GTsaauYSoLntYgPENIVgvEK6HV0huU6ErEqcdYM
/6XTEszxKOVe4fPlp2rFnlJN1Qq1PUuOsTAUapqNnvknFYBEaHOhQKww2BMqpeaq
SefEY2NFAXnXAg1gI7w6DH4QrV0BTsrLHv+uV7qzhJomfkBYp3LUuGSNfPrNzbiJ
KTVvMBaDnObL6mWKdTP5aiEYozii+wuWxk0Ss19BENx1pWX9a4OFufW+M2kGysQ3
69fCUD98PagIoNg+ViX7DX+SmEiMJiIbr4jAnmDhITIqBHc/JxA5jIMKER+Njh/G
NHFLmR4LOATGbewp7AetbqPbW/wPYZvqpDvWWYevo4AC+L1iap6tcYIp7pYq5wwh
/2QAL+2xBG6TahRdCFnY4rkYPkR+bbWrse/d03kYyYs6ovetRS1yZbKOp036fH7L
M8RyGTQUzxx6/WTMPveW683JBd8Z89VSZHF6WV7Xnh9cp9xC+/OZ7hN3KPXc4Or9
A2QliXOpmXSVPY/aL4xDf7GjJLVHC1ilA+5TaPSOoO5hF7NPd9NJBLtuk3XhN7mB
zb3G0khTUb+sdNgKjrDizO9XQuTEoZ9h1Vm7aXTEsnBGuUEzS/QCap9ZKPeUiFY4
KAPKmu5mHufP8XxeMHCLe39MkAUEbBjVm50lEZT34+9gPQIVwRbGjPuNa2MdXcl4
zNZV1Rw4IeEALOcTk7MS1HJzF7gl/vlHCFqSlC9XPJ5vULmVQw6ZeyaqFzWJE0dD
fIwqE4RPRehFInxvs75y9o17B6PpeJv+lrh/0V//Vyqcxi7PCQl43tEvgZUrS51o
xmBk0Z1XCUTGOGsYqKPdSw5Fvs/YyokHggHOjUZpJKDITZcdup7PD0bMA58OkXiS
HOo2SmNdiHzciv98W1fm36hvY1ro9l+AegJS37JADXiE/wmusbqd28+RDGjN2nXl
uQ1H6jq6CzUjfGoEWWRD/mI3FFYic6JRiHRk/76SSv93H6iS28MkrK2/VHnbzps+
wLd14Ku3QNuCo7nwsMIi6FenWv/Wy0dMVT/QEvmndpbSztsozrHjvFlPW7u1XRsT
oLApNTdlTlpwn3kFAkLPz6VOxWNhRXVRTQ/8W7y+STisWTkeOplIDNKoRXD/squw
Jeof6LNiWZ+3nG2dxulmP9VTJvhAOamSxLg//NcbobHeXAUP+03mvUzmoiU6BTqh
Q3daoiOA+hztkcOQb63HeA671B90FNlO32SFMNSVfru93YaecRytg1ZFIM5tqqJu
+rgSQPPP+y+XQSO6JFkzyVc36gIC4oW0xYixrb5LNfpgptJ5w3kzhO5+NeYQxMjA
wHs/XL1jFWeNroxqw3uMxgPr2zTUuWWc7C40yFyOoPJLa9MzxJ1HZC3uc+rT1v2n
WEO2AbSiwdhILZKuy+tbPPeRRapZYNTmk3/JoxxcCKIctNI+ILUnSHEdWD2rTc3W
ahkvFC3w8p4LentU5i4FM6JGfW7YT8dIIqqGMSFNGRb9FeO8bRWkkT3susc23sXZ
LZH5I7jGVIfiYhTr8kVeEVlsaXmzy4F+Q/13UD58xOjHxHevziKMhlIPbTpwWGMO
gCo6Mo+X2q4rLpqOI1Eju0z3+0wZLv8G16s6dmsKkMo7qM7YoJwHJP2W2By/ftgb
ELaly3pJY7ScSyJpq6JsnfrsT12wzYBapmP5XpQvgPVRwjopnBlC32j4hs0SEoWv
js06ak0Y8XJiovMS1VlW+B3SdgyrH4gIsaWvjjGvT7JZqV3ieyDjqPa+zDP477hE
bST6FItTGRVn4awWZtJHyD1NpTLHPJpnIV0w7wUv2d2VvGBxM34GDF8y1mJGgcnD
7Zsje3dEEzrIlszsIg3j8IKaIM2wcKS8K6Ed0lDNRSVLH+XgFuSbNuw8rmyqonx8
XpGKoM28f69uoEVPAHUVeU+gXNq60BTqEOFMOvxnKXc1jHSPetWzRedIKOtozg/6
p+rsmvGz53Yeg0b2q8bdicm5LbEpYvLRRbqfSR1f3ITM6/7VTn6I+jl59bnH8iU6
MdXw0ykt6FIG+ZeAAYbZaqrj9MyRfYA+i9Yx0YmxbHNeAvjLauruRELuGB31A6V4
6RdSsNua643BKGNXrY2xz2q37v9mUHdKFRFLHZMUPPyVVtuDsU0jhtwCDmmvzzRM
xP6ynCqxdaql2QhWqyiP/vWwqfWIibOn3Iq9WQ3sXnY9SuAvzc274YiBTM5zl+fQ
AWMn1TO5KH7Imz73UB3muy1yjKrThjLpxI2N89RdJQTbaYYuri7/no/sZhgimhJt
YZOUQZPOCjv800O+PTPdTdrsIvR4Me2iyQP9GLvWy5D0kREEIWXEO6BqQF/2JxNw
`protect END_PROTECTED
