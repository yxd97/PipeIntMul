`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LO547JEMpD+W6oGeOj0DeUEKBbL5eHydQkd10WcK+7BpgHU8vA8Sy8VPD6s5K3Py
wHR68ZoCf7O1XHR7dNjwVcQW+jMUiD1JHHijA2QWCFTs8vSrfv7RX1/vwJ2miRzh
tFhaV2RrUelNb9TE/Uwt2KIO7u6oEK5IjkUc322+oi6Ehcw7383OpNUabJp8/b+u
j7qVobjLFzjju4XSikwVLuUu0bLCe6kRCKDwV4CLY+HgJ2AP1VyOuo2CG/yCUalP
jOqY0GHjpCjtOTiecaS6P9lmfyv1TyMsFBDG0EDSxJ5A3G+ml3kAPNgMEB54wLTw
wG96fBEmlcqk90AMrwf3iK8d21P9rAMDXjiijCFSHk+h3t7gQ8uMbyRj7dns/N3l
BJeFXMdkIBhtn5hRUdI79U+M6yutjMApsydU6A9c/E4=
`protect END_PROTECTED
