`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+2DsdeaH/NFbco1sLPhe+YEhI0hd9ZeXM88RkEGs2dDSHjtsmaZaOq3cIpsX+dO
OkT/l62EMDQ2C3DWSEm3IBh2eiuyc6M/1cmOl2SUbrtAqfArbSwnxG3kTuCYJWAs
Ddw7d2uAK4aVfYHFl7doY7EOibgal/5peA8laB84XU49cjCEdC9lbkQSNf+TEdym
VncD0woKVb6b5JqQfW8+V2FMo7lDBpXYwNObGrm4FNK/D3MsGQQRJ3a8JdgKw21E
GYNvoZqKMmbKrL3Cjn6iNbAtEbp3f0QLrmQZ0iy6kPy4f9/Ldc0W80JPYnNpZbfi
KUMRy66covT3UwtYIIg1ki9rxVjxpPNljAj3a6i3GRXlFxVonkCaLyVosRUhsbG4
ceT38GzdlKKIHBNnEyOOMA==
`protect END_PROTECTED
