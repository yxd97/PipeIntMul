`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k0BnUd9jrlvHJAWQtxW6Cx8QGJBbnxEilNpc/UZvmkpEiePzEllB6XjnA1ngRdxT
HMMOK+AquNN7xC2Ujvm+lkX2Gbz7uZT5NkEKaYDUYI8sk1yM0Zuh0IGroH7PLKQK
WyvC8ctkoUiHPpvlnhEbBCYdptrlkH6oKMDgjidP/GJ9Nwrzix3eyMsgU80ednF7
1tn2XPOaHeihrcu0IOxkRs8D6yhe0+I8CrALGnnZuPbna3my3Y7w+cmqE3g0g/J8
67vEz8K0hzF8R7yXfJXO9uqScgsTBAgqrKlhbNwAwdvKDk0ekrpYcdzz9Y0nE4Vk
wBsiljRshS+Jd3O54PG4NFo4WMvNYAAflomroMpfq6v/09P//BuwZmUJN5YNylqY
BEdn68RC+INt3oSm3SE/SxLwrgVvHGtk3Q0nNIJAFI1fU89A5F7mclIX1VKgGjcw
ZGN14d09dEDh6leBO8LxwYDKGY9PK4/M1chMWKRuOapM9Pjhy96PS7TEp7Z6cnA/
SKsuERSghXq46cPwZA9jAViJnuKG8tHjOzO3J7tVwg5xxxrb3Gcr5B4UBySU3gmZ
kOLcBs9r1KKr1mEH1F4YWG23wQSRfOG0OctZUhlEpXvDBTQQ/Nvw6POK6AWqNOvu
YorlokO1xKOe1BdmhR1ca70Ia+Xl7i0Q2kjSyXqsvgQFtXw2Wh0cB8xnto9J/yyu
P7RQ7erVGD38gXjujvsL5Rav5ZmkwwhKl/FNQaXFG24Lrjq9YqtXcQLPadUKoHsi
s1ghVKSn5KPWXkY8VO2To0elnzIidSCUCEHO2Y2VIkF/IJDu2MK8G6lHIl0qggNi
Aneq2+U3mUmB47meEuTvVyJ0iATrkf1QkaC9C3EowAjS7h+O6YMdv7A5iO4zR7rX
LkVdu5lbKJlBxnU8KkQsySPqNphoRrtFmy7hF8Zny6TvBQzjenHlZmZ6JUAhys8z
1l5z9vbfTlIgE6QIA6O2diPZczpe3L+f9AOeUqtgRq7YeXKtSPjGc35AROuXIm4l
SFCQdIS7W7xFrItiRCAU7k4iPFhiK4ip9mDHbWbBro7U9P9EZ3l/4QnsHokMY+jy
c25rIhr59Baw04REPj66q34sNJrBs2LrCRnxNN8tOIuxpFah4lkcvD2FoSmwx+ik
tM+tUgbrgNNjLjvCInU1RfZvkpj64ss0s6JEdtlmOCZqpMS6qCw67+vE8yi1dQSy
p2dCT+W/AIDv21/H66XIkDI/i5Je7Dt9MVhxbwPM4kGnNxd476xUUIVuCJOlQ5lb
`protect END_PROTECTED
