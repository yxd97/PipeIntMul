`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWBexe8RHlpalZ4tKO2DkSyM4FVWAK2OU/wYaf8jDvT6WzqSi1xAzRLPH05Kv4Jy
/KaSBqVowPZWyY6lAeZQHMwypM8+/tP8nia09vJqmCxVQ5MEnqF+ysVF+D9XjwnO
0n25nHQUwh3eX8qOFbah7mJgVf2D/CEEFG1G4KEt1hIICD1JLPytowkCEci5ZAEb
vzrGpxhArPpCXZo8/xYvzPGdvVCeZSVReES21Cge4/xrZ5W51snd8y5It0nOWA0S
UV0sXckVb2NIELS7CPVyZ2u9yFeumJSumDiVXP2rwu/j+UMNnYo+WtKBPSFfLFCK
joOQI7j3akv5c0KMVOMYqAqNVOcQMsIyELFus+haDvWNGpHejGd2oB2Iy1X1vzeC
PxhR3Z55t94aUOLSKlbbegbB154zIJxyG85aa6LbLddB9t3+KYZMDQAU2yTPfgZW
8xH7LR1hRv5bz+m0/RMHKOeGsFbkPD+wUGeGzucTDygIuFcXxdWSUq1uJn40VWnG
FN7xK3aeIZfFckX8i6O3CUncsBXt1IKNo0PphikFY2ZLX3nDygZuS7Lp4tRCdzHJ
Vyh69Y1G3heeuj4DQR+ThGruGFHoTZZrpXAF8ZXQBaw4GWc//mWzDAGDotndDQ+O
2U/atGoBGJZ+ZsCwOBbpMxVSeJ6q0lNErjblPPp/jdOfLQ6Itug79p01awu39H+6
lnCQw4N9u/ydzAlP1TglkALNRYPa8fuA7u2cv5ZTMjRHqUmBQHJV/DdeixgGW85t
SYZBmNbs+VPkXQ0cqpp9XyIShuptuqX/9Zj5DdShs7k=
`protect END_PROTECTED
