`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RKxyEs9qy1mc4YBTy7cufzReDewOOEbBTwK31/ONwJr3yqeWqn9YjANW8Z38PhXt
+UpfHW7UyxBxoyiwT+VjKfq4aU9L0IZAOXT1DxjzeJwmin2ZTKELRI1Q5St0yq+E
l6iWX0GGs5YuYXH+3p7e51Jt3qLUNU/9RU4KxMsyEhF1DctU19YBFCjLLqoCl5mq
9x31SAO8+tyY1TDLhkf4MjOZX4MoqXecHwhq+teND6UKtiOPxBvyVUJg9SWRC/m7
tqXf/tDGtdTgq6rLgkifGRHLAfFlnxWoIkb6gYWLG5E4GfMhRLEm90hF+c3sd0Wy
x6niUAfLdymgjwKfFnUpTbcbY9au1I/vgqwmEIA6ir9ZZzti8sDF8v5efCyH+5Dl
YiChLWu17Gi8BME1ZynIEmJQcnOvUMq7Duz0Y5NoEoL5QAyNCvh6ltx3wbYcRbGJ
eQDIJ3ed0eiRQhAPKMfKWg==
`protect END_PROTECTED
