`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DyTkq/Q0i87EddJ0mTIk/AVf6I1j0F4OFSbpiZDvhaAUAUBCfr77i0cMLcMFQmha
tXTZiG0Mmx9KyG03s9kCknfN+AX148Ln4vDUpm556zhzqqUKhsCfp76p9ui8mQEG
kyl0DWvtQ7lGVpinjjohAsxpkN4YbXCrkIB/8ofjQASzZrs+EZq6pYniqROEotCs
ZVRE3VLwVLkfnbGdAA9MTw==
`protect END_PROTECTED
