`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3Uusrm4mPZVJziXAOhnkT5kcgGQVJw55nJI/6P75E/WWQzk3bnSCcPc/+4iAJ/C
QLpUQ03yH2UGkKUAIkZfJK1eokTNAe5ATEAvLHBwp3lXmjWIRhz0yIw/6+MQL6AY
coCjzTjdmryP4mInTdCIHeoi6o7HBEH7iNkMpkRdgiYeFRXnfhfeZl5ELkT3LoC6
r5FuP4yZE4m8YVq9V9b9f/Cn1fv43dldse9lvNgT0NKLbbnZPngN1KyOAC02qNhx
Cpw6+Rs079IzrVTK08QpBClI3XcuR29CxyE9jPuXsY5QfQg0h4f1HFpgbqccQLHd
r5BoXnlqMeoYRPspFkQlhUEDjtyqd9JO5Yl8MfBllTA0F/Z6uTRUlMlAZyYociOf
UmhnGjZk1kc2tO+PMMw0svpveq5dOQSb/OxConhcuAMUKNQv8UGZLurR057mQsN5
QZuY3t7wyHO86c+oQw5hShs23OJWD5ntyOE5o4QQ2FJwbpkV4ZIrsJNvK85ZZfkV
gT/WpzpdxtElRBbpYKnC4FHKBHtrZLyOCKNFmUBEWccqa7hPfh0aQ/XHIIPBlw5Y
wyQ0bDtMAmpuNHmSJFaQ4zZpFvAhCHiyZHOslFQmgwROTpmY73rGfa9n9J+IYHl0
bcm0NpvN7vUgTO1NmEYt+bU88b2+y9aiGyJD5RcyCOieA7Iq172Yto1rTuilQdNA
4pgbWZd3IWLush1qLzf55DNX1xHAfyRzmePAsne2RybOjsWyXrGr2EMXMx/wrY8l
4IZky+Ep3wyATOk4+cHWQTcmZIZGDPGOr/sBUSD8DMa+zk/gex+S/7feQtEVULFX
NZ8gkwdIekW2MwcM+Q6urHL6dZ8sdLt/yTIjV6xTr0E9eclzt03EVRSFwfzfyGLS
BjBVc1BXH8LsE3rpanaTZNPlb19EA51CbQOuN9Cq3iImu2zEDR0k4LlPpI1UAafe
UF1AE1ypeR3UzRoGOvPl/vh3eBbvzDtDeWa5rL2iRgA/z6YzB0TFWlXlA9eHq7cK
oSbSBELQ9fhBpk74edwH1sw4pXLZx8eFouv4ksvYLhOZo2t16UF/PK8L0PH1wnjz
8yosyiNdf7hy9Fpmr8Lc2ZZ24StEqUXPVFYyYqOkMtG4xGX3SP/pF/QdqLFVKYaG
ToisAVJbSnUKeQjIIQVwjNsMNStCzA6uxlywQHEvUxlOhqLr4KbzpMRSXseSYv7a
WE0m6c9nhODmORAHhRIZczRuwykhoDwW7uz9+Xt5vY1tU371WazSezDpjIXxdzU1
BJZfI8zqTrCtt199xB7kceCqQjLtcXhoueEi+8b6Cq55eWYoRpKUKqBUA5Qeldjt
KctYFUXCMArkAONbedZllYRlzw59Y091++e9D4cW7cAYqBR8P/nOvieCI5H/j5b1
uPhzpKAkc7BGlUB91wIBl7kmTtSad2qEIZTHszdjX0/iTOMQ5RRsDWMGl5Tmuf9+
eo4Ax/nmZGKLtcN2bN5LBPPQ7iCzCE8frqzTCO4LmPw9MD8EVnzM3y4NUe58S/ei
RNkPbtPg57pgstVsdFcpxlcqaoE8lBd+rNGj/MhaFBuiZHOpqdT99MU+UosaGj0T
w0nfLWXF5zsjCcEPLmeGBhRIo3MSVCXdGFj2gupP1Pv4uQKLOilbhzZe4uF4PT33
ylGB1cKVYXb0iDNpZyIKs+B74aA+fNJkhKj2UIm2eUjT5P+bskW+MfRCGzLb8Jzb
/tbHHxxlVxGmlCEA+6YKaRWC823M+eWfvVVAglzp0t6j9XpuEQfX9CMt8acxxRPG
s2AtZbReykp6nTwfX8fsuATZn02yOxhGxEAVOOVMo/7SXNFBevhW9IXex0dV4110
fFndYCjeqHUEmiFNvA5yzzhoy9BMag7l9iNRIuYvjz8teMc9/E6MK60D0KymVJNO
8E4wHp5AtRZlvmYYcBx5YSehjcAzFmuUvU1xdO+5EJFHUILLJxZhmF4sOWF6W0cd
mb+cc3tHfhil7xPDSDyol9hSavexTcuDJ2k08K1t3dOft8EIdJA+azpWAY5082jl
y9b6UJTKyJhsY4oDgxyqR0TW1Nw8hsMl0+RKTDhuiwMRin39kAlM5cF8zsgEleZn
VDS20os0+yMCHfOxRkWhoBZV/T0iDCyOnQf+EmPQxNAwdvt8p31Lczzi1xOSXvDV
6iqz6+IjoRwc6Vy742anNzReW5IlRaatzCVJ2kRQyUK0wSm7mVXrCU1PJhSydfIw
EkFs4fmTG8oRy5dSBGbQJkCMOwIY1EUdzk+8alJqKEWdK9sH/FUTl5sXGLZAEV5O
Vrtb+Z5+A+ZKRv0QNxQmHvJPQg4TNE3zFWE9IP6pQV+QDhkMPGvsPg61J7EVjiNl
5j8V70Vksghrg9c69Wdb2D8ycbtBIQLUOWRY+as+PICYvRrzQbgccprKzXqOSD2z
9Eivb++U9yViVjF4edb78TIwSO+yeluwncikjwUEKp85pGl/gFPW21HqoxvDviGd
P4+pfMCSSu/pvwpkUQqAHWXAeSUFBKb23Hq3c/2mDdC4U2iYIij/t/KBA5AW5Yzn
3XrJNrIv81DcoEsSHHp7CVjQ61Mf1Yg79Jyts818tPG3rq7a9oiiGeni1eIkMDsP
sL3yrUIIKTOcFlMnxLvJn3lIXZvXBqNBQuAWHJeYy0Xep9sthjFKenJ+M3TLCFkC
g2ANpijA8iTqC5NWYlxkbAlgnGWhaRP0ktpChZA6gwypR4nHoHiyYUMAcwJRG6Vf
C/2AaYQO3Iyr+HfrnlnCAwzmu/oJnK+l1+6Vf9S3Dcczk1oCHb4z4glJeFeOhju1
9uehGADIAEu7Ft3Ro/v8Fv8LMrsQ7nx4I5Og02mmL6ikQ+1r73I4FnyMrpkNFzxW
0JDZkcPB+KtsY2FSTu93wIfoZoUvXG0GkHZJfhzV6frCsuXmii2nwocxY+2bz3/S
XTm7NtXFd/SfLzYT1IGpfT0Y6NWq4JtCXDygbL+xAJE=
`protect END_PROTECTED
