`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c80T+ir5Dy4Nclz2FcJ3GTMafqVMfvwBhPrhagvfrjDdFH2l5G+ODcnG4O5mxnij
CKz101fyVcf9IbcvF5iY7OyhHVEUr1/Ys5GqT2IWy4BRGrjZXeAQgoDGO3p0r+9E
gZ+h7Fd3bSTXEDpqt7Jy3yk1TFO3SlnrkisWSC4fvsbI6XwneKT2vU20Q2fxIsDn
fmvXxcr4MnIdun3MnnxXanzTWgqz5BnxVDHO1/grHlf2PYm+kR2BvUSa7SZd23EE
fZ7GMZdim4NMLXELVfmLbA==
`protect END_PROTECTED
