`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHwpTpNv1Wh5H4MDCyjyY515tilK4QGIkfPAij8qqla8L9+/ZU6iWymiS5DUM8FR
B0oh/cS7Xjrvr0p8iU5V8o/+d00dyJEqGR9KivK6B5b9lAQLBQJA/UGWEMzMeQYs
6RfZe1HIuaxuJ/rAvLciLac0V8e/sKNZ7MShal8CE3oDCCbjoc1sJjxUsPYZ+AhN
6muMADVoSWv8rpg3CTZ3bNEVrhkxd0cWMkLzXV+UpxLFvN0xYGO0pe29S0cFN8eI
HKRuwaHf864HfDBF+n46rpFqu6ukO9HDE9cfUnx2QB+k2JtlGFr7M7N59BKLIcM3
111Kcu95Yg0IA99OVELWbeWIIXhRGpzB/9h76ylLcWqP1/CObW1kXLokJHj4PuVO
z/LOGRY2Z7O+PU5x8zr+zT0/7HNBZl0JwsHHedQGjHIkYmBZlGn2PyO1Yg61/aJr
4RTWLFFElzsuNmpyi7L/NRtbeaBvVsWgL559zADGpbwk6fFjD1l7BivQuvyHEN9S
Fmhu0BPJHvqrS/KZik7o4Qijpf+v3LDn+BZ45ZN74uft4/Me7yO2p8d8VjiSZKn7
ugpjgUlCjGV4Oci0mThTpVsCsXUTlDvUQc8slfKVdJaImQnSlfeCTOt/smlsnl6S
uNQixK/EnJN1+R+GVjkN//kZ+j2cpXfv3G2lQ7BkthhzNOCzbsET9uFbP6hBY7F9
uQlZ50kzFfP04h2HO/fqy9L0wZhN0R9kDM0724/MHpy4tNK1h8mdcTv0JLtu+Nhv
+EUFjGSPmElZCw1XNhpwcK13/i7CB8Sc3CqN63IGz5AHuHjOmPs/plxU9UAYrEyz
0P8yzgktgIwRi/3LSwc35BChUDT1Z2kbPybAg55RLj7c/l63de7zNHWzcBw6VgFE
JfeavAApk2+4CuBiYDiL6JkQd+5IorUzQRq4eLRQfa5z88qAhZDI167HpEOLcUPT
r1mMi2jiR5JtsFDnUCsEwR1ZaiERs02daoAUS3xOSmWKuapM+wBHJvVKra5UUA/7
3iwWOFbco5ODdeMEN3PZjaZjWJqdGQuoylmEjXNZswlZirvq6CUS59tj3AWlhqqP
/k1+Fqj9iSSdBQ4hhiYND5I3FJkmxjAZHyxwZHqI+py0KSbLxl9hEpcol2k8u4Dc
v45gkO2L1o6yZxyELLIFZSVX4qeDw9oPEIiLzJHaZbAyaL9IRJc1ZEUAOr5rWu+b
P2SLMD+TjX4eCVsfqtc+K9qFxcRYfzoETTVa0FjYjfDnq52jjXe7dR0rd4Q+56ga
NiWlDejiSMBT0o7q8dOJyiYI7i25vznbNEi6I3xgnGsURN5w7fyEyVj06jL3Dnsm
VYmufgIwoHpaF1px7+TeWqE+exqr7PevTQdtzfoJcDYdtb3ob3CI7ppOzJza2qnC
x9eIw+9wAP2eo5zof79Cy5+g4PF/OPdS9J/K12gJaoQDR1OHhoq05Dt8n1FPBLEJ
yHwzD86DpOpWcSBcmGakZGW8+IeLnHwgKLnbYkLPXAuoipCLTjQJfTuh2BBo13EI
287IBxapFRMHAbSSaskV5PVxD44hfMosXKPHCeZHtFv90u0vmsOH/VldMHmXfz73
`protect END_PROTECTED
