`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PzEtFsorg9Iq5GqIQ7oi1/ZHu9GYPqAc2wY54RGr4kFcVS7wKWpWiV6dQ07z9ROJ
2Hpf9P54pOr8pwwxI+2GMCOepu4QU/eDzCXTmzXBrbWCzIQA8VTs+KmN3MPNf7X/
TPq4RCOXPjQhfZsAqOUX09bNIaTt1D8qFxqhwlHe+4XbDvtAg9RhgV8/7QCHSj1R
vMIGaeu9YwTZApU5hwSbSjwK4g/msG4yyBb4GHzihYeAID8ut58R9O0V4WKdLbEB
Gw91Yp1+R8nHdu9LpUzXQazhsD/7qElOxc0mzEH7XyewdUKs8QlKV5W0tT2ZWyTG
gx/xzXdNOIkwhrtunma41nyVuACXRfE3a0dP/SwRytafK7Nyc5n4pFYD3EVOKw8z
qrBFavNnQOwOq/uAdANwjQ==
`protect END_PROTECTED
