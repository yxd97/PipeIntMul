`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WrFtF00RbhGQF0ELL05NdK86d4HobH/dIwbx4XrvpMAu6LRqOmU9TnOKD7pYoiUa
LQvJEsCwKhMCszE3IZlxHlrnZ0ijIcLfCHH90vmOP9AL0KpqPO/B7hUKz4zXvDqB
QQ2CBqUP/lGrfBugI0vXFYXvln79Kh4hpDyRA798lTCD87dliXMbSaPfx5TtO5AP
ebkki5Nl/UnlOO5/+6pAuHZgB8Z3//nQzULT2LkdbAMuHbdbR5DWX77gVZqMMUKu
E6WkmjXbC/LBA75rR19637rKq/khPl/eZmlJ1uIcCJL+AMS31yT0YkRna08qqVi1
M37prF2fR6TkerVFXUlga4v7lxcu59v0xRIxdGkI7MZzMbck2xy9nxC4Ptm1DACo
dbMU0Ywy+uTZRaXAI0uP9g==
`protect END_PROTECTED
