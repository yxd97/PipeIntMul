`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YuzAHticCwnIUOdcdvzyQ/hk2Hp5OsvzYGJjcfUTxMHsGwrwbYdJgXGix3Ilb3Kf
JdapyT6qUcGGUzOeRoqq3My5OHRlsoeyXCR68r9YWDwNROGlP0Lwj6pRwwMQbRb4
OWcHkIQS30pZOLh93OZ8eb2oCUJxpbnqphqjaU+OAHpPPeyV/CX1jrMk8KacnSUJ
FIW7d3zl7Wz9jGpcoEKswaEO4Al3HzkLkzre4KpEYPRdUzMpYUBym9HbyVQCPSTY
Xoy2YJ94PRRf1pASJ9ifm9ocfQsySwwcWkG5y/b34fgDUwgtf9Q7nGvVPlT/mvRs
i1qkGn+gAQx1Zya8XUYsq0P+WzvGB7MVcDm5QYKVs9jR3jJywPumMKAUNMeqHXzK
k9Gx9yLIDCHWnb3RyweHJQ==
`protect END_PROTECTED
