`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jplVdz4yoifTFmETFSQ2qxn4MMQnwh4AtgHc8qyP+p1/JR354640WBYeBGTbvz5s
5i1SGZloGqkkQMiL7SzCs43z6LgbqwSxF6ZH8ju7eaMYW4+vcC5rpMF6jMAGBvbN
ANB56uhD03VrxMg5yBko+sogllqOPoTGXZZ0UAJwAYpuIuEcJnnvydbWpvLxLAID
5rtnBVgKmiz/qsF1dYD/JZTW/U5EaDI+pE7+pl6oedBl1tlrgzIxTjr9uYAXUVq6
BPWOEUygvVjbV+MKGmL+hlZ0iY+251RVfqknmXkABTwMg9kek36CGwOirUPCMkoJ
feaO9Tjj2CINUks5Srie5ACZlhMvyOC6Ov1JR5v+285HIzrS436HTcZnNkd3uoFH
KEM8T7BrTbu1IDLGxUFRWQOcSuzpGRpol8H2WAd7LEvP97Z7QNo2WCNCGNKcYxSG
fqpyS0dRwR2kRgbls7mAwhMmhpx4v0EyXfxx4hG5jvNeTI6Eyg4pb/o11ZIoYnBw
mrN9bg6lp21geb49vmMF9/q0J/o6fyH8ugtyN8/QaYYxoPHTxCBZ3EQKS2Y8rlmg
gdgQ0547733g5VvsExPYUOAZkra9SXr5K51aFQqYKjvLovU6AfQFErXqw0s4ae26
AmXPu8WMcsr886U0kFUuOGJoizNiPZgcg00SRT4wP9G8dadQMdtBKb3GqtAXal54
C8adr+pF0n3sYpC9diREjBX+UiAc2bmLxvkE7wWBpbN2UHfN+AF4MmLg/RJaUQgU
0hfyTv7F6x6X2rBPIY5dDw6LG+p+Ox5tZEOCJM+O9wZN5VGeASlBj0tLYwlQhYQ0
ILmemV9M4q2OYRHYBfbKo0m+HLdO2ybUuePlbLWggN94TJWh4R+TKibaQjqHXtzX
I1ms6PSSRjeSuUHv0E1aixBPQcwHK8pcmgZgOoMLE6ZzLTpDcbwUMHGE7+0ux5Zy
wkwIi7lt7kkkPqSKfvkjJ3CQCSP6P/oJBm/3ZjGPmYSX3b2CJeN90KsxvXjFoire
k0d5BlYU3uhdeJaMW9r4FaTRIDDFAAuYraucL1SEUid7vbkLKCPF9c16S7rn284T
SSPjzn0sIflY+AC+OH/MEeGAP92euvUACxM7Z5hFR1z2C8tjB6fzogDPSeyg3T76
PAYnwjkYcpk/9xTteuPdFyCCSBnW77kNhRLAWMaOzxbr0qqia17rU5PWHeyUnDjr
fJhI0zqRItXq3Pt7CQEzRRIu580+kce4R4DmaphjGCxmOCMHe/71IlxW3pLcK0BJ
YKUjMVDQyAhw9OwmST+mKh0CbRNqvWzS8E9+QdzLErMRZ+3Zibq/QHiVAQi+pi5j
kxQsxd4GL/AwErABoA3ycDliwDOyJ2Ca//O+ELuI2YndNm22nnvey9sW1G3W6gbb
ny7VWtkONxO0Cb0H+Vy2lx4Gt8szVTp03ewHDm83gpMlrGboUsr87THtn9uYyqq+
ECVQirAZyX0+bbkG93Gwb9gg0BqL1JM+CHPKNw93m9fNDaATh+o2XoRKrFX76pA/
DMd1IFw7mKLhkOQbxKxSdOdDnisDdtO65W8qb+YLznNWq/TixInY7hno+oWVw5Oo
ZueHNftkxn3Ix2uvX/r39yVZtsEMM/01YXdwL4PURKKL8JLlFR7CsDVOCrEVy23y
7XapjSsaX9nZUyTZ87Ab/6ST4nVyyAm7z4G2OOZXt90b2lr6W29AwDFzHDqujMdN
HZp/s3J+GTrRbZ2FvJCXKslivIlRUP6Uw40c6ewn6OS+FybH3cx6wyilvqyYfPu4
jmYw5qA6Qka6C4fDKThprJsj+y6PmJoOXYLAA+2RlMYIPay90+VplHfnmuwbAHAO
UiFaUY1G1WwrBuXJX7q7x4cogc1WOizJn9OubOJQ/kHyfF3CPRLQZ20R4W9BIP+s
i5C/NOKDQa+rhewZW79ykDDR7oIOQ3cSDNQ4XguxQf6Zyew9zoaTiMwuPDiycVHx
G+OKyhCU/JSGi5JKnvvRT4bMWOx90vOho3GQeSDY3oJlXIFCngh293KN8u+bBiJu
j8ebu6KdNlGqPu9Igb3ujH1hu4XNeb+KGrpDUNTP1yRT4lLImG0i2p4D0dh2VMEf
qzOX9fcqi1UNm+p+ur6nPGJUUzGzEX5r/Rbu4tgjUcbCyh07NrH3aBCT8rS0Lfog
aEyx7cVX2ynYP2VPESNyLUfoidMQvkh5ZAmv5bLTDLKZBvYPZ5nYWDQchTszxqW9
LfP0OucgJ5A7aECrLYDM/1gi6qaCuOhIDkNv6kkWuP8wvxAZT1wT4G5KSku8a8uV
NTfNB/kjoLiiOL07u6QP719oXxEahcKohqTNPqjxSd+Z8USZz5cneYJczQueUSHo
228hQOV/lL0iwUlWOJHhmVnUnHbPMUxMOF78wz8gso8jOvg+1EejA00JTB/jTDWH
Oq6VU4E5KAEvBjYlzOq15FHe63VKSnCkeJKBmQChZdZmcZAtOs36bM3PEazOn4x4
PHPvozsttYDrxMWK3RgdF3uqfNM18oa8gwa3OCOMMxcekNRW2jgBePkqYe93hn7d
FvUtLy/Om2wx44MZn+3PaWmn8yLLV8bltTjDLaW4CTkpWcVdn1/fQPT0B7anVAiN
eNjky3oXcvugQ3cdGB2PBA3uo8bHzYJs+SE1GyBjMTU+TvoCMX23UMYDJCMsqRe8
BWIMHL9rgKDn5QR0tB2FeKRTzJGARDdJSHQHQ8WsfVFMIZSVB1WTvnGYU1FvqRMh
rQ6UJVtINDWXbaXLBUUfR2mZM3aE6iW2nnXacUOptxsoaOkmGYVrPYRuNsAqnUiV
dJycQx8eeevF28kedG1dl4DBle3d8GHqjN0H0mzzy8bqgC6oaEYPz0gf9oLrlkVX
zjQObzWtIiKDWlJzubeXzHTUrJIdjD6BG2sp1RhgdBqziNrdlW5sJPn0So3EykBj
go8b4kscJ3KV2rehryUSDXze/PFxPEdze4dDVDqZqITDGSNG+5l2CaIDrjRNHM81
lapn6/zCsxaPXSqcfaRz/SXiyFVrQSrUnG3k/mO1z15XTSMiinZ4BaSza8KIJzNo
M8VI+eaqI/drs21TNGMupf5DjIlhiBFS/FAAfUjqiT36Q+LoG0NSN6/3hpw0mTJ3
kRb9BOaWW0yeKdBRoAItmt06fnDj4k/ErNwIQjoxKpCOdT9PR3hm6K12Cx2juioZ
Jrn3nAmAROPkaBlPpkcduPn8kvvp04z7UuVre2GItN9xrcke8HsZkS92mOwpDhgM
8bqjfiGCRfQm4r5PEtBh6ZuxjyElAVbohdcv2VpJDBQDmYYbkfni88z7N9PbUwwk
ZveJRWstUcL+eD206DrtuQ2cWZcKcxVRH/++EQpOt4LKklWAhaOm4Xrj6p4ppaJf
hi1kUNFb2Cwyt3+nZr7SS4yefm4DXIWXtWXBwNvqteQGu+VsEsf+23oVT5ejobpC
Kcs5sOAUhBxQ4g1OWuD5p9U4QO1AoIrskgeHJoiIpHLQloLAQQNIVLIECJiYycre
tDu8HoCVU1M1AB4np1sBev0nEQnrM/lH1YFg0i4tJw1hlsk6X5osbwfrEGjtwL13
ojDTPLeH//NZ8TBn5NCygDwV8bxezVrGb5Xz7amULJ5STwgaiHmuZ0Vb/GfKDzPs
QHRpuLYz/w60ewWMm8RcPbJScJPjzb0l8dBwLajf8ZR4mdxxo0ybmpMwtAQXQqUU
pJN0wqS2FuAWqQoa438NI3epTcOh64fDzkH1pm7tMBJnr4MumLckxmsXzmry3MSy
Ra1PahEGpX2ky1ssBd8YTHJRI4IVLTZphFFnFvYHvWG0tppd7eg+k7f0qB5dZLBJ
/HjPB8dSHUQkHiUAgKBaSMUNAHEw5Z7GJYr7EASqdtC+sYF7Z56fou/03xu0YIhp
q2Qq9PDwN64Aauf3tTG0UB0BTKlBmWoX8pP8DF1NmONVsQNROWeiDQbF5cY5Betx
ZPUsTblu6zmc7YeugZV1QnFfpGWEtnQimbMq5bJQQllQXnpoFr5ibOHb0h3RmjR7
7IEoz9JIz1DYpYV1+98ZKfPFA+VGR4gzA/cIBHYdcWX3CnsQsp3U2RESYyml5um7
HTnuFs3w7X0u4EV9Gn7ARkNaMlX+DMfsZYU1N2UaxnIupfJjaZNJRLwvIx0hzfzs
tAepPOrNoeNWv1Pumlpaxd9qJIDYn+PPzYJf6Rf9DkIhX92vD3ivxAkrkDwszgMK
NLixbzNM+1dPtnvg6KV/BcqEMZy4qzfndYRdFHp6Sh08FmOLf7uVQ1PyR2CWEORe
spPf+HyMC7Aa3rL0CH1b6yhNEv37mGJNh64K8NSmC0Ov4Asv0JG8hXjplfs4+TVF
gBkcy0iG/Ue489iLI1JisifppkYkgdHPPWseHDnqlFLXSHJdO0D9S9kjBLivxKBB
+E+uhLRJFnEqvxKbJ5i2ehkqfl+LFrIDDSqa2ms0oBaNuSy4n/xF6rvZrCC/SUkP
sKWKU174ciFpg5AmbQEh0uqa7GZiKbKuC4z0cxlkq7DspibNISEu08/x1EKxspGb
kBEAN3aQFHnYlG4RZyz77sdRpQqVfUOrpWMwCRF+3DQwEzRAs3i5uOHnIddl1JK1
33L5zfk844PZoYYRysqxPqd/lJYB/HnyPMAa+R439O/RQ6uz0ZiyolzPhoXJLEjN
Z3+xtPd26I/ylvi+DWRk64jQUPem3kE9ioyW75FACugQODRppNaSldiWk4Fzgv0w
m9NM3e76rFhzI8+Cs+fmpgBlgMPgEw4sTQ/W/DCyxKb+aoWS3BtsBo4FHu3Rv+p5
nZcGtg8VX16Jt5fJTUZ1F+vby/DG+u+xWWO1a2W1aqV//Rqj/G8mcxQdrhRl8sIg
l6zvaltVuqVuprzoHRC9zKjKP0hFCWjm2XBKVVjPwrrLwxobihlG46umfDdyEvym
qBQFOYRZ7N5EwCIThsgGKANHSEa/foT3l1yKe8192OMnFdIu9TW74KK3JRRZUEHl
IjpeNkSqd6gUNmJE3E3femM/NAbPH3lzVlEtf9XMDkTBMiQ5ne2oyyUKxNVVhEXH
5dcxf9nOZSV9ma1TJvxktB9XrigfLCjD88zii0EnSw4XiqVq9Pp3/r5cal+gx7KH
u9NTDvT7r125zWMLzyDr9N6f0cBYkaiwN+WLra9Dg+TjiLDeCjZ1NBT5GNlNeFLv
+tB3k2eI+IWuvDuxXmZEpQY2l8Zt+t8NHogXOcPYPuqidVTxFTMzfleJoPBeFAOR
mrnDQQ4jbkQs3kbUQD/+YiUGNMdpMcQkt4ze2yXKaEU3wxUHO3j8x5VFFq5nwyp6
NBye1/VcDuunbG2rjvfW69v1SWm2HPyTYZXWhWxuMMJ6yXKiQ9mRxeW1I+nhjmGI
knlqQeLD6zHJKUivAc6sgoK95Hu26oOpg8Ph295yZ0kquOm8G0ASxmiMxgqtL9U4
Y5Ukwu7sx0neE5vMogT0M4xpyf89EbiOhtKr0WFW142NnUI1FsVqSNcJnoBwr1G5
WfG/XdqJfNiJFNyRXdD3BPgpPDOoMsDW9Az8myVFOHEMhXgqC2n0NnrI+bz8hcPl
KRDodrDnrOZd7VAoTepUv63//kmM+52XpZcFR+TKIQrV2hmOANC8BQ0H+moPnRMk
22VPeZS1GOBZYMZZ3onOInX9O0gKSjAl3Lu11LVsTDIs5LzXi6GW73SWvUldDdYU
g+RlQ3SJDSwJLqMlHO1eHu9QzJ8I53jl/kBbtfAeNgKr3/4c8pQT3e+fpptfJ6/k
QBDhVccTrxTArsKw+sYO29A7FuwaFD7xa9w42DWAwKAElENMmTWMaR9vPVOv694v
4UK8Flsnnfn3ISmUb72aMV4NJz0lwlwAF2HYIytkDnF8Y54JVIUBAurFH8CMr4PH
HRqtsT2vKc42RvAaI0qIvm518+Lm1tD5wX1d2YxbYuFVlb2E6LOdWwxgzVnBXVte
6f2Sbb7MApPwfTdMtUQFGJtVhgn6Mxphy4ll5Lr5Gel9e9g0r0QIBnPwjE5oaVVZ
QWrTvVLD7MhTrIzcQs4iHddVNYgVqsnxH5fFsRS08RcPnaA9U2itg3jAxH8Ha98v
GGxtHve+fAAefckTLwZejyLLJD/0AMNAhsRrlW3W3gBZWmJ3df4oIY36LkFpLp8d
5Z/MZPtBYWqHErSo4bvm9xpn+7h+KnNHLTG7FSSu4GsxkVW++JHH/vHlcuMDlM9g
t8fOJj76huIeAGvLPHfNnxHrAbemMmFOHp3Tk2JVjAYdRN5GnGi00HacKyX/KTVj
pOuVvTYiJrLp53Z7F/jv0S0pJNu6PtJOEQd1x65jNszGkMdBHrkv7VXeUj/6CAKG
ulUEcDdSD7tKYBwSlxIzpxgA+MDykmfbXhNfRNyNxsY0K27fahmzaCCHHpoxTgOh
bXZ+vaAErqSZKBSFiblmrxKdFywWWlnNGCvENkVYYxorx4ZQH07gJmVC3HmaxKuc
WUXQA7OicZOSYLo/WGsA9tlWCJTjjDaRb/w9f7vX6/uO/YFfGhIh1v0mmO4p5I02
lBz5gcE4wDQ3bGX46Jtrvaqc9bAEHL0SXQFBTSsahuGdumBIQPTywlr8BZuFn2IZ
zj0vQETAvKqfu3fvOiHGpv+PcW40VJiway0oPTF3wLubiyYUwqpyRMglqJOIVJ20
C9L+/u/LdY85tzOrVn7mtKZfAB2XJQOHDUcmCWMl17LZW2qlF5EOngQ7/LDZuMU0
bCN1Y7gqDFgcAAd0HLqywQcSNl2Xhgxa9T3oMGNraW//yOcmSO4G9ojk2ofPkw2O
2d0sVjQGHHGAe9MryyLHApN3yGWuYFZFjp0N0FCtMpX9XgkwMhNYkNCt4zkJTAqz
Wjc/QDAmcC5n1wo0BOv+i8iEmwCVuSnpJdUMuHuP2agrvG5ozPht1BhSolbTi27V
Em6q76NVWRBeexx6txmNy5mguBzo45DIqOZ7hmOlVO4qzXp3j6KI300OG94EINne
1Wx1mLA/n3C4EFEacLX6sxoAARBCt+y/l3BNgEpX9sZlqiJzWQd3CqOxbwLX0KB8
Mt103RwcO/4hgnABW0Sa4YDR2LNC0iPZAlWMs1BZQfuVOvIlS3GXNwk9QLyy2mnD
TtbbFLoj1ZdO+ZcX8XBTmOHy2ZrLV1aEtStnmxnJu+kMWX0GzyBiCKgoT/wH26vN
6CmiZuoV8DCvtbIo3pjs2p4NRgn7y1qaY5UNq1BoVxoNXmERglkLPFhXCRb1ZfFg
xKw+vtT+9rcKSx3mvPokxZvDFcdWFFVFWTQddVB3Y/RK2PCQGFH8YoeDehbqK1A/
DcJPd5+YdQ1vLXjF7nx4tuQ22k5tHd4ZTsk5eg8MwoiQFN6sVPYHVuT06iVGD7WT
/Q6MD2/19QqigQykr86JhfxGPg/W2ArN81quWywCrUpgIWM5cGXRrFWNBGpBoeGP
McOf11RVSqSfMvDR9rNRMHcmB8Yj48bdUwbfiU3i5IxCVO1SxQeQfXasrXhP7QN4
03nP5QdaGETD/ten2oZOEA4aF5iLuKFNHgOz8EaojlXSGksrfRuUICoOMADvdIKb
1UURvFmuJ720qvf1rTJGZFCdhW8zCtUyKswxOwnD4Ft4gmMdDIJyOFhdwURLq0ej
8MaznkBkzWGS4OkVH7Lz862MswIJi3kB6VVpfy2twGRXLW0GvJ0UFj58Hz7i7wEL
BDU6h+kyulEvnyn0fcT3dvjn75INY/tK2qnwjN42OBvTGIpuPIF4xqJtUFGrNkpZ
NI9ujqu1j/uGHKSvMVUCS1l2SpXwkEsXNiTBW1pw6qsMl5U/9wLh+vB/3htKwpGy
+/GKLawe+l54Jm1JixlgjdJlezx0pkhkE7+3qPOVcaG8x6/dO+IVobY4Gyqsl0eQ
Mrk6/oB6pvpKVO3q4FDWBn4JhsTN/zf+3YTGWbL086CPp9+ugNsyQIgRAWmW/9I7
Mlvv0GofVDk0Ckz/ioIvJ3Yxifq9nZRs9obv0W2HyDRIpp39F5Zh7W9+LMl8+UzQ
OMoRyp1DfbTQxdhdkiwgB2TNxzjy+ihe5OYHUe3TVHO9G1aRsUCaEntCRPNd4CER
ej0ikku0di281LHYrGZFyqXwwnOD+s0NYDX8fhcMAdPt1vwdJyps67FpoPTCYIhQ
/GGAKyrVNgXxMmjKbMzsMM9DlYYE761PAa/P+JaEudnY1i2eIxK0Cqrgoz65C0nl
DJNWy9PzvtwqR7k4al+XKPYkLTpnKizZyf2R8x/b49UVTlYiHhwfLKXXO6BtQa4s
nGOQ+P+1QR7z/SfLDi/thqSuaJmRhyNnfKsWMQO1qFA9+WCB2GGf1mHab4aCmVl4
mJY2iWY6XOSM157RLFRMuIh9Igc+PlFNgEYH7ZEIXVHNNyiv4NZ1xd4TqhOlAOU1
c+/M8jTKVP7rin21MGBAmRaYyyhxGezoAiquQ1S9XxkgEStLC0YGMi6PUOYO82p9
S5couol3FczcHRajOAf9RTqJiXj2pgJWR6zXQBCEhjMWxKm4miLR3DD2QFSWqvGw
fe0TkqxE91OQgNEb3lGn3LTmvQp15AdSfIP/E+nb5rNGw6OVk0c7qQ4QLE3DJrSi
4z2oACWaHnlp6nLLgA8s6HIS849IRqgy02o1fnDDzIFi3Cms7ZsBTcNZOxKQwH0a
W0UQdpo0nIGpFVTfyPxvwidl307uzw36YgL4zqgttoHIkpz7oYMZdlR3N3VA/z3r
w+YMlnHSIcLNnAhBChrpmBcUGMa8vEFclHxasqlJDh4dfSGPKd/lIm82bUdG5OqA
s4P/EewIai4W+Xp76ubKFiGGAHbmEcjrviQMsd01vf+Vuk3k+vV/hGb9TsS8KRQQ
CZIlXXogdN8fPI+7SX4DbesmjCJ3qkE/vxdY5Q0dXEqp4hwS53FMy0+D+Qny30zn
8pCoQ+/dh97ZFcwKjl48wegT7cXMlmzN0lj5eIX2rUJtYcs3MPus1aeE1Ags3UfX
7kjHedkLEvxIQknkmVnPhLYSe01PCm/gHOuq7Cuh2tN35BdTTmc6n+4atLoJc7GW
IbrIcS/bb9F//yXaPq9132IILfDLxEdgtv6vqFXjeCRG2Opk/NbXGdnTYoLKIDfG
1DkMKxce5IATKGVsJozdoTaKa614tW6SsxJgmSfKWiBJcA9pqNLSHEUSV53hYuZM
NB4yNtVA4qZjQJSyuKPnnx5X/JxcSLwhYKf5AS1AyPKPy9t8wRQjkL/e48wla3cF
+Ol4M/N3NIX+XWGxBG3d0ul2bVwnLRUL+dT0a+odUl6omUjRN1X5LGnD1O/f0X2T
GeAAzazdYiRVypOgUhsiWRAZSf8dB2gQKEC78udgPYa5hkkMGZ/gUwLlGdvsSexy
fnxFgQDefC10LjHHD4nvv5EGAMGVqSuJmA3JzlstSPt2VSl1wfWS6UnOeEKvY/Fk
Y5KQakPBd/TFuiKJ1bOj8o21uaYnuO/iEana6S5Rud7c2JOROMT6tGBljVdisv7a
4Y+CemUlXsTTjyLSZ4MOVlfkPGYGwucFSIxMKRFmguf/ToXObnBuworOS3zrD0uc
fQYtvNVwjRS7sEfDeGgugPi81TDnMrjf25O+5keHGmn1UjVnGLuodpptqcoU/+NQ
Y0tJmRzdi4yP3y2mXKyDLvtkpVuT+sMzVra7ozB0kAP1gVtr1UzuaOkEN7UMgJCS
nTH/cVovRplsGSWDUJbyiY25Uzv/uLu6Or1BKfPfspgm8StseeuBZ+zmOxVHNcw/
4ZxpnjHN7d7RLUaJWia6mgVKkD/PXbu2duEVS1pptDzmW+DwUcqOg6rzH/7l2Axu
8gsR9H0e/C03El+AbDyhLr1GwlhhMRMK57vRI623ZkyBSgo9Ck32g9kMFbsfJt4J
aO09maNtSRu6AWcdJWGq3BlHsdN3ID2BskVdFkl+FXgMUq93NkE+DuWUJmovzbQO
+ucIwYNZriru1KcOVxlfpMzjsKh8J1mARa7pCWAyZPcjF8q+wTI9MeGGkU4EZPnT
YoDqr5Y4QYrQymbsuO3BqqYw7eBQOoItwXLE2mSWjOaDTEmXI6uluWZ6TDsGXLa/
2pcsdO5A8xtWxmi5YeWHTY6htUKNYCAR527It4o5o+qqfFDxboYdk9lftpFNLHKU
o0GtvGPbpsxYpeaytV1bVpuTF5hOkk+6VouG286ou19cI6il8gMHdKfnpQ8N5ITF
IQQV9DShicJU7q72FSCPKNcjdaf41FAC18IoqjBQM4XBx5ABnTiMM4gtViyQGQFv
gXpS0GdP9DhoUZJjFgGI0DGQqOD+rdyUov88ALXyEAGQzLLhtnn9Wz0ZJhaiqT8I
YG8I+8uKasjbPsTq9UvP/w5wgZmOEkTO2NMmff3ceskAkA199m8/iuDjypdor6XR
UB/Zeawm9XFyyhjJL/Li5FcjNHSGu3DIZb/3tgEktBxwMSOgpf3bnu7sSYPZJmRo
/+wqObf+PT7veN1W+33GK18XYVQJqJ35V2kdHaHhe6au7Py99FT6LB4OpWwas62M
cHDyjvv14vF++RiBLQRtE8Lf2HiXKbji8hY3Ccq8mSq7G0rJYcpnCVDg8w2a/v9r
wlKwTxXU+fc+OlGd/k6na9WCwab+XkGJj+2jqVPKFf+YBFP8DngEoS0yyekXOHTK
T8fUNX+YvqTNgPsR4rDYD7iNnk1lMifagJJyPt/al3B8KeOcWOhzbhd4uCFGP4ed
OVHzgYcMQyctPYvEw5JEkUoa8h8s7/XiajKFVLUgr1z4HInfyiDaybEF+LetPxm5
iSrZeLKv8knYahDfOzlvcx/QvTbMuYyfASxHAzTZ8DnUefbeOKe4rOElea864GQX
oa6CNiidCoLF5qWqzvWfsdUHzP2TivZgA/FiBR49zwzVO5eI8fRAeZPiqUHOMElY
loobpiY2XBnii+cHfnMuXgC4ZYtW/LRHBE9uzGGbR5hrOhPMYBtc1CS1GJmIBlBm
466+ZxGU/vv95KXP5bVUJaKRJi5k0KRcjPjahx3zBiZQd9ErFrGL/jb1BAShwkgL
3FJUC2nwnoqie93Iu5KC98t9SaVENCxx7ID4j695dpe7fcxdZm3BI9lKj8tOvRqo
3g0t0DvLPNWjEY4LshAwsCdNWY1x21XNUo3va6+TFVwRKiUCGvl/trkOwHYwXlhS
EhcQLth0xULmKFTR6iqR7s+teEdc4MelaF0ICM4Sb6cgrwo0RP1F6GonaBr98XxP
OJwxU3MDpOSFFnNoXnilmMWwPtps2wyLJG9viPn/engOQruwFM56GaQu1cOdIcb2
t2r0G4bLIw38urEAC3W1VmvBPxcX3nKgbyAaDJM6fjrMiYotejUgGZ7noXAydWQS
R6qP9+PrqIdg1sQdLM2yXeIpjO2+zEKjYrCKc/gca2UdrlfyVCp58ojrBDzynACL
U3ijv4q7EB4tXS8nr2YL0UnZZdE9tB6IL/I2WpCi2qqSnEQbPkGEISL0wzs9SzFA
ZUJNOnO/XB4hSkH3maUIFPf9XwX9/+k1JE2LaBRJMiKOYqvkC0DuUhsGD5l7lxwq
Q/pgmUsYsh2yUozpEF2v+j+Khjb3QuVMMlOaXx5yyZ1dQVw1a7I5le2uvohk12S8
3FY7/pR4afigBGcxdZEZFA3ZY/9mq/x99Qehc61HMMCQrJXXaRFBEaxP5kL8eME0
A6WxUoGVQhcm2/pyA10mDRWd0aZSDvcqexrdJmXbqdFPH4V1ml6upre2vwdcnH5v
KyZZFfpNPcn0GPI+m6OSSHIUP9cTINYunxOJhdWcfJPNRatusEjXjyHzgJiAMA8m
onTemV5oNe68TXdWGZiLB5sI8LczLmp77OKV36tB6f96YLKgKOf9p9LpyjSUZlDh
uuvkjztHhj3vMBirjoCQxrqY68AwOb8QbBY0qKvi5fE5gQTnaoN+rAFpvDpq9E9r
ZTqlWgFqkBOdKJzKzIw7KRIJcsa8idMVcsIcJQqbja6WNBQt7T1oi8/9N/okHMgZ
VSkGZRzZVl5l6bi9WxxZr3/zJgvz7fn/ncFAQqlrwpVkHrMDQAu8KOacieEV6DG+
pjGDWQ6ocINemdyTwUYKymHoLsnQzruN9xtdjn22lfjKuDO6yk2KxdbjG6BNMEa0
2K2rumiCO0YaqSYHXAC9YDSyHeu/HPzT56sOGChBLbrUwUut8eZwzXNBj//eme2E
IWNXO72BI0znlYMGihWLRmf/z267l0o4ghG7CLM9oPmM6C8sP7S/rh0GoU9wm4Fs
CA5Up4/TVqhc0O/TUEjJFs5glWR93/E9VI3hB5pgfxrW1l1lrxjfWY1teH+OtTF+
rjp/onAJlYJ/R0PYPQXIAO3yLVQlyaRJw+dk/cOlJYlRpEs8bDnJ3WdY/ANajzVR
az71uM04XQnEfOCrK92bUCXfcVo80u8sLfw2IUPd+ZNbye9vVm7Mpng5kXxKnW0C
VJasbEIF+ZVWnf8JmxucZPeOEXgA9B/PJ+qc8LByVu26qs88hAeqtuSwlG/ga3Xt
nu8OjUV33262YAv4IgL099jkYGtv7z7ioYv7bxwAKWSDel+/RaNCRLlug7AvjqON
ZFiHsMUic8DkpA+yJWCkrCJ6LcNZK3Jwz0mSZC5kXS7JV/MZ51/bfmPCX54DQZHU
C7A52ge4CY5PRB35/IV9iBMco1eaXhM7CpIdOEa5zsYy66iaRitN/8RlcIWWOHwq
+TzSW1FS+w8jnT4gHizt4S9IQUvVbOARv8MhtyQvsBttHaNPSOAzotufzvO8yB6w
2ERhzhLcLOqeNdR/CbaUGLjgw/KqezFdPvk9jyMQ57LeTNORT3TAG5fOZhuEW1qf
7h7vU9fSAjBJybU/sk3H/+uWCrspbZaDHAJ2GguHLb6q8nONcbmkT4/TW5zkX2Nu
t+uhmnQ92f1U7//S87DPvKlg5IOdwwizo6B7fje/Wi1NEKzGwaIysOAXpAjN2d/M
Ys8HA3AlZJXBXY8Q+J+m6UAXlbc9QeIZrPa91iC7kGYOerD5hlMmpTzb9bWwQ5t9
O0DLiMrXi3Fu0VgQnobs+OQ92HruFLVcBUr/hIG+HeIB20QZOgDO83kCGEkzu3BY
VQHh8Qa3DN0uMoebWbLKdpGGgZh93RzP1Q3sUHQt/iqJYkKYP0MC8P/hTbHylGpm
ZXFaCAQhZKta5x23auTaNHEdpQ2ZBMz4/36oRB4r3Oq9k7a1+JU+OEs2GaUOJV3a
QWQFPk5RvsRhut0t3LpCPs3ckQCq8kzG0tOwRXazmhA8EeEASh5HnCRltSNq5Rci
4hj1d9gXGmbYtdxAl9uGFqc0pHyV/LEXJY1i7M7rjjNb4sTrSrs2+S5RJUvUyEv5
0sGVIS6c78sMjm+yg+TIuHzYII9yKnRoFUq8Hz/CqeEVgaXyRHUysj3XOnFoxLe1
/Uk/uqMfr5nY2nalErtY3p+0kFw8xmztB7bI9hCa2FolYeZR/rFwqe+8oH/0+fJ/
a+Tnz8tM7ooWa38XXUrUAbeLzqXnIs+v9JoVYfXP5biJBJb3I+T4FUh9OocjF1ex
qEeJ7TmP0rHjO3dtq9O4TVPm9oiVe7AqCpAsBg1aE/XPIPI1v4t3Y33dN0TGYhq7
QBQqhzmswI7RbyTXoS+iNJpE0aWlzeJxbUUGQxKPfQKOhIY7UnWVZ8aI5y45fCOB
fyeOS3eVsRutkTVYJzQen5P7RA2wTkoWKYgfhaF2wKQZMSoeKBWn4HnwIZU6eNvz
u330Wi9NrToPJkOxY8USZHWMNVP6QCCXpjDs9yBDNKsFY31fbEPuDz9MGWVPm/wY
uJOM09HfpuNsM8kCTD90MMGxRPQa8rmmuDxj0t3t7PFUXAqti7gaO/dLyh4pDb6x
9YBb+z1oBF0j9ItPekXMS+YM8wMf5ZdpHMQ7FV87JVeAopxrbkp8oe8U2PcoB6xa
A4WzPpxAKfqlrOos+fQJ46HXmAc9AMxz1T08rpaCTrdVpituLlaoQAy0QtOXlUtl
la5jQbbjb0uFQ9EGO7ISwSkikcx/AOVE3dST9HxaOSzLOeCNoQhSINDXwhpohe95
cJcZGwhI/Kxd/Vqx81lAk3NCJaiQbnEoDDp7gkVofzQXDSMHD9jQJIrs0ocCuswq
NyhQ6bR9QNUAr3AUEW3q4Z+S2lwuwIBCqE26ssmRt5GMEq0VuQ4MqHKfIQ/FC02G
ogkWGYttbXd6Qg42fUT2t2SUoN5o+wwxNT7DGXMj8UQbiiGaPGktN1aR9pMM56tT
hB5zRRlnA9xvCQ7j19YYkCKSM7uqdIqUXBZD1Pnv2eCAy7An00f4tSnPPa0RIDKd
Hox8e54i9wvuO4iV06IsybSGSMEqhJ7/F9H8APnGXYWd9nV7xqYp4I3A9H048TBg
S7RNq56nqrllUID0T1HFpAsfYQTzR7+iwIkG9ZczeTLUTQnnAW7ArYEdVjFYSNte
exBn2WDJqOdVh5wjRji3f8fm9f+jBRlDF7ARfCy1DaohZKW8L9BUSXcF5EprtRk6
/wOutQ4fjPKsRcQhfjF/P0fCSaiEaWeW5yq714nJkEC43TXYnCUDQzCRO86ckMCP
PM0CHQ2gJ5FPI2p8JmxqnuJ/smupTPzEuFGkflMq3jEqevZuCndHwEPlKlRTQGpO
OUWIA02c6ZL6KG+Fjgp7EXF5dpm03Dfst4FcttQx7X5TqpNoIcUQ75FKnNofFrcf
Wta63JWrGrovDqwUAyxhnz/1NTVmY3tiez3WU2oGtuGMEEa5WvWUPz9RVG50bNH0
mATf9Xra6r+jQqCDzq/+gUxz+mhG+2Y9F3ZMNK5YWATTEREV61MYJY5148zLFKNh
SoZZ+ZVIGqlOhd+C3KSvju6zCmd0QQ5VByyHmsseX+qxO0o9stH73r1zryHeMIxB
yVB8qfiXhcflbJ6KzGTX+nPXwL7bju8revb+k7Fy0QCG+tirJ2YvHVtq+zva6aZC
dQI7QylDfEFZetXxEVBxGoh8aJmUosOtrtxypzBHezrVCO13+b0gOfpz3eR67AWT
fN6mvFA+93ibpTjNDk6wFaWh8qLxbRw3kZeG6+XA0GfVgX5s2RrNVX9tHiIcMiNH
yHK4rN1OOG33RY9sYWdesf1W5l3e7cUIrjDt/rSMRP7ekzcW3ftSqMnl8ZwhM83+
5cRUysLjFv+rp6DuhjNNWXfJDMqG2hxTlpwRUrOwcB/4VQV7adg/NgPqdxsgO+zt
v2CoEaWLd38q9hNExCOePm1SCm489hhHXNFXZr+qAJm28sq1clB97/EKjnU9j3w1
lu4Kdhzz4PSB+dao2rA31uNp190XZCMRmmw6/U8xIAgwWIqkPbX4/TDznGrZj3z9
uFWCoR0tIn3cLpws204Gr4ZD63k0mQw+3y9T+A+xO+j9r/AbDKOYWAQMbF+HXk6R
nSIcnJKKmESW/iZZb/jQjMnAyixIQNx6sRZUiXnnYMO0gI7usfWKu5aQNHaIJgFp
8sY/GXjH0oeXKJkzIVCf7Yt4yRgxENTnUfT4tBIbsjRTv8W/t/8ouQzyJWAHOfBN
uknSczrc0saEcfldnxqbkHR/hmkTPMbEbr0VKHq/xKBwvZwAND65WDywrhGi4kDM
0r+azwKnt5f++lN9yofeZKKPZPfMrQHz9LBKGqovCNSOfbQ9oTUNp6Lhx4nupJv4
dCBm6H/IbDigGMiTAN0Hre97tY4myOFT0cqjwaTANsqpLfOOyARbxkOyiKEk1Z29
J7UWnc70o4ycicpP4sEpOnHr9DlRv3ePnnGHJnbHDlN/8jd+dS6KUq5AnR09QbJk
DDf9q6k+Zkp+EEi6qpjGuBK7Lck3g9PdKbBHy4k4jZsWo6niip2z8h+SOraPisrp
BA2QuOU+EH9tBPUQvzS/AA4mXbR4XG51YraPVDVznHJ0hndcz1GsC39HsjZ3ZytX
48rfdrZLUdREEm7jOvNWWb9Mf9HvwJ7izdEqAQ7B9cYt75cT6k/BUp6ic1Fpkz8X
fioBUs/9HaUKvmssjPChiTKLTtYmnTT2NTJ6asIltzLHHeDyqkltWivn91zKXfgt
pvXPPrQh7FLO6Zj+yHcZMIkm6eWWKVhG8EVv+r7hQb2DRAtxLxZEemG+0a+kIjtT
CaqN8lqbZO7XV2SdU99Y65mfis0EwaPG1M8gUG+HuUORySu7b0dKBEnGHl8nB2OY
cBQplXOLF9RQfMqyt21FPbk3C06OkxPb/Ct1iulHW7xMcWWBa6hkDukvg2ioMdEl
MCMADqYrzsHJHoO7kBh5KfeupmT+eJUHc+aR3gksf/kLoKIlBzP3IHYuIqvZINtm
VmU86gXsW9TSAXaEmoxhkaLKWd9qP7Fx2c3XDxMMu+EArH7t7ZUFMEcFJarLCZBM
aBGQ7bWIQFHBoBaKt9c/lMGNfs2T1zHQxrIWt9TwkqQ6x0P38dvuxviUIExkvgZ6
QCpQpRx6HJ1hFBoX74GO2tGasaC2QQOkr50Xf4vSQ0GarVcMFjxY1dfMuYqDfOwH
GyNV+u0GiKsy+4OwfPZ5FNZJ/Xn48tHel4TZhopUXF3duYP2o6oDKqRGMXN76TNz
+YENyQabheY+cRAV92YUKAoTufHc4jyYDc5FXsFWKBEqSRhBxdZYgXJlTVR/qWyD
GveuppdjaN1wjv3XzHy/PG57tBb5r8vh6rsohGYVVu40vpzkn7e6zZEXvCy2Mob4
u6a1Tft+Hvzc7dnf4PDwba+N8ztvBuR2HnlPXSoPJd6+llrcZPhsjBAX3mw57YcJ
G3sRU264Z5LPEM4X/9FhwN50NdUvMgHFZvPqKFI/I4JOHaVnqDnFTsDszj0AUj+k
Tak3Gmb7uk045nz9Gj1dNkJqfqY14Ej5Ss54W2PjG3qLhsd0E8dx/4Gqm6qdqkP4
Ume5SKqOVxU7CHLaIbAZX9osql3MPzw0pvhMy43/5ZakbV2/rf6Eh8NZ++4YMXX8
UQbcAwD2UHh3bRCymV/D74XnszWLxccoIK98nalZwUBJhYjMJQrOQHRoo2NARupQ
0dx9EisVx60ZlRXyhS1wk+MJFx7UEu6UKPCZh6egh7KM4hki/mdA+KGr9DyZ4Xem
WPEe4qQ9H5NGd8g0PZO9BtPZWdIbcIqUofuxDLD2QMvVNj6G8iM/Iop5PQDjANAz
5WFfth8PyKBmSJDGBouw1ON1EFWPRN2n2p659RwR+Bs2l/kSXDjb/FZ29CxzIUn2
FXQhkVqxsiidYRPJ8s5t8febqJu5I2MoeCqLGppeAxm4N66O9NRZfTE0w3XzKgcU
m6ZDS+lTlsCZsnSn5Ozt3Y3k9K0Ui3cUu83/i57/VxKUuK3Ye6xfm5mKrmxz8815
GM72evLb4VdOpRk02pkx4+hQHlwqp1q1lQ+8N/XRRKywoAw903swLVrRfjh6qiiW
TcKpy5XZmjdACMo8RnHwguroVxr/Dla5/+bX7/+fHCJqINvQXzsEiS0AyIYZJhAR
bRt4vDeQHqhfefQFadbmluIbkBVOX65L9emb+sNiNE+JZ6yGd479xTOt/xF8odeB
P4TvQv5ONg5+AEvst1uORqkhVZlwZHaxKfr3qKwbzUMq1keS+vvpIF/vtZ/22VTs
6qkOK8xA63Oh8G44O+Q6UKjcK34yVgc1Qwzu1STgpexK4M6GMlBpzQZ6tESNtah2
MEUFinoAHONyo/3LBxyjj0II8gPgNlWoLnJgquRygzxleZ/tnwXgfj6HTkjeCLjH
mcDmKENVOiit4AINx4PZb7L+BCH+BhnQ87Bi0B0hl4COjizhwSIdAA5jcs41/wK9
lvahBgGOGX+mc3Z5AFOfr9MHaTqHVV+PU74zXRcGub48Z4hlA9U+ws482ShI56Gy
Gc5Vp54LuqehXJLY8V8sCbITuXm331Jq1H1jPKSWGKrh3BolsjfSnnZ4BNwoOAFd
eN+XTXmKCsPqikBLFFQIf6BkCtds5LBeR1MqxFk3qs7JLPYInS/aRrHvfkDsKFvX
B9by3a4UR/GTFBifI+Gf7lTltxW/Jc824FoxSTQ6/BCL37slaMhH1fnjOmpNEO9y
MMXbb7429TxRJJwtMiIyw3sd8YeyJS5GZbyIwRv0rotTjIfdSJAcucQbUvgg6XJr
FrYzYtpuyoAjPsJvv5v/AAILbCUoR7KwaQ8PFi61J97hZt8IFVQ14dW99WFf7NAk
b1S/NjlNKrsDkSCEsYN1WTJcr9M+N0I6DdiM/Fof3vcI5B42oYxzMwCtXVJhf5LV
9a8w6ENJnvEwqNALSpAo6G21WtcnpuoZKGwg1XNyq8uzj5tyRnwBQhm4Oeo3dhyW
xPfhQmezjwXqBQnRB9CF3PPQp7eB50OU2FFFbEyCM8HklfkdrlFhrxEXsF6aE7yn
+09KlPmAKs23py3vl9SG8cCHT3ZMKUUdEkIOK+xkKq56/W+/OnVdNTL1P5XcR+Ll
ix2OhO87yVR1qIxOwz3Ti6XXGSIEBYJW7j6R2g95+g4/Uq4GsPfnybY9S/PRco80
URmZLskfic2ngc3EgDbPS02Tdh8mjxCPWCjlNpUBQyfCM4/VzJya+2TiLcYB3B6V
puFKgsnKi3Ve1YpZQcazfcCobxH6ag0vxCbl4vbNJBqHu4cOOsjHsb3fD7lY/HB8
kDQbpXs3JfjBo3uf1zbdRd//YAGQNCZ3EUAwmOjt2O5NaY8BQF6Jkws7g1a+f2ED
L9fmXa7NC6T4FzV06FdBjHhSDMtYWqGJQVNCTI94kGzNoMN2fJKFfycFHY8zl01J
JqhiMThX48WOI9N1ZG9HJdOzQjHo1Ne6MyykZyo6durASo4yvOQ5+RVsAcuiJXIh
WW6YFV6EupIFwROIW1TUvBTLzq3v3k934kk9EIKEwabauWLVnhlchIR3s1tGxkJO
lHK9HSTL+y4Y8kkDi2UZQnTmLhebxAH8zuu+JFGrFn4v+8CHkbkgezoRGPl8Mo4m
LijM80vUPWo2dGNNazpUQzD6D48OqcK5KPdh5+aWE5SvJotWUrT+my41jxAa0hN2
GimHdMr/TK2hpUqx7OTDOyhEIFV5EF1EIlG7XIO8KfsiuxxSwCzrvsqcRy5K6Wv+
3uEKNQaAlAUIsbRA0V02UhNYbrwWJC4iex4sZwiVgpYdmxqU0UVXW2+8CFQJ8Yc8
ldv5Uf94W4Jaj3aT+dJDj0JIBIg3+o3XCTjqaXzhCXSZyVdw/cvYGGl3r+ytXpnw
QX1ati8NitVbcq5vQH2PCI6FzDbUc7p609FG0WsN3KyoBfnnTSheM7msXuVEdaTl
hD7WtsvE1001pa+1rqNxoGpUO0uHbs6xQCvVPAaPXK/1400s3vujNx0bAXwRzrdY
jqYJeKT9rs0ilmK67ZrQCgXQcw3XN5IyAv0YjkmCPP4cUG7OBoJcav0hZ1PG9rvX
NxGMw0tmbtdjsb1niOVSimjdBxYZGA8u/wtMGpR95+C3UEvKs74lt2IkOJ1cv18z
89mUTxHBAmwAH+43IvVnzeZ72jM7B0IWRznQy6r29zzeYkakqo3YHY3Z/EtNZ2Zj
5rBaPOZCEy1O4a0TsasnNn02aWYC4waNG49+sC6n0vKziI2f9mclLeT4UhLycn5i
57YaHy7PwDDhC6Wx9uT3ZOgfTqKHCP4AS9gUt++6iCUxdj0Xy3DnW+7gMeFqWWuz
s3PxsIzrq578wbW+mvSIEnh3hX7mm6IJg7wRG6ybYSoY9TGRaGOT3OI6jG894NHM
KWrr20g5Ebu33nyJCwIYt2oN+Wko7VhRAGdJgaAesUof5RV7LJmunCqXsmp/ptIQ
yIM/c9WJleUZuQsdVksHPBdyJ8HDwJKJS+OKwk5m+3Yo9pP1TnvG7/DdY9tgaOK3
JSV7YoqV6Y911jdRcfAc7l159KnKhFVfVdfd0Bqy5T3ytsA1StJqeeGV562AYkl5
DUDYd09zz+8N0b6hnyqymWaVPcmXRoHfIl1NqQkEU2QX3VjLu7HCYp4rz+rUWl4I
8TOqR1G+ouE3cMXtXi7Do18R8sMTwfQS8nDZv2FR0edpuJ1gPYZoNrhN3b1eeBxt
xUx365CN8FDVQ5y3PiUxdIG5CmphzZ8lBgTlT+McKh821j05e2xGrY9irrl5YZx2
KmT/oDfQR1EqWqjUGGjWssubLyZiX2y+Dt7XCtgkRygVVqIVO6oBKlePEhKJdtwO
f1XexTSRI0WGW76p7y6gBzAJHH0G53AQFl6/vwEydnhY7c+hJ4JZGdxfqENVoqQH
okBTQMLr8ws03IoOm+i5dmRQAgUU/j/CidTJsfH43goqZN9EgqM80RIw0DysKsb4
xOJxpqZXNZ9Jr6SvCXGjn4YpbfIIttiRZ5Y6trT0BMcujprTbkLis+ZgNCV9FsOj
eICTA9etF6I4KdKU4Isr/g+fNynraCTb+G6gvpNzDAi5WfGGbDPyyapb8NmJmftP
3X8TO797NTA7BKv1EB2DnEpw7dxzx910sxegI1fskU7P8p0syPN45lV3VGN17OLe
S8oE7eqbGbV3EWOGilwxCHEjQkwokmfo6VOkyoTfezXyezRCbd+4Z1Cmn0qa1A8+
7O0W4ydhrn9Hu/LzVtVlEgmoyHWZsWITFcSVWr+CnXwU6HtN6cQUd1vfdw3cuNP6
zlpbQeGxsYtTzl0iOZRYpOp9kNSsebylCaWtD4wg/gBzy62YlLmDSt9dq0nTCB6X
BhgaKAqDUcH10hI7m5AzCuZCUmi34kLdHxiblMoQBr51+oPddCbg5ujzz9+rXMZo
/pCSOOQ+ibJ4IKh+8Qw5JWiNBszZvET0exWQJD0eqZllVvNGx/487FPSi3BjruVV
M31fsOhNO++lUW7+RZJbOsgomMW9Lueq62XZrW1QTQ7zNEUOy3sH7YDKK9FITF9p
LEuvn8PLtystr+b8kBVvyvsdZk0wFQqduiQMC9kZ329ne14bprxlT8iL2lGODS35
EFmwrz6aZ6m5plYCCHRDnXu+F1hG34OagkuYoFXmYiuYQ/AIOhliJVk1hjGQg5iX
XQDBjpf+8wesxKd0mgmFAkFxbNSVtOh2BNBfdGsv0nlZk7KKVBND4CBxyWAP9Vw6
QRdU5kGbSJoynb0zui+ZoGOgjEPFRfU3WYGd3jWdfIMKdNhqr/4tzXxLUFFScLd4
o0qSYUtNLUkKQOaATcHj+W0efoCYovZLtos8JrAscNfgCabemIywahv2T/fOQTzC
8C1YF003UawTUXHS4hJKXGFOD7KdhFjuKHrpPrIBPV3N5FVln+PQXdQZ2keFO4tT
LIOwRReoCN/ZheErRYxj8G3ca6eahyfaOCZgqlTQWb01pl+FJo4YGwBgLZZNQCPO
rGAkdjOrJ/ZvqdDmqKvrd8Wj6rdbq75lQawWGNOImKe19LxmaLJOE0ZAfDK4NH57
vIVV7WpBMJtLoSRxttUJOFgNdrsTWV+hnzlu0hk7jqQeMZoMHJkzhxs/0TbPz4iq
fcEU2+g+5qoBKUBlUapaUmgm8iPkHkwmU/q5bQri05wW4+pYlFKMYuWQVKJa3UEb
KftOQHtiwl+w+1LBjOHlh/MrZh1pQg4zQiOnWByRsHUNYvF+sopV+6sZAIFGvOEx
a5fW9h8EXREWM3hUDgsj2HTrysMPWwwTW/hYpROQ0y0OONDKzzw+z8I2sJdWVe1f
UK/raiPAFLvl6s7tXgNP44dRdDGZ5GecJ08W5RSGgNR8YZMq6D4/QRAYJwlAqYU5
192KiO2RFl5wY82SMmlR46u9la4uaDNNeoiTagkg+5SZk6wNvKzU3uLlqgXoIe1s
RPZEn3KYOgHCcSY8zWd0J2zzbEBagGxUm84UX0oLT6wYAj2HAbw9wwp5crTf5JCl
1BDzQ9CBiKHTqj6pZy+hYs0khmuEGDDzZ6XzkvLqQdwrSwlM65d/L3BQ8KVCqC5m
LrjbYGfBdhOHJdfRIAW6oxACsYJecb4hgxbDSwazYy9PqpPbDq232o+f3IvWN/co
XQx1MkCQ8QRYR66OU6rF+B3q/c9xtdPYZQQGE3QRxzeN2Brv3zs8+//p/5WAyXOD
vYR4s1s9Uprk1rCd70zrhZg60mL0rIJZTl5AqA893LIV1dx1bqaqspFKrym8D1NV
4vPeWdZMcitPdul35Ab/9wPHCGGVInjWEoz7CI7FXZUCuGw5lYZxgX080jq9DYgL
pRCvlJelobwcnpAoEiagAToIwlHPlvpE1a2TACWBR+y9Wv44oN9dySwCerHnf6b1
+e8loNl1pcsYlidgm4iMhUsuTxlSZ5vC2S8rvCgJxQakKlTxc4tYJSN8YQgHprh3
qDh/e2am2qi98m/FA8W080G6Fp44X1P/PC7pIqb/fVZnXmDpAhClG59j25bLFts5
2Qx9hRbU5GnxqnhHdZlKvpRu/U19wgM0zzbMQs5wFJwGOJc+J/QDtdBlMl3ACqZi
1nvPLAoWJQInuHdSiIp0flY5kA9ufZpg3Hq/KA5HiJW30CATCvky4z/TAHXrhYb7
8sWiuFM1qsqRnUc/CKkayqxN+TMOEfWQuhuy/cT+IK8IBDd6H2Nat3U7AYXzHIOX
2xl3asYHDWmePu1Vz+q4mAlRFI69yH0X1Q4ZkX9wW5LGEpUt7i9tjIS6+MNPk1VO
6RBQAJM4DOxekHZOn9ox+EkfHvrTfK4QVIiFZGj02bU4icyIRr98VtHkK3dDXz8Z
UUDsKBTjTgoID5XoI93uWsemEm8jGz1/7jYIRwL1TLFLAbcsaZaI/Chww8MLTlSi
Qx04GYN9Vxe8o2M3Kks8K8nzIB5EW0ScH4M/bpzxjZPZACHK88MBsNgiYUd/WfIB
hSolIBcKYOI3JvDyiRFKkBWZR6JGAAoDa7yP8pEsFyZfxrm6pHiQqFplwym+cnkV
QPmXzov6I/DCXX0PCFBhTtt5uILEWnRKMDF5xcdji2k+1nRB/VQU6EOCmEqfQvYS
C6fnoWVlDT3SIdHsRv6kAdBEIoNd9ZUCsRbi6vnpAlc6iAGchNqf5SoE2J/q3Fwj
qItlSxHNugO08cKdzDbBJ9seQPqQZVsiK3OxhCYO8KYWr6x3Z0JHFZrzfTGRQiTh
MIEkAamEMqn8Qg9+x2wPvfQObxBE5PqeYeaXRMrWg1kyJ6FTkBp+F/JsHHlEZlK9
npVLeqjcJ3op1qTiYBOJAIhqBGmYctancA4xrKsta4einOBi5D6lNtjPlaYtjvFy
zbInU0fy978sQj0o/2RBoUy2JgUrYoyJkzZ41nZHI2ZSe/yqn1o8JKT5wEEyu9q6
jBphNZiQHmTiNDatGX2CGqNi039pDOiX7row5CGNfA++SuoJMs7rxenaAiq644t6
QvemOHiek5e5ocVEWyda6rk5tKe2umdDGum9iwvsC7HfPrgf05GWlexwA6B6pUlm
OANO/ZCSMWeRO+YMFL6VO+T09l2k/52QIGqaC6PgVK9yIYas62v0kKB0KW1qoeC7
mHzzV5XreTVTxbAHvIAhul9xtHo2Mi9wRLX/VWLeW6bfbmETOJON4nzG9CZkySCQ
6uywLWLhFDhmiHK80nyVr7RpkYaN4rI+btBUffbhdBGHmm7bTD9mOgfRP4UcY/Q4
9X3G1K2GymQe7jfTvjaQJI66UvoPURXmr2aNTzyzCMYFgcW8tSHuaKIhHpu3bRey
uBcmYFKdsY4wsnH0Z0PykUj3/bo9RNMjmqeS/1T57jNAyrelbW6BvcXlIZJLCbVC
ugVnrOpbR3bmI1e64nCAsDjF5mFggU6PAypK6P+9yD4I9Iqv5hSZg/oYy4TG2rtW
UZckZeHZqK0CRhjsFHGzi1m2KvGg+8IvaYWtiEa883X8Ewcf6sqw0ugElBMdjDNd
zeu/qDJk6WcXaYOOHzBRYV03JYRdO/DCM2QWS10/oYarP+S2dEDgAxnVwhjkejCC
N+h4rIT6vwFPo2Nt6EMK14YSjHBQlhoaWztIcdF9VHS+WdyQP3pTTMNQIt540fYl
JlzAMEcDL7LyL5lkFxK+xc4DkDjUadnu+M6pSu821iXk9A7jNTFiK7WbdsyZySyl
tSFwHFQ0PpY3w43LkFdsvotfhezCic81X5ZMqDeZJo8jaoa5eXiC6RWebPURhyGx
XhUbGl5cGj6DfmcyDvtze4FlYd/5gfGWB4qywMcQ3EAibvTyzes4OiD7vF/QFC8W
3T3ojNq1ojje8oEYyaogfuCn+AY8S7ZJEELTQzuONjbgnvcy7OMfR3KdNd2IgVHb
7jl1mDOEap4z34LL9C5vz9XGMILyIkgolk2USQumi6w15IoVsEumu36b6AhX6KMk
HbKB+m7PbQJbbyWHAhF8ReOiXWl0bzyFycl0/VoYW9ZxpirJcduAyIhNhNOT5mKr
/+qdgtz6q7KsT7tgNBuXT8izxUJcR9m8w8dhHWfAgeZwyEolYabATN6giHwDbUf2
e4KDj+rrTIPEdGb3ZPJSgEl/q4TuKqAiCqqOQ/sSR3GrzLcZPAMGV485vCM47FQd
ABOXQ5gwpYg7mkKXxk/ECyPsOrkkQzgwtuhCIRiE3mef+BZzjScEY5mtfhnvRDxG
P581Xj7rL7Z03bfr/R7Mwh2+qnV4HtWI+89f9PXFCiyLDsiFKE45FjpHVN5uK2fk
YFYk6yVtIIyipbP1Apt4ddMLRre/xZnz+MrA9j4iJBWtc1ZGIyEPlZlD5cMorGz6
3ru35Jc0guakPRwcO2Js8mGlnDSGZFDlxDSgybHOeVdldabx5OTeaLW6Z/Ufrj38
RBUmvmOrS7Xia/UjY98d6UxMH7kUZaat/aVXxFjyYouKsE+PWqVDCSDECUxuvJWj
K3qTrhZ2K170Rn23WWgNiZ10ATfMD4ml1nRo2idjsQHhQgWVa7xjP1ZSMXLmIY/S
HhtBNsEXnZoAQwCOsBZf5zpZNMAGQr/Ht5iLujheZZtivoT+eg/AiylEazNh7/2k
IrS4q+Mvm/MJk0Z4VuUyO7FcGyA/Dh7zGTadPsVLJo1UQm3JMRkCD8hmVBr5JYlN
9KdwTG4PAbfkB7+n2iwXhxIPBaEVobBDdpmuSgaS72qwKI0OqmdX8eT/OYHXkjMd
N6E+/4CpPoWpUVrLwaPhmQBMKBV9jYHpeW+/zuoBpYdx0fRUIhVcZxaaRR8xTYTq
3Y7uoSSEJJzt6IsEZB8aDAAyrgKTQ5ioS+HrAKiYTMVwHqDmv/30aEHO1HCJd1sU
1lTvV+67dCricapgHAfNrnlU7ZjZJjdM3GlQispIOQI4NMElZB+hzwOuOcvB4Fuz
5gKOajZDzE2BfL5hBrv1R8QrzQVjG1eg4abwEav0ULEk79pfQsxRLlTXi0Mr1cvd
0sBien9wcwtAPF1h63PcuzpQZPhDds1KRMqb2uK5rX9rhFbUyjVdUTjoJ/37vxEh
yGrq/JR2P1fJXUxphY46qIUjDGSRP7OZI44xXYWRECWzuA6zQU+7T4Iulw+BrJQW
KLmcHlXk17/goBeIP5Bs+xin94UXL/2UmOgZbyJQT248jHypwlPKrdUuEUGNy+AT
NgF/VuLvPiRX5OSnjE2qfJN9iAs3VhRCqcTKFH201d0eRAVeO5NE63AMX8PNn1a9
UWdrsfane8a4UvyXTdr/avjClhJeU3E82X9nWfbQjt2kuSQybBTNJyM4Yy6jLrCy
Pdtyon74cgRj+rJeKwG0G1QaE/pEdDqHpRxG6YKG3S/87qeBAA48dEVyFzqrWSar
GBINLU+ggGW/g/ejW2sfBp7h8ugkKH+w5wNwLSxw6/a7dqOShKpSHuSQ3Yv1m+p2
evSPn5Tvae6MxBevLyvP+g3cWF6Nq1kXP3w9ix1cc+nt1QvrVMZbseq4eoAr1JTz
ION++qNbGYPK5X/y+Lz5JUvg66WZUM1wAga3GOL157cqPimWEsa9+xyxL0xmjPUH
ejg1UItzeG7aXeO5gP7TBVgnkvl8BMEypOIC6JRzLU5ypPkewxTOs9XBs/q04H8u
narV8nS4p7tJQO5XCVblrBai87QEUDT5Gn/FTtq3WJUNZ8kw4gehiG6wmccRsfNT
75CGuRK6BIBS3JpNF9M8JYmc5o9ZxS9FNlDbOB0dOvpBgvUlG/vsvPpnnEUnIYTI
erjIDNPxK0o+CrtYN/0C4K6W5HVsP96K64FlWyH6jOZKgLnEheU5bO3JEzaf0lqd
3fZJ8rL4GQLNKPKAHR5tgbAB5BlfQQwy5NrTjAU7+h7sWsxU8IaAqZ3vG9jHxsjN
1wYDOSSaNLjiKWhzLx1WUdCqHpgKtKW5voI3HNXPOMblCOQZJOXn0Kljn16ZTjM2
iBgKtDJ971fL2BcI5hEIZC1BokrBVNarfOLUjlbSknFrNyN4fNpZ2MHXkF6PDqHc
YM18fNkXiov2HU4byO4qR9Qv9MQ9EOosx7CI8YXWcrWdpNDzjOhlWEwQ+UUP2os0
sDudMImq9I6I987y3ezsvac3DPDLdClv3w4M5Lrtxl/dJWycDCxQ+MwXgn4JBz9r
GTZwH9/Oh8n7eEdM9nENYmxZM7rCuDaAqyJ7TBS6SfupBnZCXYUWyhdRROYgGYrN
uT2Gq5voH9AKs9x7CMmMqDbQlwqT7kZxxAPWE47YFLCAewFByFA7es7rqLvM3EwX
iXjubsIjlwYjDgeN482xztUyYXq2uJCYwafj2eiodp1UjF78XIxP3hKQYZmOYH3j
uCdCSEwq8yYB3dC2Y5fuFrui02RMnm97zhSZ6vjEqU9/rk6vmdaHbfVmoEYqbtm8
HjjpLXjqqcdAP3XAJsjrBIyecmbbr/okiG5s/z+gTTDz+EOr0RY+Cp1+oUaR1CK5
BBBvm6g2EhIyM4JlYMRrjM97wuLvSGL28kf61PwCLk2805/mJttA8cUFHw8J2dXC
v0uAayUKCGIweWS6CRjeYAd7qmGqygvhWJ+NkdE2BXJ7dPmukE08r5ZWikyfBW3p
3rnxyAYyqLoGuO5Ru9audhL5vFieI3j800bfG7UDlhI+QPwrcagXheJZJx6A50Uq
OP0CUb0Rc0momQ5EVjcqs9ZK4lOVYtmcQdkb0tLs9v1iempASSfNiChwbbmIxyuO
MUCn7h2iszJO/WnCIsRlZbkeUl569daKvq5kcio2d3evY7P2Ci5+UkvDqNbLosr/
N5hdx37dRgpzqEr3CCRX5D9tT5gP0OpTbFSQo9rzbwWtKssrwvDLz/2oEpRuZOTB
+SpTCyGASeecjlWsWqmgFsAotMzP/3LNeMKsO7lR+SFw75+S/92KMuvX0f2IAJ2M
etTbskcIg5jMB8KiT3srcsdRPMhMNU9N9EHfgX1yKkmHXPR9A714ruiT6qMXrHLh
bDyzmntH4xsa8DUkwE14VQEH1e6QByLoB4M7+byC0qugX8wDysxJ2gwqHsWZTZct
vulcZx6zMjgtntA9UxemU6NgOKJ4rbXMS514M53gA+/upmfy3Yrw3XZPdfh/UUJp
+xhhI9WEOfY1ZYLXkDnVT8Y/4EaMRi7hYYIJBp+bjtGWlzzXov1Z68tbZghYuwq/
Gr4QQS2mxpmZ8UelGQmUoo01Mn5uw80MeN3AF+YCApSTig5qV2pC75MjiXSQafUX
dDVyg1tCjYa7P9AHoJw4TgLGkPK7nZKP++KowqCOal0b0WpEMPp5wvl3xRMcLrQA
Thkv4njC92DRdf4IswpLgiTZ+N/aBmVlKfaW8NDxcGjk/dw5upMgiK5qPtz29d/l
cNAea9G/xI6+s5c30nVHoSl4mTaQ1Z9jJ92vWLZKSCNzg9sa8VhPw2z4lng0Jy8c
1D9Lj4aB9R8eGx/joaafLAyHCDef2tmACntGhgv4GStVS3HCz20D8eCIN1Nt+Jls
BMvsCyY1LpJIDqpLZRwfxJ076Z+zJkmVG2fwrJ9WnxbaiHvRAmJ2FCyKh1EelBnc
K7EJHqQWx97fzLUSCSAhFgRilKdN4J7jpSZAxZ7rmxr4ovFzVK0f1UIrAwiKXpO2
MbKkwsLy1trTNvlJwoVkgcxrUzm9t0jkuHS3JxmmPqm5ZyppSGK84lrNBqEjsqcI
R54TMzyKh74NJXl/JLSiqXYooOjeyyB8HPW6geWom9+dWJSM+IOtAw4Yfm1yARUf
sHPA7YdrFyj+JazzkeDIdk9kMpENLAvdGSruiDTfkmH2jzWU7h0aLQU00/TaXFdT
yHx0pZ9D2l3FCy9ygB9CYkoOYMXhq/ADDg2pmrDpXVWzrjM/u3ApwOOJ9GNsLETT
v+FZpD3SMmwkgSm5drGlgSGV5DnUOPA4gLOH3KqG3/itGXG9320HHK80R8fOrDAj
VB5UypHbW9Ic3BFnfu/dQT4MRsrywkh0/zNlVQgfBCRO54YMyF0Wi56KuD9/IRns
n6dB8Oh21LYQ3PTzVDa5wq0ztgNzKH3TSHUx3iQsIILWFKMU745Xl85gaUJE+ijy
jwF9TQl6IK7LsUhh3uLPev1DgvS7//hxYQ/roK6tvm5wmK2Dh7YkxulcEfqcmoKm
zdcOxsn62+IYgAilUy3WbB783jx4W/2REdzvlTvZKqdnSnPY0YEaH3velt8vVYye
zhg8DKGFEk91SEcFPBIIiWXraHZ3nF3J83VjbYjBjFEJSdNo6J6UKz4zH9mdEnHj
mnJKYZFsMIgkbgtrNAHP2kd11sDUEsy1f1VHwj2TXGK8ZY2vAMQkcCA0qIF0tm8S
6Ok2HuEPstaVbzMiJhNQzHkWJR65gGnFjZlt6677iJuJ+15S50ttaf8OJOuPf99g
Im8K9TFT8r06GrwUlNmKuT0B20thLAfc24MOKR1hYU2amrVtS4q6a2RupY+PY9N8
hw3i5rWEiKvrE8xRv/rDzdV7/3QEUNzRDVFz8UKxLll+tUgGji1DqAo0GzeiCpgN
a3c8Us6XcWSjE9Gi8fNsQh9l/5sJoQBqyCwC1VV9t+fwajIHOW3dPBkFiXLgPA6z
XoTl7b40FOsHOjsddHJtmnAB+sYAaZBYWXcGF55jOclW/qSzeorK9pydnP3IsptZ
LFvuvqc0T0olnLCALE72W/y06t7EI1gnXZwDnqiEfKXF1yWThWqTs+6i575hD5Zz
TzsbYJrjcqqK1rwq9FY0OHrbPqSr2VArS5HB/K9v7+09mbEItmE88ecJBJhZuFMr
15AIENxJ7wvmYWnrOkuafUt3RhZZjIRIMQcm1cmyosCane641k3MD5AxolyIzJYy
zU4+/N2jEy1/SwRWGm/sj35v4Fwm6pPyz1BwCdXAHjkIMw6rRH12FNszk6+50cct
HhOsEzMKmfx6HTJbvUfh88M3CK0fy5IFd+zAYVLAI60kyUzDUOxsptKGa3TU/84y
LjA6uGOClZdILReSNmd784n4PLIj3ZTFgF84bDc5gLUosjjgPyC/8MYtV8vH7s2N
ol721R4ye/BliloFeQk49Cm4Y3XyPWLmHwmqaJ+uJcewNRRARb/zZ6VVWtRBq57g
D9pf+RIrFhVRhME7v2++99GbUUZJexsNXagiWElcUoxASxJ1w/SEYELIp1aLP9bT
+f1ERzXUUUycphCdP7Z4BChrKUX3yeUQdsIKD143uUGbCA0g6Uj5FexqfMVStW1m
3yN1flonwSOS0iVryR7xG3McqQCI39Oye5rhYPPAOb4TeNTizthDKZWx7rgjPkkL
KWFjS9oQgKkYWaUXPrkxsOCKW4zofgp8mY32THWhvPylDEH/eq4YRVT3DF2uHZsG
Q6YpX/FEL3Jf4ase8tZUoU7frJ+qibBUpNVZVweEYir+/Omm7frtS/1K1f51q9zA
SoXDpyWC+lVxbHtSTAQJ/bEP1Vq/Du28CJyvVRAzFlvbVekMGYK1DP82QMr+6Y+Q
nsajOcwP1OTS9poXkXnKwWaMEbcEXMPIA3hpOitg5tXKdOqaJ9qEsKqBMaVY/aE9
rE/Qpk+5MUbut1rhU0das7UD7t8CZOe5ezyAx2sKVpDubMcWioYewYICroAV29NE
EBFkHChecZU56o+KZduT7A8/wSk90Ek45aofRFhSdScDV98mqtm5rLm1FIFmYQ5j
w5avXNr8qjJSBv2tDHsaNzC6AJery78IZ2numyfXi0P0PYRnPkwIX8LK2rFt78t2
WykyvftgLegZsD0VpVAduBKgRk5WaJNm1/QZGt/UkWu6t6SHHFrQTIu5fjsrXJ1f
UmUK6GbKjLzjl6DbfzeKmPCXtyfrKvR5WHLQIudESgGGAGrwqoXysla8wVx8Q/oG
B+0ZXCmBDQ6FrIc8Go0VEsGwXDcRKxqBzr2mSBQ3ONO2ezb5ONPBz5xw1vy3EA30
CPL9GERMXqFObiDguxhWP/BsvB1wBdiwLIUV4KawjC1ktuNYmf5DR2E6yauyijYk
IVekIUooN6ExR/+zGBKmoK8pe2BMmtwyfqYMH/LKyjcvWfbWP5L2XJ8ynamkP4Cy
udWatMb8OoOGtGiFdQJ2Ryupv4UZgHmWfkScUEV1wHihD+Wlnb9pxWAfVQmb7s2R
JhV2buCrEpO6/da4/xIpFFLELpHvmt6OPg2qExQPH1IKoGYuk1i1lYwCIt7tBDl3
1GBCEqRtX8ejLFcI1UzMfN72gqWe0CjYt8/WVmgVEm4+sSGKSc95o+n7DSUwiWgP
f5JguavMvUZKhkU3MDbuVT98wym4KcDEXCJ0Xv8HLC/gqRsiichzIwtt+QfpVcdL
ln4BndX/79aNsdmjTNC0zuZdS5hPpnk1nJMmBAYklFclyhJNRG0dqLErIaFPWYTR
6xvRtx6YaZ2Ne4VcpJv2jQE6uTEvBbrFBRhVAFg8kEDnB2QFX5Rt6aJjoXXvP41U
IR8R8oWsYchTwLshoWjdKxgSOUzPwnWKUC3yMRTM51iKr9GoJLyFjjhjVGL+YW23
ycVdpwl9dJuwNCvZ8nZDRLhshzSab05uQKXIlaxwI5SKjh34gWxdp79cB5OFw4nr
qs/6kuuuxl5NRn08YYLc/q37KMooFtHrLQ+y4NnN/l22z1+nWe78GPrdhjfN5ocm
mrfZxkhk8dEWth5JzjskL/jGiUlYChXnvdfL4d2TM4jqmOyQmW69Pxl5RbZ1RROZ
hu9OZL69R/nbNUBNnhXZ3OnoPWPdUStdIgnvxhTdlFrxCuGuZ+XKgBsp9Xlj3jMo
jHnMn6MOk1tmAlprGxrhxTvAfAI8r6OvfOctr3X4vsk0OQBbdf3jB7HuE19KFc8p
Oh3c0vSpXS1ih8Gd4FwK0qYjXQiPSozR/J8r0qVK9WZMybM0bbVSHIjAzjnP60gj
6NtJgL8twOS7ka85MZzEEA2KBpzlUE09ddkiQUXvlectTfjyVyPKxBVC8HbN1eqV
W3vPvzPcm+CiXgOYs26X9PMoUQPlcqpN0YlXPY8CSD1RupoLtn487nnXELK6Z4CD
CqoBWjaHf0WAt8HES3Hb77qNE1mQ0fCK0CgVQcFhKF48JI307SeXXZcHITrQTrCO
1lEpy0B+nETIC/XqgjXbCTRytq1pgs1lLxwoQsuQuaiUkN1VczDamaetUGJTvEIp
M57qPuRNa6oaLWTanGlSGWYmD6P5mgo6/2V88Gs0kJrAnWoyY5oC8WPG/55eG+PV
PTitpHZfgD+BJZ9301SwT9LbZ5lV1edZdtsrMUY8pAjA1Fu2lnqIE+CxnQBqvDAk
vRufKsJqeKDDq/NaIhXE+W//rCrv+pOc69kkensxl1pRa8lJY0s1ocxXL5N3hhuE
CuIFrbnZWCfwtdkpXJVCDfPiqqoy2yEAXGOFHW4jhDY0ifNR9SLKomTw8Py8tnl4
c/sycV710n/6LEDew5Rb8zZvisYPzVUsnph39FwqBEt8jSsgg2b4eZk4Dq/Z8i1i
zFte4rGatUJOmbXeh047tupJ5NvHE03txyQ7vRQqDsGua9WUH9AZa2XJkcTIMy0t
wog6VnJMjJzYioLRsAsFcmKlLnQ7HJIAP2ZJmXEkds8gqATQa1c6nTw1d0NugL77
6L3U5ln+ZFUPo3+wUmEsHBfKca6vNRE/2+oNGfBA6TtiqNT+KmKHLbLcRp1+bQnH
w2klzRKBB91AdwzkdXvEeBZJuLMs/YTeiMvSmvhual8CvvGBb2AJaJC5GHdYTsnn
Z2fS5iaYxNXfJ61kxA9Jk7S8+G3TY7wPQWrQON3OBlx8LTbTrk/qfMRDJrL89F+R
IRMWo8PqMMwZYxs3E+LzBP0hDhxIo/EcOklEMK+GqC8gbvBbgUvHR1bPRORIbjCG
eWBuSlY/P1Tu3cvuE6HLkjwZP3EHmTbD+iDBn9rNTlTdGUBx7+e447LjwzWRwv01
yA9uWhKmttpIkKHXEJ+WWCPAf1zhj1TnXyKo9fyLKV88oqtyXW231qr9kYatajfh
h/jglU0pnjInP5uL/rKRN3HxQDhrQCLEE48sFTr3t7yqw18VGHa5jDwShx8XwWfB
W066/wUl9FmGbggWDMOLhbKrc85n68CCaROwBevAyl+HUd3YuMwMsFui6QyyHhNO
fuEJKKQolugB6KF+DVeCeDPxU8W5VDrN8qzzSyL9yqPM8LFyxlqlkIamWAZidTim
llEt1JIgXEWlxbyRN2qjF/lt18jzzqOoeYftPtXwf0fIsDE5igyzulhFdwJ1Rkqw
alCMGlbNkidFvGNM9ba7+LGYZueq58/2fGqNLdFgNpkVB1QylmSwAV0IHNnwnEUP
Yo0a8mBu3JGMB2zsE2OXmXB5PrlEXMgCgq97yQhqwpYJgkq6CYQ4zcicjLoxME9V
XiMdlpY/X3wU9c/rWYrTwfgoEglj2oLngV1Mg4dNBNCm8qDRjAVIC6XDradfjVVY
Rc4VUbKLIKvG9pp+bpj/4chIgvdZjAR19kubIJxBwo45acoS7hqEhlq/8dIUryQN
venDoM5YpBIKC/SETQhQCHXyAKGIBpse4Hc+s3BUdq6ASjpU1djFpkx1WbTVz4U0
Tiw84nzxKmRhwqPS6fAivhDTAJAbASsZgSs7Kt6lSNmSjPuGvmaAjZ7gj2FiBl7a
rsvNeqwwA8mxbsOxIpJdLBTT2vCGF2qJ24ioHZf9xJJdzbl2JNz+ZKk98pOCVfvb
omLoSXwhcY5SHVi1Uqfm2WgwLaw2PiHoxTJMS0reJYGnzZhtr1L7TfwrTuNAXeDJ
wKeXRw84fWU0noPLl1Ed/Q==
`protect END_PROTECTED
