`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gdO5zWbkeReQ+9Ab4Wo8nvDev8TKqmDptUZhLinqaf8qcWOgzuLqWfQ40AkiF+WJ
/WJygZkrS8GQ0mkrOFl4W2HYpIuwkMHs9Wsjen1sQPHe84av4LyUMXrNfBQtY+Hj
6Y0BYiZN8U9hci2QXofF8yKCreWTc4dDdI4FbJsnQId1zKSJdHwL8L87z4p5od0Q
49zFRSTrzR5pJ+gvV6Y5yS9Re8eL8Q82UGunYA94dLSZBr09t0HH8a8ZlE05YJU6
ek4VHQgjCF5DQhhHuzUPx6plzebnYhYDnATOayyzyopstirFjj6rWzeDB/QgNqLo
VqSiiooJ7Wn5Pa3N+5IoRw==
`protect END_PROTECTED
