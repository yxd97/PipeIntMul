`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5nWSEAMAERzK5o2VFQgjLBBoPFTFh3gS89DIrHkGsYIbR2lbgFGvWbnjT1MK6Lk
EwedEaqMxc+yxhop3lnmRdja+aFNxBzFJKbfUe4ZijJc+yyKyN+trEAclVow+epX
KRCwlJidgMPoZAo5272lx5hf7zUFJ+OSdegiTkhhw3CCaceQwFoMbsUE8gCMyNxB
ieGqOuzLxw8cu9+/MeKe3Un8PPrdaiRBYhXX59zvtoP/57PTdKoFTniddju7SfEl
Ty0t+EtdDSKw7l2LGwjU9bS/KUevAocA1caME0aXi3obWXzbITGyXV+Qcoyk7K4Q
kOTfBnvQdLyGtoB0ODWO6g==
`protect END_PROTECTED
