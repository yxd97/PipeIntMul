`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
suk1Q0KlGqm170blctPeztcLeZs8fSJdrjxQEq1h/DEozv0TSQRRFIDNetM2iSZs
lqQe5CEYxTcmfGzx59jSCqTAwkS4+hdgiaopEulUfPrQLS+X8Q8YiYoKQ3w++CRs
9S8EIk1EAQzaqmQZFR7bMIJKvMUryEAeIGrU4eUKlo/uYkLp1+gLy1+bBojug6Ay
fO+/F1Agep4z77PfH9bQvb4i0nKXbYV59TSTsTKl3zUwkIZNdTi/RwQEuz66sKjs
B9KOhpKPCQZxk9hMo4aPgJjZfZt49LIjvm3pXGtGaE58bnk6idPYcN/k1JLH0J7V
19ZpGC84gwrxQoB/wYDfdwTkOI9ZYiQbMiGLkkZ3x2gRbDNvLECiqDZcTZY+2tkN
`protect END_PROTECTED
