`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0cVwj7UgDMtljdMlSw6IWFVWt8BBScktl41iTbCTAzeWCggSRTcmcTg3Ch/US91m
Quv/7LB9JLWTtaCeVbIZkPctmHCjCQU7pfEMU2wy7FxCBIvzHxC5+Pmef8M4A6wj
o4zros69aNQoJBeQxXpaSZYsa9VuRiirDdq9k+AmyRzNa58pkenQm9R5wews6/Vh
Bd2sDLy7M/PBurKLpb0FNWxllNSfffIHj6JBV1X68EeZW9sCVUX8v790bO3T/VAA
auACOGzYnN+JfU+5nuLH6w==
`protect END_PROTECTED
