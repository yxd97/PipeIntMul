`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8PIGvCd2FmI76cnaePLSWkHe2efyEU8AbfUzkGZPFsPeoB5f+HkxwUoLd+xkZ0aw
48cq0Ro/J2iDtEVb6ZdyIcwCsljAjsOeSj2XeeviHC0tzFbydObjRZPcUed/N/eJ
McD7DJ33tA7IvjYM+XGOy/JVp1roB2IgQ+oW9IbcRjpl3WEiZv7CcB4HOwpyhwM8
QtHJnRbcdA6mFRyo4Yrn1xrE7f/stKO5r5Heaa9C7XP16S+DBkA5mDF3fX+uD1G1
wuK8u/n0ecp1FIgCvrSKGgoSrxtyepCIwfdJmM5c4gEdrTBEOCtJz+ca/CkJ4JXp
qfMdwfoO77JXnsGhm3Mgt5nz6OucwWM1k1yoI8K8w69yFrBXRF76/YOpvrcWVT8y
BJvBDXc+yEkKeOruW8sJNXbOSBLW/p4+XpSyGa/mKh1R/f8Y57S3fCyXyw/7Hc4d
PXhuCUuzKN1yU7AYbahL+NhIFJFNd2M3MTV+UlbkBWvR7/2WWkIpvKZIGFYuLse/
ZLzy/NO/QORIndtdKohMgF+GfbXrEU0VKvspguHdk4Juz4joV0e1Gig0V5CWgI6V
W57THOtlqpscItC5D6wd3XhgcXhBL8sKfKejKNDof7ZaLpYHlUoBa5HYiao8soCH
WTKDzQ4DAn5qJYzdJ7L0e3XpIYntNTU/0/tKHn5mSNLAzJW8llcr+DJbcILGslm/
3dWwgi142nr+q8XyXNBlpCk0nhThC2Bh6v4pIZJLPAJXFf4LEGeRI+ldkZVcimEB
nCZUjvZe5l7uWWr/aIYvQ3RgPHnZvNyUZfonXNuDljMRWV2Qfg5b8GfUUH8u2MP8
9eAqyiXDiIwh5wUFsJrstGgT1OIZDDkl2WvrQU3ReKMzuWHIyG25PXhM3rZs6aqE
lGtPKOSwZmO0d/YM6zChspmiUgVqCg//cCBWJEYGiy9o03QsJyC8K9u0v035FJuC
QvP7XK2r4s0h2P5mhWQArCVYy3JXnGThtl0DL0s+9DfSRtk5wpp7PfSt7oYlLudM
OwGPYSSv4gKo4D5/P/KWLABy6r2ZasJ5gQXjqe44MS+3YykDPmdoHi7TbQzSbx/e
pd1FBJsgr1tmMllpC+PiBuTy/J35e/MxOErimJT/U5L0KFMPQANqQ3EIgqIu7Rtm
g496waWk8LNxH+jOhxmD6Lr0nZjaVFokPYOHpaRMdfgJNVyCKbES8bcy52v8tyuj
PHs0vIljG4awvSpiLe8ak2GB7q0gB7rXFnKu1qNl0ZDoMwWQX/ZOdpUko8VaI/Tv
Cy/tCuz4dw48zhH5Y8ZIcEpAwdrWe1DmBnahRZN9k5EXuzebOSHuPxzAMf36Vv3v
Min/sKR0PEOHnCflIiVGkqHlBKf0z0ZH6H8g6Tw83SNYfvYdne1rkEk1fj2/ZtE7
bK/dOAfMoo1r9T2ZD0M9AUYjzARoMU4N9iU+zDW8W9ByEwsL6WxbG2dul+q3yt6f
GTXcxLpRZAeP4uT366p/XgPSBY4fzONBaPsDMleAPxMV9T0Jk2jGJVP2T6fXk/2E
0EQuPSmXSUN2x2gyhJvcwA0jNKxgWHsf0LOJ2OvYGbIoEvalEpqN2J5i5wuhBjSc
eehEr+UWOVRYl2ictvjnq//jmCsRPPJdtFh0HHeyumYb0h7ilNhXnkTOxuOC5Glm
ezdYpzex9E+i2LHfc4t2QWsxT9AMyERW5cTS59HuAfukvhGr2NE+ZVDuOUd5nw3L
8DIiF4+KkgxU0t06Dde6sG2kfH1HwN1MIWA88Idi1O1tnkOaG7RSLU0Oh1AhDl94
4PLTNjHie/J09Rhaj/JAa0NxIN3nzDtNl9PloRULGM6Mwb4n9z7NXNtvY4Mbv2ik
iyzQWMlu+FD85JjrvIi2cvfaRm4ObES2SdhvRQfnSzQRCSr1TOt/bzQNc3bOYZMc
jdpVZ5pwzcy4GMbIQaUNpvHznOirk6QbGGVsSrJAIi1fm3Om8dkdw1sy7KCXStwY
nmGzCIvhysf1jYUQe9RXrbVX7ag2GOapnTO9SqkIj4jzOYx37nzECsYWuwIoVL8t
`protect END_PROTECTED
