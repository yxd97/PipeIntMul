`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbf+LJ2ZlQCKB88Pawp6jd/6J2pCywl/r/S0jrKOp4aB2DNbtxw2MJoDb42qWehM
xP8WCDVeJWbQpmHu8Vnt3Qn8elxgJEiR2XjvTqlo0DyLNZboUe1zjQhVIpLTAnVa
Cv8gtrPrxSvq8sxuw7Mq2vvcizShvPaq8riLJp9t+BlxlNCoaVAn51RY3EKZX2F5
R19QH6wiMkjZHUJMVLcerfWKs5vfVAveNeXY+HB91w1c0mLG921JA5uajCaz+1NP
PGUmawLXZveQ5ekgpOM3Onur7q6PdhbJKpfif+tENdCt4LE9mYrTsCNYGcMLPM9q
M5XyPl/zgLmeYYFvsJy0mgsHi2X4wTgLYUWIRsEoN1+e2kctAzVxN5CD1KbIzNsR
htxswhUl2KG5ulBaL+1/2WckSP1KLfYAb3I5nVJKo793/6l1kYnYHZmyq0nDzgl7
KHlAkJto0jDPGqEuGEf3eBZYHnvLoOLKsbGloCkIjSSRX07NlZGaIHZqiVMzkNfG
oBe5REbWiaoi68NHGH143LVrV5SQ95aufiIRHHePvVzVpk/GNCyIXeol9glbkTs4
qSHTDeuc6R19tyWOWRgyZ3YfA5N5fqtpf4Fbd8GTXZ/0eCj+y0L84wc1PjPHo4lX
m0XuaOGxuxjdv8RK2CjY8d0NdwYLlxIrficBF3EPCTY=
`protect END_PROTECTED
