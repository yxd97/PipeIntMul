`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/H2NYqiQaDRDlW0KGYY1Qn/4jsMu60ZRf9ipBALw6sIxCC/AhclJCM2DMgk6Vi37
lqv87oxNmCTTIsjLyUqn9equNYavzm/1lTFWgs6Uum46zmOf+6eogCLjTwndUuR7
SYe8XHpwXXNq8Nj6OH4DSsGphIqNr6D275owZvoPRp9SOcQwUG5+GvWye+YqumPh
EoKRnyxeChi9YxFbVz6WIUGHZf2guWxRlItSBodq5JNWsxNSaBkZT4wHl4k9grp4
tPE5KedmZ2DNrxWhqIPPnOF5H0EYiH5tt6HLIJqTbILimqVBaoKGBgkN7Izaglpt
MXqGyN+tAYyxY/itmDG/CnwpiYEUJmVDB+bwvGTh0UOjl2szIfUybe5zW2+Shdec
xlHihr7S93O4ScVQrxX0cM5parEfOtqSm83v8Wagb127Ecdmn6+bh5Sd/csw5jPd
st1SKsaVs5MU5OJKkfw0OijnoI/hRVpq6ou3wmY7oiD97OLqGiAMeWQEfz9c2y5H
m7B8t0Y6NcS/qflh7RiqJS4JNR5zQ4mNDu73qq25BDb/5PYd01WjGsE+FTjMP70p
eCuhnIeFruYmLxy8GMDIRSk4y2PkJevw9X1IkSy1SdJ5Pp6wtQuLFDnTCtH3amda
luxKD8CobW92U0f09ISun3Gj+fV7GROyXqgDLxp71tnLdQu+IG+65MCQ41ty5I3m
jpIt4LuhBX0PUFU/gFH2C0jZ5CEg0XEM4WDh6aFBWuae9sk4xYKF8DcQl1QcbD12
5IuLoflZqoIaovqhAvgwMpYRhziLGaXow8HGTc0xgcn1rgDLKfpCDVIvAYXmH0pq
SBS1ZG73O0Pe33AVyx6ro38HB1NFfpFc537sKHrP2IZwUeT7EvAOPvYIyDwdhSZJ
36SbcZ8p+ea5iFaK2SWiCclTxRsTySb0BBAVPk5trvIPXDomd91uCljKM8Ltvxmb
yq3LI8QS8t4SmDPKIXMk/goGGoh9RZgV93QlvpMWjhQY+JrGQ7evZmTXoSLtWImP
4orAom1/MQ9/lKgxXCksgemLcfBILog773En6mkNhFwJLCchcGG2hNwP1cWJJ0rg
VaYuWkbts8jJRqDv4eQK/beEQPX0YxVCBJah5P2Wr9WvnBPWWCbegGt2lzaF3A/q
eC1g01gNhgp47BowyrxmFOdEGdVrL5BHxsLIyMX/oPbcL+D9l3zjgGEg8UCcBED9
iCjsTN9YXLf6Wtn+jW2N3GkHgj4m8iZDt2StAS8f/Lzx+8wmVOXy/yKytTc0hAWc
Og1CHn101Fjpx8I7qe+Ylid+q+1oahxs3vnScMkZkWxBbyCNO8J/EGwYW4ySB2X5
RHL8qJFk4r9ry0C7jPpW8jOFLKIU9T7VvfCtVwEiK06KR/OaEklA9YR4bNNkPzkB
R3TOFvGOzMI4RyM+QsLesUjVksw2+3Ur1Q8sOg8KXgI3IKykEeXADtVmAokHQZh/
iorEkD2B1WILKjfS7EdoIw0olKpwyeclVnzV9HWTYSmNBoUWdfMYbgKwCYgqbHQ5
LGT+qU+cnu4cLQ9qFTJ+8OmA6RTEnErfoDqs4b//6xBssV3LCK+TNSRlc+q/iQeT
iaxml8SPqFh5aMF+Kx+nNeqC37ZZq2nTZbIP7L0N7aV9lMCR8fTEgpGGiK75gVFO
Md1vA8BtdfjOh1wz74xq5UR/TUEeCSuNVMh+UtkyM854Y0bOTUrf9cYXHEhtZD8C
wTWEds3a9BqtxGGMRA6OPlHJV3v8fmlVY6qr9F1tpQTicKGNjkCjHJlDnoC7Q3wz
Fh2l8iNxYCiKSZ7/SwpZkF91pMbupg0KvwCOMrZ5pwCYSFg6VflJy4kq5CI954uB
oFQLxtOFV0SkpYURwhLI81f2cIXRQEIRY2a8HpBpOXXGI/Y7CRAMHv64CFOWYWrE
6h+fOSMFVWSqAasxIC8n1cYQ06Ny9UmugUb7w88Xo8KsYR6iTh3PbT9Y4PqovUy8
6FQGiRGy4EmaH+u1JjzzdD7lzao0SKQ56RUrhWpF1TYxhp/KAE31k+Zxqm7UqXQi
e4tPhylYjR8Gha/fF3WYP4pQ7+qQt67mhELCoSDVM0bJG0YdUv9t6gyy43zST9tr
s3MafdQfbRokoeEobukNE6eH+63yGMyR9P7uJA/rUM7NgSlJ8DRxjwTwmRN+WYG5
3ZCZPD+BMmbqg18pH8rdiI3qiDfBFcrYM18T/z1u1TcWK5q8XFQccDsByIiaypS8
YOEy2O44YvdZD6RIj7eQJ5eJOef4LZsMktNlbzOLBGAkl8/ScSDYci2yrN/6TypB
`protect END_PROTECTED
