`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NkZIPQcGhPU/5mtNZxZGE4eCxHK6ZmzPbkUgXuRFATabVq+2MUQkm7639OX/bKx4
dw7mf3LtFoO7TtElznl9JcM2DkWVbVpifF7hsYWtOKrHTwBEgw7tSo9phQDKhcfN
1ruDCWHbWRMfBFgW5qkZIIkQMmwJ2B31r1mRQWRRvDzOlqRW7FOr6u/qeezAY9ZR
8GHYmL4Ka4ELDWlv0/rj+hDLh7HOndBGeZV+L7T9W+1AtdaZlwK7himZ9SlU2Cim
A2ofL44zNppIXLBAHvwKduLu/eFFCPMTFC96jt2EOQfrehpu0XHBgWFwHrQmfeBN
InDXvXL1KPQvC1djKNcXcg==
`protect END_PROTECTED
