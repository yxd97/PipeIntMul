`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gSxrEBaydIEGhsL/G/QXy3fKGQzCuAwqi7Vj/9Q3Tw8je/VNAn6abG4ad7tnq42h
R/cIF32ZcquW5HA2xF6uzuvAPEb21F4gW/W9eyXMdvJxfNeiYhSz9HTuUfeZfxio
PjGExRQGumFWq9zpQ4s/6PsIQ/GjLjWtSjdm1gxisvXcjzVPJiTBT23PqkTVn4eP
XPZSlAh4zXfbNcdVyoguV53/A6ZbPUsRgllSe/FvmXbEKfMNXTRM2Y5qGaxIR7XG
Q2TBI2byhdQtSmbKMPXG/o+3u+hgaH+N3ouY2EBgY4x0FQRZeYUJE2QUmD7ohk5/
njAoHgVvTTMEttiF1p7obvXHtMjQmJ/04uLNst+aMmr6EFG4okPhcrP6+OX7qR+Q
YNdmYNGvAf0P9O+lIJDyYyNokqqF5xuwnl1lu3gHzOUH8NyE47HFAyedtPhNajPm
BV9t4oO8ta2ofdoM1ViEtdx0QQFlJSmCWyD7qitqznYSwEi7SusXUnd3aDlwIDoT
`protect END_PROTECTED
