`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1fup/BU72OUQKBhncThFP1WEUMDoED5mpo7GZWiMAw2xz+1+BEILaAiYANapCR0
wlvf4KpQvqfH69GwylezDIw+NbBQNvEU+izWSXyTW5k5SEFsm5IBf6D9ProBD11H
uAAr1etq9UkoLl47dIXpEYtpqrHm25Tb9M6kO/3jOdTOEuWIuQ97coUUht2JSpZh
l5kwp2Z4UutNPEYyzdiCQ+qgWkPrdzql9Z8usCURI5IhwCIkXgGErOZDE9hbfKCQ
e0N2o3j5YjpgDjX3uJZGMUGbwyNhhAZPP6XCnZruujgIvJfQmLugNxeWDhpBhrYK
LmOUoB0F48jQ7s+A4s1IFP6vDJVBMrlQ3GZulhXd8Z4KFYxX9RIOOk7AvKfaJ+J0
5LZfuSGDospyF5PClF7ikF5Sg0d3eKvcn6Qk9qEtgqlPwPsb2K1Q/TES3GcatNdq
1mtcndE9KJrTcwiiTmnftVGiqelS1IhYFki//AB8PadKvXtTlgJYCTlwFrCTupRK
LFU8e6GrcAMgj3S+sl16ig2L4gB8FYBRzxilOAbenfzP32k5iUPubUJsk9ekAI9A
+s3ER+upKSS+/YNy6oyQYOXL/WMkCbbZA3NGuyMf2tweWUwwTdbovk5XhG9ldrTH
cR6lHjo57sUHKsHt7/WhIaXJv3+v+KJCo4LUD6nRQLeysSAZFsaAkSFc7xgU0Epu
GZA1GcXstHreSlgWbPrDMFkuYeTCynDmrz8u1SdgLyapD9iNClCfM/0PssfD9H63
0kRhYCYVgTBxYVpYFEGkny107GLDraouUao1na3E46aIaKGHzv9dJryzo3vLip7G
6yZAq0eT7JudFjuKL/vXoLqgY9DOaSr/iJZRhetbBjduqyOx6pSWkIRTLn+AIjkc
hqeQ0Cejk97NIbIWXidgrIGNWgImug9ZJWleNBoTk7MFGChLluDzdE7VcOw9XXjV
i3L0NeYfpq44pZ9q2yDw1G1gyu6HLKmcDwgUhbDGeEWGT/ZCTijBxzUrZ5MFdmI5
slSmF6tfsi7Ve8f5VaEAd9psJnIt8zwkMQAKxgmyVVrNTzHIflVw8KhPA4NUVA+F
8XzMM5h4nEBXI4059uw0Px7nQ/Q7lNM3OCBg7sZ4KfIvkJZ5IUd1Ql3dY2Ff7lqF
fVyVUdTgA++xspRD7aFfDgprpYcEmEoJFbsJVlzjs4f3YikOPDU7J3ZvGL1BbkST
gJcgw3nOqVZWB7Kb6uopc2v6fQ20Jgkvb43GtShn8hPbza/ljVlycX3i5YqVxt5n
MmxrOakmaWgx9UA6YEr3MiDXFQhiJq0UdOqfI8RclS1ckb49Vpa8byXc0fPBZzY1
p+4PHMdjxZxYqC0rCT4OXBNOipQaUxdfp8OO9uT6oNwbO1b4q4kAIJb9Z7M8Anza
V3RoM2onVsxKBbNCUBq+DoUV710LnGFWEsr2CxcYIdJLlceOqLJTFrSLdeBH3wJE
AswZ+DuDlhpHjKSrWlvl46U9FwGiRo9xyp9Wsi15aDB+wSiEq/6hapn5uf0s7D2C
r0eikTcdwbSu9iuiEiEqDPY6W1ykFAXwFUv5dGsHypjOyq/FJJlAEVitmsGwypyr
dpKhTJco0ZEV9ubokWfFw3c36HnZObGsn5Km0nfASjsmyWhdGAh8yvDE+hU5djRH
us2l5KLBag4TxV9cTBTuxRk22sV9HQqY+65gj3QW4Esz2gRaJ6q/Col/7zwJYMD/
2wCSQyRgug55Ae4Ug5YvC2Kg+nAetGqknUG6UYTFGuURSYo5HQIU461C8kXEiAdt
7xOsOoOBmlH/+6T0OBmmhiXh8+EcXIfTz3QdSJg25FB9Vkdf0qLJINAh1Y2DwucG
mc5RBbTODc9Gwo/Szol/vRQRffPfM9Hkjcr2L39vHdBzw5/gkdbSeM2Ap8s2CXN1
nkgGcnXUWYmdnJKrwt2T6qzXmxusM8KiKNGVqWisbe135UfMnCoPip12v1O8ht6S
Ez7yJcethlGuD1ZM+kjLLoZNu1SbRiMPEBMef95c6qYPMep0KowXhtrVg7usCcOg
Pfw2aS/gclg/6n5aSrxHcHv0bFYWhEH/vRrZ6utqotfIIDwPl9wSecwA5jEWPr8v
tzgRwne4wOjhXLvXuMELfEFXnMtyKIo58YEcZfWtr/EQI6sGSCEEuBp9m2b7ADec
5qZFV7TV8zsVcZGW8TlQCIXAnrKgiJ/s/ZL4zQvBnpz68LL0hDSp35ffNC1R6VJf
pZbN4C+if6CihbBXdzMEG7RKYqjZxyXktYJCIxTd6UVlbeh2SHfVn41OxNfDR9jt
FMhxIr9vFaE3Z53iaQlpvxVT4D9bG7IVs1iVr9nNrbCIpZbBZl9EniDeLZoGANAq
HjvKx3XILm0JWNJlNRHMf7V6ClCZkWn4nXpEed+5YJTrbLi+DyOmqFBlqlrlO7Cm
7mAhCJxYVkepXSucTj+7L1AkSKOwZpQjePisKGJVK5kWDyxocYZrqWEzrlcAznl0
aBmPxYcebq86hgH4Y5gqco/170Go3gBB2DqUiLmoLNeMxYsyzq2aCAAP3iP+Mow6
G8p9cTr6GH3ECZ/jG/KIAZobzl2Q1WCqhl2V2PUpASFw8ava3s4ytLlCFGdiFElL
l1V5mfFeQTgKEbuDHhZ3hpmjl9t8Z8kM9AT+ZgUV2LvxXyxDZQcStY9e2tWdIa+r
LWqWJmX4k6/tOJj+RMymKjFZSjLhDS/IqboxhhZTzFHTsTucEybCv4sS1MlqU1hn
d/GiD+9IJM8+bulIwigaA3tgmILqOWiycD1qLwtEzbXmAyrM5m3QW7p2KUEkFJJP
+Y8VCsICNxhgGuiY6Uu/FUf+fY6e1nA23GkYhM+c+ROEnIMgH5fb8L2RXFwNwf+L
g4zMRPcJD+pri0cWfIoyXfgoAsVwGO2Fq6BFjZJRP+DGaPnRlsGznVNp3V9eUbbi
b+VXl1cR4lm78+Pil2f+5FPs9pdKbp+RGeAUiefge2mBsUgEyvyTHUNF5QFP1yYL
/HOGJn9vVrsnaufnR5yf0l7r+2LkM99dzd3h84tz4d1dL5ZKOZXjMvpZgY5aFv/i
pcbiJ6eDBYh7EhbzWjHzaMy2SwqHjbxJhtdjN0HlxmtrBooFgKekN27kzspnFnpL
O0fIYAo9QWwGfsRfmbLxjoyRG9nCnQzhMnzg6GVpoA//Ir8MdcZJ6GG3hp/zTKdf
x4c7s/8DBYJH4SrXE4n+9ixqABzSS/nPZLChtsRp59Eaae3WOU7QcICTJ4uv/a1H
g3GHVNyV7NTY2buFUHrdgDa7e8AYOfNE/MbYW9LXjlu4t8j1wpq74keXFodu5ju/
Zm/5KS4CBr22QVHczvxhaZ0sjMuTblRtwAry35fWTD7ODVblhHRCRYKHpN0Akwe1
l78dS4yacv8tROWk0EYEN0lpdJaNT/wzt+5LPtrk963a36No7uaJvAa3R5/cfGsR
dxf4hw+rt0wF+godW+ONiGOYY797sLfY6SBrgE97kYiSYUalfvDGWKOymdX6HROd
M62dRBmcFYLXqUi2Y9zTP6MbFr57Nh+MkUbwvRoIEQa1NtslXkvw6P5Eql+URZuM
gEt9qUt6kB2QXmHHehsmJd4iZuDRUzwtw9z15SerNO+OEbALE9rOUTxii5bcFBm+
83iTioW9MjAjN4T8IGR9/utzgOqQvjMGqGYX2/k0U36RaRNQzF6FzJh6vZtX+UWi
HrQ7ct9wkxBXwxm0UibhlfvPHeJ/tLcYIpQGPpUCxj2cDi6rDB5aPfPTN/sS4g97
t4KRr9Y+zlNtgee6XKonAgZO15UsX4mDIFJWeKtjNiViRxBg7fdL4DRdp955B581
HvRzRoEvf12a0OYUHZQiZIh3pufOz17XeqtO/UpLoOKQvoZtKaoR3GoCMt2+OxRk
Ms5kY8XmMO2aaotvRbpw4vAjiFf6irymmEsf79D2lfJu+BrnHKJ0KjIF05AxP9b6
PU7XDfRejD0vBdJPhAvRgBSr85ZOqlbbd1C26kzzPPXR1vQiQyT87Juy720QyPOD
todtRDXtXGEeI/Em3pL+xDzw++Zd+ISVfIubt6CEFgBLjKY/26e/PZbQbQ5Tc4fF
OBo2vkJqD/hKYMATe7xG/BjMzAWh3hDbRMuiZlqtv6A868OJmdAPVYUKfxY/0bQL
8J4rA697T/lN2GtUJ6mRXePi9s4g2Vmof2GRlWVg+Uew1A5VR/iwq5g+FK2BdUZc
jyC1bD/1DCisMojJSAoXTRURNnMaLkk2qrjvVjJsro2tf3LPPosS0i99i4U+CrFg
qheoiqwc851yjjtIvMBplpdE1VDFotQSPGheTU+9a82X47NwMk4G8sQwzTsNsP83
t4s6ADFChrrbUyII6JeEJrK1+STAROPDaDyspjRnx9RY0IKn6Cqf3JQ0H+5pYcaB
dahr1S9yvLaUMutLXnQ00nChwkLA5sFXwn5vdCpJuq/2clq6X10STcrZrh+ef+V+
DUZsbRpc2Pcr/5yFO3syJfPTqBparf9CzTMMtm+T1iCXmcV5rHojO4Zei9D4iXqL
DIUSAscZa7g3L3EBSDR2Eu78ocNXUQ9gVLIGVZmP2Uu9bMRB0e65V9ldmD+ATSQo
fssaYIRYG2UHtpoNpY/szjaeZ4eQu3wWUrO50o2/qdKWGfQu3t5xOmHci8daJZdl
bvGomVx9PSdBbg1RneLZOMipg5iNmPG6N+WZl+H9rQhzozEfIr+cqdSdxPEG2c2P
rIFPKj6r5bNyXDn25vHnRtISlG+5e5h2YnyM2I3HYH5j76zVd5LHKFaiO1Rcjaw2
SqCvuqxxPjk+hnKlHZTmTwGw3tJWDV7ni+icEZHmLweGlfvJbo7CgW9Faw2wD2Y5
HcR/7C0EmRLplbf5d13ArBSqYhjUQaFJKgCaD0CL+1wckx9pGQfRFpVPmm2TCA3b
HUJSGKxOhX+WyY+2YjMhc+6koXiFwmlzJN+Abf7BcqcZGWvx12/NUMW7rJjhTyQg
1a85uJ8XO9WT8svK+k+SiRY7jeULL+l6TjUICO2AzXVi9Fz3Lk7dBur6+BAd7XRk
NHlMss0d8E2lOMF8zi7vf3Iev7mFwuFuzibE7pNo7XRPrd6Wg2Qn/r56YUWJ/POl
oQfa0SieCpugcFxkMLSWv0E7b9cmDVd6lk6i6MXg0tnfH6jz71Vq+Seen73bqvH/
Wvt7ww9op6DE/S0sR7OVyXn8gR0Lldbkf+wlyqXJke0/7q+lVUfmYLO7XVOYx+yU
JCpqstLGgg6quPyG0JR0QinW+6SO4d3t88UDDlSn+mSC1vcisfQeTaeEQXkidZw6
fp/LBK5aRndv8mvIxXVe7yMv4m6tlb7aGdel3XAo/8tCATwziHpfbllfwhu5qNfK
Q7kdpTOSLwPTjIKk1k/y58+V4I4hUNnl1Rjh+WAxW206TCM3ZiVAEwkk0ZVrpr1c
J6Rp77dZAI7g3QK1r04i4G7ywVquOMTj0t2t6aTqnQDudN58lOdB1kygCcYe7FAJ
5XR6HVDaM62Mmu855N6Hn5hT4wj4ysnh+lDpOfRpwnEzCXQh2+QEf28mDnB2fUFU
b/1XVP8glu40ZqasqS+fhD8+SErMO9HLanpp/x05H9ZNiROx5/DcKli8jFAN/Riy
d+GkYT5kC1IxZ+RqEZ3R9MRTCryDsC38MubJgbvFC3zL3gUKLZoEu4WAMlbbJCaE
cIBtKi6vnMM9G7rwCEiCwme4/KhiOK6aM03I/AzayhyzGwRSyMf+HiyazINikonG
Bsjz+QqnAb0zkS1pNUp+YbYBayx9dEfMgn3YD0ngOjowLOWYyvdPIEUV5HwXr4y8
4oY7GrS4B8bQizJJnaYBFkNSyPOvks7ADkhjHSIR8Dz6puac05/gtTi+arK63r7h
MpHtOdhcwicjyJbkF/RWMFVKqLWSuDMsuLZG9CDzdowj79GsvpFeT0nLWZdFFMOa
VPZJgiQX4C7zdliEruUdg/vcFvZ0+cvnzpvTRw4OsFqEdJJcgWjkv4gT+0sDDUyj
OhqI9I0no66mhfwzcoX5Q8v0f4qlP/Gi5PtPTwQb264VElvYVZx4Irwrelk3SKnX
CXz/MbbOYWc4dJI1xHrKSip1TUYe2uxBg7xrinoOT5Je8HmnI4+965QGYZil3yNr
wnwUAVXgV29gFIm8g2ArkuqUlQ5fhwgVZ2+KWfJOOxL8AL5pX7CggzPBjwoYpw+s
exjJezEaxFCC79huxdWATChDXwSO2FgARW8vuYNR5lEEn+FAPsnACGlocMrAVZhF
aDut7z8V/GFp3c/t6tmLaqdxxVUxopqPlog79sBzMSvaaztoc6idAt/+YyJ7uCF+
MGQwQiYEtUOGuKnfvPUlUkhlyh4WToWw5KzfMoxUGTTqZr3Pa3bGlWwa9eM04Q4d
xeNsZ92AYihCcAWyEWegmOdj+hsaOJiiiD3dOwJCvavjMz35ED/bfzILlm1X9yvo
zMo9wCpozKojKXlB00Op04pGBN/E9RsOk3eaJ1nr66q6IhSR5wOW9UO9vk9T4DT4
tBOOlr0bjqzywe6G/9KKHMX4HGsnSSd6bDaTwJWJ3pUJ96bmxoqys2dBRx8GTZaM
ax4bRKgXFHivdImUIO8PcVzCXGeipgUot53+LoXbBKph79ksOVVJKa96H5G4Naa9
kHh3dDVZzjr2d5j7brQRpQrlsyzRyf/I3lY5leLODUjZU4FutkBBvnnopZeblA8v
YGb6uJlWl+DQwzqUScPkVenOGuD6DVnwuXlswcNAwQHG1/FiQaU6fd3XbSGv2ryA
YRHcYx1s4mQT8uP0gimXE/fY2k18WiJuTtbyoyajS/HGeztUKI4fPXNUv60YyLHR
MBgw7rjYO4AnP8E1KNH4k9FmxmAvzqtm8NAEUS2qDa/Hntz6ET52Xjz6SIMEGxBN
XChV7i3wuVxuQ47o6dbtlK17K1htvAaw2Ka+XYyIFewZCC5S7hyqi4BX0yhaUXuX
tWuIv727DE9+8rIe0vNUFGACzltKcuoplbIYV+qZueP4NwoJWuSXLB9tKxqDe7WK
5pHHg1UlWzZEUKUFI3cTfdAeEVynB+CWwdOTUbFUYpMalBlC/VLIYUwPepPfbc+E
4t2HkK1AuUefEcv5buxSmt7A5zSh4+HRCPI5rkF/ExJX1fsZvyZq54F0LsGycNXE
P3NXoQ+dlbwv+7dfhq0dBRazkZZH8qa2/ZwtPFyDNf008TcxxkLLhZd36euhpD6P
1/lEUq7LPcO08I96Eck6B3/NgzjVY+3DAQhKFwZYDGUS/c5mMKKJ4GdE5zeZLjWJ
phDGIjlHZO7xdS4pnVJUjh//B+vJFLJ4p7YISClviIkZzchhXfb9VGG/fSEgSvhx
m2hCgj3egRSDGQ2FddLydoNdn4RcmalROTwjQGSo1eN3638PwPwaMWSDY82QIf5X
fXrJHbnFXglY7hKp4W2dBvcdsT9wQwLukXHPndrlSiXNh4E2I8YQViFLaKIuyZHu
mH4CPaIxUeaMRjPkKDO0iUkzJigaYW09iu4a2EqLc9HCCGolGBsAn1mejn22RATn
V+YcWe2PEsN0idc6WVKTzPfPA4L5FZ9pF4DilPT8VwSovZjR8Z7vwn63hhpWLXc0
J0d63TllPMXfRYFTJ4YKoIn1H9ZKEqcc2HRWRw0LJM2ycLWvGfDpcx5b1Sy++uVS
YB0or6T1LiVgAzFja5hjgySTc64aHLz8O772OWEaDq7Pebu4+co4M9SwX78W+RVT
k136+PGdpzF+X0lYaDkHpRU6ZUT6xeDLWsfWpmvRthTdGNgoEjSDFvDV1Mifiwy8
uHir9+lkoSTPUUvJgehYNaVqIKToA2g35JMc4eIebE3Jfhda4S2GPekrr5s5nKZU
M5R7FGqKH6NgDJDMoC60OX+L/Xsp+4OKi6XuXJaCmFXLf2TjGcPlgayxz308wHmv
5YM1j+f3V8SXhA46Ur8X/LhlqezB/z/t1mB/nqxzyuVq10Evy3hHaV/qGBBpW1+8
xOQG64SCKOz8h3E6uPs+SIZ9XwBHxMvKKwuElvreH6uuHnd75Apc3NgCoFPZu9Kc
XXc5pIQGZQdzz7tc/fM9oo7qjskLJZtLf2SPrKwgQE2sH3N1Fv3GgOVAIXzJHI9h
V3KSgb0o+0AEFBsoZ2DgHQXjLvrfEkh3qtB3ms3xd7zQ0M/f2CzVnRSSbUGa/aSt
t1TabtB0FwBAyoZ6HyGcewyAgK4LTjfOOlFkkWtT5mIVIMUhNh5cEae6ALUqquYY
Si6NeSzWIWLWugiuQmtMo24nj/xYVZVG2eLNlR1/n3nLslaU7YjG4ncoWnxyM6Im
1WzDVYS1oTfKgKlJYOehDp4kauPtmMgS6q8YE0hFHVPF93V+1NKZfQ21BmqRyekB
V7ghfPZ8nktaNhM8QlQzYSVVDK/nEEt5PbPcn1PX8WDflHTbphSKSss2yoG7x3MJ
WTUmVd0r7KHvrfbKypP6RSzTaJ4ZX+JuDITyhPWTO0CasdeEsScj51/Q7Wj0vfaU
nzm4udNDCaaTNR5JpCyfCcE0Q8dUldva1UgyDUzdsigUY8b6om+9vjTymNLSpO+N
USG62Fc7S8polvlJsLsJWhoqjosgvAAp7xD83l3YSgjLDMB7sNfeI0le1haVONC1
FGjyCLYwvf+aaM3p4NwTQg6zchaKi4N0ZEj7K223VUqUaiQxMbzpMlhxcTy8Fq8J
ysKWfkACsCffCcn6Gfzp7rmP40CFm+Jkq7z85EDJgZ7mCDctGftNnQNs5Lzow775
BOddz3G0h8Disu+IQspkE3S/oEjHhgSWaER9EEeZkWzcokAyvuor/TYWkvRNYMCY
mGq/ksBj1YhVEfbS40GiLkdtf9ZjXGNoes1NDXjffi9n6CVDEn8oxWkRLD2s6bcu
whx0/aBKSYWOQoaibHbTmfE3wj8DGf6liMAyEloyOWepSI42ADGBfjY1E7VI7Vdf
GIwg6t7Y1H5Tr34Va1fTpYkKA0yGCqGnlLT8E3VS2m8/0ALrEZ9xLKesqIJbVoOj
7e4xFNGj1dKMSOmqfq4UZwA3H4dW5HIEYERcNibOVPc6kZr24nOIesnAmeui+DFL
I+rJ5qPYyqpQbPxW4opDJxFyqF0bsPKCNn7yF7LVM/dBLSKO79kuyDfcf+YZi05i
KXlS9dJWaLBIYWwCznbb5xqmnv85Zi/XJPfiTn/seJIm209hmVs1CJyi2vFAjoQT
te9T+ZQKAEsx9Yhsd9CK+j0vSjEsMU9NQdYNF4jlTI7fzu8EpQk935Bk3aLZ8zdr
0/HtxaHFwzihIofuOWtL4QLlsbiOFSvZKk+5U0TY0VvNKHZptCZSYhQRgY1shnso
Y86iYxKOKYnv+prWUmka3NV7rduEOkjjq45An5Ax0nXmP1FdeCLUNMpx6t8Agm8d
LBWcLDW7wP5PVCDv6Lw/8dJdwrLpEKeDC9I6s90qEuUkAVA4MxxXoY52QNoYWbdK
bozlZG14yT28xvBPcubUQfgF3Krc2LH8j/iSaJDW2vfAabF2vLd/oJarhjmN+mM9
EgYqIptXmC/4nhWmJ+edhdbGWQIPUHsUM9iHAqB7jRPtM/wEfVxvCyD6dx+8+a/3
1MwKVMc8GPwplLRW4/aIsezJzKIcpPsWJVeuiz/C6GrWSOLefhWZxPxL0c4Ts59g
pFpqxegxYd1n03Alh1NyUT/5fYFU3F0lgTQRJH0zktHpAHd5w9sWhjBwJZCEgUjJ
zVQEv/WmXgFxF5GXYXsmQfb7EqC44hcG/vAh5XVOoQYtwAbaivMkqq6SpSyeGP5o
7Bmy1/ZjB63O91SksZ4qxRUiywziPPDKFbfLteK/0UeI3wZKZ7+fGrRT5D1zW9JH
kzWTwsGFeAhkjVr7AnAlkMTdXIoSDPQS9qFPahRzpxm5Z3gv23fVBXy6u/c45LK0
DtpHiptz7hx6pN5dw5sF5KTVaFXs/qTDcT6AVW7A8BDLk4WsArr5VSzNwhqrwY/6
DWiEtPjLTuLR4EFkJDwU1A==
`protect END_PROTECTED
