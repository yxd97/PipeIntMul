`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KNd7iG6vIoM/aBqoBLyPy2ISQwj8XZhDPPUWNWEl8c/UMmcZaEd6uPBZidLipxB
q9vf+Wh7UB/MW3kSIiZ4nWLIWlZ9gBB2zxhe+DjCaEYmSlEFq1lUhohMkXSvsO9a
eDPvExvjOUzeqi7cTuiS94BTwdJ3d1Da3XeO7PSRUIHvM+bVqccHsM/PAntsr11e
hFpI4hyRTiMd0gtTfKOhOJg6RuGMpz8Dro5G7wGm2nULsQM8Dr15J0/NQ3ITnvw4
SxrgJzWj2xugWhDoVkjFhXxzaxm1U0xAWAwf3fMZS9IcrD6nvpdGbFuWcij3QXKd
yblAMC7U/Vzozkcrxdm/9mD8l9nNZwamEiN4vQ0s6gU/DnJxeisNGHKvvCLSPPnv
jXHIdm5S2vU3dzwMwNuMmYHiC7c3pV7RZYHw9NGMMoUD78NDwS9K9AQRkbSxrj7o
o6vyzJObUTpk6QSV1K8YPKZpVxCLUHkQ0bOKtO0oaEDEuje39hBwlRNvCkWDQRDK
ukHwy5eH1/8pxPydHOG0npgQ2ur62LHZGs8/H8qwteMRYkIXouPbvl0koDV5OQpq
`protect END_PROTECTED
