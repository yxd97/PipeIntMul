`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpfDXUCwfbGbRJvTshTFMEwHJjBRoyeJKGoT+a4zZxNN8c6pQKaW4N+t5YIPUpkz
Q3LVsON46jpMY2OZEdOv/TH78DPbn1KT96kuFgMNYsp99rsXoKBhD7D0peaUXWFY
pfiMWjGBTHi8Sycim+BvfO8Em3eL7pM3hzgkrwv3KmD1zoQEZsMExvyXPKRHXmM6
cBfh7otz7L5Xebwx7aySVGMpTdG5xOZ3+s8IfIb17TO80Kiu6ocSefjKTHJF6w3u
9cM/DROcJ/WVjLxUoOx/B841PLevb60x2iaX9oLA4VDeeB34eHbU695aXuM6BKJW
6KZeMfi9o0jFUQV2yp+xDaUx9DlAGr0un7BqO+0RZqprSqI6DpnDb5O+0lZcz5Dh
/kekfMQpMekYeuxyheILHogBCQx+y9pZJjGqqrmerkjW8AqcZ/ciPu9LmkkFH4wO
1Apt5CDm87VaORmFWq6w7gDCebltG9jnkylj6ri8jcs=
`protect END_PROTECTED
