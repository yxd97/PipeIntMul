`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CpZBx3UOaTqp7bQb4+0BG4JoUBLs7gNzydVQbQu90egJa5R6+VxOBuNtmgwZbgxh
bPGRgmhyrpuFOQ2LCIpMpsJ9SSCZMGcgADTbeUy/krQFHEvh7D0OE845dhkCgol4
gncPrZQIPqHTQ0DfAHFxqp75rapG5CCvuIds8CGH5x9LxFl/Mnti4Mc0c5gohnUQ
g1OJT5eO9tnylFY5xbLXXsMJP0QosC+YrWF02l+bojCciQy43QA9Rz8xswLo6VLA
+z+sDuYOX+qeBiM1RSwJ3j0lvx3874jtAR4aPxKJewbLgabCvJXp0giT0yCU+jEX
wIBaHSGeFFafJRyfyeRo2P/lC3DrDipH5ktiIkimrbdDllANOZf/qp76PwTqJ6tH
faEwTCYxQglaWbDq9y2NFrjczNgREjgJf2iRNay0L2dSIbeo+Kus7KPrxlLuSu3x
S8ggGCoHcnF5gapCIZTjo/PUE5BblRs6rlyJ/gjSz93P0eIivgqKcEtSQepiVqah
UPyekd0mCfF5qH//3PoHBzvywvuBbCJ+9vRE4BNK2ZyvAkyS835aBvx4CwCj2OzH
t+gHrvwg6uO1VCxFiRb53uSvR6NNuRlD0p1UABpz4/sYfNUj1rf7aiXq8vNjn4F/
MZuznQU4xt41DEw1qnV2yylGfpO2PAD0uOhHXQnL79UMqRnzJnXqL0hOnew1cQBa
cB9ovAyzUTf2n9cCC8WRr1PhE9hCFzIvsOs/joolEvkUL1C72rNfWOqnMPo5BQwG
Z59ipVX+MXEJg8WrYibFD3QcwQKlKiKRe5SC0HSQevY9ADNqM1HcbYV32EXLoyQ9
JhrrFg4wlGonTvMwZ3lxquKvwDWYexRRlGv6spW94R4LOUHaxDEZ1Qn/FMxDzda6
cIVDmt9QnEqvqMRWjmivdFX/YOTpd4piGwbTCeuaiGo4uQ/1iYCfFCzqgCThW7Hl
fhRHuzukBcixLbM3mffyqbNIG7+Xilw24IQ7OZNoHk4w01k7vNWLpR0cjaKKz1qB
BGB0UKuP2EZu/0DdGQobJuInWf4m283UdDVTgjXDkGtBB65q3ePFXnGfijqXB77O
4oL18ntFQxfPyb01sfgUgvR/k4tLe6kxiJg0aB4behELaOrCw8ZFWv2zotQaA581
RcFesluCe69C+MWXdlCq6TtB0latEqghOddDExp79x2MT5U+f2eHlelNhiBiGb+c
Do9/mQEzDkYuj89Br/urUA93mif9KOCSeMoIlTGsPGOTP/R8eHUDiWurwAS6gDUG
iUV/CTSKTs2qXl8eXLx98ijLuquKl9gOpZUFccNQJQnxrG6MTC3HVZ7lk1JPhB8+
lf9YR9aac8DzXbx0YdY/XEPOcQXfcWIlLhUDoerhPXpMverSsVg3ju6gbylam0Il
mJFTmH2qC+nWMlssG3ST+izQmGZ1jqBy0rsOWmjNrw6M2H1o2qvTqwR1T8ye+9MH
JOEU3a012mAstZoZlXCcUay4nb9h/T5DDSrtqqc+geKknlicTFsdRxqwuQTr55Hz
rATWqsEO+Dg4MfaKSqbG2+G4hSNdCBqnpnJhZkbCLcsyv1CAkxOwWrL6BrYVi7pi
s+ZQPuHfxgRfdFIAs8YuaTKxPHErqIoBYinFquewLIsrYudPDC2E+aDEbut6fnzx
UzcMEVsRwlPcTQCt6eKmKA5Dwj1STF2gyTy83ji7sX3VN2NLeXQQAvoqFGB7RSYd
n/GFWQjeXKev5aiYVorarkzDvBMNdbqS/cW1aA9wYyf+rF+yaTE8/rfXvoDnLXsg
2+CYtnF3UYtsNMBHJ4RoRgEoWsIlveKeefuLib145QCSG124NW/gn/DeEyIehlk5
ZSZ3ZfWfgp4f6ARCHMRo6a/kJkwCDXS7Berc/GSNObw1ZEVorLbKI+vPbE9Ob/j5
zAv+spUtoKILmEr7mQ+6/nIKMBjx4RE25Sn2Kyv5c4hdFiqqVBGwIrKj4txo1nGr
PronpVhZI96hK03ERWV/l6k9N5ygwKnFU/jKGIWJEOh6cedmtBEuIhCT52sFqgHX
ZV9el1KTdcGmMr1j684A1RkphjL/IsjFgRMrQJ2bw2noIEOlsPQn+hE29pl2UpS5
qHZkfByfXNtbicprdY1+yxXbujiQfuuZN8/bpAN2ZOl+Z+PgK25BoXzETojJss8E
3H8XWD/fM9u50TNlikyCoAfGxlm9Zg3lJlFVD6RgqUIJanGg11rmIUIqHdTfXm44
xi5rt1PInCDJtdlXZHGktOqEH7uwI1mxhJ5uPtvBb18sHTIMC5V5pJ/hOjzy/jNJ
y5OeLZpx3Z+ymumAq0u/DDYOz5QZ6gwStaa3RkpObjz3agGzMdAUX3tVUrPSFnh+
EH3fEW97bfi4VaaO0gVZOlSuuWO80IZFDwqQlcM/Ss7PunJJkqAV4iynPy+TE0qe
YodlqBrP+4sN3GgCBiVT08atYZwbXelaeqYt8mzr14Q2CrSf0lYHazUu1hpUPDj0
gJCVwPtUb/NsM+5n5f7FHh55I9u+/GuAVZQoVj3MWeQ/+0pBJPGxpORqsJtOPCel
2ntpj3fWY2TqBfrrce4vSOiiLugsCrhJoQ3SuYn6g3nERoybmYpCFfw8VDgm5hLK
JYSJQCJBCDEZI6Yiz3XWZGwuUFj5YrSa5ssEvUNzqkHhP8nGUf40LqxJ/z1I53IT
HUUkgoQXq5yDgWP6TH8jx6jhtiCBpwCCIODwdQa8SISnGHeIWiFW8OfAuP/iu21J
+rsCs6xL6gkT2jfuUmb7BgPENwbAKwhXqLR8qaZQjFX4TFvIiAYyVziMz8K038IA
uQ1h9angNNnsBVMi/BAutEqWc/gStQmve2zBOW0gQTjGhcR6wzsujJ3ljCbahY5F
ftzVuDTkwiaOgROOdNw1ABZLMkipydWI9PpSTwQbvO/m4ql4+SjWqoAndVbmka1q
7CmWCNPS5fY80GHE+x9cKqyChPVQLMPbyhZYq6uBLg7DdQ0qqjZWNhplfiaoC+Wp
1TXYvYl+xvmfYkVZL5vT2SYUbkqU+sEYOnP62xvQcWQDlwQhAngwEFPuJvV90ULO
zIWjDo9labew+YoNMJgOjXJFjQhEdtg7NE3wzEi8ziw+oBtJT6wDJ70m3dfyPAnF
6Jzo87zjpQiiwBz7mt22wuWArzZCr/hYu/wbsrje3ns/jaC0nrOTiM9UnU53U7Uw
P15nbgk5T0NSHcYOJIo1YmHt8ugxzlujtPz2TirYuaKt1lNIKb7RtoJifj+sborG
qwHGTsoUceVvuO/MY7og68Tm0aplFAK/oVhCvIEYhTyD5aVjLeF48OL8MsGLAIVL
CiqQUpxan/QsjiJRgh3CQEGf/JZziAgV0kHPLr99HTihJmm1qD+z1E/injOPJSkF
rX7f9BtB1wz6X4Px75vB3ICsgqdH91I4FyaiCQpIoTbX2VgyyFP40RPTF72BUVxL
qScujw8NVzKCOzs2K3wscg==
`protect END_PROTECTED
