`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9fTPMQWb8S5P3+TsWWHdNAyN19m353mf6FRhQFfpjKfwTFep6MMAYQf9W7utzmLW
9FQPhhvIXjkZ2TkqqB8ktJ6eWowOJlQKO33nR0a9SoZzk9nZook22/n0ZhhGrgPk
37xb/tqidj480pAK8nuKf4o3mReSw21m2cM+kQX8LaR64pjiBqwLrIa+1LeSiG2k
odlARB2cLYq9Itlw8aoXK88Kn5YU+62qMRjjrVpnZuDZfkyj7/S2ziAhaQSoiuL0
O8dE3FIlc+ETLeir/UmZLPO4lbGDEWpAVPoMeRuEbzCyQr/Gc3W5ZmKjiWNAHKlt
Rnh/PvR4uLA6TPCwwXWWYiw4DGceFo2rNs9Trvl8EJvIWcxZVIkLNUddqDbdyp1M
OCHkg4KSTLw58UdPMqqIlBVpp0ZKO4CQ3DF/69kHV/2eR4yaB54Sqy3XJbvm4u9B
SSkAbEmRHxzxIh75Oghx+5M9jGTOQMvikmwp1ngTkXyT/AQylpMo2KkLn5dgFlaF
xE8kuZi6KHHZVbiapS5c2XFBQA3nNFMwBxRZDfNY7+eofLa7B/rVVlyq/g4jZLbc
IN6BSEfvsefjGIb/A+ygOSG4Su69EVUjBHD41ROGuipXkoBsG0FQNG0DNpYTJrue
oiqanjmDIgDE3EJo4LArfgWnUpEJtC4bbSkqLLtATNjIJsIiCk2IkpXiVkEeKC7H
VxOc2NtN5uyq/DUk+XMD3Kr89HPykHsxckcUXxO/f4Uufi/LICqgl68UcWMTSaCI
Ii23HtwbcNck/FUhEdbrQQ==
`protect END_PROTECTED
