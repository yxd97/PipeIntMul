`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SIW7NqFcBYyV5fHYaOJseCJsPtLF8sl8svIosxR2JZhpzAzlaBgzGzliSGfzRPap
eR9ynNokR5oryYrHAXiMQOByaOQ+G9/lADTMvgQR28rmrtvULDWCQVBOBUk8UtTw
xqfgdK9LpRPqjbKZiHpIvsUpEVkPV0lL9pSOTmHCURv234JY5VE6oybSswt4nV+U
nrnJbOmT7JpeYN31db5/uUNS1UlOuKwej7gQAydrVVaC4GyZUGObYlssVlCzdzdJ
7VrlZHh037FVIrG7P87m4q4B3ONkthPQt7tzN0gzVIdNmGi+b8qe3+9+y7BVA413
LFZAFEuMLTVBVXYKoIo9f73Yv93xkCEDLWLFP5nOGQMJLk2yTobFoNxBnSn71IEp
rqrjWGA6K04gETtCcWM+OsHeqA7HuCfb4NFASwS2tgnSd5JmURXX0udEoqOERVxU
n3Te/Lt5ZB86n6bTOneO1BFoF7m/sgC4KBImvHqV6ZMPs/W0eP/z0a7k6Ug5Dcmy
V+ivJ/RM0exEorVZIb7HIqmNd8Beu4/9vZmMj0pAJACJy4nKbALWQXvoKfRDrC8D
lOMXWTJlmNa0G8cZbVmZ0e69ve99VOUT46610y6hXlOcBEstp9GRoOKAz67Mmj+F
NGbPb5eVvxPyWDpPLtExApvEeeHlYCj3z7mT+ay6izrVvb4Z64YIjR1wd5D+tHue
clqIYaMWqKcZDDSXxzo24bYoCCAzQ4tmtG0lN3wGkL/wItj9MzyEuGaoThjBpwGQ
sW8KKwiCJ1u06PLv+Q/9SRb4SGrXpnx5jqKyesKjonFbKj9BKm6ifhxbe740n5pd
HMMu+KBTzZ3EeY2wmpgsVlF/FmoM/HBzpgk8STqiu/AdVvVafTn8dizVvtiBpO25
r1XEfkiX4coomuL0klF48Rmz/0DTyLjFDnI7qJuQE8257M8k7riK4cBbm0OxyTOW
yfYRl/USWFdagFL+uH3QcZ/GWTBaXmt6YwnHIZ02X/SkY3sX5fGBlAsU4Rdeuhi0
nfJoQ78D2A3UJuX67UMTKYIJfwqe7QX496HAmrbGOS4N5BwhIgASU1GqQeKiiQL7
ecyEabyomjBrfNWhcyZBh34R2kuDO5qLakgVGlURUuT+20wX43V1H1gi5O7J4/+B
qc3mpHd+4aQcuQd5wOLwGAFKXg8nBksmbH1gWCgpLqBivZW6hmu0DVO9LtUP2Uym
YcYn94Q2e83YV7116sooS8khDGKHAqO2FgSGRE8POqEkZRnSCbez1O0eSAzvnfz+
7i1LJrZy88g+ua98ONeDro2SQCYgY8QQQWIrUBscZUPmKm54uwn/LX6SMws2NRd9
n8qbjBVYSN9HA/CdA0GVOdPWti7MnrQITArmoarXSwPJ3LgF/yuHBdjvEHzG4Dt8
5uruNI+3xNhO5DBEeBQhoyk/SZCDTCSSOtmGCOytzA7X9V/4mWy8Lig9ItMfxpSv
BVzL8Xi6RHiNn56ady6enlDwtxcyuoFfAGXfDiaB4EdLjtdbRo9ObfrSvPbfhCsa
7hAgRFQjbsW1jic2TThLlxiP1y3uqjwAI1sQjoYm5aj6lp2FS+PCWC7+eQgoDVHO
ZxPi8t5P21Ji/NtVXVaFYK/n6ig08t+2Ub/8ntYeU+I=
`protect END_PROTECTED
