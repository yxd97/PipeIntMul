`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtZkmBeORA8+I4ExrKsEwDJi8lY1h9dT23g52nOFX2NlXzYhqT/Xvbo8KJPh+b5M
+gBnWVwDwUzhc1t8gT+I+5DgaMo4ofH50bxFiSskxBXOWBRFS++tRxQ4ENTdJcXz
h+fAWLrrnqB4JhUe4L808NyehFN4jWMOO0PNOBd/gmXxSP2PJuhGX2UFmrb9AoSe
WOwPp4EHY6MMqFaCuDHhN5WtJQF8YcvY4NhTPwcbJ9qnf1gs5Thq3p+Rz5Rsr4Oc
Dz32/nFzJ6gmnY5BMGJFKuG8qoeSiVdGYR1OyS4y9jJRKlcNgIt5g0+8Jfn5iaxp
5bjcrw5OMN86+xUOuneThzyouQOfu/NPaF+3HaWHHZnJ/VGXeylQyWXoXFV+tniS
h9HdfnlK340AblaQEg+NPrwCViqBK+HPkELPXCYNhDsZth1DsR7sEkmMAJ2JXM01
QCUAVZm2D9yVejsB5BrLRDxQRp59/+nMp2J0rkhmzLLqq1MoQTu5d0CYHaQQOHxE
`protect END_PROTECTED
