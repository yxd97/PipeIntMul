`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V0hjNJTD0G7CU9QFsprBsH4RLSRj8+5V75AaFqJbV1FGlA/DttpfWUsTvv0ADD3V
8NSe4A7ryB96ek0HXS9WFwHgreWvrXmmp5+t7w0OAcvxnDQUt5lgB5t3IoeKsGgm
tg1TRGAJznob1CIj17v8jOd2O4euWwpl+diCxB5XljpzzC4ZG0k/ETniOXPW/7TR
A9uvg6PwlDzhpdMFcHBv5Q9h+BB4Fu0+es+0xZ/F9EHGNt7wz/ckK2/Uxs0fRSOa
0G1aFfXU6j+zg4OOG1oJE1NzAN6YciKrDFKsWKGREXzLU7JO9vqgHyqV/AtOn0dO
Zq2vK8E+MzeTXAqRUcS25eQ0BB32pG6hX23zbiNz8HaxY2LFqXAKwLQGAQKpTlCw
te6El3mCtKqj1hiHacMCjop/2ll4nICsDbV1UEIISpAKtrkA5ME4KW8zfyS3Gfbp
iLC8KTtgcYPfkDW97zu3xLfk/x9zm151afRDQim6qz7f/UApIF3IbwEnqELscIT1
gzP+AAeBQRyhQaKOtDdovNXdlJlwYISFG2jQiLvfiAmi95NeBqzPtJU2EKc20DoX
Q0i1zkjwkozXXpqXQs/1AYWJAGVOAsfqLG0JtuVvUcwW369mag85Bomi2bRSX7/+
YQ8qLOucqazWSa/qhUmgxT9TbkuLXroD49BczIowLzC5YvtO6gDafBFU3S4Ozg1r
n6rTh2hvnX6x7fmQRCtg+v3RAEQEveSYzcRNcKtXXwx5lva55B6rtPP4FunR/W8y
Dyt7Z4YzWo8d6DNRVLARtsvjbvT3D7/Z1ddzDgISbb6b4YqoS9L1bikc7b5S9dp6
SXbjquhzVBzcy1PqNM1W+METq/JJ9H0ru5mNsL8C/rO1+7FYFCJOCXRPMFvqgJvj
hf/PazJhisAusg2UIaBnUkyeXjszt5BUAaM8u5z0gLuiSUwzFsEt9hYOvFmnlT0p
bqS4rqI9pRMLFDDeZ4RTNttnGNZlNpFFxIBVd83z+YLsjvSz3+HojmX9oEk23kdD
/rP9cVNZJsBeONVxrLNqwsB0lgv0rU8SN4nikVZw8ubB1LAi/VNqspkXBbA642+0
bF22QmsdvMmvEQ8pMUTgkZsQMpuJsfuETrxarYEDj5Sk1VrNS1JpGFgnKGceEixj
MEmKm/t97LMjhlBSZc/tJqBt611Zw/ikFwM1dbLuxTql3bYx0FbdqqTghVAycqp3
sxbG3gSjo5Ofzbvuoc2P4ABJvBJ1HqsKXLNWECcJJAsbmN+cKi3BooUAaGRHlPxH
R8HwOIhyxWXSiKKBZNVuA/VPkFtfGKqR039jKG6imO5AW2D3XoKPT/TCvpuoRvBo
2b5eSG6oZVZYdp5TMdBWD64mHtN91j/XappTnjQaJgrzP6HvpThbFUsGOEGfHFIe
vrrGv42z3m+bpo27bo6mynCix2RrvJV/GI5iNFlypyZXenKzfGJ5Wkz68/B1LZbX
hs0CsvjLmZi0NdtO/rqBmHMH8XI2QuvbELhBMWf6c73nP76d48v5rZgNMiOzfM3/
ek5sVlSOOQWAIjOckELRmzp8d1UhsAkZW0O6yfwzuiXLOriKUtdtfrrJHYmnMxRU
wXRaG/2grjD1Pr7dz55WOyXZy6oHmKKWvdhK7p43Su9omcmo8bl+M42VHmD/woZp
5BCFrnquJ9nGgbgCJvA4qnplSGp69VT2qvqGHO3pBA2mMx5tjxbcSnrd1E4PKj7n
A6yxK/doJ3khOKZqME4yKAblLSwzcItBNLmoh4DjOEX4YHVpFZvJvLPlSr8rDRMG
KV5dy3eRwMcjBBUZ1nc6J9VkJwsC11SFbgLlp9SWbUGzoSkURfsdJdoRVgpy7hip
3FyWRD739+7/R7W9e8S+/Y4lwMQcYu+tA2bNhAIjfBC7p1zy4z79m6s613YDTpp/
s+rv7Kvg1yVjR7VPT5lOUfAMQn8SkBZClM97ki1Y+suGTNKDGv9Ba1LqH3zIq3f4
2ET6kxxuq6n7zUA6kB1uXysZvubayaf57PmiV4QenD4cuk1+2XITi32FgDe/CJ+e
4xgCHLxVzKBPqVhPQ7x+aw5VdwBFOekilsLuKIE0+UlGDH5xhz8ibP7a3W4nzzMa
ttE6S050mSYyJYUzXWZT/H2TT1+UjrhiCTu+6mnG3fvxPWCFAUn8x7aXs8sdgV9w
NbCoADmRAvYFuRSAXB2nrHv87dKfG26u2ft4HwdGJenTCu/reBmZ0BlA0UlAazrp
wUdR3gUk7XfdoC9t+ujotqiLbSQh6aK2OhMcMw6ByONire2iPXzbtKSfyg3p4yU4
QKk+ye6ZQK7Rp5fBuuykcMUhXEmHfkwrDpMFk2+bMQGcqIcJ3lMkuAPphI1m3uti
hfBTTIyeEn4eXaxwr8ECx29Oa6eIOCgduMZtCsZri8bmv0DZXhp73Fg7fhIVYmrN
TvVyQULbRWNHHO5fTMGhnlU5UDfARAs8J7d+yZ3+qtUBNoWrLUrSPFtDChnXZXpg
HAZ0KlcY1wpXzLcIMHcYTRI1Pnz9HvyfBBcmux27El526N+4yZOo1U6FZHLBqZjH
MvJ7RYPoPJn8UbrN7MLwx7EoO1DO9nqvD86co1z2tGdQiCZ+BB7dbePlEBxJTSpN
kO2mJD5iXJ/7aWvYWdK9fJ7rIajJ45gtekuaCcsDtzrG9sZQZVGtiQcm8xipUZQ0
ZJv7iD5F2oIviZcIJhMYNmPWRmFo97w2aWZMzUxjYwVHCk/SuAWgr/4F1SkaV/F/
GUCNWYPcrb5VtQMV5DlQI5DIeSIdrJ/HFk8qNFz6yArEUrvUwiSsKFXy0EbkqYHA
RaIindGrG0o8lfpLmRhtklmrWbH7dVG85DZG+GshIJ6gYkk2bCYXB1p2OLncEt3X
1zeLuIuQmtHszUTxv9A51pgRTtJ/Fvruz4yG1x49xk+GD1AjqKXbv2tJVJlPDfVg
hoiZqEMCGzWFo6WJOWmcvXiJ3sRIioMCYAsRuoMJN6o1KEKxXwClzKd7fcOfpGar
Ydm4OrG4E1Yegm7uniqtmsspfEy1Uo8KEfz/5w7JWC9a2ZRuQKV4/Z2O1ZYbKABL
rySPl8K03MVIplwJ4H5rt018HH7Dt+epKuByu4MA/xvSsqJKuBxiGC/oQ+YcpKIo
y2UKThUTNLZ0qvOoAykU9F6CfHlF/gmA9mBDglIwtQr9y2bPE9vIbg5QQ2qqmuBT
G//TI/rD4nYm4031qsgUHUogKewRUHM2RK6lFGWggXFoP4BqeXdPUsNroRCTN+OY
T2bQM6gPtmxbVgUdMZD2M7O7DdP8jG9HwhJWKicUM2TBRk8GQSP5soVLeNLp+JVn
D4OXaU3LS4pN5Su4ELzbz9mz/ep3cO0syvwCmexpHacFn3mGZzsmYnqWAPdbhzmQ
/yRy6B/oKnY+Sv7qMAytn2xisbPJQLjGUs6PjHmrddzIfiKFU4I1DrxuQcIqQv0N
W2FCRaDDUFk9Fl0Meej0138Jb+5tb54vpCODiBf1NzwfvPaQsgQ1uj3vngXRXn9F
Cm0FtU3L3Cvb2NxA5Yc4pc6aDOVB6tZ/hlOEDR+UhS1atW1yoKGDNvU9qkFFkzdr
pMO8zkJedpJC8NsAR/3p587kzvjatlRQf0ubgbP+mCOHN+1RpX4y1/AIGhkXiN7E
krARrKxaeWl7I8l2rKr1GRvao1BKt/50k0QN2fJHIvO+kD1FQiYEMwQ0PZ/lezN5
zP3Hkb7Oj6L9mFWz+OnRIjIL3/dqLzNabZ1xyGaOWcUkf06R6jp+NzLFDSgaWoLn
3tVqduvk09hfd8sb+HvyR9axzM3gCVH/Ic3A67S2ihg3UEGJyzfzFj/8sOJMhWZ0
vtuTjn4+GsAjooLOEz181NrGorMaUificmWuT1gO4EZzMDygWD57T33aGSQnT/qB
XRmsaaCxu6r3USdiyB2OGu9tevukJ/z9J7Hdjk1HtaxmNAOkG1+WCq1U61IGhbV4
bYA0N0QwTrghyMu8JVn3WHiFSq9ccgwkgAIuub1z2FjF2Uk37Snt4nReAfwfADTC
noi1C+FVZWegj8anOA4Plrykyf3LJ7jVjlNZwgKS+iXwbRAfisQc3PrWapw3L9OK
A842LVPRuaTPCdo/vCxAmaDuF3hq592vsxz9m2Cci0u/rE4W02a+GCOCEhilIHhE
5XUJzvsWRsTRHic5KsJaojycc+LbpuO2WbL6TrwhQi2nK/7JGyHf3xD8LwLayxYE
hTABtMbtneYvzSHidEa6JauyNzO8a/1K5Do0GTVlObxeuj3lc6VYbXwfpy4ASXx3
wIzPWld1kc+icJztn3HwVV4658dShVDV3RqLQO8EYN6+1uHyQ5xc5hjQNl6miikx
NODFWpkTcVnihGUuI7UgSnqcESctUEIOIbO4hf06hilnaRzm/zL/ffucCpeR7Frn
rZfuCwOh4cye5QDpoq5jd3+suf4HVFEVgLv7OJMNDYLWXsn3zh6oJXKI7MkDDrbD
EkFW8x9fnSrE0eReEOAumk/3vWAf/zv04nELfyz57jQtOAHmYSk4tReTk8SnvWKB
Ui4nqkPvx2rQEglB4thDG4umBC4hibfh5RoaA6Op67Hz0kNXdTbpN3/I3AjifF9T
PLmRKeKCQJfb6XgPDXQNxoSju3rBV8Ka6TM8iUh/8ZCyrq5jJVQXXCrY0TpGz0eZ
TyLa1pZiyRsMIePb5Kf2dRSo0lK/pKatILXd2Emv1Fzlny7TMUkugFIqpbdpdOsV
CPiSigefsyT4rDnjOOgNIHsEGPQT9Y1KKLI8ZWoFKgPZheZlRx0z1LGgrMH7tsbt
IxpFpipxaTbTGGVxZKCEy+Fxux9Od3s9xQJvw8Sha9YjT6dOmgFbALQ1pJVOCj5a
x9WvSUB8ztA5/3V66fKACRFyBeZBP/Af9K3TTNNqGbuoJfcKiWL5ncmQy+yKAdSS
VhJ0HJdnBCPecyRZBpI4oC98AGR6qWfRqWuKUL6G+OaBgzQNjoBzyiyx5LJVdAWX
WJqymVoEJveaZ97TUrI1i4pQXdO/mYNniQzSfwV+XcUCIr7647gItkCkA7vredHU
VssvXbRTCp/V+pUwZU4uwdlnGcg4PsaWoIfC9lqR+tP6axo4rS1BTgO+k/7zHuzb
6Wq/rh7e0b0lrmIP930Uxr0dr6bfzsmPbEzENFlLZ3tVgqX5fbngSSdO1VOndXzS
mDyCvauFsC+FZm4zZzRlfvqwcOTZPybPNY6QFwSZek6G8/0jH/h8zH3w2cqimrCO
qT/RqfbqFYWhRclm5HW0o5uUGxx4Dfkc4O6TbQiLDRt/yUpQwn0XeWYSA4MhetZG
wE1raEDmUNYmUJz491a0exn3NPieG65rmi62PAG0o8kwsEc4x/VCjTe1t67ebbFj
ruY/3SgoVHJIjvYge3Yr47YCrijXmyRpL42slUZTRpoOdXBi2ah2ZYMPrqNN63rl
/sfMCG0zfNvX8sqB5j5Qzl02APUPb4YxTEH3YKBqjBpHpgEJ56oET29JJYiGKeaC
rH4rknhCefl2JVYUcmiBX7cJVP6QRMm4yFDiFVPG8oJqpRUN/qD6r52SfvjgZODG
c6awCmPq+ES9QQOeLa/f6NMHq+iSwVE2wjUdTFBw7KBJ7tUFAbaOjahgHiLNUUqg
WjhnhoxELpcZCPpwL72RiACWFLSILxJWsMl1Tv4MZwwtarVCX+PlsXrdMJHAx+HC
lxViRV3TQMiQMPsMT0501AEgYhRF4//f6RL1eP62xQnxNYXGzkqI5KrOMoFkE+hL
cD5w3eAVk24ikEIoDF3MFAzAGUHuSPnCAQABTIo+W1OO6is55wMzygm3MLfDUE+Y
NhJQIHe/l3oLq5g3j0nFfA5d8lWMqFCbSBzi9k5ghTSDhdlGbFQgE90Ql1BIwSxi
bx5nN6VVCf9RWv0CZN6b0D5s5ScC2kXoR9Ks6OP24aRVkWN/3dcHMEjZILf8t+lJ
zcC7ZDNcDPnFPDlQy2xuVHuJ2nqeeysxwZvrPmboFL63R2LqcXmNz5DjV+VJtIhV
NLQTC+BKvyMKvsq+CK3CORAGFZquCS64D1eGRaelNN6ZF4e8O1h3wqo5avX1otDj
40A+1XCsc7e0PC81wVPWHzA1HofANgRcyBjqx2WeRMIUrD2wRMhXcA2IcXxHdat/
r6EdxjB5DUOI/eezIcttKPIdi9GeWx+BL9jC3r1I9/utZZYihRuCkXuoRHKuLk9d
/GcJZ3gn78iMxWTO2M3jOXX99KV6o6UHpwUcbdrckQs3OK1GrhP6IVfCyoSVt4e2
p5OrhXUx/hyDGX4OuzTcdStFrrkZVdnrU0kk0CCoQLqwJIuXq6VkIye9aJzc6RuZ
B7B7W8Yg6S5AeJRknzicm6qmYusTTF8JTdiPuDiErigqcNpuEKDOtmT8c0xs4hbA
IhtuRY8vzJz+/LX9TuZOHuouUsp7gKsE6YqnBPs00ncUWh9oNZ9rIBFwm/8HE/vn
n6fOpzTbhvUxYxqI6URRFMRhB/8O2m2kIlgfOGgCDXYJlAghaZMs4Vikiv/1Tl3l
CwuTm7ZMaGZ3mUB/3nWL+zD+VYAj4bDgz4skAWpDXg7B1+y4yf5XjEC9TfRHS2mq
V1M8v76YxL6cR3UgJsJyzRLZpwKZ881hZkLhDehxhkJOtU3JXhSiwVbTKlUneffv
TmBSd/sFNy2FfoTA/6ARHGz+w9zVEDJQo++EHwIPMIq89I25+WsmLo5bo9MYrGT6
nCwe67jEkTcorWtelR721eMPQ/ZIje5R5rC/hAvL4dkNJGf1+bxYy+/AwHCzz6gI
dTl4Sg9LCabkN+cwYawq4LHQ303Yg7LALirl2Mea8CjmuNWwwsmXrPTNxwX6h86D
QaiGfHTgm975uYIEUzJm+X75T4WA8SgTvx1SOtx1HZrUBbqfVFSAl0kZ3XVPEGeQ
DVBw9kz/F93KdwDBcQijVA==
`protect END_PROTECTED
