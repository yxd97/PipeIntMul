`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
udHpJ5o5sWf6SMBKHLejRiADOqlrGtL2Xew67gt9YfaQEp/wnl5qxxyZipWyPDLv
/Bmcm1047iZ6deU3qL9kBISDEsadNnmJ3pRQy+YdP0chutGLApli6Mz6jNFJIvYQ
0fpySxJh65hnwxn1QQZqTf9l6JrqjHSOC6kLxtbeGhwS3PlgMhaeqB/G2WFVRBTs
m/uCaKXqdtzOTRBNJjvyY06wpxSBOMj3/u676LWGemE5gpWQQmu+ywySxga8kW06
Gwtz7O4pfEbLNn+lo+dvUUk5SO+yAH71dRQZwD4RcquVk+kKkoMWccYv91Lf72FB
`protect END_PROTECTED
