`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/ZWPeNF5qotljXlWYFAYP1yK7pmzXn9YYI8piFm/vM2Z64z/MT1y251ASCj1mwl
JUZqWmaxTyJIe6fhCX1GGZqH0gthCcslmHTEfvCN4v5RqDE3Cw7KswamK1fQhj/m
FNoZhi/cSJQEGnzKhuR1oIuIFOfgQLQgGxYKElj9BnGAwf0gxEw/BlsERIyE9O3U
BHqvAURCb3inzor2ujdUMJt9fN8qbClW7BtrJWAClVFHQ6NMrogm9iZcxEowfNt2
09FO1+yzqC3ujSYQcdfaTiazJNJB3JcnpOPmbgQ1SL/pTbm5cBrkeUVR7Izqov6J
`protect END_PROTECTED
