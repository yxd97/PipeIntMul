`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ep0OJWMSGtlJ4xh0jpjYPn3HEZzLtoa/HyksnwcYQ8Xfqc+vrJz64RpaQm/cTsaD
GyvV/TjZJATSPxfYpASamNNJXj4kvEhMHkqdgsahxG0zXqAeGwPN6Y7zL8AoVHzO
Yc5n4G6bSHFgGUQigwmSResJNAOFL2LhTqXf7fFP3yHu6V7Ms+5cx2gSRzkDceWG
Z+daXrIYRVbuNaKBMYDJE083BArwjgTUyhf8D6/Zle3wEGOQNOViL0ryV6QJtVUw
fdNmfo8fJYeTKV3xZBLDdYhRne9jqKbv/heWez/OzPnqPRADzOw0KK3SlYFYrybV
r6LBECF/QBe5w3du+MAxE+m0d8CuD7ksfxBggGcdvFAQOAN7kaNVCTZGSaG9/NAs
+ftfzHzQnAyXrEBI/CoNhGiLu8EJNY0thncXEcIomtrxEaSdwaftQ6PJ4yGSKonK
qB6uqyP4tj+kXlED3m4qGvpxi4AFVLaCRu8AWiBg1FyyEAqL5xcdCU/p1xdTvWX7
2mxQkavwxpQ9A5t3pluWr/dYzoQ0a/cUMnmWFr6CdklMs1B7Tpvg7dyTywJiY61b
kCf4rca0ZI/2bmW9467OVLJDYdxeBTS1TBsk3Y3nadco7zzugKwiR2vgtB8xqxuE
gLkrqULsIZlHiLmjgkGHSH6APEM3JkMhGSeYsNx0GeeyTQ68bel3X6AU5sBUIWjV
YO2f4/6XBUST07OsqAyEA8cqvcTe912bOnsWnDtOiR1ZM9HC90MX8AktVHIz+v2A
TrxtsyQtRIEyItH9EQ1LKUAWGynZK1QEAFfdHyp/20RGIT7BMmIG7rVI/i+xcWIk
I0iuQiBVbsNKAJAKas1al4DJl4WQjcpMaJdmQoadCIqmuvKxyAzi0V7yo/3C+8S5
X7To1h5LhLzgUVfzuvP6vu5LZ5n1LAy18TwT2ijFa+cNCVk/J9rhtvVE1CVX92zw
myxt2zqt0ynVIBjjBUzdBafbftKObHHe3RuBipYcCbEKo4Ql1DLG6Wvko0/MKELF
awhmr1f80EekBia7HpdRI8mG9MTI1R2IS4Ld5dCaRdfSoEkpllPNGhSO1XMp0CCN
4xg/h+cAvw189B2W1+SBvaF3kizGZJRJ5IMSdgufg5wuyfyQay/PmmK4VekeL1TK
FKgnZdMcAd8XLc3EbnZ+CFmmNVXRW+3g7NkmpZL0wzojTzxONx7L1E8aonT2G43t
ojc/rWZOJl1ysWZZ3sbYWVYSzf2KXNrfPjeof7t8A/pBOxynouGb/t95cFRX3dna
n07Xh+94cshVXItb2+bpE8ZtprgmWGa7nqOh/W7QB2/SlNcGkxl/a6q+wxrYDLTa
JpuGCvvCITymjCipXswwmdbRlDVoeV45dS3CmXArCv/2903C39SDQRvgDd+ts7bW
Y4wcZ67thv1RGNlo2f9dvWyYy++swMdh2YwiY6knSUZk27mYbHonvq6yiHgWzQwn
tiBgnj8qACi5PmFzBCjlbarEQ16ymjAexdHjT8c915Lv/ginJkDGIP7QBsaKE7DL
zCFg65lTqLiiN/yjNKxp8V0t/Y3eMkPbei1honZiXjSOe5e27F80eKMjDqwVSg2o
ysJ8E50ICf5XTjTD8RT7VHYmMd+ZDPi3OPj2i2ZFU2xBbHua1v460hWk4ZNQ7nhI
4bwtgWhEPsIJHqNysXxb15oCo2mBCYO9adCqqXbI9VqyuIKoXfqhyEQOQEn72q2k
MtxaHaur5I4322e+TUUeM5PP3hGaklxaTWSvN7R5EZ5DuKRBmCAakI7e9jP8mpQ2
0rzxNg7XMt9g22hkYU+Tkz+uHKRdc6BNtwFc7TeW9eFqcMnk8QmAwxKpBhVQuVAt
5n6hd+5Xa+czSU894PrC4AnPWraZmo4s8eMiaeBHx1MqvPpu52Idd+3OpvsyV0vh
RgiWBG4+5EQqreBZGgnLJYUiUNEXmYlNJPwP869sTsxgkCyrfT7iQ4pzGj6WfjTh
1uaaYWtWT6igU9ljIqALOe10asOpOqILjF0CKueekHueoQCyDc1IiphRvkye98XA
BipCu2e9l10kGJCGuof45PYSYuWcmKOPgOwTtKMYAzcxJe/ja4Z+rhHiPRoAPoKL
R02DQKRWOf15y5lfoA6lwddCD7nTRZV44esuoxRBbbbQqV6pB5g+STB+efDoK4HB
Mf/1sVzmlpjaIakDVhocTXQkq/0OXNiE8Yzkqx7yrlTEAzD+wXJF2823TsdknVyT
B5B2eNXsIOb5OgB21IwFvaBC1JWKmhYcKlYJSbZnpCO3ONCi2cavF0KuKR69NpiP
ocAI/eXaMNtIXjXb7k2Bb9lLYwJde76FLz4f9sCM3YQ6MYZE+Ny4v4x7V4x7z3Pp
Pe+QMUjEneLjAS16cDWQ8bxY7sefANicNvzOKnUW/Lv1ErRxu3sYjfSsM7cEplRv
8eiitDIU1iI+GcDELE366RlJsVaZYPBX9o2/ITOGqnWcDgI4m2aZ+GTzrKTeu84W
QEmv4OqWRPY58OFx6cgzQMOur5M/UiRZ/h5Gf3Ossh04vsb8tcctsmKusntVl/ix
3TbwOEtWZG3NKyL5k76vPoypLCoHj0Fl9kHYOSYa8ECQdLiw4eBQu20WD+CinD+z
86M+b093yTNhAjCGhy8QIJAGynkw/xi7MZws1kJ+HY0YmfYgimijHyCijUF5+kLq
ZYT6MmUZZ9P0NVHUNNZ4TOm8Fe7LhtU1hruR9FUNt3hFoPRn/Sq9zk4Y7WbaYRfv
rrZNXC1DYB/+FE6ZLMEVgS3SkeDPSxB6PauT4KLiheuoMn9+VhZp1ejHtMiwli9S
FDfRcqoRJOsfUFjHnksnFrq8EExiLNim5ytjjeRfT4t8BYIzvyDefwOybFbH2GkK
PNZkVgH2OWmrz37Yy07wO0wPTfPZpKVe6TTyw70SkgYyKB8n8E3k0EOr76hLA+3B
7UGtIaL2aiYjvxkODZjPZprW7voevAu+qrPUf3lnkM7WCrQjgAppjoTi8TZxwPSt
hyceb/ajuckmmYRdmR7IZ2upB36ZvW65RMWPAXC5kjLholPgOzuoxuDgZQFlL8KT
0xiVJ2CQBxKwKQKMBz+seu8G/z41b1R/batUt7Civg3bFsqU/fC+rfpwQSNexFqX
n2tTiIZs8svqD5mI9zyu7+mAEyBlkx8MIZz4QZDIpP4EHgLuZ2XAPqnZTVmG9Pmv
LvPjxC9IU9ZgUl2NtwRXk1bmgGi1drHFwVCzyQOGIvwk+zvAw0t3dgSjrKId93BW
6lFyz4w7M5fGJtgpsnInB6Sw3wcLoAoqYVpqetyCxchd79gAwhr9bAIlj0oQteg9
gvLuNCE8ql2ox/l1jvKEnq5FWHMCc+QVHeVrJONM513Xr7pRlp9jjj8QsJtV0NOK
1JP3Z/I57Di8qzpjnGl0XXyPxzTRvtWySgcnkZomUAI5FdLP43j96+XQqTHR9Jy9
vQTyg/Vaa5BWw4HpWC5A1X6lLTdRSYcel7xDd2TzLOcOanmmq66rW9PyP7HlnjvK
oI+go6A+rHzCSoTvUGOPBTY5/QqfRkKmMicT3ZEK4098u8p9Ed9uaQawMSIuGyQP
db4OvCXkHwoMpkHtNq2ZgoHN3GMQL4jDOMlqUIEILabjgAH+khoKuik+9FU65uQm
UPGOr1jvPZPIOW+VxSJUMZncqXy0ObltgM3npgeXtCo8GwtE1p2jmsmGJuuPBCeg
OWOERVSx+wxJ0N7VjN9uzBMrjRcEtEPyOMJsbj2E6zFkEs/BROyeHBm5h5DTCJTq
H8xKWWyfGRj/A9ltmhznUFTs4YRCKJdVJwooc1l7SngviznGSpVzpetKMThlbdnO
6MqYONmZi0APFno7r1gnSdCVPos0VPNs2MsGNrrz5BFsFX/kHXf6TNq0jZqzyX/s
rqb/gpKwdfgG454aGCDpJtutC5ZyoM8QI4yC8qRyc//jeeO8nM8n0rQyqf/FW/wl
xmF4ghNsQeyrxgBnZSIbDLBrrSS90mWsUV21K2p4Jwv0MKbBRR+bxm+1Rc1ukYtE
tjGf0h4rm9wfK57eCIayND7RQltSmcvD2P/c4xOCPm0GTn7XwuRyc6wgG2YAZb2+
BFRbOZ273/eg3BolxL4+VtbJUJ6ByCPpBSeMLxGQRuR+RG69MliN6KNQQGb1LiY0
VgnYHeqYx2CPAaxEoq+PXmZejAFJTukFARZf8SX9rkXdGDzigoEbPdEnd8Z8RORu
1qdr812KEapBeIzaMxJMVbEf1WE2tT3RwlwqVUFw8tLj283GboBT9Wx+5AJXcMGw
I3L3BeKV777S7LmreAtEGzdHUrTb4hOKkvd3qBlz+GItH9QUQthwxiKjvDNFwCY5
67Pck9Vza2renWCfvx+zlh4WDghEEHDrsy3Maggv5xgQq6eO5bfP1n4IxzJ4eCNX
4XH4sODfYfeYQy9hGB9rik83SphQIq3fF1ghoNhvuinvxMMvA/9TseuFgDBZ8/3i
vQyTnHty/RZVovux4+WXUJ8CNeUf75g5AhaBcT6CkOfVTF4xqfgABK3sClnvwa3j
vfm7Q8AkG1CZTOzk5Q9B1C+Y00IxysNh+JtehaLCTktoYaAQSaXyMOvu2vloNTUe
vJba7A+rImES/WZsikCFYrbYTIGkNCAArCJSxjhs/xRpx13Lhb0fUBoH36ULJaMt
NmQJ+qsjT3y6w2SGa7+lY2i/Z+X++GFsEltNwUBUWRZrAjusVmqEWUkM6QzdALdW
yoESZM0LxX6tqiepQ/sDeBOGd0im37zOsx+nz8EInBgvk934b19QUzDcMVCF6P8W
sNRyMpa/NbN4/gHD/DOa4S8spQBFfIZR5TuIzNuqHE/JDAMwCaYQrD/tWYyV8wo7
80gIC1kc4QFZfUAQWclmA8P5kYFqIfETGWR8iXV5PCUyiDYHXN85quhhz8jo7f1d
JsXsYyTikFnmWxW6d+1h15VIiFn/cEP3ycqdnZ3JZyfr3pg1lzXu5mOMlExD97Va
1FWJygfGWeJU6BImSF7ODVDswuQWahu8NzMKsSjCYZsLipUeqYBOBm8nCF32rDoy
D3dNyMKhD7wzHXYThUcFaGUnTlv+r3wlFrBKips8D18NRZcUn+HGLHbvrZ5yucOg
JM1biT5EbsKMzdE6QOq5yODcOAdeJazS8WosmQnOacwdfVvJNebBtemy6lIXwv7h
Zwmb8+JRiSSRbNulf+8Pje9k9fRsKitYuUmLXujHZ28bzW+46y/rsY5xr/N08eig
NtzYEyjTCpnC2jfHnTj3pMiqTGlrY1GQEIUsRlnf27n+VgWoK6cEMEYBr35QJYkK
o2LKVKg7YIRuCodZQnmgxsk7SRNv2Jgm8OrpeEcr5wfApXMrPW+DFKo2ptmu5OTR
H/q+KnXgFveCTqoCDX3n5ZHzFCOkVfeiMOpRRXvqZ2witzENSbYApyWaGNDtdwpT
8jR6RgT0cVmMupkVQexCnHcybBSh1j1QadT4Lz/CctxZq5wp3clT/Z0i7RbO7smo
nS/LnUpKs4tbW4GEKWeL0w5+JYQ5XJ3Vm6HuNEBjvzh6koc5AL3TCcTtEVCG34Jo
QKQKK3RV1vFyz2ojMArqxp+Xu6wvgGyAXcOu6JS4X7kQsoPYsP3xV2OdvzVaNmIK
86hb7lff//Xdc6EV1Av9I4bDVIWel9cIh01OWOFHdrfo7/SzZx/uyGn8HWOswlZq
KOnAjpuYnl3lM/VTin7Kd8Zp8yyZ0wksmR4vGpYYFaxgQWIYjBG2vBFrb5UmoS1e
xnFAnYApo/KK655aUkdrs4AmK50SoCoMz57maAZuQ73rPgPU5astqc0vhPAzxnmi
h7WnVbigWOTlg2Jg8aM3M8VaAIre+8GVYf+hRdBhHnhGamwcHhDW2ulEE4ebkVIf
ElDgOHcN88ggGjMHSQjqWqsbgglj8Xn64YTib7ogYW7uyA/8g8IJggbGXtXhWc0a
AlRW/dNwE2BSOritA1HHrCAGw1gh9ZlOu16oQNavyhFiFpwur05RjtXyRUdsd/XD
tyrzDVWMmZC3NTOfKwdTM0hCx4lun5iRVtx58SrXEaa2kjly4Snwai0dpdoOpQTT
jocOQxYGo8NAdzznyetWdUMwTyx+52hkg9efIuYT5gnibvVK/zeeTIOcxvdo01/e
WmKSF28+b45YRJcmBe1pS/wN8N4c3VtjHogC0jkK7uatIX55wLyq1Xsvrn38BYNj
wG0XhoC07wE8trXjEwQfFOk0hii6Wv8AV6HsW4W1KpjhfRR7bNXgG8S6QlUQdgkj
TnPx2TyiSaMm5q9/CRVjiZzMw9JjVp4Jf4iWxEvN7cm7te8Hq+5ZfvlOyIK7uR0I
1GF4+1Nlx+2UILn5p4wVHu7STnOxI9nSRahTKeSjxLIRmpFKHUgw1T5uPJej2rvN
Q+dZJLmr5eyPDjlM5AQ19kOVx4GZEoVpYdRjdxqLXvK+YY9KUH3SAEZZd2CT1xOI
dV2WZ30TDw/Rd8y/6q2URNJB9ZDNYmZmYk3meWU1PZQzk2oHrMmlBiwY91a0vu7W
/WCG5vU0NyynP9bdk+uKeQ==
`protect END_PROTECTED
