`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+048WOv/ScoAaH9wKVWFuzKBSKJMSxOoYUGfo+yikDnIvaGlOb2/MZezYfBpP6f9
8j90qoxajDFvMK9k+WszRG+MrxSAe35hvnqPfivcy6c/HRa2yOSFbvcQPP7KecUL
KWZf83tj+4H4OtFM+RUsH2QSkD+inapvYAeON/JUUibZTOIXMB+CUZkIpGBS5Lly
R+NvXLdrY/c4kF6ITOoeiEyhqfW09+o2oRS2KL8D0YebHxw+KRCTo6nB8vuEOGx7
RCiudvu9EmRwKtPCeUsBqZrh9Cnvc9Ch3Iwp6vEkqw2oUOLXLmO61TpzN0vvoZYx
`protect END_PROTECTED
