`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xv30bFpPLkE9Z14rBljNy1Nji3bT+9M3HvlxX/fVbl1JK1c8mYgJ6a+G2xuPRVoh
/c+aXhBpkaPh7JELVndU0WzVLp/DiaBV7t7d1N2GXaBqgNWjXHpk+Z/IEwGUqabJ
T7hloYscxVp3RH+jktS5bZ+UJpG5s/AN2KBJ+5gMEskM/aaj6imtt0U0rZAkmJfG
djjIs2AFoU5jtyBU1kyTML1icA1Q+GpbYOzCdfTvc/08wtE+kl5lXMjaKYfQgn4I
nwBZ0fCj62IMbCT8kRgd8OBUw5tXxuzKFjvTnh/bHzAipsQbN1oxmpLPLE0ihLn2
ZmAZKEdQPxkCy37aL/igl+8i9i8T2dn30YQtQ4Mj/lZnf0L1ip/5z4Giwajtc5m2
4WL1QMBeYRLijgsglPsqZ2Zip2XrDIn8/HLUmVGMnQx+pcRJpOqImgMS0M4TE4XC
2vvL3AJkUbmIgGpFYR6LWTVTK3/1S0FpZlhlStN6id5kJD37S3xmuiuG/zCwQIde
NC/4BKCWDkbPtCwaGGrDX9jQ/mvIsNmV1HPKGm7TLH8cSCCXHQDjUtLCLyljymsF
4NUYbxEwKT4GnTI5DrzSJJrHGdBj6WNbbSumAkSp116MnV6N/ol07Wg5l/BcaOHV
nixL4LDItvroZ7UUXpVgp9UA2BaVpbM8v8u8NpgqEVuENi7pRHlmvCz/MnKh6OLJ
/ilpLfYNMEdhIaFClxbQoy7cHR2Gy1n5qeyVvxfvk4l0c5yn/b+s+0jcFjEjU7s/
6RfTlwHqcySfaJcIibULVPV6Eu24MFVknw8Myn3yWZPvvlf2v0jKkywxWXSmOsXm
xWNzcUN8Nbc+2CSplA9X/d9IVRTkSdQ2vjz0mRUTCv1Uze5WW06iGqyx0U+PVlXL
26K8YdTet3hrzsujthbvTIzBlfsS9/qZ1CMG76t+z7sJZy8bTFsvZc6sP4UoFPRJ
35QPJZrFrqG7jDmAcCr5zB19dEZHaHopBWME4OopakAd0HYxxJdjmhjAcihQCCq8
HCOWWPJ7bBZPWXUa8Wy+3Qv+NeRMivwZu0mVxxTmrdOO7zYm4oKOWpP8X40NvECn
8wFZhSK5/Y7fhxKm40iG5xY7ICzgdgciYY/NtZrK71xGDYhGYXaZUgLuasjkZbH6
5PGCxayKkp+bRXmwxyUEpXYcqR0PAj5KyD6btYX5D8L9KUPaDH6RMRSpVfV4ekYC
0mQZqI3vr6vo1IkURoLimsOPKed9ESAaWxMYCMxhaR9yfSQGiWrDt3euCLnTpMDW
+v59yz/30JHRV4YRckmsEg1rzxBAGxnlN7Xuu5tNEgkRLRRPouPaR3ggPeSZWUnT
MTqwaZq/GR3I+UeMWzdJpppF8YhH7lgLE3CYEaDl31PFXNRaZZCJazKU96jD9nQy
FxIDcO3/c1ZWH/3oNYs6GkCnQeRrVlmevmdFJmVPXrFjIh/XZaMjI5f4bltoqddc
w62hRII1qZ4+YbDlqoN0hbApgXjWCDGe61dqZQ/3HTI74ASvu9MyLsW0Jk6lNeGJ
3lWYpYhlvh4E6GcegxihdrvWQOKbc4E3Ql2NldN419hpzEy5DfG14/4a64bhk+6l
jOKkzlvWNbr1OhqYVm6DNLb9en/QX6HQGBHVoK4r5XIXhcE1mz4MNjfeQNQXPSz8
nuu0raY1K11KO6fiOYznUHe+JNRVGmBTb3LDxNEphADwmIXAkPhDySgZdZlbD/eh
U7mMpOkejuD5FoN2DZ1IE/qN3PFI1OUD/USvMu3Uj8GQPTX7pdP8xtZa7c+QvZhC
3EvwfhcGzhZW8bFXtVowCExDdG8ajeWGqW1W2h84vWh5hj+PtD5E0vK2VaQcLvxq
ZiyL3AxYsYQ54u+FviQzNzPm7qU83VOtyT7CkDMTN5DJxrXbLew2c6QD6EmqO4JF
ddWjecDwb+TPZ+2k+qCtZDnkDCrXvUeieXsBoUg5XovipfKJXY7mQQbi/LzG2KIS
0ssKCH/KDi5hQEnh6jgVVhvPxGB6ReYDxkQybw4Ak8YL1b5PRImONfEynMl7/Vve
ACGUg9h/AikvWcqofvmY2NwcK1Qc0zheaB0lFfgZVGWUG0UZvN4bu//48JYRvBYs
ib0nHcDnpyolMPL3I14AhWR1h1k5qja0ZWUfyP5J9tI6lG9UljfaiemY5UMMQEdn
Zys0fmRZ9oUBuhQaimkTLlqWWG+TvjGSS4o0JlykfqVDgFMQUh5X2uPxtgJ7/4oK
WO9lY/GDYrPwgeZBSOU2Rtym5hkxKFOLnvbD+mam69fucohiKEnxgSFEspNqHiul
3RUqN9K4NO4p8F/LRTlKetm6SdwOtrT/djw+gQZsNntQ/ZvwxJi0HiJbTvtkjTzV
o+GyZLUkBbimXRRfi52szKLPWZRI39Qcc1kCgVei0Cn8ZsfzI8AAqmWpYma2p+eM
FRNT1vl6Y5eC/0hDHlYd/0KQiYq7v5x54YI+JClITThfYG2Yv0nUjGvXLT58QiAo
eeAILZxGZpXsis1rM42oZ+j8g7WJqoMcTjjAFoBCHAXU9gExIuU85Ou9Ty8G2q0x
/L5kfQpwZ5u1hLCpoV1g/rYHDiMxh1hbQ1tLYfPNv5SX7GwWDYYCZyCP0kEAMYai
ibIqUHRnddRf6zZh2idAfHmEgiQ+DZewdqLhhA9Ge+WtaBgDrUuEEdRAqRzS0ZIi
e3wzsMhIkZGtDvCLvUKy8NO9tXarK7ldvZCEPmI481xrG6y2i0tuLoOWMkYepJoV
3gPe27Cnxvb6R3XBXXEhVVYHiWrCDUeCNghLbjDMYg61j4dmNmsqyA0+j46reFFN
8GWvgkLEtsCiIWQFJqsG8FRo7OpC2vd17xWx/0I2wOIQx4An8HP0D+wFLYlHG3nK
guEvoRHCFz1kOHoAGFu8cZEmKWb3KdoK0wFORYrkc7uMeO/xctQ5EsVZkG8W22lD
Zbq99u/aF5IjEWyPn2RkxLYm4L/fmqDcBBffTCTOL/PtuCQRvw9BqmVNrutpY453
kvMj6vn93lpA1KYcJ408yUNDJ75fk5YczVUVh7Vf1Rpf0ai6A0RpPhFnMpO8uTJa
OP3FzaGCZsmYAKHUgOVC1CNLByyhoFVeZ1lW7BKSs3Q4xyoMktuQ2UQPwFuef7Dq
MqtpQWrcPIpGcDM+HlCUFIo1p04X+y5tJE8horbE37msdSvklDKMu1tTYDrujAKj
zeNZv0iL/QYvOed3bgT3Ae51t6G+e5CVq4qIZ0eHZfIXx2dj3jmUqNOQTKn5nOzV
7WKMFHrMh+iGHFnz1k40ETIsT8nx60CSg5mJDjJ3Qh72zNf+Tsbda38XeWqCsdIn
reZAHYRO+xeBo2cdXQXEGGQT67vCuax/suatgjrp6zcUVl6Ak01KIzifQMsmGkAT
/dHMb89Bks3G01OGEmnR0vxsmfrSLsnzPAzkCNWcmadXPJzGj1QQ2+86Mth2uklY
LxGQccZ3j2rsDAr9qrS+HSgJJlMCyuhuPcvnasoUShGxuQiYtzkk5FXMlwE34szx
LsUGe/RA/tWWfYZDu4iy6Dokqz33wJdsbSPdwbLKDgtYU6nFP4lpdIgqh9T7Ijnl
6hC6K+4sQ7lh6OfkasZ3aQgqP78u6Af4UhGhiyxntdVYQa5YDpjDcD6W2mmeR698
obWXIaF4E/CSJD8l+wK43GgcjIh9/X7mTOS6EnUgAWA+oVjgm/F5YyTqcCHPzE+1
y2BCNIpiNicJtEWWm7sMYA/ibTZi3rVBMYcUZpEPD/C/0YWBBlXiQey0LzRD6fdw
vaxt/zxzuORTnTMa6ltPt+NZVOAFxaKXF6vXuPAR7sXX883VHytvovpMDdTFdzb3
b+OZPBFtTMpSx/J36sufMMgV+kGxae578786i3rEOsaPXkAiYGLBj0zlTUpPj7ui
FVABOLDOqPKilYwn/2GVlg7T6juYbUkF28FBPq0KSy3MNnkgRD7c/GTtZ0tw5HSw
NrMR7yrhy6qR1euolu3rpaUkmIeVfJMbjhcRVHppzSjcdw663YrblHCmrU24Z+kl
Z/CkRaEaB1HHdW2sca+c0GAIxzf8Cjiy1/nJmVSm64PHZL129Aw6bfI8y1jLncJF
kpSQ33BzX8gLjc0bSncVxgXu0lBYir31FTpsPw7bPRUAijWomEVPp5xU5fhQyZzz
uOOj9tEjErzfwlhovyGEv2b8DS6aQn6lQHPCLQxSY+cTxvnpkMWynafNtHuhO8sB
PthO906WoD6uFzsH6GMu7Cs4ATKy+EprKcVNYbmQGMFB6IH0fL4QCTQaXOYcml/k
xnKfVJ+AL1AeG0B2bIA5IVjSLOqODYjdq0ESWEhShe+NFeu5S6By/DX851Xg8zeP
4l9XmO3Y3uEXDn2k3buLouB+lqT+oYAb6wB4j+Hy64LL9vE5sNDTfg7/IXxbwW7q
Hjzx5MfZ2SzcSSeuZgkr+x9+wVpM8wTctkM/zp0eoRWPC87kx2Vtl65xD919JpJP
eZvqVu/HXANPJMSFkE8OS6w9M0V+d2O1Lg39Xos8Xjdj1uuf2a+EGiJCmqxgj/2+
cJRbt+HpW9VKGZEQoRw1gN9zfIb5/KtlDKpEbTE1joxYNf763z0GcaWkQOxp1P3S
9GPHLxxwR2EiE3BWiHhrcAkV1QI6586Aw08gV5hlYDblGvw5XuhKILTaPpuDFCgZ
rn55FHlu59HMi/9hXVcLYfTeSuN9KuXUa3YzzkknZC+FYC4L8csxxlAlLrW5N7gN
FbcX4gjnJhTR63TebWrJOkLA6/uOoMEzUmXWrfcINIleM3Ij5ZjRHXSmLa0wx+K4
F+IuXeg4FbvBTIn6pmn94cVzus5iRrT8VhrAvc82ra/Gc+M8LPzr9nmBGMIxnKDO
XfnMUnkAPnM6Lnez23tEc+bMP0EIy6jEB1nfQ9hfMQNs495oU6DTjWLC7QSiQyCG
BhR8z4RNscN32WxO+lrM2Hrv3Xj+zI9JjhBEoWYzYxaI0KsFCouoKIQ67oqXas6v
OyQ50erj6Cgu6mLIzyL2IsnlHu2gLUGKIh6ei7fRAEvfNuZ35mhtCam0rVWpPmWB
vQlm9MLfbBjeCQUvJZByYkLM+ok4r4yWCrbEmsxvOXIVqq5ssp7JbSWfYCqhnCNq
MJ78rZ8bXW5RAOIIxYllAJvRc8HHRF9rBWXjxR633QODbWb9b28Hf0CwaARW/xw4
6fPYHkY/Li/5bJkqex3UViSoQIE1rNw9SWWVcH6pv6E2cO16tFCT4c0YwGKpyZMK
GpSp8BnF8ZPPIp2TydyL/WiOC47gLsTewC6aP9YHgz9jpHUmH3o9BsdViu218jaT
FOxfyjmWqz2SmsDPrr1oAMihVYnx/4da7gwlA3Y8CTazET3pJSHZoJcJceD65O4h
nYQ8bxTCZAzXkp58ExCbfS4+i+8d/3AjzQUE886MoewEEA6LuDZjd7Y13moeSMWW
VKfarzvQCKwfbBD46igfezfY7PdO3mxuuvBpF6XWpnCnZhOgoZqp1BHDo2F6znkj
SUPxU5f7FKrPMl30QkMuevf9eKFVEvedvINty8Ul1sZN3X1ya5cslRtcRVHWuG9F
kqtzTAJi9z+8Ii3gxMbclpoePI6zNpG7U6KFEAtwXiv/0EGtqCOv/ma06F71pVHv
Ddq3f0pklcH1tQbnFfD1jQS9i0NC9WlAXYHi7YNnncSm4rxYRkutJpIrMoQS0nbV
rQISyZyOV1DfaqjThcfP2OS9RBYVt+d74Nx8gfKMIKe4Uxyxw1PqBZh3mLTQFMN+
m0sGayAhSuH0qAqcUmIywta2dF32S1VNQ5BZrzq6Tb/vZOIf232uIxQI08Ip759T
Qhc0+61mxIDHmC1CxGwz8RX9OIKuqxnUtUjJSRqiubYKWpZURVo4TYlTBcH3VQCS
QEIeY4WjD7OwRTP7weKQr01JlhuaP0L5A6aky7gzDQrMuaCfnkfKiZL4uz7eZmde
2yZsnak7p66OX8Ixd7nfeu0m8FtA39KATKYU8lrMHRTZE2OSkwKcBvIzrKe+1xXP
uakBzIDSbfwaZi2Fnp09vY3pzOjUzCEatSYSX0Ge731iY8HZUkRmYn+gI21627bB
4/pIe6YQifKLxHKjp7Nlfa7VSv4yb/rZDiPdTL82UR0AyLGC58j+U54vtxnhDIoy
onIUGXzZ+ai8hOe9Gpc3J2tHFcPLNEAUaZYRmXNrowjuHJiDIGOtuvU2iLiyhJu3
gqIrW/nBAjCfzp3gFjsT33VfXt8ikGFiVCGO+q3rZf9da9sfRRFcFGz/4oX3epsX
U1l7q3GMbBOw2IO/m/K/iRaWK87vDBfdS0izwXfDOvKp+nkY+/pFLsePaM2pk7Mf
z7wdGSajN/Ll0KYEAvivwA+bi7XYiiF6+txVuAA/297IGAHxSfRqPXawN4gaZib3
z1gQWBC32xrMRQcdOwY4qez1cs2R/ICRFnsXE2T7Q0hVeVQ78vKM5SsXVPAl8Udn
AaLIF9xT88sUjxtL0y/0intBUg6lugKVbOkastCEFpp2d2tJt3BB3EtD0xmD8Gek
Q/5P2Zi/+1Kiw/tD6UYZYE/PoRTFHyYYOL2BvgV7OhAJ2cSdpFw+Ybkka8Roj4yw
g86IrmOu+SvlpF2KMXjQYsYOIeHe2jWTUIQG9rne/LjP+WY5COnoO6JrGNmUVLMu
UQV+HPNuPK23BU1xhGQg2+AWQabJXuPHssvsBZptFk8EYGU54/9Exv+KzmGocDwE
cNe0npefHhToC7iD6T6ff3Yo0uSg0CEM9vrlULJuHYVGMqRloVG9q+2UfkQuT5d9
vX7FEdNp0+0gwEm5vh/PQDPHXRjr4wQf0UGl+DESbMW3ffPFj2vKbDMcl2o3q8Cn
rBL27PsdwFFMJd8w40YNAygOEtvawiVaMqDasDGd8awYVI5c8TA2CAQJ6k5Us8kM
vURdE4CEFm5cPG3/mGkr/nRjxdabChEd6o1pJ0uoGFvAl0zfqusET8smLB+vYSho
vAdAWujizeJbCxIzn2fv3f7yk3VZSAAekIQvsrbijP3c689ArZANom8SxWbevpC2
dMc3pymURn1ZZjLn3hs8lH0TvHy8L1CwRYURHn87qRYxk9oOf5kRawI71uxcy6D8
ZZTeJp4CmYT/5CgEqYi3LtJ9FziHBWFDEW9Tz4d76/lZudJhlfuT2bg18wlMk3TQ
1jBx+dOG1T7IBLGrG6IdRA6EvjeDY+RPaoIj24vWQrGwPR1D0HVh2yuGDVS+cuWZ
F4DCn1Djp6ZXV7rZewu0/4Z6Gh9wIpIseJ49x79saX9sDUStEY9bD/Srx+KfAPTR
d1whtdv4oHQ4PzsID3IiOenYz73hO8K0/S/GDsYQCeNOrH91JoSUAGq9lBzdlhi7
LjAf1qWzT88MGov1uvvNibIt5d+JZmnu8xoh3VO6j+a/OIY/t/4jHfDZzGPhL5lh
/SHB6+CjXt4JuPA30Xiadrb9MOWTmFakrOKmKYBSS8RYzIanfK/HogzTFTGbI+/R
vKEUlVLyh5PE4anrlk2D+tjNRRq2LKnWPH+XQSvtD+2CM14QJSsdT+TzygS69T79
raUxMNB1EiTGZSowvEpYi0bpe2uj3zRl9EjACJ0ndTXXc76hUdQP8JEBuNeVNjMw
P68HiLHIYgpZgXUf44dbX6C7l7EbCHH8OBvAibsOxAmhSDPIhiWt14xzE2Nfy1es
XMwaslEgycfbB2IIRHBaLXu61ffkayk4VWXUX1zAu7+LYY7hz6sQCWK/qGnVmpq6
Ohoi9bwIn1/gNP4yDcAGUACrUAbatNvtSdK4SWv9g9U2YS4rJoMyKokZbPguuSs2
pfNAMaMAqOYckeNMqA9fXInR8SV3ejjme2e7h6NMyneLqgDALBevDEp4L1YLwWSx
TkI1HuYJybggVcbuFEjiV+4zrrYl746pCFCzBfR3RimJJ2fWSPV5+UEchpNH1AvD
03iuLANF32FSHzyc1D9UwrfF4iH3j/1kKj9KW0xYb+Dq8Mrbq7mm+utCAgHlGBBh
eVZjbuKZtaqgTmw9fKqVCqxOfkG/RvC2Laig273/UW5gHLTBTLFGKSJojEg19daO
1cbwznq4YefOZfwPc9vejX3KKBlLhpNinK+zc2R88wTWZ5zWnGeBHDdZi6bEIJdl
3rUczKqUP0reM/2ia1gAP/E4CUsqVeA/hu+HyHncY5iQ9TeU0WmY0o5vTjN0mfDz
DxjJNF3rPZZNgyBCFe4JjQWGmCxQR6AI4U8o3gZ6Tstl4ejKcwIQXkBS/ZHvAWuM
2oM2/smTgM5Mfsos8jIgW1cVwodB/rtVyiBUG56LaBE2Cc4ugbdAuzIEMeBdH4tz
bh8gt3q3kr3iju98ovn+yTpJENT+PzbpK7/HQbvAeYKWYH0biGoHyjcug7pRhbs7
MScf9VFNoFiIzHBO1+lJUvcPVQGvGP+Z6lwY8UqCSctfoNZ5Wdyj61DUJasvai+w
cPhBdOM59kJJAp1Pr4u1+wj4nTzF4Za/SWhayuUuD2gCyKyXfDxT3oEDXQgqjlFE
VGIL5X3bAVg0hMh1OLEP4aqDZhEr5p8PxwQIjB4AWSS09SjMRP2QDG29T+kz+G36
H0zUuqBtmWRXuA6EHpja94NUKncBkqnsWBh/bF7ae/BCvgU733KhwOI5IVKozB9u
oL6aSNxDp5T+T1GaVOYxVQAM8OfNjg7tG6qOXa0olbf1h6YomW4IiNcRei/iI+PB
Rzh7tZP9XB6Lm0rvdX8Ur5UnD4F0NL55sOxrXUMFJK1y85T9XPaNrxljiCZrxr0f
vcDaSZtt/JXW7kPrl4ZVP/jXnbGkRv1vUoGs2n5D81iVodO8fAKZz92c0StrEm9h
7LrVter2eEXT6pqR8zw6Etg8/KX5Hl+CG4tBhc0OoRKDazoHLz6N26J5KxPYcxr3
uFxzkQE3XDrz3tr3kpNfFVz4xLn4khWKvuZFf7X1CzQ/RYZGfuCsdv7dGX+ET6uX
k6C7rQ0o4qtZNfSODi2Rk8SNCza+r/S41jGqIpTa26f6qxQXke0cteB64URXHicB
VairP8SHK+bNRWtG0i/SvJcxWVOClFWbVPaSC9stKAJnhtPPOJGsZusCg6X8VPzM
EqeWXogK9EnZh1G9rym2tsxfSeR0s3aq3Kiv8aojOuMldXcxp+OqtmBbHvYl5kk4
Dqcuix4Ma3jGs2AMPQvK+7FRUg/+/mQ0+03Sr9FFrMRCkJeVTZtqxxYDnBv5z6GB
V+3y4HPwl+WYsgJjfoSf9LQN+s5C2+aQyAtQ2ELKpVyUJyX0U7A/rfITlQUm2F5p
WsU0BoiEZjTJj+Tqsb5A6ZPCkv6cSrc33w8nmSjrI3jYP4SGE5xPmYHFb01t/44I
GYTfFxwl2zeZb4YMSGBn50qYmqFCgXGLGa7fjiYhzZPRXqRdTuwYAzwFt6gk7NH/
SxaVrQkohzPSMaplTMYsmpY7A/g+GFQ664iTgLgYQSjyE4XrCl2BmsmZRty27DdH
7PR1Uwn5KTddVt+USuyM+rM7kSHqLgka8UpA54BSTemKLN0C2o+R1i3Skl50IjOJ
OPqYecCqQqGeLHSWZx0b0DvMBgge3i072Wu6PCu0eVdbHy0KPMf4J+O/vsnJhO1V
L6+wh0giibjz98cw73YFyc8ShWJvXpXEACWKnGs5K2GNbyy0SAvX7s5A3TLE5gRT
AjskpnDVa4ssYoQpbIqVsZqNhwLGyK7c9fu8H6PjEcJwAYEgCnUNJYrq+xzhTWry
LNxWLVBDcFO7Okvvzs4YMzOAjuCs633SuEkzrMEIx6cKUBN3g5mJrtHTGt4Gwjnz
f5qsoJLmtnANYfsB/fC+ti0BXc/muqovqLyZMmg9nTae4n4VolLVbRzUEHk48cx/
q/9EFzibtCAmk7wDKhlE+ZsOmDwia2xqGjPTd9EPWBUR0XH/eElCZlDVZ0MpVhlZ
bnfUZZDI6DtEvdX8ks55LQivdf5E2JF7QF5DP/Zq69Se7stFO+6Y7XOtZl6NJjtS
d4Znuxl9Tv1dFCjjaV41CTqQVKfBFGNXU5iiGkpWZxIbFqIa7Ed5/ysPus0Iw71J
iVjdBqjeTxq8zKAwqmud+bG7gtWTbetYChyrixhVsniwblvXOuXwEdOF3cV6AGeR
0LZo5dBIiVg1Poz1az6KDbAMGfETFgtjx15FByjkvMs/7zd2IasABDPIJE2nq/5S
M6lXeY+03OecclC9/cRjPnNoG3VoUEj7BXvue2gwgD2hQWCWkbw2W0unpU1DkbnW
ySTDb/nsT5gxioHqUfpkU0eXtWH+R7n1O7MhicUuOIaiZqlflagIv9tbw6hri714
+phs2MzdS/gFmHE/0+Au5ABIOqo+3Dsvma4mjc0zeQoUhzdXSxAqyjN5ICpKCtWT
AKuQ8/bnzqdfQA88H18MHcg1VTsRIjnNJLZVAtY2p25YingoGRH485pNUExKswnK
kqahB61C1Wug5bNEuaFt5+1C0TCspBg1pdk4SynlIBps2YUyIUIgGpC6ClDU9aQ9
PJuTYgSLyB2pH4J4Hp3HyfQnJnVRXDYg4jEVEEXCpDNdb3XDUGxZNeyQDijmpzjO
sZRmUh8ZQizLea8rwuqkrq95L/iRUJqWgw3QicKnaVXt+wkZh0XsTP9kBnKLa3TG
iS+AH4+eANzzhQYOHLYDyFxadq4q7MLjI4N3AxB24ubEtaH5vy39KMQ/P6JfILCr
/IIXzHjfm1W/a2syjNqtN6Zoe8+b8L+hlMR2DJmYj4VO/phkdV80V6OemYqijVUH
HhVPkmsvMdkyncl5vngBQzvZRj3NoSg7RwxQ3ID4maCgfW44HZPjAZhzkJBbcZA6
d6q37dwKs47aSsECFV7b1Et/QRgMt1EYdFyNKbYnIVmZ8gtrDg6YqSntn8ynDuGp
6kVWx8v7tx0RLAV0OfPfXZpbtkt0ljOk94ZCmP4Th1KadLfKps8ntPwZWlSChkWZ
n+fHyUMRQrHRNUmvi/pCOBPC4+RRWegxnnMfqfloZMaBsIG6pdzx59Kvwe3M/6Wu
Hws1hFwF4jwoXdr610SvEm9qAsW6RMtOZivSJ7YIBh0pqZua1Ue1v+GwEeXmNRs1
KSVt1cvtt94w5gQ/VIzektbfmY9NOqFhRFYG1SmfLnmKetMhu3+2XCHerNSEuXY/
ibFVrIVPgOoVvKr53mqFuq3YA8EndpGWbuTNGDC3XPsfIXD58lxAr69sKpvI/W5x
ZAkrfkIiZCOknmCdrKbGDKiTHhjprA/6dkF3toOsH4O5wdOS/VTpdM0Zt8kgBC10
a9e99zdpPhM6wcDljWvDQcQtDS1GB3uiq58D48N3A5M3O75AVTW/fsFGmV8N4FuW
NB01eblJsO50a5wkfZ+68iDWDnPmI1l1GE47XM/PsYzfV2QUiEpDziPOsIVNMVta
HLLacWRXWt6EfyMgEO185PmOLUp+YwJI1xroVrCN7pBGAXPGz/bIpu+OCs6gWFw+
07Sgq/sw3bUSOxOAa1DhQbtfdc3wqjgCoaCIZn1RpX6wkgxO683Lnp6tYiaaeK38
Vwb9WNTlkdFWBhQeaqiKO6nW+KvRzOs0XKy1Beazk33cFNEgZpn+s2C+bHOoWiEN
zkbWflcbm5RfRKAggOatv2mpsZz1pZJQMlr0wHp56xsgCnoLzgdCGKPlU+y+iRFh
1tcpiBI52jFiDSoOGDXLAYefYHie4TR+zsib6Q8M2vZ3b74E110aUHlM9410OEr6
/imWdLBymMSDm/KzOJpJF1EJsLLeZU0g8dMNno2NrzX5RpmqAl3fESrPshwAtl34
hpcoVsBDDgaEqUU7YTz7MoCtbCoqVkRqN4YDP8DO+xsS/p7ulbHj0JammCAF3sOz
9GGPxRkkzwec+rGTv1RkLnRUdFNO2FIuwy3VCM4/vp2UNo+FPi2NH/IK99GaPGQK
dCqfMkjkp+cyoesvPCuF+rtfTnJuRqaEwAHL3ld3+xFuus4yHjmd6gcBb55afF/D
p8j4gxNiXKDWG6KynLs70YGuUb4XB1fkC8AUvlOMwo0rzXywBrrhgKgXJjMEvwRf
Ijq/1YSw6leXTfF0vhlMGdP01Wx/0YLWU7NhxC+MJFxVu0LdmSGGxX20Ox/9OzGQ
d0F4OBN8AnpLTOHlcJvB8UkdUtTAwCSEr4Ht26NLn22vb7FsX+uv+zmPfCdaf9Z5
3fDxTSjsuSZv608ypQpDbROnpAJt7dw33Tkh79Drcky3TBNtX9eq3xsbkh1Q2/0t
ESxJ9LZF13DEnrpZB5CIyNTBymKfHLf2ubLuUalaay8ad/0zy6blF4Mr9Qc4+NyD
GhWRb4fq9qNQZI+B0sT5Lj8/ms5zavoZDAkNfqon6sq6F08Ks1IS+CA6LnaPYLLB
FTPLV1jajCZPjO4UOtsDjgOHG9IQmiPAVFx2oyevDJScm6Y6AjEmg1o+DN2rkqy6
c6g7nppl8KrTNXqv3dD3BZw+t/zJvCIgD2YsKW4ihksH3pgzGhrijCx91hT2NuDO
IAuuFd50bqyUtqPq+AkBvNZav37oA/dVHt4ABaj14fzhHaGekmo7pUWeG1Kk/TSI
XL0ZYPgKw5TyTzCrPZ2LN96GA5uxq5UKhKtUPG8KApyhuaaFt4IykDbmwx0dPj+g
+YWyarVinRxF3JVXHAl5pVGq61w80F6nEmYgjaadigMyiV7Zl3NnD4jNQ9yhL8+c
qZ6wyv7PlY7ZEdN4NXVpVzyPz0ao0OAplrJlHj2tUUXSvIKuzkM2fAus7V1T30u0
sKG6yYIhpNyKzBMlKacVg44PLbGqj8EG8fr+CnCh9h43L3MnsoqiW4DemR/6InHZ
PFcldowM0IFuYBjWwK7RXUvGjnf9bJE0CMI0cXLtHLmZKq0PQfyeM2iwkE5b9JRA
edKTYf37P9hRlUCdZ4wPm6ykjdBpLBlbENH9/iC6OsqcH7dvy6RgHU3T5ub9vqg9
lPixqb3kQ7lsbK/UsuW9DYzhUa3bTuNd74kn7E/zvnYxst3WOF/Q6VnLqeuT9Xsk
yl753DZUaS874ZbjodjKAn+d/2/XlxXbqkzVh9Q/PV8uMnlawvsxnJbhAlwKrXYt
naXf19QfmX85plrvmHgrFKSawWBn+Xh8TgJ99FAbvJ8QWhelzjY2y0LwfEDb9hly
2iDKfsXEVRU+FkLurZ392WBtO65zTkLij4yXLbFv9tk8eiyEk5Qkvw/fQ5fEq7hm
EPJr/ndQ0d5m8+0dvxDOaSW+EjwWGsPyWMBD6CjJHXvs0Qgdd+pznNosWHWTTjZe
9f5wxXHubJ+KRHZZ8Th6FtTSeulUOfPQaZG+AQO+iFrb0LqcycfVYSLgcGgLJCRK
DGb/q31xGzNK/ufgSQqSorgZACnUTxbo4m5OIkmxvNnlYO2nzx1pXAA9ZySNMU6l
/eCprXyA2ARCG2F5e6mhHQlh83sa9ly/DY5ruL7SEuobDF9/7zRncuc5KKQE6hKF
OB7yG9HrcWz/kMM2zUr+Fglv8AEPuQFWnhYr70J5VVAclQ2NfzzBmc6vs+zuXwWn
ElgPrFn/beIKZTsLEwSgTbHbD0MRBG2xmfy5qgS6T3C+npXSwnRaQ37XfMxcHBnh
3G9Rt6TVoA4wI5e8mMSgRGoroLmXHXRnVVAF7O/+hpp6K0oXNZBRFXg5Nc/bg0n+
K47DHL/qmlJse1h+S7u8xALyECnF2B4+9dgJz5PDqb0wJNQDSnTpamTFfBUx9opB
EBvESVqtF1xP7Gudm4Hf4viaocxOqN95ID1c+BsSbiM3pPvDbGo4987h5e3NB78/
qkA2vShPKVRlOxeic4tysB98I9WlZmu0WF3QNLNEYXYeKOqBt+kmkcb6+0/DLNke
1yn2HYxzn9XlH6PzIztB+Ek7lPBH2iG4a58faR16y0N7J9F/ezmk3mjlQoam1skz
SZP//TDHy8SNwOcpKmyjWXOGlCxKr15i6npBDd4IgMHtYKhxmNO7a70S8OZTqhnC
EIFCFtjJNTbLA0PY6fsIUBXIh7VZTSVH8ACIN0GUPVjeLL9H6nOchhFr/B0VNx0f
vp/LccQTSN+s2cYryeMC2CfJi6sHlFAK4wsAEzIdE6g7HsCwRaj++NWov05jhoFg
QCqeAj+DjwdR8j8OaHR5EX10xEIMsYq4+S5bS6w3KW5h8dFYQVV4TPtox3usRoJr
dtixovzEhzMTuaA3zfAKCUVVt9FORimEvGsYZBO9GxVFWWLi4cbFxo0mukXPR7Oi
XSqzMNkBd/B3btX74TvTPTs4I7fVvvwFyuOATSyGxb4Q9UCUnCrzGxeMmLE51TFW
ZuLsz3RL6ach7/iX0w+CDqzlbDKb6UqibjTTi78U556/mM6eEltcNaVVIw7IOj/i
l8TewakGJk6kvqZIp4F0i/deKcxOpTIA+Lj+2MIZo8kjjwq/lnqDMtu6tCLb5dx2
WbZ+BGToavI89FeJnGkoFNs67hhbBmSOQ0j1s/tNjZGTZtL2Wl39wGboOkbGsBAm
jDXJgVJmAjNteuisGUqZXg3GJyYPu67im9h3lvZRUI5SBEOoFYWFOjmuZSjGTmj7
PXMg4mBBnSyxkbCBUjucYg8E16PgPZqcakl7fqiZ9q20mprCS0KGi85QTNNVRFmB
K+Mnzctx+pxvCXFXeMVHn0uOgMdkHMNVDHXhlyjZcloUpi27IH+DPHEeqDeae4ie
HIj4DlGUm/hX8ZAY4RzaW8K2RbuABoQ1kwEgVO8v3X8/EGtsjHvUr2Du03rXY97v
pz6eWEPAJjAp4bSpcDg/1ftZwXEY/B3jOXbkiVz0gvRucy8jbi5iOX5RcPv6FQZM
LsWQwW03M7dgT32tPLFACnRtA+sG5GuTTJoLZ40Px7f/chu3x2H3dnWv6uJeACsq
84z1wQqaYwmV/vgML8b8t5uomZRdS9Pf02QqGjI2VdwTYKtpKblOGW2fZSUpCp7C
JzNc6iD5aWH3sug7VZ+k2M8VkrYQMT+Crr4s9LFxQSHzQDJTkyvEOVmQt0xPiJNl
Iz2veiNvLM35HqWpKYQfdagpM39RQex1EtBUSKMFDEL0HPCRfEbueGpXYca+nthB
ofsgmUdOjRcXl0QIlGx8ZEycJyTzxcQwNn9PO/TzqopQkM5XedGfbPrzkWXw5ISh
ULlLPaf4BQ4GtgPVhYPZaFj8HLlt86qeaFBHP+LyBrUD+XdTFv4TR8QYxWd8AJLH
BtLmGOKHrcMsY1LIM+R+Tc9poymMIKt624U44N+VLiIj8v6mevutKqZwrm2FrQ/n
a/dddViedYYdoBw8nEzbJXw80iJo+Xbf6neZBDsdNgLjnssOniaEcPo+SZcGxDdO
vy93Edd4pOfrD3bf/2SPF5g9elKtD05y5vAWFy2oz1hfi8wneQlO/YqZEAT/rojV
/PJzdWIhXfLQ5EWkwADl2K2+l5cJVmn/KDs5R/qmy3EaoVok+7hFyL4T9D1bu1B0
0fMR68krpmP5Uf0o5EtFT3eu7GXfg90paG0QaZRsTzaUU0bNQfo9gDFj/fxKRDDF
PY4fq/nx1aHQpZvi33qgCiQ1OkGYm6ZaP2uAscnjFETpOcptRkZ06E+5A1MNBYj+
NtQxCiVn+RryZFaRFaC4Xtp2IPvhZpq9XzgHLY2WbpsZWCD/D2PLDuiiFs764VPU
P28g9mPiKK7MmC8BGsBF9PSIa0NcetEb+BC2UlY988iciKTn+wxk5C5QAoYq6rl+
dx0M1uA1FrpYMTDrRAuHnpS20d26ei5F8bKB1F0HvdPlGGXAItEpbNHZOpB6Y+an
pyRfZJDgdzBz6gCouJZVMJnh/KmPEubxeay3zybb3zHFzYPTOsUoDfMJPbTjmxoG
rExRrczL0h/jkxv0HuFfXJqlmm1H9vbXu8Yg0Xedx0U6SIWsBza5xVtGSoSRv0oR
w1h8BaJGmIW0ka7VBb6inaPP64lPn3kskr+bMKrXR7KNKEZz1iPN0e3o1C9iAzJV
p/BYyu935+wojGSl+qCwOgE0zW9mYtPwDtQyiIGPhpYTphDw6uTZbd8Fo1Bi4Jh/
NFeoMm5A5xygXUBeP+f8LJIWoUHY66lRHq8X7GPnSzMr3HSDTQWR3Cub2KCjUi2G
iKz2zq27UM7D5sJS1gPk1qS4TrL9H3dJTSNLIk8NNlXgrNWW0qgX+0b0piIPrmQt
ZiQYMX9ARjvx+DOKajGKVkecpnDjjbxA/cPsZ4wOzMxEqj0FeVHCDsKybkhwRCQs
GqjsM4fgSA9DuZN8teyYJE94800TuJTGR8i0Be+B78mhY6Kxc9S/c2a50RWA0FRT
mC43CSbQ1XI6gBoJFc2eJj1owzgSu3xMV41n/ntGMyjL+ySP5Ue8pn1eILa05xd9
AhMfBvFWYEmtRh6GnEDZoqKweC2NUvJNXKZIvTYcFUXcrLFZW5vOeilHSRQ3XwLx
zFihcO5WNZsg+dipMhA8PzSVqGFMGWl89l2cYtvSGLN/+TmIwGunm6f0K0MFYBVF
iwuYznBIvFASME2p5HbVoHgjkn9uARWSgmL0rWnR9UdcE96iD0Z11wV+CGJgQ4hi
/44VOLaSNPXAwkAn+zPHxM2NWEA8m8/PUoqpT7AimDm9obszgDSt9M3gJBKvMBHy
c8+LL8XJ253YwsaIG6R8zMi7WDh+2rjD6n12b46ReaIGAe7SLNxBwODdk+IT7C/R
LM22A866KGSHlxRegN6TkzoVi2UEo3nhid1R2yfmoDNmKo2IahWVQPzWXT7WiKGV
SUqFKnMgGkZOoNBRH6az/jpxTD4EjpMestiuODiJaSDcWqNltn4nRFuUcpt+7VzN
d7OExvFtwvhCoQ9acCJhoZ6TB14pl8Szd3uGeN1Lqu/AsBqHGb72bfFhmiHXPSQm
vCRJTq2T+hdNKibgzJCZiuxs9Vv3XrZ0zDrWqf4tY8w0EGCBe9DzMkDWxHDv7+bi
nsZyqAkdXADsOGXl6GpQu8DOcsM4nlyVMLRPB9NxuuJl1eSCH+RhclViuIDuoVUE
gvqDD6PWYZrZpbyW6mFaN73YgIqUarydvkVOp9ZVo1q+JqhdoalrBzEfTUTujKGp
wi1+OAxzxbBNVWFQ254GetoFt/sU+fdev6OqaacqNNIQCHwSKJgB7PUBKA47FdJR
WJXflh2lii+6PJNOeAhG54k/JBUnCXQyX3Mq9aAactEgLOTaGCgl29EVorokFwGr
pIomhUAW/dXnBQpVGiWwy5K5BEDo0dxQEpdaZu+gcd1wt97LnvxJ8tUWd8n1jcXL
83YvuTapCQZUhHPUOVDkT1NfOIMYoqQxJnIXaAMBwO32oOK1EEQE7h2zYHrAmkYJ
5EYwFdOw07jGrVfgBYeZLuyt8XUINJz5zE+VOMaqDXsoB+/r/oZoJtrhPLfpLah4
szwutBB81gs35qqhLpePbBexS3fZNBVrVfTM2lcaJJbC4axCYjBT5O3NaPppkyGZ
kEHEhn/O0jpN90+KIkyRezq12jibpnnY+nZ+plEoOGPrcTfP5OuuWAsDR41JSjV1
j/RmeHKu7XOZ4VeDCuGFdF8/dJnJKNcl1Qe0I1+8H7PcgQxfn15vlh8QnzrX5sSR
cW8J/rXDh+hFzKDx9xVermiDk+Y5YVXP1h9nzDxpxzD7lx3SS0VihaSAOkjM68z0
7NvZSE4nMhSaPfoZa6MJCveml5c5bsvR7d7SBjj9bSlKMwczVpuvrp5H264iImsl
YABL1q6jyMwT855Gcv8WAjxnqhKNB9Zs8+YftaPrBzuDI7O20Gjbf8PiWOCJlf8q
LnM/ivNPzD2BT3MyaAbwsNU94ISdRnu69vspqKvAlc7SUYk0pntdhk+gIZdObCN1
aSm3wZ6lVaTdKUo3lTttjajtmtd9ZMLXR4d17rOSU7/xW2tZPMc1/U9sZ9ClYnVJ
CUrjzZCE4SVgscLv60BYYtFcRcYJmmCb7RDOdA27xplgF9RLKmPYpC2KcD+DSaSr
hIxIj37xlUq0rnA04yPhcn8EjvNXPp4lwzhXgeLoO6n2YoB0A/uC3lc6wXTe9XRr
ACAml1eH24B6I4v92cUIIucOJyfsENdqifaCLo72Rjly7OsRgyYrPEE+OgDswQZf
9JF2fSwcSLjoHi+hCs2tMp8dyUSw3ZRe8Wtjh5mtmThrJmi6/XxwQw+aGTHRvz/I
IrGrwfWCa9VjSVcsG/+OFsCIJDSh73QKyQnO523PrRqEOm11T/3e7BjsxXigCcNU
dWOKq7kjYaVQv/TMdd10KKBt6AfcxW7CKlcUhLON7cqdpeg65e5gujPCAbV/5WoE
Lsh3brqLCVeErd37Jtk9NJ8kq6rWBsRk5bwI/VWsyJjKv1EbLmeC6/heKEUavhFU
PhMsP6RYY7mCpDDYp155k5IOupEylFeaQVdLCqdX3i8FAthHIt5uqyUuKdDfhn1o
klb8Jk6ouzfbM61SSjCPo+Up9Exdk3b8/FiglRuq+ixVVxfs0hEcIr5O+pcXb25M
B7Qucb+hsNA/ZdUZkJO7PzcOlYdKuwpu0jXjEQwPq0AZY7J0iRJdkEMX48IeLHcN
cjDbpzmaJK62DU0YJlgZfoWWcoNLpqlW4h/1Iu8vNKJrSTFflQ/eQ0eKKvE9L7R/
yOTj/J5wSmwDl/W+rSablMeyu9YD31qeXSnOkUekGboacdZLC33fYjuPMHcj7Sl8
ZGVKSQKhgxF53TN3MMJPeNG+cdbQELQHShwE8c+qlj73rgRbMFFyyCfMWoAgmmlX
pG0u6O33qMaCzvaiXQe1PQxuYd3oTGwldPt7RVakNFZgW3izNg08K1p68gZoen9X
V6lOYZUAZkO3MtXa2Q9mCFdfPvXIrPJiw6+UQ4XXELXhoLs81tvc2cUv19RUgOlK
XZdGLBroLYzjh4A3MtgMCW4vSRyx5jA50rbhG2urZwJ/UiXCXenNoaE/jnEkCSkq
++IpQwhpsJ6OV+vDSBr4zd76DHs9bFQp/TLPAO3vaH2rHVqFGW6KVjGkmFMl0uIW
7vdBPJzDjjsb1tErXgTisH1xO+z0lCPyCI41NYd1+iVVoQPE7/V6A8lfqlyiCHXp
kLW0FGH9RBj2JXD1J4K/79QNRCeKXgbunGLYiBfoND8cq23pUp6kyWI78U6jSun6
0FVI4Xl6bGWz5FFVt/qpuykg9cq27fGEusT6XAlV91miS2B4KadQaYIznOU2o4hP
2oBsW0u2dg+i+/8Bk8ZXkwSvzg3aR8hABiXUsp1nuunvFCQMFhxTQbsVM4Vu8Kmn
uKBYyxWwUwqT9/7NlXi8OISsukVemP7tts84ylwvE/Le45fLsz7lsr6qIUtQVQYG
rpgbqK8uEEvY6mcLk50rk63BhpThMZDuxBrmzdbVfelIfarpOZ0Nm3jA5rW2YeNY
OahcmbcZHxmWCMEwkE57ISw1ScWwWy2sGjY4UKw4E2boeqhCPsVcP74mve+k6oMz
9rLKR5bIfdpE+GiKpeN8wkRRUFOXgxZ/5OPLiuroU+wlha5nA2H/QlLZlotl4tHr
+1YVby1UKAFUWf8Ir6wenVHSw7l0gI5D4kbOMMmJN9I0f6kdvSiFF8gLlSjwYxe5
LPdVtiWhfGnC44IdvNHc4wEnTehFbDjY+hL1zMAunqA74g+X6nV+S5fudV4T67SX
Zs/kK+pNSV7POtFYs93x0z/6msZMBNX49aqXLQfGTbI6XYFu3s54E1ocYIQ0MGAw
S7TRYgTeDmZfCaEO95fffAMW0yqLt8fzsDcXeF7O8YCHGryGhdYVBnbIhbqQymCn
b3bb9GQbo5Ynj5YnRU2Ielw7QhJsliEVRfz4jNKmViqnVm2qYFUB+UbS+tt+JUWZ
P+zRsD30fFWRjsfYbp+QBC8Jp1v3fDJXYenXfR9L6kW17m81qzZtp6qAwtBO8xq1
9yn1Gc111fCsFfCK4qMaZkOUtYv0TRWGpl73XCHxbwwntBozb8ZfxZWzMOfxfJOP
lr0ASG6YM+vYBGwAxtkMP7f0D5CTM3rNNEHE4okbR0B6x0C9z3wrJBZ3DkFuEMWr
05n18l8Y0M2pGkAnT38oQXMn5IuvgcOw1yBxsb1lcTkLgX0A61lpSfULLpeeNOl4
kPGhXOX/CWNCsO/sk6FQnCCtjqgIhx53MpMy/Kfyfaeij8zQAjKJYUHyzHRCtJRG
Jb/PR4/K/3ojmW0+V1deyIJPM8kBgGDy9gAAjPU0q6+h33tiyO01M1heVdPXnFFv
xCSsxPvwqFh0GSM9U+gk0TIf1MGV1Ou3OipMDcexL7xJfWCdRW86r7s0mTwF/54W
+SO6fgyndEbVsnvoyAz3HnE5B35muoDSHSX0n7B5FyXc5IU9pmxqiBjygFC3taDy
E+7m5b76Phe969EK3e83uQPseNwGDgUl1EkG4S00Und4iBLhOxSXokNs7iMKPmtT
8A3J+NW/iPH5LudKrLd6ZCG4Q56OgTq3qmvZMLeurv6WVGMWBVADiVnEfkCE2C5Y
/X01BSKwj7F9rt/sPXVIPryihZdkPJ2vaROzlXGNj0QqL0XhO0e2Rc7MdHMAVvJe
NBDwExO3AjEBfpx9tQ1k0C6R462NVBtth2Ogpoo+H9qGzYKR6Pe4ewVNT2oMUC5R
FvCsBHVQUso6pUxvExD6/MSZvcCHkXg1BTzRDVvyTfB2xJQAP3Lk5zu7EUSBmr2l
A5UWdSP1WbEAcSM2VYO77PzQBjuZpY4Okjtl/hc/hxZZOrL5Uf8kGOorOnQ1KgVX
t2oS3IKW8cBTopQ2mWhmuo9bEuB2GeO3lOXJOI8LZAQ75fTFvgabr9IJEgIfbloJ
yonQhtSzFcKF84nuuN/Lude+XoovUTI+Frbbk8db0jG9jFQ4/aBD0l6Msd1lnZiX
oBdObfijvgtrIIJVTJjkFqrz7APk1xNWUrE6mIiXxb4/hDdAKzMrbyUsC9n5A9Ez
sqT51BblU94qG5UyGd/tZaFGRnaI2B8+ZembA7l4vM+/pQzMUHhBUHw5zub9eDOa
gGPkQmKzcPa4XAFOsTMUYmPPbrZa06QfTsV/BTkzGBpxzFxBwUMe3EYuXIk3LB8q
edCEVYwXjUFwpXmpQPtGy8f0l5bXdiUwn7abo0Ze9co0Ff9xtTude3zGjdU8fJ6t
l92ITAWo4U+gUdnCtjNIvg6p0BBQvHgIYa31hCrct8r57Wu5I4U+cMOQX49SSl5y
qILIedGFhnS0JNPjd6GfTh+xgt2i+mOl4W4dA3XZBVeKdiLEowWN/OPa4NtLqvM1
UpqfKiGBKiWyh2FwdsYdVkELHWeMGRx6jbPi7kflzEx05k2+mBC9SHsxRX4eeq4N
/4LW9fTqfiYMb6q1/eklDRBAtJW0NZWWKI5PGe8tx2BHb4X3yxtpeDkdkB8sXNfn
S+oEdQ76qGnC4AzA5bDxyrXEzH65tPnhrX7p6oIRim3Dzu/OpEwYpExo9jolYhqo
C0sdL1u15PzvV7utSNnkx9XJBARNaybr+qSMXbm6m1Wx9+KoQOqfzV7bxqbA1Vk8
HMe8VPaVNmHey6gDhssq6rgHQS3VDeL6JeJK9uYe8oQxiZjaU52QLBhXx0QeHEKr
OVWt58IecaTlg+cKhdjzayhwA++KT2Z4ShHs/PXMcpC51fTKWctPGUuQ7O//4oyN
9WnaPSJQ615H1GX0gcwkWp5u+5rE+NnuewEPr5QFq8qDu7jcJXCAWFUu7zMB9+03
MIGNTxibb5zn1i4PrNlZ2+p/k/Xz8b1sE0JIQyTea3nV4Q2uMdWNR88nr2MhZkT4
zjbcb32EFE6CFgmhq/DILBubC7SKL2F8Q0GB16hYjE4j0QV3JmCrRJTf+fKjc+GE
IaDh4ZIuyqcz9pWOGs+kf16/cJglL1ManlcqohZK3V3qQ0IC0ghhSNoBM4Rd/8N5
xrsreuucFXvkNcq9qI5wRf3RuM8vOOkkLCSfsurFEuhT546+rJ7yaLpcO9QIL0k4
mhfEte6gT7hhL8yRZsTZyu4JQi5d6fc+pRT+9h8cOVRWEDNQxXqyfAXIU+9wiJof
3L+2/iK75U04SoO7Mb43THx8eslDbNjs04THeuUbJcHHmMKrLbQGCmdHq1oilKs/
y5TrVfCDXyO1ciXtvQRyZDQg3JjtduczQ7iyYpSkTyJAC9WBO6S74kjZnInkr4kj
NmYK39xa5CZbHSTe1LLMTEva1Up52DhCIdQplR1yRza/w+ZI5DhOWO0UTs8x/UPu
MD/hK+1HgU0HdhfVbz+08Zo7XyAkV1lV3O2wNqgEekRqlGEegWNrov2S+m5AMi3W
sKOgeZjYaEzJnHbtevtC7iKn8S61JgO050lARamzZR/Ner7Q32LOkQYBe/SDMTkL
5Mx8zG5MfIZe078BUsDdRjHNWYTgBm1Gh/FLPYdQitGw6SW8ymQGz2T5IEZvlmhv
aMvtqp2rDUo/GCxvUvqRb8zF2mmak3HvQehlzHK2TQdEU70yA5E/d8Dm5u0444sM
tkmsl6ifYy12+tEK4Gy5vYXB/sVDUqKQr8QZEv7755wxO3tEiDtXKuGfzUT7p26f
ISivIG+773RkwtCAfOErLPxzdAPSv4UtRB6qiWyTGvLo4300IhETnmM2Br3NsSBs
r/Gkha9E5KGXqsjCqwoJZjoQHf93n4/Opdpu+6ZstYrK3eD1xlXELTBBIZd1mp+5
QXxiR7ar8z4lXbw92sPLQ/FEISztcD12dbl9zuLBrZcy3qarKpEouYghWv14tCAL
RzuYXRAWRAJW3pcoAFstrCyVoe85sEEgh7Y77GKTg2b3Zl97B67gSFYpbXpwjDkh
Urb2/6h7qPfv95vngfBIq7bLtGmCIp+DHM9ON1ddeNgs8IFwQJrG3+5zQ9w+DmG1
pLBdFuoyVFJSeqnlN+LOOGQZFCA5YPESHKyr5tJ7E6PfrjuDzUHTm9aoyBMWWmF6
LWpkyQKLc5XjW2N15N2+NPaMIefqWHuD7U2pOsyJ46nwtZCVXSpn2mBhMkLHqUWH
2cQt4sZv/U9csoTlzD7+S5FoUyJ04+7+Pd/tjHppUsUwGIYBV4LqmujcXQYkJ78/
TEJ9nOJ4TgHPoCNCIanqsQzCgFEzkOzt9nuyTfXgr0s6fINgj/svYpLHAY1zIbkl
PszP1hyYopEyt/fplXDQ+gYouqXDTUrGVfQD4xQlQaynjA2xbN0NuaLNW9aHbcs8
EYnYAvR8cGc37r5Ivt4g1nJN+ln0js+fzOxkV0jgoUz4m9h4XAUvhqCtr93qcbba
258THPXPzx24ZP8VaFGYhWRqOY5vt5WoR3uQ3cYOYX748tgTTLR8XGf6Ob16J1hk
AHGQReP3ydMgqEBft7ajt2UCAwPzkrPvBZoxL1iVZT+h2IGhkrLQBg5vh2FBbhe1
gpHPALfhCTn34a+wrXfHGHg1qq30CkiVykeGnqkbvP2kfxHZeqBKdjquyOX3L/WU
U6BnhoGS3C0hEKFDE9uJFH2KuD81EGwwP72Z+vHRabwRsRRRYD7ztGwCheeACCZa
TluvODQn7db6qMdfSTDOVCbdmgfiQWRZIPDOXpU8MOvFBYIjFLEtUAeskfdJ7cw/
J7IiNRRrIO/VSwEiGE8MkjKX+B9rFPSxBHqxqD3g9JJIYtb85aSFJVVw2/HeYxko
T50TLZqj+2sUXTDMmF8IJtq1PVLMRJbt7EoSDicwb91T1cXTj5vDBvOqai3hcfAN
UCuEMPKCD3/2e0vG0UIJM8PRLEAL5zM18Qnxz3yBGEZgpjt34h7RyUdbRha7AW4N
yveQXcLm18G6HlyTstXJZIO9lowzUlcUZ4CZ09dA58czSc/2qzoXoIVbOZF81EyG
74VXQpHbcKlHy052mAwmv15YaEs5PMRAKM+816xo9tJi6QC/Pn8e6wD9dt0tDAyi
szydkGhzc5Z6AuC8s7CwmQwvtGRs1udmrYqjmLKeU23NM0Y8sBLwXzUc2D1QYJOL
kNrfSvw4xDYmcgEa0M5C3CSy1UhxjMtIyno1RiKNhRfAENbBFbXYJFGy4e9WqWtq
vGW93RHGCbTSidfP/OZt1fMAjMN92ZbvLdU+hWUvg4O69b6gzmTP/QCEO8mR77yY
WcGZSvawGJMcrfQdBuh+9OAQBEBRe3DJpwv+/ha2FBxZ2ZmlFn1C61VciolbNolw
+FhvWIUoxd2j0i+1vjSofLSsCSaHPxpTK+tQyFdlmv15EsJb5hwX8avKDCXaIC75
aFjyty3glMq5RV49oyYwNIsKogURai9NVg4EojJbnen97XCdxpLxgU39kx4TqzbE
Zq08l+zOHYZOE3tvGtKRfziywtJ6ZovXqmpCXRVnwXaQ0AuvKQjJuL40scpyvcl4
RsiKMYOpVmC6g0s7JXPbIY/81tBEU4AEiYv0cRZF5fGdfxcNQPcpdwgyQL0g1ORq
cYT+ys+8QH3M3GZLIHJrOKj4Bi+y9/ylFV1SosQ+LSlgCq9550D/LrBjCwbpJuAy
NQcFweC+KVXF16Afuv6bMKrIcYhXf2IlXNnzExuFclyLlvqoeQ/44q67ezxLqhu2
VKzBHjKTQ01ZMr79zxnoKjxXFRnKJcgkqqRkBx/ydITMMJuZ/TRtlSo24P3UvzD4
+PmBLmyDDhJkCwkYkhqmcBFF8z9HbedF4yH00cx/wUdIweMO7iTVHxPeMCmxWyfv
rsSAlxA3VGP4t64at6g0WCxAb5+w1C50x9XtdHa4YnsAFAyXWZc5djmRoGtpBPR9
pDnF6NMcdCldQjMcbp10pBdseOUKl4Y/j8p54XrR2H3LavaKcDnKYuFhPbytVk04
K/UamUearzqnU8ACBox3jKis9WkdsdWjnwc0Bx+lVqG8Us3M7zNf+th9QbDlHOky
zo7Z5PAnqBRsfbvccA0xis1GhC+zLoeDUnbcEq5rX084UgBLH3AI7GHaYFP1tKiy
5n0X1gZHmdOsN0FinpEJZltDJX7W6gpSnE+/Y7uVsfM22jggED0qmm/7bQOQGv7r
Z9wjwkCMKJ7A70ymn/U/GPECirwGPYqM3LzfSyqem4izSitckeH7icojTfMXbKjr
B3FZJ+V8nPwbBiw+hXMnmJ1GRsRq9ydrwbK+srGgLvfZK4rZ2wsIEPlZKJ5VgcrR
CPLLS9aLXhArzq/qKU42OVKOUv8QZtwm0bTyq83vSY0KThuH9KYYMmYgH3u9xAA+
TVteM6lCHXQjv6WnFc4kqW6e6MsAkTwL/Rq4Xlg3kNjkbmLMivwUmanDPMh6nJTz
37gOsbAHLCI9WaSdIGtCxJqJiMVbjnRWiSm2x+MHP/3zBxn//OnZUlabyU9U3Tpl
gAhLK5lIeYZYPkyIMoj+OVgaTTYynK3SpISkD6U6SAChhvfd/uIy1HKRPNjMOZvw
F+s+74iuAsYNs5vE6mDNyVbg/Zs6Ts1ZLf2zvBCRWHXwlUrqJ6kvRcZVnNOnnxc7
kS5JqTvta5+uBQWRyN0HJxGF5AhE1JDlsGtpSn/m+WfYLI3xVeWpZFOAIEgn4hEw
wGP6f4ooE/cliMc5Zg894S4XTFaLaR5hHtLYIxdv5NoKUYJ68fEymFWEEtIZBkWN
I0atYDDDJa5wT7lAv/clCYFR4uxF0XpJAJ5bh5FTeLLh4Kgst1ygEho665nayles
akhBviAVQrImCKawe0JYAzvqMBEUpXkx+Tq6ybma9ultUziJ5ZDljWeR/ISiWKO3
wdgg7d+iG9nS2oxEUYIo5sJ4yRQVTs8mOZDJKjfbYJL0u9M3CeUHuV0KgQBx5IUU
PlBGH0gn13MfedvwxrWOYIcXwaHgZ6bwr5KzJlWm+SHvRH6D3OXfyxE/7FweExDn
OnOSEaIf9iNYgTLeCLNekL7JNGMfOmDVGyXVHXFgZqh8N9SfjgPO+UkEHuQXDKLG
fQIxwmmh+4AKvlHhMIX3mzYWRMQixoAHdYpr943CvC343GrClBQKnShMYfsEcof2
l3wbd8piE+wq7B3GE6VxIxFh8ok3aibT1OgjhGx6OqyD2pltFa+QNEFrzYOwnfHS
IDeshA5IutL+nhOxGQMf+XJ7XDkz1W+jN0pVWoGma31ELuJu+qCWcyvFATUjmCan
ez4wf3v7AX208WOlrajxxZn7Kugy6utz/iQeHavP/H+ozCLkG3oqyqzIle2fZpeH
cIInx42h5eklYYwldjV3nwH+hKsTuhD22U9irHQp0npIeEBWQoxt7UFSp7iRUJ9g
wPHikYCDbzyJDBaBv4zui6vyBEu8hbBobQgqjxBSDTRxHyT2FWXR5UF1W78/8Pjg
r0+NgxdUtZlRWW17koP/xqkximr9Us6uR9iZlIkwXdJvrAKUpxh2phwGczoldeQA
Niw0z5BvdVizLaDVuZNipfaz5uAapXRVroYcJvhTZNwlt96u+e5Nt0KRAzkuGFkx
nsDeGBGojdD6iaxmxT8VSu9Sg94ZkP82zDMKqjsP4e2pPaJhY1tNFMZrlt/8zH0G
/G9keKJu13jlXPcwNIgP+1SAh5qmSbxBY+AIBaud2BkLU6yyqIe/3f2DLPm1f+5X
nUhfyBDkL0G+klMwY01dViA6YgcuVrTcPCTzpUdtwjrBEz8GnAQOarclQieyy74T
rH41mwmNU0mArg5sb/EXOyUXd98AiVAkOHdlMsiLZqo3VpxT3wj2apRlYI3/ORpd
GDhQ3LDL8yV2X0bdATsVuX1gcI9ZvURrddgFLCk+Dv+TjyAvNDO3N+sCUaVWL9gh
KPsSaiqRbJZ0KEYH2zmJj5B1GoiDaKlXjA5g/pPfM0BT2BX/mfZD5LhU7iTjPlnj
uqaN2S0ffOtX/byup9mcczxtoMUyD+2jTqD+n94gxTWYHWzahSLb+Kj1oDskY7U9
SKJoMx2ijt3zCLqAN3ENKlSHCnxcK9oBITeLwKCsoTsu8lvFWEx7YG1YSNF/lJ6U
ZsJwzgzQOjucJUuAncfZz1R795+/rLWvH6OcYGYn9u86U8weKfadLynG94ObsN+J
qlMlGXvvslIz9b/X7pV1y+8N6UKH2IMBdVHD+XV8b4y6ycOij3x6NHvkx5oZj1MZ
kHI7Zv/+uoa3Ro6uZxWXfar+dItLyIpzBzGFuf6HSMaHBii2gRHV/qA8YKsmpm0F
QZVjddKt7gOHcGNJ6HuuDYkxcqE7GdLH4v2w7uJN02WFrmT+yTn25mwVF5KpLLXm
pek4LAoyQGNcyomThPLDwMRlei24hTl59bvLSGzRyPVpRej7BNi37fJeS9ms31J6
diAOAJzpc1LlSqPCEo4gvjzY+UsVGEq/t7vcMswHlib2Q3hb0Efafoonsa9B0EXt
vqRSbinPnDuXKxWkE8r/OzXXruNGk0Nl5dRoAhy9+HY0O7uOZasHEYfniLl2AOwk
JckNrByiigtYbWs1Je880OYOZH/SVJ5K1LmpyNgvFIA5/aH9/MFUGH+hIovSKA70
0gt6FNbVdXfz8Pgqs4B9O41lH2UTY8u+ZM6A2sTRUDj7FLJh9oFsXRaCUDPFfW/u
eB1JryF06UCyWVHwf0SrW1pNn9PKUlYaihDhHjJBKs3Jg7kzJ2nOuzLdtl55IZw0
jGUBYG2YdK84OEEpOq6ilVsnyVTu5EnZ5geXxE5s1oYLNY1kGIfdxwUDZpb8KUP2
Ozq1ynoMMS5QoSTxe5pInC3hTA94u/HamGO/hI2GP2qzX+OeVRGnkjKpCzo8HJUo
ugDtru2cBlZIQfaY7J3Zi5z+jizhee5kah4p5YwiI9gvf90Ed8fdGArsbiKDXAN+
gmgrr9ebjMdLSf1X7Pk8nRa4c8bv5FwH7nESPGDpyD62+dFf17AMRSpwtbApOW4w
sRbFVCVKlBWQrE48jI1hkpHN4+CLrI/4wIZ0HM51w+SEPK8JQIHP8GdiS1cpfXM/
FPFD7fz23m79fvZovxTcknFhgaA4ehy4GCm7kJAEbcL7ujOAAZ2NOxrHv/T/LWuS
lEWyjKhwUDZbNXIqkp/5WwmsRMtwSk/u345hPUqAf0QBwwZXbAWaw5UXfRu+/7Kn
FG/2tg/pvpHfEvUUM0d0KCfgSFAngzqzjwxd57iPBvD0YlB8/a1O62vGJwvmFhxQ
aC7omQzItl26cTd7dbbcS+mcVQY/YSqpWfmJFYElBv+wJvpIi+4ha/mksFAzbfnu
3vpqOSbEGsn6qipgfI6YcRrMGjkuPPYRXMbc3eUTxspqOS58m9IrMvXRh1b/TAnE
YuasmzuF24f2fFNXzJ+xlv9wTcUl3ZzEaaDMfE70/GrUMr983lJDlDbvhzUOYcqQ
1aXPcLeLezSvmPiXFn97AS1TPhhWcEaJMNcvjBZgg2db16qDpqoyt8Xi4Bu6/80N
HqN/dGbl+oZ4KogveId0FzZByijCfuU9ZsB1BMa9UjDAlxdq6hI5b2bvk/hQzy3n
PbdPewShY6ISnmmxbY9kkI46z8BrnZbJAi5rc8owzY5mUutAVfY6x1Kj3OC+BMs1
bwjIK/YEAnQNWOG4Z01vMqXvFhKJv70aq11zGQZnLbitAOthDpPO1mXymZIkrxcc
fU8sT62yhcI63r1Tbh6vAWWMW/zo2GcixO2pi8t3Tg8=
`protect END_PROTECTED
