`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRY1RzQOTgDW9EX9R1DBuv+y0N4c5u+wdFi6Sxsh7Zr/7nPYiliNSCRffs7lFkMP
3JDcEdklU0gL5fW1Qr0r8MtB0vz0p+dI0GRbY1WCH48QyZrYQmJarv3rC4odre9Q
/sYzeB+0bcwtxIfr6g1p9XBIRMWR2hf5/aW7GBFQEWlFCmBiHCnPLdlgUpOG7DY7
xCbt6V+w2oz3pKrQ9DpmYlEbH/pZF2DBXflGzj/XB/uK6uKliXI3Qdgt5UaNN4b2
vnQBN9D/eV7ypZNd+TJChA==
`protect END_PROTECTED
