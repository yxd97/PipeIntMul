`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFaVSPJcOgPetGCXbqhM8AfKZ9P0YJPsxG8u5eL9+u/1ewvgYEGyedRWzsc0m3+j
2cDGKCk8lKwsQWf9abXg84dFKAn6xAGPYEH1lg4Xx7/3214/cYnMDbKcYIvgJN89
TRrMJcVenmNcC8qaeA2cbZ0jS7cxmOZbLlFnKWY3DeylkaEIFMnnOZi0Sevyoyce
GTznD52UhNfOdpff1EHKIzUv3sJe5B6iJjNGj8oGh7tRmUhl4icR0FlQchwbKi9l
LzMmKrb/lv6EfT+0fOkUGA==
`protect END_PROTECTED
