`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uteptFIrkwyruCxVXujnMD05TUIBUHwdMGale7VvtdctO+Vfne4OApwUaS08Eqy
VKj5Y4acjuS4lSvt5EaSpqd0qM+rad60NwIh/JVV899QmlEcYCovZpUi3QujAszH
TwjmBFrhnexI0KRy9wI6OCOQTCPxOUBNKV0/bB0oqn6k6Kal9gpAHxtqoAhFf92W
jBeIRUdapTEXowVd5SmEUfd3u9FpMu51baZt8T9ib7XRGFnFfm5808APf15c3c8x
WnRiasd2/Z+zIMy9nq/69A==
`protect END_PROTECTED
