`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GpzZgznsHjtwOn4AzxxrO8qBFabaRu03dgfXpjChRGl2uU6Bcf4ez9rO93ukQqo7
4eOKp0Rk9FN3nL8bIIUsOIFQh1qpqjE69kQnH9T+IcWb90bZIByFt3JCNZLXt+WW
XotUqDvex4adXHKfYc1xF/Tp6wdqMDGtOboRqsIVEYevdHonTFcGRvSyyRNnBEGx
yrwCM0xm9j0ptnzaxZi2dLB2bI3ZLW0cjz8qXDmb8BR1/GAI+ijHhgrYFx3YtR0i
o7djvdDumB7EFGBFwZ67AM3FJcgaDKOCTakY17CzLz9OVkLF7O70Yoc2XbtZv4kW
euPlGqg3m3gT8PezlRaq+EbbZ6NpMgVcHDYY1ReftAwsOnWyiKsYPQLGyMGQ5uBJ
wPxS5JMEgNPZE68DlWJC1pyOL5swNqG2pruzHUo0afqjyyk0veukMlkTmZaPzKVs
Af3b1IxOVJJFsVFLxwRvIsdx6/da30j2BKsY224WRkUQs7UTFIgC7et3zLKA7msK
fAcQy7cpWAfh+uAZtmSn2K2irxK/vynCEVYVLdZtnvXgssa4ETN53h4/r5NMtfhh
/cOgnOwwffKnbudPDxDhJLlJGVdExPK0H3dKAZez00NTyqcfqYGa3Ui/4v7QTKOD
dAOIXd9rb3U2Ngh/IYmNFB5iccjXIcw5ItP8Qt77ChIAADOjcqPd3LjGYHr2Wvop
4fBZkugv0RzRJkqeQk3kSgdC6V5bEWBkGC7d8I2CuK8vZLT90S9JW1LOUO4JG2uP
3PYvYpIeKykD5F95oZ5U2/RjewIk6ovNs7k/mOr/5HJL9TpMeljynHTfUp4pzHU1
IMrbqUzPpMae7AZQruJz0cFY/0J2spnP2hOphWBebNkcZ6/PdXZh/f12UT6m41P6
pe0yYYqdCO60I5AXCLZGPX7fVhiflHwSmq1Tz3HJ0O9zrO9jjsdMxKr4+jx6xkz5
cwtpkqvsKhoa06WmOEe7czrXXJ7TvEAwBUrU3c02I6YSKRgC2rS276C6OTHkWNcF
mGRnF5iG4hTzVvhWsYqzaSm+CvSAfhY7Zn0rLACyVlGwtD3iOAdyyxFDbDOVIQUf
GmKfP6OIq1FWdJZJw0uQrJTdt6RBZc7tYupDLYDo4GcXP4t6URWjQz99YRexwVVt
6R6XjjC6qWT0iCCMyD6ufN8hQRO0fmI6I6NQYBhUXUiPDzlOaN49mR7+tSuYflY+
KPvzvcZEjBXSL4GM0R1VflAnF+qMmH/bUnpC6cRwJIW/AxFD41TuM5by1Og1CtHW
F46jqh8Uh8/4XQaQozTfqFILVm8Kj9IuPuWFpIfDYbW4p1EnA5r5gg7r7OdjFyFX
kKD04J5MAg/I++9aEPK3QqcBhr1v/h8ofh1cJIrIyQS+5NAfShcWqssAnj8VqPzm
0mHJFQQdxzNXiSFKduH79TZbVT8HfcfDyO36zYNfbYV0+ixBOzh6pnJWMBrMeArC
Fm41HRxB7fPBGhQemyfOn9UbZ+cgPErC1LgdxaBwOc5HIgqqycSQ/BJqK3q1NRPY
ieOgClYcHoZf0KJ4t1RoHa6eRa9TTsOTuOTaY9XUL7f36aw7AX/cbaf5F9ixYzyI
/IF+oLULCS3to09hPVkE+bccUQr90DfhTpAL6mMOUH4n2KEtn6YQ4NoYotUjXgjE
Br71NKnVvas1BEg3ObEtVanMFzLA15Y8/pPgcKd5AeaxT+jraKpS7QitSn4CeazE
Ic9v8y18kN+QQIRkOAQGYaM7XUuKmRRCpwHhNVVayBSIe+7gZq4O7PBWaM6PpC7O
QepHgJx9rAN2/OLP9ahIXLMSMBFadEVuqqcAvXjzOte5pvdxJ1ubZR9U4VO7wst+
EjVPhhkk6SqlqIFPspb6g69xjp/H+/IUel2DWnxDY3w/64ulA/xLVaGz5bFPfcCZ
cHzs7onPKk78U5bMIfZOhRLmnmngPBsQKX2jm5CAjRqY00Jzoztlf+M/DBh2+V7r
HTIiEe7gZf/pdNMUdemjzvBqUhpvAL3NdT8ikLrtYP4yx8AsEdIjWGml7TSTCUz+
ZRVtt3EK6aFEEE2AaTrwI2ZkL25frnYgVzkCvIGtVMeQsvXrzUbDl98d9bIxXxYx
UAPzJIn4NS6SlmWd5vkD2B9wVY9/v3FUzCl4pQNTZjCBAPqJ4Cm0xrgQUoyGUKFe
trQs7x8F6utwehvgf+aOoNK1WApZ8mgQug4ENRIqu4FFsdvv7Ry06onzlw3Jjybv
cktEYUCNvRR9lJi56L6epfLDlYL5mROraak25pKD2zBFbLEZxKAhRh2xijdB0s4/
mWaDQwNn8eCeo212Cf1H77EMKzI3r4ZUSwRNoM2YmRqJyg7etST+D4tsQ49jmASl
0gX1to4ROHPJFEgWwdqDCevUmCctf0fhn/IIE7M3RALPMz+CsdAmPP5FPvbFoX2G
iABsJxk4zxOkQi3HvxBZU/vL/rtcMa66MXQ/dfqcKWeqT6n3TuvUA1vsEbpwYOhV
aBBsxVYM2q3fwZnijwNCLPk7SVYSQ8cosAB7UWJp8G0hfzxFXZXIajrjEOhSiKKU
FJXFEyGX0G3IcCQ1n2uHe4Dw9Pple/CeBU03NeMfh8neNN/Z4BFVnyduVyzmRmXQ
kFL/E3HRZ05FnrRdJASvwohJCYylwtq2d4D37pDViA3LgarcCt+VEWJr9/41VTuN
Fjbxade1i08hk65Z7JF9CVsSI4whO2naFTPxUoaD8Lty/bqw2REwLIeAek+XQPbI
pa58UJPvdOSvGuV7L+3VP26mu+ddm4sTG9I3QpMEdAfqv+cwfWGdTwVEizGMQnm7
feGVscSP97/7rFJIQ+/Y8MjWa083MLQzZXC99+6+bsInDFO6emNxA2Mdt4ujbmci
FY/b6/mMDb6lNRMnoCNZVeOHOFWwVKitW8tpufwjaOx54TdQdcX4Q3ihlsw1is3E
+4DR8cz3GxsIyeKXyEzhV2yhlVamMUKKgSKBPFJxjn3rrIyW7ZdAXBg0vCmHgMAI
Kf53ztMoyhEFA9leuqcgKAieBD4fmn+lKCQEsuHQR8ymIQSgv28v67kFoKs4pq/R
bcEcEEgxx0ArX3y9MetprT7wVstTkL+UKsYIlSjx9kKdAyEtP61EVGvCsMu1K92Z
mZzm5KYCwVQxoRMMMAwAp9C823OO1yJBtotSElL3zbEYu61S6Ycwvs4WYIqjWJTc
dgzagQoyrIF27/ygUPzFCdNV3HCv91k53lwzBDmsp5BYsLcVyuSK/FHb0QsZrcpE
jujwtzEJZCU3kwe+RnBqowLGt8krSQIr7z7SO2nJsnT1Gvndb+yjTnUnvY3e+u7r
2Y0ok98q6UreYmHhu2ju+1z66y9Z9Dn+XRmaBs2CYz6CkfC498GMlm+3M/nxpWls
Pw0ASqa5iFJLk4LqAX17G4mt3u7zpNWwSxbtt5VFSp3PxcQolyng7YLZlkW7fWO5
y1SsJTHzOiCGURaDS92qAg==
`protect END_PROTECTED
