`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDjJKOJictJhXsgVn1zqiV62dIsyPunI5QOVGwzxDNh25k0fwRwXg18P2x8Hdabp
PCEV64xqPzL4oX3jxOo1qxi1toRtLGJrHwk5/5eERDhxj3CsIRnww87u71cWldBB
jWitgOn8byKW/NwkUKYObJK8imVfhwX5Ly5dTcOUhCVB6LXbp9bt3lYWsAjGw6JV
3h72zcKByFYZF8Cpngj8iyXD37/iqWB46mYnEFxoFeUHH21A+hjbcT0a8GsCgsMv
M82E4pVH87SFf6e0NbmkMpL7Frc5O3hexCII9dtcx7QfbMj9K/sAIyX6P77FZd5K
VL1SaUJ9lWjhYSDexYadgFZzzQLGtnlacpTue4SbomPLzuU98IoompT7BSji78Ci
HRbyOiXHD51AdvHVofG6Cg==
`protect END_PROTECTED
