`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iERq+0fdUMP4WnpvsqKLiskE30DqdKdc4lHXvTxhrhbDkV+3Vv8jFXp9Ja9AFre4
eEfCvYBAXnxY975v1FYys0xwF7EiPd8LdSqJNPjM5aO1KrdiUqjAYGvFj+Yi36sC
bML5fyhpPnkULs/jS7ggQxfYv+prEq4H4BtOCmysuwYa6PfIauaAASjKwI8ZcsZS
Hc+jgZcVdlWHI/XD3D5qO4pjqeJSf+mighQBlbclb7Ma27KdT2kk4/+QmAi31Lp0
UoS9GjNcj4semVgkdIigDxxfObKLrvuLZy7Z/ZqVWSbpuYD8v1Y6oiAC8u9iPMY5
AethsDLKY270uytLdEZRZYwQ9MLx3VeEsaFog+5+d4hYY6r3Te2YADI74hVQz/NA
nxVktsB9BzfwCq/lxUj/6MestAzwqt2Dh21diUTWFgSqXnVN2soCpdNY6+Z6XJEd
mpUAKZh8atCGCjrXhFoiWfJd4Cst/X/opBCHDRwzfJAGw+d55BQl/5mcQERjMk/3
1+zJsVWCFDmge+qWIF/pFBaJMopi60jjU+k4ga/2EN+Kpnwo5aGVVTM/ok7YxyUV
JbvKx2ZfVk+fCnIGACBV1CDKLdHsbWG1FR/0ox2Js0CWAo5/ZtwpTFewdiZ4zC30
g0x5mFtoFiMj04SYMcP9oKANs2VigNE7zJDLGt4V7a8sYyEeQL2gkZoDZSljPrAq
XRxt+ImF8rSXX+vatd34Yl2rk6DRFQhbAkfO8Jo8RAHUxE7VxvSmKeeQojCyl//c
PSFCPDtHYhbhqS70PC9OdmeFZbYzjJtWBnAjkQMB9lueC1sFKnhW0/sacGPm3JpS
MSZ4WIP5Fnyjz2fCmxD2OsfJ2NdL8sxQw/ZSggpTdbY=
`protect END_PROTECTED
