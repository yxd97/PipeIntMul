`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/Q0USH1YqVvNRXMOtTi7/WPesDa5NN3QZg2kq5YapHjFLi88VSlx+AZEiQ7cwDy
olgLlNYDLZ28iS7yuv095+ioJbqSj93m0UNOnmtBPWWVGZLUZjEyclY1AkocwGgC
7EhYvmB6d3GRa6nEDgknmlC0ELe/ILgz9QQ/ZDB0A61MQiZXHpd0XUxG+VfWYKKp
zarVWm61LrRR9EV3B59RbOkPKZDW+CmgP3qYwjWG/Rzw7oTrzCdHHSDjN2M67u20
gUGD14540V/7EYENl3BwkppDPoEweB36RXBRy7hVn+wuRSw9zfEqLO7Rp5qtPRqm
8CSWZ89wkqo7bvW8aV1VvH1ISZLXz2M0J+/6czrZaV0/wpVcBE22SFChWp+XUVwy
gFxulHZOsWBC3jo9WoYD5XrJLO5Mi6Bl+jjJl5vdCd83iZDzFwpl+mtifaT0qKkN
CmBjLtn6jCC8XkA2wtf9IA==
`protect END_PROTECTED
