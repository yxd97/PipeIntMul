`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
peumGMyudDiXwWe6drmxdaR1GUD2vImF8jlnwzT0sPSfhkC7Sy5QEtpOsEOoCjN2
Lr+d5xrt2MKJ0dxjGGsAHAYbMdD23VYh8qQK3ybTB4zHggLowbNKPHDRwBGLjfFM
j9HqR2b5CgIY3ekX2c5ESbDXEzC52yTVJE1Nt1tgVjMJi+/583MhcA1V4Lu+bHb6
75TtQbOyRaP2H2Wm5E2AckpYTmUrkoD22+D1ceZ01ZNk6T1bgHYW61+1pcGq0SWZ
K9p/0lDMnvJpiPvEI1cLWXKlNKemvMj+EsR0KM+9IVWOCpKbHcRLCzSUF2LCsVdF
H4Io4jBUGDhgTVMAgvkANxgo2F0/0Z6dp3xY1ZGbfLpKikDGPljJmZ16xIlO3CGK
QVHnKqQ1Dmo39a6waGAg144CLadaSzrg6NZgLDT41lB7AWaLKTt8mA9hUYdGEdnV
4jG7vO9SczauHlT27XG52kQ9wFMVqkZAoooOS6ue3DECr0/6kP12Pp5MbXS9SvuH
B8Gb6pckIxGZHnwR6MbqaMSeLxLtu5Iufkghza5eNfydcR+d8p7nzvPZKZ7xetkV
v1GXY1Zx1g1SLoCQrUHhEAyqMhc3x1s7a08N2hXQhPBmaXaYIHbwzCC1UZoWz7kH
RYXlQHGH7Q5J5GA9JZ+/T6t/0mY1snDcWf/P+YI14O1D8VW3BMJ3SLQwO5huVvn+
4QdLzIb/qfb/U4oxYDKtzPPc/6kxE0eGfIqseYVRL/JfcuROkahYKaufVEAYrf/Q
5LnX/WoAJqByrm++Wy4aZ2JSzG0ELfbZFH8RwE58js+uA7aID7aVw35sJ8NkwLnH
ybJr1HyrZoLdGwDj+0/ij6gI3AEUVXU75H36s0VqreQbXuz83TjD6Vgr6Qzh1ih5
+u8TQc7UfUQLNEQ2Fa1KSi8Vmmiu/DN08Bn1Hh7N/lKS4K64rEEJisIG+IaJfutW
jyCPGlFTeeppg26X95lWXMlkDyKR1+0v38cno2BWd6sVpkE7hHPrIRDLPf5ZsV3K
HBgdQqbndEke6KrPSxnWIb8gkDh+Oc2aYURWCdm+MnIUIcY17QdzH1hzXhvK4VGF
Jyl+iXt/2wpfRK1bi5lkSOOfccFg5aWM9Lpjr3h1t24sxKgH/TM2GCzOe+S+3+SV
+iUQx2kfc9K10nmIQraDikO/Xjp1pJnTj/e2M+fOoCqczFfKEpBfVrWQg0c73mR5
XrUmsYMjG8kcUaXLMfkv3JKPJOX1dPhPMc4YZhmGmXwyq+/55whjw0NuFuSovQs4
N9d54jHFE1h6FidLYpeAd60Vgslo80NCsqCamk2UtuLjZSGeCejnzH1aQ7nQpZNN
acvA5dVih7FUSM9Z+HZwrL0jw6KArxVBIpJz4X15ClrQKPhiCPUBtCZU+LQKJS8N
+NqOVX4gXbFeC/FHJFfadweWbYpO+zdO9PSceQRDE7AlWm2/OVRR9dLSd1ACAggX
a6eGoucV1kWow1W/tYccYVXua6QrLY9jB04msCda/czB6A9+bICJTnxxYudlxerv
x3xrj+0yVidXxrCwUoXyOk9kipXElg67izKgavc1nQ0iO6RywOwJwsWnzLXYMCas
/8s6kQ3Otc7ZrDlr9Bgq6D1ZI6XWYvQNNPttV8qXNAl/n40CUWcKBXrqvz0DgW9A
DrRDaTFw7sJeZRxGkp9UWM7rjgbtNzLM/43SSQ82VDbyMcJU9XzNMESf3zay+0Y0
dyEolzmL7N5pEtgiSNdclT+ytzBmh8dE0YyIuNEfNnDqyqtDhGd7X8Zg/CGExk4s
0Yr+xvMSW1eULE248aLcR2XdqGuLmbA5XYr70xUqQeBAzoOcgpFrKB5AxrY3l+3I
NV5Yt150hxtNE3dnzumXKbkwMuyEt/otUCuCE3J0j7wtDC4JGbUpzk8CYsHEMQOk
yaqRisoalV/4IQxRX/HCUVfhJp4aaeV1UcNcNu8ZfJpbnyKYv2NcCMSMrvREgtYy
RAylrxBNG0YBTZ27smIIB87nmCJyvGyBsVNI8NvbRB0k1SBWH/XkDEtwbnZ0dqzO
8//T8kICfxgXg2osK4vy668HonbDtQPChMx4HD25+QwPk5ELxe1JLbQ7gRGlcMBx
HnUZdllZCULaq3sjLPNC6Jg/w3a0m8nsi3N+h93WxuZCmRsGtCe+eAdAQ2IeQT7q
KLrybE4eXIZnXCvq+3AYyfW0NKEzGjZztWfrLxpAkX/d45NBrOCkJNNA/pPI2ZoH
eHYU7xbFI/za6xpRvU/IQO5zsWzuUCUu8C0TZXgco3O532YFOydmfYYdnAySiayU
i6G1fGRyrMrtT+8g82IXfPJg+W2OZ7dWQ153bvWqNGic2GfVDHkHsFuY1i7LepZI
tPD76GMT/maICPo4GgeW5/MbJqz9bOFDafrul8U6aLJwxdJWMqtCHq8EF/yxNJmX
AekXcb55NdjvTQGmFXmn1nC+yFxXKhwA44CjeVXnePqbe8dHyzm7EC3E7+Ac2Bfa
wSSqBHu5GtiOWoGPMd0sVCxf9G5Z55esK0Dsr7mjX9nK7MJqJtVLKBKXaAFrYEAd
3msyRKHis6IRmH9c7RaxEwultoB1sG9LLyk7q9OLrjHdG7A6kLZ36qLkJoX3D5qh
/sfROsgHGHkZaUoc+1cZmKqLCMRiBFvANTKCtt30sqBEvpIEJJQuu3awJIma1Bey
hET4zwZKTOt0GkH+Z7x5bWXtVgos3ofp8Jn5cBUaN/wIaAq8onj5PkF/8/Ad3RuN
fHHlctRTIXagZ268Lry/+fZQFdflsjsOFHwwEF0c/BHEspoMiAtW05aU+krvk98G
jNKCj5lXTYcQ9JwLEMW6Wqeim8tRT+g+S00CNzBxXwLe/+Z8RgrKr/lJgh81/TEW
E+dZyPTBCNgIEnM4susCKLMAm/zke9ZBUvi3koO4KS8d4irl646mBaPV97MkPji6
pexdx6BHnJ5i4q01/2yxIOoMacXEuIANSRxiUtrs21SbPcTd7MAaGHxotkeDiCla
0vyCb/PKUYU7W0Q7ntAZXLHs4XcPMI7Uv2jvUHRn6oUzN+Z88FtDkCDIyJ4zM154
9BXrN+LAJq8HB7TUjT283Tl7J844wSvoIuj7w5VkYFcYCSqQGAbhMDqgMbeYwvkB
tjBpWPrcG2s1fgElDkMO9SwNrdGICewyXkp/t+QdQsSItblKicUm64YU/dB7kaCh
ExE3Q4OH23iuynHg/jbVWRauzmFBUI+KsFRu5EkLwutKrXajyZ1hpRDvOzAugslj
hj0eqjbMZTPcK2nuuP6GW/2YnHHcaWVxW6Y94F3SZUXYKxkoRH6FXLEFipY0ZfkX
jQRVd6GMmiPbm/lT/68/Je8bhCiWdpGotSXh3sl/TCEfngCyff5Ujx2KlYhmto/L
kt3P0d1cb9ZnsXjIxzitlpJa0s3pCcg3ulGxhAEMmjiLmWl/z8/JPDC+j4bEcj/N
FtqBQ4uxSQMnUtJJKZ30g4yvkjjnZEqE70yQWDSIhE7Evl0KyPL5PV4F3IYKfp/S
A+HCbtfEkUPqtdPTzF6b2wK/VcGUlPBwQpxINvLQzy50zS7fW/miXcOP5ekc6uvx
+/QTn1Kt2uM3iD5kna8AzXdPFeYXH9NJk8fA+KYew/mJ4PS13jFcA8axGEZ7B5/j
JIKPrFOpkUungh2laor5ocZT8gDVtRMg+6a5x7iHNSzy3Jp03RY1iS271EcXlKHy
t6ApDBKZi1ymDTintvApc1ghpk91m+a/FGmuwcMVihhHrTtnGyBNp1MsDK3LQk71
JinK/+Bi3Q1f8VlAWhfo/zfr4YpJZY/ngb4FdiEH+qwvGvSovDcRgl7OEKUbWMvM
345EiAUDm4ezikYLo0wkpy2DWFvjHuQMkj2IJCeylXD3k4UuA1OXKK3tpS9/qJ+M
JFp+NiP2e2M6a1pdOSfl/eqRchaDyRjqWFwK0/1QTW6/dAsK1XhNAA4FI1tpvyOc
hr3GH/5FMHjDKhGxw7zRwbA9kaYfGQ0SzycSCo73SIHGEGNur9vLVWllDwNGJYQX
U21GvQv+QMbRk/FTJZ5WA4JCiMWN84UfVSzLtAq8GSD+A/vRd1CBHBzB4HctH7FJ
A8YWkXOeWeZ6H2lF9siAKwZEkx8g/DYS/LyTG5a/SQnZE1Jaw9Xcnbdl72TtfLYM
brAaAe7AzpNgzBf41vFjINeYl0/XlGB5ZPcUhogIy3brZIhh5D2S4zd4wEu5InXL
e38Fp8GILofiDB9pPEaxLfHjE0u162ppW6cz2hVlYwkOys3mIlpa9QsFSR4mrzJw
kpMWz/O9AfPy/p6mdIbyJJZ+e5S3VycfPRi0I84vTM3G913ykrT2IezHLZ6y6+et
qtoYaqrJKN85Vs+Mmh6w/LLqewGTpCf+QCQFpRG0/q7jnkrx+52q6bHPdYkQ71TW
XtLsEqMDMBXUjq07Dh39/0D5iALu2BM9gWGF693vAg/CX7B9es22hQyjBRYA0ICn
OwW9wx3OWC3873bdu/XXtKNnF6+tZ3BdtBSvBWXcM9gHFQCXmWv4cPm+PBaSP6zC
7Dyi2L8b/Nflb/8T3zecEkntygy2l0QhUGzdcAXpzAUbLrUNAZ0Sb56hqEcRm/KS
xcfUgU7WxSl2S13xGrSH1YogshACqS4+f5+Cm4e478pxkv5S2BPaxy5A4yEkNgT5
VGhyEenJ6FxCsM4TjjtqorDm3qwf+2/xGstPW7ss7KKFVo/j85jigjFEFJ4N0Uqq
tsz8BNzqR1ELuYCuoMIToIdZ+w5bndhmltcA0SC4f4QaOGKFjh8XUTjxAEJuhX/J
jTSUOBC6dnqFvdlMJQnpisQMSPkm5mJR0stid1LD760im/M+6AaNGqYbOSpUXZdN
JlUX8SZTJabd+CSHkFQ2cG9e1/o3l/Hkma17C4hFABPLljk3I72ulvD6EBsfyqBQ
7swQZrZWxis2hI1ps90qguVk6K8v+Hguc+7U5FX62oodDLxHHozHF2maZZZO+s4N
yKWVWe2abp7aBr0nNZ+Z8U/k0Htfg+iuAgG1XW48T6Ztur5p5kZmSgf3Gdr34cF+
FZKJyeupXFBVaJoZyF0s1xCeBh7GD8hhfmF9ntXs/yFYrgaQYC/QKbztyWT86D0j
BwhlOvcmK8VJVQKNM+s1TMToOT73n1jrSWvKK61/Ll5PERstkwP+96RXabrsJKZD
JB6sky8QLwF1p78SBayy2+kL//nS/O7vVYiyM258/802fVzFZLH5UC0kKczCXmQq
/CJ6zqC/Q0bjecbjfh5YD+eJJcjBrxy5wu82k/hVxipt7QRrz0Eeuxur1YNCTv46
kT49hIqxilEQC69JpO0vUNLo/iq3PqzYmVGsivMgECMlwZey/O8jSj3Hrme22pi9
WSYL5nO3SoF/wpdqIFnXBGnps07NgMmxXAaLd00C43jUA41hWRwnq/j+goEjbHMG
y+zvDMEWk98e4JWyDfZ+dF9RLmSkSVnqCsDxEiyzjA5xhsvWhX0YhAh+bvofYyeA
g6FEdNSP8qNBtF3ad3F0lvtH9BOEBBpfDZRfujt939mH49Psm/qOCgpOBhT5ez1x
K4bCCUnl4VPtZSPK9Rwexb0MfIv8P3v874McLp+TsqPDGdSb3OZQw6QBdS0FSLj7
qzFgbYDgeldvjLAAmlACNivhhdNjKmHQPxCwq0LBs11AGJkYoEXvNs6XfA+Wxjd+
4C+b31HZ5XXRnQo/Ry2mpxap8JfFdnUwu08yn/OTswJX8tDx/Fuv7g9MGfocnzvT
845DT4rII1mHQQFHi/vUyCFXYUUvdqoPIQuVpj0aJGjQnhC2VVB0d9CWGuOmthX7
uz1BBuXdQ0krIh20OV114KU9NFu8f0/sQG/Q0puI+9DMgrEAhlk4TzhSmarw23Sc
C/YgMPY9eSItykhY7JkOnJ6sLD0OtFmXwbvm5Ur3li5D1jYxCLIs9UfaFVLdhPJv
83TlqauuH56/lt3hPWR71GH2cxuy31Mha/oycNFa7oqCOyWdBayqHLuYcZe3oTSH
M2btuui/S6BTuZ/4dAGJmPTaxHHz7lFi/UsZXQQ+3jG6zSJuDJrP5yMWWNTfIZPH
/2zcH85nHIfMHQ0Z9BxOeSXda4OE4GcBezX35Q+ytkUkfaVc+6539UStNsS2Wkv0
8gMR+1NsBELxshUau46zu81GAIDUcOa/BT1NEpu9anpKOndTi3f42zvHTXBoF/1H
xktS3NUfPGZ5l9LQ9sb8QLjAsrUSJ6IFirgYvEtRgRlc5IG0OrWeJvlFHWgzctZT
HfDmws66vVQekqg8rwVFh58hiNLTs5yOjKHaZvKXJ7VcSkvgaoP0kQVdQkObqnUs
Y45RuumXiwPfYmvEPh6h/8dGQHDsY5CsleRVMr57yHXhgzwNzrtGp7Q5ucoZO5Ol
2d0tv6p/PxV5dxDOe9547I9FuWTYbcsD1Be16aRMAwFWS9ffHA8/y9viF3mXh2Nn
VFZIVk7WWpyvkRlhoVBLGFjvNISrUuIHTg5p9EZlJ/RRs1fbmoHUJJJdyZLVu3OG
8YVASKuI3gF4giCO2qgqZj3x9ZAxhFLjfzOWnTH+YkqzgJYHlFCyAs5mqhMBLvPy
XpimnHheGI0C69JussfYdFaDtRtYKBdDqg2hjBHcr0zPuAIiMNMWzdjQ/QwMQGfg
BCYzXBUpjC5cLMZksi/NGE3l7Lj3DF1puntGw/WgBFZBbMNxJ3IID40qJrzXb9JW
P2zp0UKAxn3cNX9WWXBrvcLnxgH90OhTjt1HZAbh5SBCreRs/c6YIZVLLOUUV7uJ
91UebvmxcUZi8o0UFCUS3gS4QnI3PHjkpv7oE5HIAOhtWYSdJVYCyM8i1V4KGG4V
pDgqd528LM8/yDhoww2Ka7vGEWbMpWPcAUrepohWXQrqs9IXRaIq0sM3FeU1KNbQ
vS2T7VBiORbGM7zSQHwuWCWrRMIF853kCCUT9CXqfy+0msZTBOBkf5iQgwWb1EY1
tZtRdJ3aMwhnuH4gFTfFWATN7/luL+vO1gnIY1E1i7ASPl4mOiHHNbIw1N9ZfnEq
R2OLAUp6PPa1xJBjESgyPxyjcO6v8IRBbMfDeDC25YBELyatnZBmeffW8p5ctywd
pNMtQI2SFNnukveVpjLPqlGCPSPzVkk/ZaW2KstN5+cfF50r0tLNVkr1bTz+XlsR
ap+jLnP4b4D4XVZiFqXrfbX65gg/RmsfjBimZb7BS/papxiCB8iW+Q5TQnXEm3hV
CHnizGl8LWQAqhafGJBt/hqdWDU2ar8aZnuwjgpuhL7IrVj85tq+I+lxc/xz7PZa
ef+VLV5fUU+l10vE6IJ9HrfNebGl2UPcB+JK+RRh5kw6n4bqgmK2edh1F8dJkUXC
5EctzrmC5QrgHePNqYUocROSCA/78xHBjcEmCdE9HmCakr4ItQg0u4otJ2uwhT8i
vuGB9uYYa5j8JqeZ8BANCcJA/umDr1yvQsoEGY9pOKzGOYESxiqUE9o/rw9BC0Lk
mwxqXAlwTngOQray5zk052c7Xjoszel2iy1HSv7dlhG3ggraq9KhJVIPCuq4Uh2e
UJUVJRQm0VKQvrRNAF9ki9hlmjH6DTkmzZIwkey94hFKpEb6Ai7gJw3p9uJXKMgv
eKqFAMiMHYb6CKi3P1nvLG6/hBMICr0S7dkKx/unsCMecKuMdWeXANeazeTd9F5N
CZFIQVuLU3j7EsQSe55hTyojWSakeAWnkt9lbY+/dvXXHKVGp24DRgNbv9qJ307F
nRit/DLjz69DCAtoaykITaznLBMX/cyJiqme+jAiYW7TnimFqsUSGe1A/LiS1bUK
Wi5jv4Tp/4RVa81cQjCq90MIQTKQnunVDnH++6XTR6wT1qKqre/BYAOaNB4AjWUR
K89LbmOB0rQl45JqieTW7u2IFI+8xMdf60VHPv7XsBWBN2Ffs68wxbATrl0XPxrL
M7Ghtj07Med/pM8eA5S6tSTLa3Wg8il0IVahzm9mbyJTcFHIqi67fhq9C8nmHuG8
jZ8HPR1fKDMK2Tj2guhNUa+TQM+L/fpbVe2hKSV9kjbD78GxoAFhTwilZnl/Qa8N
c5JH9o8h3zABd63xguumHssAvl3j+KiHMfX60i20erF6Y/+36MzGdA9g6sGKdadI
ivd4ssa7jc/i9MUMFY+hPY37WX7k9p79Ecf+/QLlp89O8lmE8GF51Ptb2HrRDXvP
yoqzIGjU3C6HT452jd0Dub94qFJMcXNzYBoMPPq2rQ4bftzpkKn6S2fdkU4heoHq
hdMDRFvlpnAI435bFhwdlFJ57vFrJ3rxqKapQ5WEJx45S25OCg0ToyOVBVdrYud2
YPNjP5Dvv6R5QkOe8FGFfN2j2bFKNLgubdTIKYudEZ/CQKuPEIjP7TXcUlCVRpTx
KxfOEoUfdtsIWEJNwCwLoFvjExR6aBMn0QF4xCSTF5u5E7AJO9IpttQ6RKoDMA2E
AI1neWVMeUgChiB5nWpTndVXC63Calchw5CxT6nyx/WUroTK0hCDSeifxmGnC+Wv
d2zKGWjptKFX38UN4KIGuBby7yDmBBWiGC26LdGI4Ub19jUU9Kmsb6RMg2bBmPsE
0jEKwGXeLTAKzUe7Cj+OMbu7GT2MZYsN5oRRZ94YflnE7pZYTOLt7ET2Whixc+Jk
T1n6HMW8Kgod/GXCpgfAppeBs9xbVd+tVFe5bpc+neO9DkgPM3GAs3NX5uJ2P3gI
1JhxkESsAuY1fO1UpyA78fEhVhUNvgj5k8txvtmduYbQalJbgqQJtdzn1hnHbAuw
q5f1Y7fXzKw+IBSl6PSiMtCfFvy6Wdg4Wx9s1JFQyyYG99/nBr2dg3nUPQYgJZlf
acxbWxsa3ZTeD7UifYzHbEW8h4xsJyJHzA4KxXZXppQr8+BlVtYsD3wLQzf3mq8S
6Tr8m02RXFJry+zsA9gpdanrt3hyqsmOU3k8NN00ZWwRRPAgk9yyk2hduekJXt8i
3QylRmT+g5Qe1XzqRaa4Ky3iHsDDPknAReskM9hctLoJ6pSIPhwv31hBeX7vZaOD
CdRAW8bDHXR3HJjkEjgZXjqLG8e3sJqqmDs4hiKavD6lKbZNK7VADvb0cXgannDD
U2LGyumEaJNPdcAAmfs2Fm9DTteqNm8P8O2blH1nG/gxyN2hCxZPYEXqD98t3Uzb
FPTUqp3VEXPLBaMIgqS4dFTXx/2MpF7GG80Fh5B7TamT11S9p1YRYo4Cbu5DvBjK
bKF2kYIo128B2BvZRON2YM74qJNWUW0wOh4RQv3g9FCrjWQ7RnVxB8RxyP1VMXdN
aJQairlj9Zb7GU3V2RC65xllb/7rR7/aIBpZSokrCJ6Nc7lPGndq1qdCpPmSF2KL
Q/KXt9duCKoklM2zSSOhFbIJazy32a7RIwqw0lzfpxi4kknJxMF2oDms978YJ57D
DsksD9fBq5S8qmfFNTY/34xVk/3TE2lfsmiM9pdzOnjPyUv4wyjBzqtvdjw4N3il
z3FpTkJUdoMlmXLOZ+ZtHQQxxi5UEtYXbj2PRla4a6aBchVsy8qFa/dc32c8a6bl
vVEcV3nb65cdQpVU1FGbBIuDdW/oUbZr9k6gWZf0TO08J0k32SQ9GLxtR2+lAPSV
lUe3MeSGelgXcfKN6sWBjbhoXT95HoM9rEyJczJgWo+dg1E/BMg3COnk5QZMM922
8xTukO2lVQAXVRnGty+0i7uf0oW68idqrmiaBj7Umeu8Tbrdh+OqEl6W2odJSX6t
221E/Pa/e/VeaD29o3kpUnZ62bZooSY5CeJb4+ZPU3kXZzBZGl4HGNbvpmYGNkC/
Z9YrJe+8ac/FehxJlxPpEhcX6EPVwdv0hWSBF4xLXUf+L1CVqijatOdtTAyZkMwl
cCxpfpcFIOj30Yg5OKSmHaayOgiilXS7lRg6g+PNOKQF1Hbp42V7nBOzUs1cqgOG
GZK+c/tB/TwvHp2YTDs7kKwCp3c+6Zcj1HXy9mZfD/Rxu3pCjAtRPz6F40PH/kyg
zShTqRq4DiXmlDkvoluMFCZtWGLTZugodukjfEek7ZpsRnx/q7v4O0RBDK4nCaej
thnPYE5v4t95eoA4DBIiMRqtcDTJ+3lTSd4AG7hOKfyHMYlob1pbHgk2FTTaU3zt
S4p5M4E0e4D5jYaEd7A0XLZ0SWKyCIivuHO8YVYEYsHpWOLeKByXsyGQlHKWQu9z
rVG4TXHnVmbF3hM3jDuNYytBMpgyIPBmwG4fhsspbu+YPlSV4CpXK7r1XfUPYF7S
Muh1z6JNcUGgHGuIBmQGKL+aPKOoMsQych18THLi3OVdg6048JJ0Ax+pKgNLfBzE
wKcNWYsZhimjrB8hUri1aG2jJIFJ8d+Q6fe9h4I3ls5+ytieo+Shv9xMNOXzxrC3
qzKaucrOzNkh8F5f4pcStkdlMAgN4B8IQTfh+cmtzpw+z3EVgewswcjqFxpjZr4G
OAcgEKwDt4x3UqYW7r+YOD9vwG4pCRMDrmoQkSWHJe4MQ5WQMtJGvzgMlIkG0sEX
JetuwCHwl+4VvSX2C0XVOojUSmuXS06DAEMbBZeYVZ4TE9Fx0qp6Z2+TxlpyXzUm
9SQQMKRRf/CPONQHvstOgYp6gBFtoGwKjtgDcDemqjj1v8aOhHXPMx9OKcesu8Cg
c5LxUQTDJVDtGjIO45RFUyaxIghB7TiNr4AmJCDpYNPUi5f938obpZE4UE+UAuvE
y0vV8gijdAUqmOuIarNQ8gexI80aBguhy02Ih7A8Da/Ta4znozAbD9SHtWNM/ofY
2fKxdYzeodyMKEhc2NFWd9JEOw2i558cELT8HQspYjJJ4NXoVLUsrgTYU6meYmXA
m9pKj4Q9sZEv69Tt9K4A4GSpnhvWN6VSQePcNFOtOCRl9W55O0ePVqEDdSPTZ6Fc
jJOYE0bJHVVJCqc5cTOea/WAa2C+g9OQCISUJrzTey4r1oSvwCyj88NjfhWKTsju
VfIg2yiRpry9hTrHt/rKtNBI51JlJMZcJ1eveX9892Um523RDV7cmrQUBojsVNeM
skIfCkIoiboPCbfjD4FzvhDr6Qoroo84dhpzXV5mAOdtP9JYuXHFzqBNYx8FiM3y
n5a72L6Ni4i7nkva2KieHqK2sqbT3Dhbcx66rqTP4EyqASZxy53VHJHbLLuGAc68
h1seZfX+LDvihbn10QKGsAl3HY9fJ+djRBrCniFMonCUu1bhalCKu2P4GkC6jEA3
nNT6hW1e4uwGYTGTiNE0aaOuST1MPROuMGStwgWnZ+BOX+hi/plBbPzaghrZCdvi
8aMMOElk4YH/3ZRV+liO/K6wROIACufiR55gH8Kmx2yPL80hEJAMmAs3ySdJJ4LA
7QbIiSTEnxXfA7tSfIjuRO+Cey/vxGFi2Tlk48jSWroqts4yvDd94M87I/6rMUo9
cMELBCyFdDTgOuvKHzdszqTS06MgGHYb1mW8RWfSTImuzC3rD4w1ziENZ4aQ+Ppv
WcZxHWa5B5q/cgMQv9LZrSciYdJ4wEXBGE8Hp0d6iByOUeR/nsrUVD6MUcbBUALt
mWFYwcj4wTIn3TqZP71XSWTVoPQPva7rUlvEMW8EhuIaflVSsGGvP5BujsmmBwb1
SJMMTWYBHGM/xQgnZoqhAajTDCRBSNc1r5MnczKmjZTmf3pXFa5kGMAbvPbo+/eS
gDGhusQu2vvzGVylooIVNnktNa+VZ7YpHTC2FYwn850Z5P8YwXVJnb5VdLwH3jbP
LhXuvfp7EuM8fRzKyV3duWX0H76YOQa6sdLLkLizwtE=
`protect END_PROTECTED
