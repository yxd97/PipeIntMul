`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4X74HygCmXjPiyi+zKPSSKZUPEnCnJSw2wTr+nsXWtdg9rUdobNICy2liCO8eKB6
IN1sm5Hghvvk7u/iioZL4J8qFVIVpY0W9b0CoypOtKN+eJvGrFlFP2Nmollj1QE/
fHJgXfqoI4OvpQ6b1klpxMNAmFHIkO5EFuggiAvwyfnnaH/zEJvssV3gS0oHsn3e
v/Z8F2K9Wub9LxpMyPV+BOEs9NsnwGl9UujJM26gkNNJKimms87f7ocxsL0nsjKx
LJlPlyYB3dihCgJgTPYxFH4lOZfNuiEPuNIjQL1yHbj3T189ACaSJuHAf07CuvUq
rDsde3YGKg1YBMjPlW3PMXgAhSC/tMbnfJ9ilv9F3wWmo5DSjukFtzJihl4z34HU
`protect END_PROTECTED
