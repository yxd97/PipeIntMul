`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UbFg3WDa0n2zx/vkjioEWCUBjv0DYevoc6lGNEXLLn93cKbaapmrpFKi+TUbxlji
WK+SVDYQYyukXS+OHw4lEd7oRpmdW5L2KM6mBW8gWWWLGfcsQJ/b8hL7Zb1gC2KH
J3GO3sRBtUGg83QaT+L7yS+RXS6NlL6Z33Fw9jcylJpml0kA2pjGVT1CICAuEMp+
oOo+xyCLI5YHnddiN59o+w==
`protect END_PROTECTED
