`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LyBDBIq2l0FD1KNE8anU1X0+q+OoFmX/FnNI1C+vp0a8OFkIymXtzkp6up50vQ1m
ye6AnLu32n4C1/EEu1oXMYUDt6MERT9YkW8wyVBab2gJj84QTOUFB/er0t2XPwn2
9CL4fKS3AsldfyVnClvcZ6UJ3HhxReazK4EzOCIetuvnlfYFE39OGoyUUaj+o6gQ
diDg65zCZDqGOH+97ur5SNq0kv86ZJ2eNTiw7kAlSjp2D+S05zfrXTn5bfN4HPIw
VUIkR91/HQ4kALCuYr7llsedBiDFIyM5JYLJ7WzaM7TdRlotl+nmJJsuN8Cix3p5
PKa9II50NAVwuR5RQbc4ZpojWcGXDutMJxH1+phdgqevBUSbzCFzOZlNv7tSP08y
197ni+6sVhOT824SSjFUreAmjW2ruyXWhafU/1ygU+GIS5pFJ6T98bYn2HDMfCVN
FeODzAP2hCxujlQyRV8WCDno9EN5o0QGlcmu0esm4sdWTY1XCtXPPoWEul6hkG17
Q9ojSSAnDsGtYKspUmFdOQR7R+bPMIYokIMvC6Zt8B8OKVKdbhlsL3HS56Gvmsn/
8nodUQkBMBg8BcKtjFs2H6y3QSjHuH0yT3J75g6TOBMKFwVumLbabmOwcWYcaw1z
uPCUI2YpXR17487IaXtEQtyvvg0e4x9z2hEnAcyF0yedaruw6oEjq2tA5DGZzekq
Vl3FI8JpQ3tcnqkOcI678Acd83ZLLd9R/wFO7zwCgPwr96rt0KacmNBWBkLk8Uye
9YCVMfGUfjzS6VYf7LO/K9EmmGQH5032MdwHypt+MGr0FRniwVoF0ryHitK8TeSU
v4OE4iAFXqS1TVuASfLSs6wdY/RHt5xPjTfoqbqsub1OkTmNPO0IUThAOC3y+77O
Kx+8zKr9gK643ltbWB0RxA==
`protect END_PROTECTED
