`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJMJAqLUExomAPL2zQaDknIFmhzJxFIE3pzNpLOo5IJLb51J74NyppC9VXUPem0d
tzKeghCTiYZDY5nJiPiM+Tkgd2sXqL3h88Exe2jgnCluCeIy0WLynuzrjmUemD11
RMk7R61c1aFtAqrJvW2ZDz4edEAfz/poBPjUSJJLw84U/Bd8yN3YbIta99lgguMt
ke4iBS1WMY83uoLsdtA5RlRW1K6FsKejrvksl6n+dZ7eifobqPeLqphMaXP1SfIb
ZU+kDjxf5SPKvlMyMzbuO0BebNiGtL/54ZSkZz+P8mXTbGOMbabOy13BlGemH8XU
rnTVEHJvr2vo6xpBfkLAwLybuxdG/9n3rIqUDY4ybiZ08s5RkOLRFN9IgJFdb/sI
F5193Thy9dlQqvZnq3cLmQ==
`protect END_PROTECTED
