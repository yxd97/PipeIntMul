`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/Ml6ZkfejffbMYNQGOGFLdZOIj9+CKp7UjCR+A9DvxJy3NGC47UL5m2fU4MhWAC
Sed+/1/2vjA/ukVuGQusHC+cLLFqMTrIZkQlrrXQkfh1+G6LsCpVpoTjWsAPqCC+
qveBRdMY/Ai0LgcCbgfc9rANP2s5tM5yl8iQTTKBECVmYi2sNEj9TUaa9dT7ptpP
z4l16NUDcYyOc0jpqc1tIyFIRkTJ+VDtZWqauuEFP4HtljEu/IciOMTHnDXsJttp
dpldg8cJpwM45RyxM+kp6A/QKcDf6WnI3ILLanf45vpjdIGJRPGrjwz6C9OvBZCV
Mt2CmhaHjRjLcd1fu62SeQ==
`protect END_PROTECTED
