`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CYeczjEFXD8FmaVTR+pkRt32JiPvRlp2MMaSMCP/Udn4c+w4uqcuw0ZJ025h6pp
7XgbvmXk9asL9P+5EhrtO6XPGLU4czNxUqtz/uSfkQve3CsG8w+3nlvDV9Et3Lf3
u4Jzu9HLrpQR1aizEb5df9VrMuXd/l1c5gOe8K/0BR5HHTT0uNXHSmdZR0B5E2ph
olXmfz2rpfWDLcUm9IvfyhfnFxE+MvIY5+ImnZo68sLLlGreW9Q8i+uXUEDZc5lq
yGNSowXq73BqeY8rLx1h+a2wBMeJ3+gjaTBWeqikGHIf7Ts7l3OXVl6FqwLokgrY
l2YRPpyXHZX8zWlTjZrpwZCOUxaz/hwpXjIoS/VpEeqBqix01WKhS0n0d0iIRJJq
2mDVDYD50mcj9/2HzeB/ZJqPJ3t3i3cU0UMQ8AtlWs/NAdVmyxMnshdiG0LVrjqW
nsgDu9xjndlXjZkl81SEcCVKoOtu8YC1wA+UF++RKSt0yAXOxP8dO2f7EgYYWX66
8Ice5FDk59DOlbjuFPClnr4ARfb1ViSzMuqolyANo/9JxDle7V+fXlIl6tQOTcjz
RDUHQ0HDNKxaWuUyif3Xm1qEqeri0KbbTcQA148mDh9uZLf62p9LwUsxaKHzHDg7
B28Lnx7pRQf6pQqSZv4hiA==
`protect END_PROTECTED
