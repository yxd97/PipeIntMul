`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EApAOY6LFsgiywMuz5EqjKA5A3O2csVYnmS0xK8sYaoqxD2p+jl0Q4C10iIbsmt/
dMJBa71mPDdDNaF2PfSU9ZYOXsQAVkxDF0NdJHxpe+glyBnEBzMItO3dndDQQftq
ieEy/l9Z5UyYJzaG6F7jwJ2yyxcOwEOTM+Orl+p+Za3AWlIgYBi0+qmHU43Ttx7S
FrvSYYqRggGmQeyo2+Po8H5AM8JBnbMZeMVF8NhfkRAt7D0O4fyixcVgC0R9KsL1
svrB95sdLA7fDqXR/LlDsnQbsIFBmnYl3HYQd5EtvuFgHlP9qELk7EdRaMbd3I/r
w43hrJk6q0u8m4sa4kIv6awV6BszJTyjiyrXK7t8rXOqvCZ7H6KJH2l0znN3gRM+
loZQGvqpOdIXg02T/TYg6u3caPoGjRKs9fUU62HKwCxkj6M1MB5wif/oHWl1MOdu
X7AsDmBiH7kanW/RrSUHhw==
`protect END_PROTECTED
