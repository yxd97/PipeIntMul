`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhamX0RC4cNfjgbD/i6+mcfDzX4Zu9MqgSirMG6JN91bsIivlNO6yS2z+T4v8boy
CVllQDnR3L8Kx1mfPmu8JJ89HJj/QEm5LmQ5/3x8D+zEDCcQ9Dj5QTm9/4fS7bsr
7CfXtJ4Z3F8eF+zzCjaj0stbh8SCdT+lTjuIHAI2T9SAmgcK0Y+R0fRB0CUoOZzT
uuD6ndEpBJxqM8gyPW4oatMXgqchVxAyjSGk4ojb0H/UqcGE9wEXwSPnwKP3uspC
SHLVzuPXjHqsWDy3fEjihLjM9hGIU3Au0qOzsVeZnA2ewDwCh9p2WY4ZT/wINRJn
oUpWBZMgWivz8RMISq8lQlygZiT1MgBE5h94rfO1Eb33VepFlU0DCf37DhA14TWO
akOYWQgpycNyQ+VwGY/swHl43z+RwK3Iwrdf6R5YnQYvCOVI+SrdaVzI8jNTKw/m
LZ2m4OYO27+CEyK+2t0tygdDI98lS5BHtmot80cIyOCZ3OLTOByO6Y667PHUJLbb
gIvHV6qjD4P//uJK6TeFllGRTrdz40GGhufJzBAgNRxl0U8bYwacOP6kQ2g8cMXv
mDeCtVcCMhrnveccW9yfZdx2eS+AWg/VoFG2vFoVbcIfV2+ZkT4rNCjKWuXAAIit
j6m+e4YrA+0m3VPusMTdkYe7+klWcL6tEinlMW1FXFo9QvhIWfSqWbOwADuGfpKg
m7FD861x9Mu3fhpjxzMxLNulFB8HeCJ4690iA+QwU8zSFGWUNO5urNy4OnVbRmiR
lch2ii/tSFh0CprsOlqyRBEaeudYSiHfb9ZBMtsZpvFABYzLn+gw8zs/MUzISZ62
Az1scYYWQQ/iNivchR9ScYiyxxh4xqqziMAAuQddah3wFJSfgbTcDVx8Qo78g+m0
H9/zTAEcwE9pYknn7z/0nw==
`protect END_PROTECTED
