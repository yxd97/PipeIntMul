`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3cjgKaabO7LZ42Z4aqgex3Xn08RkFyp8Fs6D4v50/ChHU6JEVVrhOuJNt8bIDnnA
H9+/n6xcgXp/95TA/myS8yVLgrG2X95stwsef5vNWy1olkm56vQn/CLaFjoPjfVz
60xdeXBzWGMGh/Jevgj0GSuVZt+3fF8ukv20SYUfDee21vVHwsX2i0tlaLb+i7WD
Bf3OETmQkyfrKKyf/HRk6lsG8mRffyQjNa/HBzN5W82z76ECZZ+TOXfHOm58gkNh
gmubnWWx189eIvKpkWwqmMlhDxG0c7T19wiTQR8XS2bDpiOqdWL9OuHr+4CNbEyj
zKJ89n5Rq+Q+UoYZZqmaI7AdS34lH+WidrVkTPhNkI2G2kmxKKUHdTnizXxnS8x3
2gcLf09oyQCSj5PsPelHPFQP86wbvP70P4Ot6P1Y0/1JODQcCY1iMhN3CmKEfoo1
clx7Wh/4OSU61GqUoloNZEAuypNjJJoNfwdaJNUfdS1btueFw7MSrWNszS1wvwbg
GW2S3NbcH2vqj/jGSbBQtUHI43ukKq+9VQelA3isCbOPCbhn0gfpNHMbIaCHdsSc
pvflM8nhB90SK4p1yvedizVh+nNNblmgxIZwevNjs/uuhnq665tlav6wnsCO8ZNB
SlGmBhpdCeZ+Vhi698k2WsF/SpZioQQlu3cltvUVydpDTF8Ia/gXAWAIkqnzZFaM
QOGp0n6kTASba1Ua+HN0oNjaOAjplr/DpAa7m49YxtZOiiLdZQlAIC7TPDG/8hQ3
FzOwPW+omuqRKr51iizek2tC54SmCVPOBDROlFfu23wNqxlM8kwlWV7iNwQOg8mL
OcGMLQy5PBogSx6+ubulOByRVTFx7qmiSjPX4/iut/I=
`protect END_PROTECTED
