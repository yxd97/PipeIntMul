`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfM39I5VMWzuq6irLStSTTM3Mw7dpdklgeknaA2oaKW3Cf6uZhPKFYzm4lHTMMq4
7RhLJFGtLqoJ0glWoq7L1NTMQPTrToFyM29li2o0oCfwW/DkaPlWNrdxM7sECB2U
aetCdxFBUEDguda6OdpSWgsc7J7SsDWdo51WeaqsZ4qcbs1Aw/hruZUnwCfJeDA3
cbrxiaS/bonmUqISaOAc8tEP8aLmQFIa+PWSBM1PBi3+ks2E/7E4Cl7Yp4xYs7cC
oMbErkAFFLjBQIW0qqWIzg==
`protect END_PROTECTED
