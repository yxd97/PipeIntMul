`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ktU3qrvlBrdKwKwCXSJytHFfh/bzu+KWac3QudmlZhWloZrVk85LUxOjFS/3QvgQ
nEuXKSLsL/kTd9ouCDaHV+sukl5uEdMlfx7t+5bPatsXEmdUOrrXq156JaMSBZWX
8coH0THP1xq81Z8XPy5ZTwmvxSGH8wbFQmKqWIKJkSkxLixVRQ1xj1FO2pQWPpva
Sug62F5afOU0w0SqZGZOkkG2cLj3t8pdVwyEkjbC97ESJ+wD3P0Ao7xUM3oPiEXk
LrIZ/VApPjyWhBLI+XN7P0jKwQlHoI3mUxSMVJiDNvSJ5DzhQMKCLDGoAu/Z0DFq
Q/k8F8HURQWEbxgSzfHfXANNfCN7vI7ZwxvzkvX8Xu/A61ZeqYNXrwEFH1QCCa2N
8ExX4LZOz002agohD+8fllh4JwVqTpu64Lr30bS1lf+OexqAe78EXxPel4Hoq4dU
dvibHpMuo8sEhTQq+bJDAQbIWvaWuKLaWmWHUho9ddzUKLXvK1P36VjrBJU28j22
/TsKPtfKEELCxgDl7kf/9waKPAPXWw+iprUovxcaC3DFwdG/UDFJISrV7GL7//V+
uZi/h86B+wBdDTZ2+MzYFdC6z/LjM8aRarh/RKK3Ulehgv0F6bJfp4OZDtelnhLR
aZoLuMNWCnq8QiUasdjpIQ==
`protect END_PROTECTED
