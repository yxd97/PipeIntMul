`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uW5Kk+4HQINaFl850bn/eXJPuBOeY6yzuORCErhgfkMXbhQnvQZjB+tn8ewK9nK5
rMuAEJgmRTXlodt0GB+HGCLvp4Dz7jnqDn0QtYwkR5/yuptG7/9Aq2Pw9m8+6uWt
7egQCGhm1tdEZVCDkNscseyWkw3lvkz8HQCw2VD3B3JyDCm38IrL3Q7+n0yuMKKF
/epECQkcnQO4EGEuAb5szn+ebMZ3vzBNjqVe2WuHcgQaoAyGhn5ESKjaLnr7cuTq
/SXEJDSKq7sSNq016Po7ReS5WPXc+JhsiiFZAHmF0YBya4ONAp4+rly0UXPNFBzY
fv+JuPuCVYC7u3rDlM3l8puoOiWpRmCRimwyw0U9oNs5h/IABgZ3jEjIQhyMJ4O6
DwUViP9gwPyitS9plp6AC9Aql9seuNnIw1jlhbdyth566zieo4vt/dMJ6cAIvjNI
`protect END_PROTECTED
