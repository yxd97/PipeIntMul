`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFBNwJNIYFm3skZmtivYdW/IbCRQm4EMENY6tU+1WOAEr+aR79CbganoSoJCKjMA
g4+6RPrKyvmUXIqwq0gBFiSjEObF9usQ7UZIKNiEIKDvl38q6nWBhFV2DjQzuf7a
gZDSKchSFBVZRoZlE4xH7gQ8p7u+aURg+yKbsXrLwgUmquuoMTLfHF5M6yBG/2e4
fcxTxHZRJ5v++Bvv8vQ7bjR3QNAKAk3lB1BLTf77JUCe8Ztukoh2pLEgrgnPGSUv
hgNzgfLh2gA0jaCDAY/UHEJ8xjUIkNSYZWvph0FoRqSoCETtDxJNsdKLVSz5LGnI
2d5xv72wKggriq3iUi68/FqR8fp9PHxoDNBK7lssGGF5l/KejqakO5OblmA4Xhla
5sVUdHEaMHAsJE6nbhbhNdOK7tnL51UJ1DetVlzFXRs=
`protect END_PROTECTED
