`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTfcauylfcRWRCfO7ugCpe6o8brzVYO1zja0rQqDKZsRb6Z8asgzfwQc+m05b2is
XGRTkiEzmhFuaathKYpK1ljiyFLcYVYNp1iNh8jG7bCckHL50IgVxEHzOYLSG3l5
mNSUjGKHG7dpmB9YmQ13p+FIxpgBwZQTuipdoLGfjFFYB+65KN/csOvroDcchqOx
65ARCU7/bi4SI983kW42bXDj5WQmG4g/YxZR4cO940hcfPoXmMAWRFSXxK8PJJf2
dFAqZMhnckSDAwlAu0iRXY74ZgiI5MQ5Wti1gVMm5F8g+qYLJ2mOZH3r3YNJDxV6
Oze65cIgigQSZU5Ze/+S6x/YAdHrWz5Z+hWcSlcdcwQON28VU1IS0KQrtbp4Y6pO
7MLJ3GmZg19pdFXzU0E8uxJ2YBVtKDkvF7DZqGVkF1QB8dyZKucou+5521eYxTV4
9lE8/M+k3HgiXeQQGioKmICkq9ac8f+iGv7pAy+Vpf0Mt+ddpI9d3qeNTs09Ch/3
UoCXx+DbI5lROvvDJSkWMrEnhI3EjNzGyZLa9pGGcDheuTxcNvtu/vaBaiq4qJYA
MUKluoYiq0dpjHt8W4g3RnfdXM9E3NouZM9o2M8qGWN40p4JEtM62uEa0r1NLcrp
f+eTdfXSnO46zraE14B7WZV2Scv0MuQnYe/2n3gEFw1wPTiAQUtF+pKE4E5h5emd
MsSx0xV2Lva/3xKtCsraFaWlyAm6IT78tmhwtdOK980=
`protect END_PROTECTED
