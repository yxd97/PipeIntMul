`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4P1dLZudVnYOMVy6vc6WxxqdAvlyUwt8WCfaajafvOFuPNLfPXpAJxebFze1F9kp
8UmcB37t1kZe5tZTBy/NgK1i6BoXa8gKH2QJ2YM6JXyEBpyBWWH62DiMcNuEQKoO
huWVdg2Lz/LvrlNAoB/Wy3UmcxqCOzMVBWeLf0d9+0NoGJZUdn6napMHWYBPpR++
d+mWHj9nzI+LDi0Goi2Q+1wIl4r8FSZEIFXdHVc5WHexBYZDV/PntRQviIVU2XG2
+RomT4uImGcKf56lVyMWVKlRFtl1sXQzybCSVwB/6e+9V+O7KfSlFMC7QpU6z4A2
09UP2phrw2FKRnx/lIrNuw==
`protect END_PROTECTED
