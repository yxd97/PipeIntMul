`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c/gVTqB+FOQAnBh3mevrSQPoE9ZqHDyFKpcBWmnOBfQfgl8gOB0ln8ePE5d6HXIy
WaZmlyPBU9S9MWsqyNLesh5z7+V0fCSwLsF29gKnAiqsOv1v7bnHRvCQ2dwYci/e
NEe+I84nyYZ+k8L2CalpEIuVKjQfOsOa9meZS9QPPkV116AzOgOGyZdn8uObm9xA
O+i8iK+xMwn6RYtACLhtPObXEGaLPFLVQj1Bs48cVHDKv7oTcsZOO2WTn4KN68Jg
kiOQOSBJ+13YoLNpT+VjqyFX7DvbGB97OizBpLXXg1jF+31ZqUMCncGkzneaVMVS
EuJgXGp8k2muo+tfCLI8UEemM+Jcmv3FMkKDBhGevqBe3KCLrPOAxn+LqwC1tQJ4
SbuApRStIKHQmOz9qnXOkZjgDblQJO6IYdhorAxQaYaTEWVTxvyuYIrUOwKUEWyn
I+IMGTUskCIlxodB+Pv/BWB30W31X7hWCz2bdyhz68gjQPP1KAtzjr/qUsR0uih2
DYEBnXuBY+oVwcVvEM9+oOAYxhme+uFtFga4ud+Wqs/g9S442OIt7hYZs0mBLAka
wieemyVNWk3QrO4KMFTVPeAgqI6jvwqR9Lp2oWnDTKbeEg1n7mhXbhAwpEA9z3Gm
qCHYbMGTPtZKcynrfwzYXzm9jmScxfwUuTzx01+GTUalKjVKAF+oY2SmCNdm6LLH
S/3+iGPIUhYQYEOmaUTlvKdVjLl9jiBOnlLljkjJ6et5UMU3u1d91BjbzAwj/8eL
+6rS+Ig8wUssuW4dKUyXjaz2X483bcL8zJO82kaLfuIfZur1oa4eEQHS+SzsibqC
`protect END_PROTECTED
