`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvXmQ2FbEg0/TsG1BCX0axGyRPk88ovuQGl68Y4jCpPcQTprjVsm4JoQeTiQyaSy
K+AjsODGyf+5Spl6y95CjCfCNcshUND2VfE4ABJoNUo9z2NG63djBE9M2jc+2cwV
C9GWVzTFT5fGqg1eXx0ngVYzDw3DValYk3EiRxD4DVd8lTJxjgdGSD6D3rqEzhqK
reNglYLfTFW9yEJ7LG7xOoyUFPhDSP451UW4Y1AjHnU4A0ZkUmK8xUrr7eVbPlqb
Ucc/BxwgtA4SFWw4B10vQkpkYv5NQkAW6nHzRE9JloPr+J1t/fuxaPFt1LgxQB+a
F3r0ukJGXE3uWmKcUX67YAgpf2BV+UHBlV4eYw+NqctsLNf7vaZ5/RXeZtgOXKDK
1ZyDuBvy7x1lkVlhshucXpFD/BXfOKYT9YmAfKj9tw0GToG7IUoR9dvRRN17huNp
CQnOqxL8AfjTXpnD90O/l7FbsoNnBv28DUNvQt1tr+kJPJd8pjlg3tRnW7JWPooR
GZ7Jhagr3tpTdTjTqSIxWl+CVxUpckjuxrgTm8I4RKFyaKV3fasQrPnD+OfCcAIm
ij+1J703LnrLIHxp+UMVCItrVHTMqkIiunqfvMfjDtTFOMW/PfNbdJ5xfSC77f8d
y9Co+kgdR9JEeLH2Den7BeLI4CzTrpRjk5aUb/X3YEJd1uojw1WFdAR/n8cgPveX
oFb3uSFSmZzgOdfS8hqZcQ+XPeWfpGmZ8U1/JH2+dBXVz0VxQ4arXt9WjshOYsHH
6aDStGE5bsPJU0Pb0Ubc5GHox3DqW6HOIZimabBkdf5CcngqQUwo6fQmB0dl61Tx
`protect END_PROTECTED
