`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zcK4iTVD7tNfpj2zOHU7Y4lQBvKD9a+JiaihWulrzgJ7XG+wUOgGLb6Zz3WCDPvg
Mx54Yylr/XWdCJkJz8tBHmHnJbIlZlXpgkk8vKFbUewaD6GtZAI6lpfm8vg9jm2h
sAv4JpyTPOaRSMP4J0V+YbusZHO/o1BOSSwWcmsu7OsRT3SSF+8M31qFsO9dkKIn
PaxA/SAQHQIRD6C20k2EpI2uGkO6NJ7timcmg+sgys5IHa/dtk9FBBnZdh1WmuXC
OLqWEe+rgvaAQfPN0ACHdqONkcHs0qYylJHj5dyGvaIeJDPtMkfRgYFZzTgdl6fI
kVQ9mDOGxAKYzspyYYUkqyDt2uKUwpRLmF3fH3JTzxc=
`protect END_PROTECTED
