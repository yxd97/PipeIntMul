`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v72zvXBOGkRMUXQZ6+2a9v3E3clAZm5scMtf32OrK7dSoAp1e/30UUnmSSSCc7Fl
CtXfW6k8krOIDdLw5zXTW2fXQo83bknX2cQ+yQ/U8Xlz2tdL+1yS2nEdnvx8M27d
3jhyDgdfy2N8Fy6wnUARbU8vqCG458a+0xvec08egfj50yEP+uDq6oWctN1WAN+d
VPAGuKUSpxKoEsjkAnhwlJtU7hiTAIlObIEkZIS+12gYcCmwzO8sIat4hGk+AkBm
6B4fRhRxpANxczJrpWllX1u7F9XC9RZSAD17NBC8+jTowIVG7LcewA1mvGlTJqdN
MncXn1l3OLsR7IR2m1R7uxQzxDywQqkxClKm7WCnIORhom72fQQKQjIzyAcIYANQ
2YCEUiNUzZSoufqwlVlW6rhceIagWVx0RKwMQQZ4SfVUtJUm95PuhgpXA1M00BPG
L6zsNOKU9Re5WiFKS81hVy8jIMsarfdh/WadD+ltg4u6AqYWFfDxERKTqVuN3sh6
GTPdOZa9FzYNeh5INpmLbgb3UGG1Gl9C92LvI3KpnSfkUeJuN2AGhQQs0pCCQcUz
ESJGQrh6XcmGuWdFaEqY+nDrToLpunIYnEUepTNyn1q5FHjjP4QjWqA4V2nmZkKr
JCvJHDkf9ZvTex/IyV9KH8GL9g5PCfdlSMAO6Ud+lQ9ahcAuvilLXHJwroirZNSe
IfeMzsM/ZBkrjQfl4OsHuSVeRv3QqpaU7H8SisvPpWfYh7aEz3sUksl00+SS/HfT
rbSDIjqRh1dYHbJoI6+a5Hamrm9vsDbTNBqsiseb2HfWB1IR+jfb7qratnoeDZ4E
FORASEJ6K0YR33cJCoQtwCsv8fuOI5coqL+GRdgypDVbQXOBQC+tD2VK4j3fziI8
awKVq7CbhvdTEMhwcVQA7kPNVVNYlrVs6RDxQE6Ebj1bkHZj2Bf3Z5CG/PH2kK3Y
llXxfvzI2iWi1he9fcgacvXnGdgsP3HTBs1bpfqRwct5mNI3djw95J+77Emeecin
3eW24gQgMDztYQuD7eckhZF+ylsLeBBd6QM+eo7KqDHif3bTK2+vaHBfmj+ktoix
Aa/U9YX+dS42r/Q9rKwmmcvHmSmHm5s+TZ2LGrDSBCld9zyvmxgwBf0zDKl9Lsrz
9czkhGxyJFkAB1p3Va5gAv3RWZ+Cx/JUsjNu5QCyJYXY3VRNAJoh1KJ4FPQry14K
N4btfTDfjoFtxbDVwYR9cvNyh4GbbGSjnLe2xpTzODPqmz9U5QesleJku9neHs8p
d+O7o6sDkBsihgf+tA3N7D86v4NfQalglCQY0G065xpKBb72AJJa4E7zsSoJFwB2
sdb8RIAEgYmtdGSixaKcpFlwU1Px+/5qqI7Vp7kO6qEHCCaI9dt8/bNLi8bn0TYk
J2/A5HOzQq2PAOhA6riWD1H1jcOiUwTcaeTXqQ4d2F5zTwa/QgoZ+RzaXHGJ+D0O
WgVpIh07hV9XqWKWFTJQDXmy23bwH8fv8zHBgN5ywofFQ8rWxYQDWYngnRWDJn0u
`protect END_PROTECTED
