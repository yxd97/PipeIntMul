`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NmvMehuLkJoFvK5XZLJirEiao9RCNGv/ixjZTe2CcCX8by7+ZCTu/gea5ipefI4H
4y0phjJZs7V3M+lDpQHyGyTJ8+aYwRoJdGhkypQmlLprMdwWfu95JNXqC8Gi5pfP
2GL4kZnnTRT41mzYp7soubRDMDkaEsEplGwSyR85uCv7jSJdNyJqYikUkk2pfHmb
/0M++dP4lW8QuF4vfqbP5aGHXWQp3xqCX+PvZ5kgS5Eq9D26fmag6YbRYMNV3PqL
oMo8yFuMvqx05ChEQS6wnL0iAIriXGAVcIDVEUKYXk5TqHRHH6PjsR4a8sJMiLl8
upelfQgt/9qC2wggmDzYzA==
`protect END_PROTECTED
