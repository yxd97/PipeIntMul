`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nManvteGyZPARl3K89loTKgbFhCWoi/hx3jU80N9hD8R8mauYl/u49B916cMEuO2
3bLv30qnFVL6CikYz8b1e6URN3yfW47CbapZ+eLFgXRl+qWWb0h6gcjFTAA5D8rf
7ASrrlaj4YXDJLN44IP/es0rGGDdvar1mocFnMmuvENQG8keZTpux93f88idQafA
YNpHgxkSaDKO5VtEQVVWJmL9r4bYHC/XtXiA3li89XikYDRBmgiZIQwUH9ryNssb
9wyT4gQL81SdQjYsJ1QRe3P0WYr2qYgbUGxzbGgeDksi5PlhQoFvZd0NYuxpNAX0
B//DmNi+rRAW6GsV4KNajLWWvuJu4LTy5tF5myWrcYSwMGa3GxLGZA4owR8MVfqC
TaRkmkbYEJmvxKNKFouPCnFpATxVAlpxeKD8VeWAG5tsH/M/yFk8Cm6+RzLWyHgR
3Xmw4kND8reg5dqZhyZZ56lbXh8l3MV+8L+x4NTlhGJX+74oJBcde6LrQKqnagf+
PTYNavUcNtC9OEoQS9A3YZAESFDw36UQkjjLLNd/e7b/StEhMUODD55T0dcJjbbB
9qGpHg6PPuIDo7IgTN5LXYYkiIx4LSYXxP5evNknYnQxlbbsewXjX8OGk3KaAa1z
Cn+qcwwqwuj+w/gm2pbP4l2JaakOFMOUy/GcL0Z4TXTLJk84TQUkrJbk4UC2dG/D
6fkn+3dM5EcrBKWpKNuYzMDlvqIuZyZ74Io0X2c84lMpIo18lwWuNY/2rh+UDG1F
gBEYXrzKNee5NhKKrSyFNsALoZIvB8+hU2TZQAIDkgCsLvN070D6EX+hgfN2XiyJ
QzoZVQZM/wUPTQFxmOjlg06lspjG2+6D8MmjzJ/PjbKEtj8xoDhkE5fSqLfXmY05
TmisaUSe9n7CTL+E4TCsrmPkC1CWItLrhIn3ghutyiwgh3BS+zfCFEc8+gE63E7h
o8586EyAj1uO27JHhVS/xQhADPIS5Qg35fdPSNoEPAvJHz7pweOQA0Rz3YcDRGWt
/McUEYWGEkIUkvicuCKcaSehNeR7FRouPbF2zu+JmU/Ug1QdgBhZhJTJRBSTlAyi
x88qMY3MyPZ0yYiiDOaoLEB1R6y1nIbnCdZOyoHyb62530NH5V8lBmDh1AWqFMmt
M0XNs40sqWg7kL2bpnsleBb5wLdRCbZTgJhhipN106qE0MRqCC70RRUrJFwSuBOM
nyRLBdd5aZAsK5QEBgBnds7kyg7WEys6JrHtBBaUXNpfHw2N9mcWTakt8EcqbEfs
mbEVjubdVAMqqXLFW8PDc9rEGIrllcYDXxChQSb/brdSgtpj0Whblgg7wVT5PnRX
hbRBLO1Mng9ft1vZeRMd6Hgf6QEH9fT7NMYpxwid/3r+Oxt4I1M6fJKzK6PFy72R
fqNyV19DklLwVU2lyzof8oZVWLKEsR55gN6TnM9B81h8BBil5bXhN3qnm5Oy7yw0
UU0+eEzpndLMxIRY91oeh4xe63IbxXgM6FTHijSZoWy14Ap/xL04JI6/KesqeYQV
FXKeov0p7ZeDvQC6NLEDigx0y6oCH1m9DGejgvbmwt9EpkoeS+EsJzVAOgIwgu0X
Xde1jNNaJndOKCJhHC5i7nHRB4NpEmC+Sgw1de7awpl6LWRrjAkUvigHOsoKLMnp
srQLaKkzjq5vJH6MlUJY8F7JpsCXM9ORBO/fpCWruUR+F3Iu2C4bH9Tg5y8rSuIe
oySpy1nDNmBX3zev9m67HsIki8yq2L3LGe7p2s7VNaI7qmHxD4UNdTJub7nJWGHz
u7hM34ayjRnkaxZMQ/WuRxUPCbIX5MKVvPGkKB+A9Hoo1nnYF+zk6FoA315jAX8k
cag73sbB2cJhz09XZnZoI8NDEKzZsDx0Vhs+1sB8zVvCzpEmX9nshhUk0YNoAJli
jbXB7WCo3gctl3B0gxzsPj59/li4rbSCg/CLPcl9egKsc6TjjlCY0z3vdBYUtKwE
oKgSyrRTnIXg3brnMykHW5FDj0fgrwH3fOEaZy04YFeN6eE9QkoKag2h54t1/bib
nNWs5CuoHnv0tUtTTEX3XqsulCCRaqwCMy9QAaCADobqDENU9nwy0lCAaaOQablA
BVWjOcpw50pWAtnfbXWh681QG8lsa3FhITIApBAMpyYjNvl7iY68eycipNPFoMev
8kMZMiNUKfiVlXe1RJaxZ2rIDzpAhw7GmFHOJviWfdL729++XMj/9m5LQY5Wz045
t5JpuwngFChkMwDn+v2n0jo5cX6lZn4cVqCxWKwRAW4nfek93loiJHEOFR9T0VVJ
8jXGpW9iKJ/zJcFb37B3Frp2E6Di+5p7op51GYwWMNrJYwJQauFWop6JU+mow3+h
fixQISRPvSWpfeJZKFJMXWESOHBhEd4oPEvF4QmX7D7v+skZh8VgOYitJ0dcLmLM
LZ9wlMF5e/mhT+LXF3pPwTrmwG0MmxllSaSbPVipKbwiK5kBEDJ/pu44CCqUXU2u
kWyLo0XcF3TQXDWqU7Cryioo+r/N/ebU9lssEbi+qTtdC1KcteZnbiE0JQk8uHWW
u/mO+mnaP45rJftS8JZ/pRnD3n/6vYya79Vc+ZIOrWWy5W0F2KLbCq96CKKrEADa
MhfQBT+KsBZOgYDpLNoJ2gM9RUvHKNzRG97gx2PyYYCxc7pPUSWsxJRGHZaR4hXH
FQ6YURwUhPIeiHn8+u9iQI0/Opu1guOknlJBFIdZHYD1i+5UMzSlWFlz1IcI60Ul
jph5OY42etXvsxAtaT9+SG1hGTIYZkRmTe4N9gzQC3CxYIrNIc/y77D0/4hHGSIH
QXKLqSDkyaiQCG33a1029bi/tHzbI9MHf/btd2GCzu5uyBbb5eBs2BTXbg1JtSiX
rsI3vd5Y2zpwn3QFAEesoQmi6+HKVyZ1gte5PA114M0auCMy3rZDDsDii8TL8mPJ
ckr9GBus8FxWq6axpy36NlNVDp16EJE5GfwrE2g4kt852peZGPTt2QWHo0h7b1oO
OLrSbN4myVHh7ZuHv7QTm/94N/PsWxOiBnpbtAH0NpJHOwXK9Ni57/MXaL2pv3vP
Tyb8L3TGeMHoz16Zam0fbR+iJcseJdmCjUU3IidpE4Bi06ywydVQAVw8ExDlyKjA
ZkuHM/rwiOKeUaUMEW5b/H1nas0IGLRRrrgAkRwoGIFgzVTwskXV33fAiXKonFXl
DObl61LxKjDrKCjKyAnEM6ddmC7mXFdkHcD0x7E3eJLQouhw/s5ReweJEPr1SU3w
4cszAWnJmsxJ7bsQUa1S4mBogkSVHe9oqxcMh/6wNsYINXoKSSIJEy6uIWgFiP7n
jCq8PwbxwwlEWpyiZ1HjlREk3uLqkDvDrU2rrec6QSMOUmn4jhNFKzO9/pHhOxnp
0il0hDN/0bvqmWfeBdkfgKL5p3Ijz4gGxHRJPtCrm9UJ5SzrCz6a7FbKdjt7hQh/
mu1aXzo1g6zXHowN8ja7T50zlhypPx9r+5rk0o5so+f/QtAWWTNz6Mlv6DM/CVl2
MFDOd5ZAF3sVQRy1OnAWiP/FGEeSKsiD65qr4Xo6oZZW+29Te7nxa9gm7hJqALQU
dH3InLP99JxBW8iC9Z2ZTzsxecxCr1MMTPZaS1SdwlH62X7qU+qM8h+wwyEV2fXj
e40dnRb47V5vaJCS9HI3mZnym21PUbJoSwwWxcJr6jnd4dkts0YJ4vMp7PZVe7ii
8cOF9qA67zh8gcDemv6zAw6N/86KPz1w+8KVKjWAyhF8hQ7xjirgIMrpoOvX5CKd
VVYpLcCutwaP65hYGdFzGEplHvS2XcjUETawTE3Rrthy0dqV2WPGP+R9UwQMcQGt
ipUVzNpRTlgUQb50myOwkc/63G/qVPrhlYmNxh3qW2rr+if8k8Rdnlh6amUhszTK
nB8OF/m24CFJben7sqAW6pNsPEFQlpdOrbwt/+qm8nu9SnUciSzUKD8n+59fwZNc
S5mY4Pwff5IH32VJ5OzbabRP04KBLhe2wMGQGoQtuQZiv6FtZfWNNh/BIorCrqjz
BvgWLX6ALRGMCM/LtiJ+A86OzijppAqHY9+IV0zONFlqNxcNvGMyjhyJcaVW3XkK
W8N+MODmLlie6bxPMJh5jvOaZXgKsm9zbJcqD0DjmO0a1Nxskan6nTnZT8i9+mUD
uPY5kWvQmIr8b/7Ae7Ge40ZXHKivISbefdKweIor3sZ5hQANTHxIGDGRdbttUIoA
e7eapXxh9S2MzeigmWH0sZWa2qnlnq3vCKBEMq3Y1W5SRobrQkPsBpfSWdkPBk5/
gxHdK/s0nhwep7JvPPWsC7pfiQsXaCbyHF6Ez5dnZVQlvPuUgRgsToSR14pHKnoE
CKUBN3VFm9qvvQzYladWyN2nktMN0LSwWs+/Kh364czGL2uzSdHQVIWU8WjbTC+j
dMZmx14g5HCSQAHTbIsyaq95EDI7gcyOXsa27nAyFOwPwmHfQrEtPx/hJqrArje4
2Heh6h6UttVGt7M0rlFjIN4hmhHd+rifhTpBGnUe2e9W3ZQaqZaPIR2eBoy+64ON
Vi6qWuGFbZlvgP/Wll4tlPnrBFIU9jILI9YQFcGFh9JMeLmdMDEPN5o677DQzJxg
pjLbuWOBQ8swcAwqcOlJkjrHGnmZVEvb2fxMZuKO8rMVCt6GKJcsmlZy0Fu3k7c7
m/cqE4vRdv36Qt3tWqDgaKO+HcoaCYPDkh1WPGkMB0SCFQretOZq2mSv8GVMXROW
L/6Bf2gpZTOfLo2tMf9UVmaZuw0l/p+MZkSkTaeHkUWCGNtAixGsIN56AJbhV2gz
hCoMu8ExBcqpJI8LPxn/F0WqWLIQS674VjwsDfbQgX54kWT2busSrNd8rPgQQgDd
nzZmrcXdyiNj3vlzFWEidOLsY5Gcb6XCOXqhIVLeBKUMEp9uqiWNUJUeS7s4uDpq
/QfhGveKLyPZT/4v5HiO9/bNHLZ+lg4Hx6Pm3Ez+JtqSt5338hjz/18L5TgQfcNk
/U983sO/XGnBhOGD6pjAhKWvCtsw9i3gflrsY5EQJSDpCBUpF3dHzMnmyvflQLrz
OsQk1fdJhcTNl1CNDa5sU6zjX84dqlPimFmpHHXhISJqwUbIERoY9ms1LzgN/cEL
pv8hXXnj+6EzZ9l2PKAyrN7hkRoFqYxvjV1wwcEgE4vGsjrZ4CRdfqqyvferflb6
+0OXWIi09zePKeGul3EXemhF71sL/DHJiEBVzhEfW2tfxAFedFic8ilV03M+UW3A
fBiLRTgagx+VtWUAQPCnZRDgm8HVkB/4QoxWY9XiUPNP7SU3yW8wQAvJYYxOfvbB
HLNVgNjYS3vjV+gSxYEzb4L7c19/lJJ61vAXLw2/hUCKhaDu7q5nKHu9VMSscZcX
ygwi5Em1+pVV/o10FteADitVXbjOcLSuJWTYNVEGcvojds6/+M8WZQuqNMT4364E
jFiZpVqxDbcKwJkKJgStlLyrLl+8JLz26J8G9Y4jR0Eju007oT/x3MpEjy87Rv7V
wWvigrTSb79nRKty2BOCMAqlxIp3ndj6odPHabHh7h/R/lIjec+xMg3wTMU4oqA5
+Z6qCDvhSTnvHdakl0085ko1xMAsctGJ7iY/425vD8KFQeKaVLcFrmZeEcyvvyMJ
N5q0LE+G2pBrCvfioQmBJpSZuNaEjMNZkfUf/XDLeVkCp+0pZ8KQ0ip38KpLU/EV
1GRkX5fUgBeWunW8Nv6PGlGQ14hJ2Vz/GIJSmCzahxnu/V9yZTOl58mKXcwkPD9T
WVjiuuE/tnm/RVecAAzQGNxuM18ZbX6QBfr1VXojtFqMJ/d9yTLkSgCPyvuL+kUq
vovuUQu75TQPjykQ44jy+yfe1ShHrn+0LWT8efzFRdpvzc8lOszxiWtWcLqthag4
v6G5A3wbB2kFTYHduCSRowfSydEdkMmRighqObnQes4S8pISA45jEMbub0ug0lPT
KWvER/e31jgF+oJiZ29T3zIFrW9CV5yaVVR9KkJagTguwC0MtvfWxZZ1ulEf/GgH
rEGCJNULJ1hJNJG3QKKEGtQ4GAjC5umOj9u5mtPoxdUBKrUX4QY6lbghsLeagAmh
He02gA/bJNrSMiCPUo7Ru5PyGbOZRDOiwipiF/QY3utjmhSz505ChC3xHPQjRrjw
kSP+vgn8Acz9bNW6L8HcMD31p00LDXop2TaG+S0ICaKAqALfG+yfvu1uXnPEq5AG
EzyEMWdPjp/I/WL7sjV7YfRSIYwUigeTTt/Q11bR0tndPkNEpQF0beIrGB3Aiq0m
eKBWBXb53pEhqyI7i+qQd299fniuagMcNX6i/gJUH55epayaWy5exvSaBJ4obAGd
m+NtqrKTPYHjhLX79M61xfDvxTvZaF4tJtgRxQUB7UoApp7oQF4f8I2CyCFrQpBx
DVY0plM3r8o+VV/EYh+DaSgLAzITrbZu9wSf0JAUIlbnhbgtdsCJrrFsfH0pkPck
zqnag+HSwjaI0tybYcpwZNqIWmZX2Vc27uGNjauxZ9xfrTTJ2LTRl/VeiR51VC0I
FyV2Ey0HtQhxIdZaac4Ho/sEEj3dJk/6v2ToTooFuGvWeU+R5hw+tfONDXorPqeV
NoPhopKuvFSeIKd4JjV40zDdzlyMexielQxHgWcMMm09iCzeoCV/thjmE8i7jAWf
N23d4qo3BjI1dqCmncr/z0r294K1WMuWK3nNvkVu9qg+qWSQR4mw12QaSp+aN5K7
ZV2BB8SfKveLGjbg5Go88ffVozkKW9WaisgEXPs8kpVXtkeiZ1NebL+0CyeojzFu
nFZm6XJRTaDMLJEXDmkflkRxmLVxYaGmLasqGBGjMMLYv0z9WM6RKGUqSwFCa5xA
u8sYpC+o/E30h2+xctLZB5LLB5qTPt7rEu8Zu6iBHEsOLaznOvUH1zbhv0NX0lBM
PJKP8B85shhWUZg+5FQ6Eg9a+7T0KRPFa6MMt37bjZAnvUzMjEGYKaLEW6ypBOE3
P1NSQzK1gJdRy4rwePGCsubk9DD7xy5hqRVICKgeWn+x+49RWwekfNP7wLr7oktO
lX0KYye7DKMhmpWb2Hy4wUIjvTJQ92PFRVkZWbxQDmWp/x1tlSu9Iige9Xkmmebw
N7rHLTSoEOGfuptT7Q877gcwg2ew2l7O8i9Py/gZKHd2KDWdXFdfTuDR72Zt/u+5
cE6JEaVC6wxMCZCP2dS9k6Uj6NqnPTqVUg8KiQTZ3/8cwPuDwvsYNXiUB4oXi14Q
rInrIGI2sD1WSURq1bKcA1UK7/kT3hIeOoLvkbqu5aUzgaoPMO5iI/nscP8ET3E2
VUtuXvFB/nSW2ymWYqN3dvlCgbB88cjMdlIw9fmizmtTJ4jA20WjXCSyqiN8rrwf
MoHbqb9uAbn1lEDwGXtGhm7hh80JIr6vvanVdOm749J5RRVW50OuB5scXq8SqkWY
Iqi1R1J5YakrST80cDKbv2LGgN5/ouSPQ7w5aCWRKtyB+qVNhMIfPO2NtoA5Y21/
zEGlgIuk+zX4v11nhE1zWXymVqRSSnoGX2RLcijMcOvAFTyv3MUEWVyONyvgC8/A
qt1DE8VuETz/IUzWUcJGNuPOIKrXEa1J3SRcNFQAO2R2sF+hjk22aN8RAymIgOSJ
T+b3g1z0bIikHj4A7llhkv73RwpH3JSr4bTdmE5EvvmxSVGFst2qQZ40CvxE5Gx/
YbDC1w62UGws8PuIy6rJAONz0o+zqgE7mEZcvxkOkoFMnh76WX/MLHQ2I54xZKbt
c/48UzbUb8e7XsEme3UWQWIQZuSnWH9HTeTJCCyCJYMGT0ft0F/WnnZZzWJHsPZV
PSf/YUqfmCgooA3Y9C/V1g4VdfVgUyZKHHeN++KxrmhM1eqKhCcAd1cX/D0Shj03
uYCJTVskbPN1NbD6DE69vG9CBymEBWWe+mmW2q56hTMMfbdjQaSmYZhn6s3b6EX1
fCYdzi9lWue3b2dJfv1PWA0gKUIHQrh5ZZhJeRvwgWodCL/P21ykyLFzZRMXKn2B
UppycMLEai0rys7W8Vf1DcSm9bkt4kz0xLm/UPyA4RaFLtsflqtzDjUjihBo32/f
6ySU/3FfDrisdBl90Djaqg3N1i7WhOI5/PaAzNSEIHGMT7Hn1VNSDeDXjdDQL4MB
sBgwxR3y3mNvKMH/gTyTN2hmtOFtVVsW9EMRj1ESh2gRIB+XrjFCxDcReX/SJ3/4
JW7y4AMuRS3yAZAPOgOVV+Dyvc2+iouSBNeUgs4IV862Odk6ZradSzb348IE0pu6
EYHoKnB9Y3Adp/0b38qrOkofdRJc1X1RqdGEDQZaZ5HM76yYw/0nHUWn5rfGH0q/
PvtACuuwAwGpEJpTgF1DQIFT3Iy9h7sN3K7+mFS8BY9PApxneTiqLlL5VN4b/CfF
wmCHywanl2hsdVMqCo1EFrlwJJ4kdVccbk66/0CmSZHpCr6cWUpmHazlwZow4BTn
IDnrugtTQGCV8ZeKt6I3BfuEIRdUEEYmyvHTcW88sXoKB8DM4CmgNLjYYpxAlf2V
9Y7yv1yyhp3spRLgv2AM6aeuTREtTyDI3iLPh8YTh4JRq9PB9LIrUNCp42IrlFUG
YcTSt/PtFmcAfAA11rJ56EVuqamh+NLD9X+wBNzlsbSd7rxXlZpenTKzQjiSHoj7
tGvQ0ZNZ81mdvXpVajvdeQI/hrbp1Vj+FtZqD1d+3WiRmblsq4q6s0HKPzROGlJD
p6cFeqWko3Ra3U72udwUmwXbTI8vz8s3YJKxB0KVJlEi+ITeOBcFpb4F9HjVNBJh
69/vpfOGz1JGBVVk0IHQLg==
`protect END_PROTECTED
