`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
auuItsUH/Wb/pYlNusne90ggkqYM3fJxDWIvajudTKUiX86+hDB4SFO8ytNWu90J
0FjSEYGgsx5IYhyEfEjpIxbONQeqQsdtGGT7pAEF1ObWsHDcFLCMDS6K6WkT1ASo
l8ialGd9d2bFnwhSLbMkX67BOT/lJgEIgRKW4NjWPDbICLOS6gIFfbP0jWf7Wfhy
M0CNaSiwLnT5hHGibV3dW4ftjhRvAVNQG9jXzmtwFuQblcl8blixSxrcHF2LqXfl
OES3oEC7UaJ0jRpc1xRzD/YDeKpmzrl2VATTT0UxFHniNoZflnkFdbcsNmqa+Y6V
XJy/EPUIqaoKdc+fAYxxkgHLPFPkwKw8avfnlZIx+YveSRZtGxBUhYgbh9bF7GCe
`protect END_PROTECTED
