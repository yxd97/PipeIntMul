`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tV7RmvLHHTuKJHjEwerMmC1abiuPYN8Z0a+CG0GqsFY3K5Lh6q5OKrKcRJU26YJg
4Viz5diM8dEXYp56FM2XghtaY29LgMtzGDAoGALEp+Q80p2ZRWk2ZQ261tUS/O1a
3EK4nVZLM07ED/s+8+XUwbjjzJadVf1PxBeYyVMC+vQVmGVMHA9632EPBWG/HjUS
qVv03fsQY6thLGyRigmjAdOBzOZNezqIyHUUsgAx9HVuQB8Vi1W7+OoL0quEq3qZ
xBV8FzYYfhNVthrOL2Zuf3ISbbsC6yFWMeCxE5T2PZMrXz1cPypQsHedYzfQaHY0
UtZ9LlIsGAG7mZNRU08jN6EQoB/pYRlz14zhiKt02T07/Y72nO16jIUezsHdfTk+
wgmojftQNsk983mb72PGk7nlddH45ds9S/8g1rYugfYq+vpggSbnKU13Qe7dur+s
1r0bTTI4YDYvKQ9NBH995jF4FpSJeer8de5ykUA2R0UULBcrTW0GU/ugRBcZKO9e
W3O26TkFG6+Ic5/1LDtrdx7tZyNx/QAAj5qKeCJkkCr3C+slxQ2TbcnH5o/m2pNt
RvLPF3G/xdBkr9Hsc3fkNejXVjrEZMPWB/tuWta2GTJwLiafhm9ZTtR9Lk83mMy7
A+Ja47Qj8j99ht3OGfQ8tjxj+hkDfEZTdOvUwICgw5XfstPzeCoU2qcrxHhkGckD
vpVxltPU3jGsReWcXH1xL/V/FDNtLX5Qo2Jf0NgdU6NDjnI6TYetDodRb8lBzBct
y7xj+zbHNR8XGuOP8Je7lYX1rW6+gRG3HQN3kkMC2kTdhV7dBRsvjcLq5oaupaTm
E4GkNc5oDepMa3TtwDQgQ/i20843ce1d0DGcpPAhZaBdNlwhfQz5bkjntwxjFrHv
nh2VjqgWuhp0Fqhs922i81K6xZsa7cvlHcMXdBfi5PpQ+5FLG2HvksxVFG+zZdys
XMWhHuXVVNFTZfy+PLl9I8oyZPfdporytkpm7IFASFoncag5tBwsAf/AumD4MEJJ
G2ERaBMPii+2UOwqCC4N2zqEHdK5HR6I1XU830pQQBoeulwNjmGiQ2ljMZ9feZ5v
RbhoRHwSXyVLp9T3gw+uRDZOc0ch041KDGqg17hnGzTaTFvmrLlFrpJo/CJlVDl/
TB9ROqNM7xErnjvW66fNVxlpSCptX1KsxTXHMHgL5MratbWHbFyj4Hln1+ovrmgg
3YuDcDmGyA/iWqPzs3IqoQzRyA8gAcphDYmarnVIGQmzqxayhItm6umu+M8oWMoP
PDquwSzFlAL3A62SHGI1haeDu/WB/t66AfuxKaVbSbVLmHKrFFV3KiNiBtfk/V6I
Lsh5Dxdo4cZx7hJ3hjMcLGl0Ut0RzQCxbupwmKZwanHAOe/EFf8IqzCjOKaYFKX8
TK7lW0nKJzBcly1yaD442//IuqLUOW/18AxoHz0mDQ5PdewbHru6N1tjmOHTyIjH
DFf7S4DEXsPDrlewdaR8OwxsOvaeqVmpQmlGT6/lxdlnCEjwzBDAb2e95DZbMPH3
op31OSppZLeomEeZXMnUMF+hZ1FTDj3WvNBN0V4wXFc1GzcYSE076so7dxUFhCox
ym737HTadws8I9zWYbaFaMjnj17mwkonTcvtxK+K7EmV7SFKIOUbJm/XaVx/bfBK
dm5ItmE1I3JZjnmxMkw5oxbevVx17OkKK/eaOO+DzG7w//tUvdi4+euVTG0NFNeo
iODz3RYr0RImJM2BJ6yiaqWjFZMPkqyJr8ZHiK27X0j7dk7vUzmdOViRBZg5MSxH
JidxMed6AWJSUyzsTU9NzEK6QFkqw9Y6Eyd/p0m8sdweYFSIcOlqTtNe7vBZiaIF
TSLRQ+hZuUBBMgvAcbeHtUguAhlbV2kXJQYwi8/HV//yJAAFYhSHtFNbYZDZcehp
+4ijT7oQ3grEDg5FucPFhovAoWBhPYze3H6Nzeu511dP6Nf7e/X1CMp49Ujs+AVp
H4G+B8pScVHFYLjFqXvEcXTi+BXl3OJVlHFAqUGfKcsmq7lPYb32H+xjg0VRj3GM
V5h96DCyeFjyqczhkAEgw786++S9KzAr4dCIkxnFlWSs13Z1Lexe6Hk5qkxmnJJX
NZZ0cXfV+3jIgayuoslSFTbVBB19srLFDbZ/cAa6eTENTmSlZbEVifRxu4c7q872
gZ7p7ZqFF548MgLO4RK82BeoXnceD0JUj9s9d2uCgaCIo2scFMEPU7p53zirIIwe
OT9GTNcVZPc1oUWlsNU1nEmFBFkOSC+mq5P4w9FRZQKtHaTcImbhyLqF8/Nl5L/F
55UEbDhoU822Z9U6TO3FdIZd2sBRzAizSV6GfSSJ5rz6btpYHf7aLFg3h3+YFKh2
YJ0qnVt4kCdRIFKWCTQwMii//leWJGZG4iaGEuIm0QL7QXoip9DQIPLe5zHEGRpY
2NFQYZjaSM91mEfedT8ppczHCu72aJD2+DZzkCTrIVDswK4qJV97oWZkQWrKJSdS
jeMs8J8C96kH9VCQa0XmRf1+kElR9quPyhbGEXPlThtR4Bq8mtxq7BvtN8Bb7fkr
9OOSdC0tl4Iedi2TfRJKN6HApM6KgEQ4z50fuYVImVGB68gadf4Sf53FkKorSvxp
ZRRV19nneycMhhUPA8f+rQvlkIpwKV/j7Q7fggmcHSaRHfQZNmKdf9SezWzy5LB4
d9+vRXz6dO7MhcJaBxMgSM1838DWROaqPVxMQ9h6yjt0k+k5hH+YvrfuZ8k83IbW
l/bXARwm+utU0VtC1N+dfoTMX0UnDENf8pUxQlnJjbTgvwa/wOogRKL59LeZLUMs
sC1duBDAXw63JyoeE5HAyOil90anurpFp3gtLqjTeQ7adjkgTTddgIBzmk+tIkLM
RKq/xTDf5gShaDfOSUrWJ2te2eW7Tu4Sp2+4D3Pg5kBG41aquhpYahS4282O0WO/
NzAtuivoujnOhQCDKlgRFONNmmvekSaNaodi/+bXRuftsxiSHeXSAMVYARBYhPvE
FLKGAxKT4bKnpmLZNrkQQhhrFaxhplm+N+Wr0m7EwNBNO/I3L/WpUjq2AUDmLj39
LF4g/mQ6bjCmn0Anh4kPSBVqXcg9e0U3tdEHGvH+mZkL3xjDZs27WusciMdN4zM7
SaksJ/63y3cpurLio2UN8Cysua/b3Bg2Yd1jAgx/OUuopaLSLMkmxsgLdRyrseXW
TliV4Y2EUfbXxuA+dIu2BNkwMxCjN5nfHN36TWp5exaEF/ScspRq7SPYEcpJN5VX
9CVXd+Xiwk8JpxUpqQSiUoLbe7BK2mlUNvD8q4Re6nTu126p/1j6/MChz6kWtynR
Hvj06yeDDQUfezMhHktuFuRuSU1vZtwFR/FAySwPRLCqleuVXEHFo/Bnt/0zaHgm
Bqd6d47SgQFKTwunHgrr+cT9wlxHlx+ukx4WNHaoy7EE07pNg8773UVirHo7GoIp
+CYJ7OccViZBPD745G3lMh9zcMYZ8HMqzizrYLJskQyS4ONdrnI9jPyMYx22e0Qm
D2bi0WBOHk3wHDt6Ftylvljddo9tiGwg/FXLNiJMQS4Q0CrxxAk4I5Ft5mHAaGW7
96b0uhdZPXpU4hiIbqug4etSQxRriD9G2hz/4WiVMVsiY+X4LIjH4YRtWQ07w2Ww
QcMfdWPyDNxj2UGZuKL43CzVLatSnjTPml+SQHc6Axaeu8fGVR1Bi9vowYq5Nrhb
2wspMkzh5WjxEr4mPP1hg2qZAqUys0mqhW1tZKzh84g0gkg2niJQKn/cEZDMK3Um
zbWtjP8Ea/Ul6LsKecJBqshT/krkpTzSXKbhwHrQTx62OMEAogiDyUiLOJTDhwBG
8V/taV7O0FE0QrC7tPGtEbJnMgKbnD4U0EfZddDnPD/vG4qu2f4UEXmJc67V/PkO
A+B31JF1pb9B8t1k7RwEKbZN3peiLv64rTitqfoQjyVfI6Q3Jc5Xr9DOdirQJIDR
oA2LQa8OlX4zXGu47+WD3qIkxUm7Zg6Ow3tnKGqZv/sejuaA2eY6RiBO3F/sVval
TD7lXm/95TsexuSmG6ojvj9TfxZqhdsjygH/b7oZK/lZFS0+SCLLvmElSHWR1cfo
hLDpdicRrJ97WHxE+oBMDseJHs2oF05yVbogmh/rfX0mdaChJPvfUOioD4lZ8N2T
wDO2zYSey13/OM6XIsMdaUmbT6VOjpN1rwSFZiRBS7uKpr7Mxwv2JKZM0UqfSRYW
kBaOd0NxhiBkq/CCGN/x5h8XQMnux/+pZrne9ihzv8bChmYodIwFUvTzgIw47viz
VeoOYziSACMI8aYoazGZE4Cl4W2pjsbUR0kOFp6/VkfWDvLADOWTujM3SG6RdN+l
guhl13VOzQyllj7LKVkDXkzio3M1yEc1RQ9O7B4hAvX4eccS0RyCEUu5azZw8jH8
kuzDxoORe4RkQxtURozAehE7ST67ep6q/0aFPYHUwD+zSob3qESXBCU9Wfdvrt/+
HmxOrpVf8BVowRER3Xd95qGZMjBLOE/ExQtbzlmQtxk9M8Oy3KdkmsMGkUv6uqSG
0Wow2aMPnwGVU4P9RkKtiunGfMStqsgePZAGrQ61vclemf8tyiU3IW5lPfu1ZYT0
vSysP5o3dA6VpFtSkjGP2JeB6HjIdFRw0Qlxa2CO8KDUxxvLxKvCSzvYAdYjjK0T
LO6GkAj/mC2Rklj4i2lp9IW1uDABJ36APfGeD+tiny+CmHV3nlXBnxAcmLfIFW+V
ex24xnn2Ck0sSyCmt3e53zdkXpoKGf3lCC+RlHBwf9fbct2Jy8GeUJTHQbAHf/yZ
H310SliPC/tWiCRsqrRfmKhBM3IDFJye5rqlAiCUO1eFmrJnhwWkZGsbPIlDbKyN
E8GabFlMELxWfTAiWMe3MQlEc4isC36iaG7GCbcBkt2KO1jr7+BfysQ9gG0R0gQG
6Q0VFx/PxwkmuTFmjl9f1Zu9tEcRCLxtfnUWt/251wDVIiG526RhWDbzpywL7yXV
d4XHWKAvhHd4aYXtbB/rwQ3k9g381b/P5C0JvWzVgPySP+JFXWZO2ITQSx+VDprf
/T6jyy1LhzPkF2uTDn2bNzNWl3rXhcPbXC1ZEJ938MCsQeCK1YiWpL1GQX/SLq5y
WXiy+J8WS+9MJuGzBwgw3bvu5EjF17FGB4tAap9NzVPf5ZXBQIFm002dgC6z8Oqp
3CeBXAloHMuk64QWOTEi7Zufg2fhJwdFWZSgdSjnf757V8qZAEw8DuGs5Gr5M5tk
FD1ZhfeJ8hmE5rDA0YZfaew1YjXsSBVv3W3+knwHfsUJqNzjbdQcz0yv3T9ejjHz
oppXHfEropOBrCsg/clpmtz69e8F0/WQUvMZmioBAgK5RnwSvEu7MypWSuIeZo9g
ywdsmJ/0lvJDKGFtMF+tOcourD0iBO8A4+4WLEzwSWqADjK2JilCEINE+faakLgL
XpzwpLxXMrP1RdmMTCrP+RLfxBBbz2hTnBxkgOqX6qXgf36FedRdk+QJ346z8tl2
mWq3oyuYPQTOXEFX0aF2lMHU+/mc4dkFs8l7Kz2EnFE1AM10NK1NN/xIbA/t42GW
FzigRbjTwpOGEBSO9+Ry/KnUlTNl7pBx0SCZAMeKCkg7g0PPJSbn4UmvmtQ2KXNp
uF7QCyKBvkrgtVnaJT4Y2NDhwwI6fLUne7GR1cBg3fgkdOdG4kREuIqeK8q+ULu3
RlQNRrg09PR4Ovl9ZgIw+ge2ShVF7GQKKDNp6gLdx1FenejAXECj6a4yi9rdJWtg
gxB6kgA9vy57ZJhoiH7CbdTqpLNUsNGn8KUUXncOyV+m3LUrMw3dXYbHg5Cmm5lF
WMhscgzkprxMvkhtww2vIeMEfC2FBjx5mj0BwXOtKf4vLxriDL0EtEgsuWoNTcDM
rQ+aVj2iw4yRDPVv3PVJj1AqkX+luYd2APHwLGxVMdNV280c/5KKYdDGf33EGnIl
PhdBSL3tWGP9wTim7nehqlMB/8WdxDRgU8AolDThIzn2vETyw+sh/609bgqTK4mB
/y6GMLXApTGNBfwXKnY+CMNtOe3spwvQdPZFVF9Zz85yT1lhL+GPjEZONawGcDy9
cFvBxacRjsj3icO5ayY+9fTEzYXa4jhhfv4sekXnz6zfuYHYFd3Hs2/Cb60+suyF
EuW2nNY42G3E9bIUSBVjoKLljVH8tDsx7SKxAYFIwYxRXii3jNnSnDi0ufc4fILb
EPTc7wrby++hA0Zl84K0FH7MwpxhpC3Mv855ZZz5f8k1b9Cr9Kb0W5rQZwpSMQQT
VuXVQsTMnnHhIii+n0okm0KGOOyDQBk8cZftq0NGg8QSpbAZjOlBBZ2LY3lov5Ew
iQ54W2Jsw9+ggPCa0xYbypqCxTsK+NT7g9FO58vQmkkCP+0JevQbLP4uhhQb4vSe
/p76Gg+ag5hmYCqbvd5iR0lVfU31jU6dl4hkKmrp/U27aQ+ubcSh6DoLsePtZZFU
vLirbSOB/WkN4an0tBcvZhpgtWHU/pO45+xZwpR56Wcov44wwnOlFG/CcKWvN5lO
1HzR106bLRpGjvFzWnWjgubKb6Pts0mUpjTJtPyV1i9SXMJMYICRN9gReN+SoCHA
7wqWZteiZMRjncDITKQwt210UhmuORCWiCmEAS4DR6OIKoTEErtKCR5dWtDp2/+1
1/Euki6K3vuQ3Djd0z7mgetboseO/dk5rtlJaA5pxU8BHsLOP4Afv6Uqwe5CM5H/
5LkgxMZ3r6V8ZWezdqPx8UXPrt3zJ0cRadj/fGv976hVTr7jlAS7odiAOAQyspY+
G6Aoj6PC0uNAabmmZo9LPyTkxpltwe1iwpA6yqMLiPYmx3qc1Ca050Mnxo/RB/vJ
aiqn6PpK/ipgOMZPTl4jFK5Zlg7RdcNHUsRtDQ9P8MIdj6Hn7NJPduW7KdnY7/nC
vcE4uCZOOMRWysZe8UGzC6Wk9XpA25CyhYu5ub/zRsDNRSJJWTkxoAhv6+fgXZUZ
x7zrXniwFBIl1FJRsPLpWf+e+5KGHL/x3F11pHlvbepd9WkfE9q0SchhVAINpzp/
LniigSfge3DhB9LaHqtWyGWTxvKXVuqmhgPzJfyklmphHRkCLMG/Un3A7E+MaAqo
sNfr1OHzWbG+NkU2GJuYRV+zYShFUWPi+rjMWMSO1aONkRhpr5K+X9IdjW40upzP
WCTKvMzOfzVBbA+WAhAprC/HYsVCS8skZ+0fstDCwlpgZBScpELwMhSOYBC3GiEF
Rilb5bjTA+9DpKa7NRpOGydXTxU6nTkDr/8di5MT1tQCZgiEeXziwh9IFjpAVq/7
JMcExqMqqH3OIYR8rxBpKwAiphTmzWLd7bbDjFzkeRxzALgA52D9rVgN9Fa/8lCG
52uLoVliWzigyNi7H48txkrs0nbMzQOonIc9XeH2XHdWrc1iu0xyY8tiSOOFNXkG
+/DHpjXXSgnAcKNs9HCnIAflBlwgW2H3XNj6KZS+3jPMCS2B597UOVN8JtLRbXVx
egMRkGBrbUeMUtUN4IT2fdR4g2gmnhc6E4qWYRzbPyObL2JP6u9+f/W9+kLgymWc
r/0W6IDpEa277yCpeXIX0bGkSBn78EUypFWzRqZm/Mkti43+CHAWiiVJgXT4bpfR
zrWxbmiUemgMmWvXdF7lhpSkMoWKUnQ/MER77Xg0GavLHtCztuUqBYfRxgAPoL1z
eoc6rvAusjKq0N5wsiVnHRNJY+YTLzMkWx6lXDg3S0uaOgmV71xxWRZ760T/SEm/
Ex8YVvGYPQzS0UF7sabwn0/+kp56RqI1ft6opCDBJ4mJo2D9+BMK8/Qej7aztAE8
r4v3v/m89GxIIo95j4p2WhX4bwEWvtPF83iDNMUzHmHXjRrIkARF3lCRIZ/QFQlH
YpetmostXKHFOCprVx7oQKLQQ0/nz437iN500M7xk28AxFeCa6+CUsUYABT0ATcg
02KB50CC6gWB6QnBE+zIL1sGmHquyqJwLXn2Im9Gbva8K45FIaJydvUyaE3eck69
iUkABdAjuiv7ebl2AUiyrttNJzfvhKk3DIviklr0pgGEl0wG1oaG0yPKF+czomCq
DlvzRI2r0OlAwUXSFhqM+70K7T+7bt97LIJH/F10V++HpgOh1xlDADKHF0bUwMuu
v5z9Wgn44QD6KqqXhkO22ikfo1zFGZ5tcnVu7eYXkFvqVlXI/SUIQe1AfwM7Wcr2
pCtWft8jxjfZR4p1sQQDUSjXoWUcPgVXLELL7Y2rSiXQbU4mSDKgHm3zyzVD1HlV
/al6j7Ix7TOvcphrXmA6iaAo5iXfH/LTr8j3DqrpBp42luaHUi4CBBNC/JE71YQt
AbB/QuwCG2NOZXqwBMajeFBVCSAk7+v/8JcmLtJkGJJjaacX6rF9z33/5Re0+1CZ
2jTxqnZJBXg3itzTex+5FslQXnHhl4g4m6ZSz60zRWylazO7sXzjpaOiqqZqetmH
eheO33KB0S0Eu8JBT7g6IaHKQ81cd3Fwz2b6faF6lORNGGPL2O4x7VT6ognHOgAT
cKhuL2JxRdfAwvI6ha75n3Ve0fkZet4ELjBGVBfMfaW5YNu7skmyHCeX0K82EU9M
DPz2hAlIInXG3oOKfNLihiy9kk1xkWqRas5cVAG9al+bMtdn3Ch4fYl/LUhx2/zE
DequXfHyo67RVmZJFWSKBkQJJ4a5Tapf5OBQ0ddEAYyKqwQ1hy1kVf8imSu1c6tC
RxJim+YOzplvSchPnpZ6DzZRLMsc4b5X3pxNdUgzOZdwcv9Bmti5+qq3lbo/hY2x
c980mOCAC6KNWw6Um1pocAu02A8u7NWXgFK9p2FnKfCncIiL9cuIL6dPS8OWA40H
RbgdpRPcOO/tIPfqQ/FPJmyw/EC9bzrDNXT7yocXyQClsRmLPwvmB5zi5GgA+LhZ
peu0SIv+mhMcxrPWIFg8GnmeGTwO+r+9GLUKRjf5KJXRYLAaADzC4tL1tvTYQi/J
Dg03GbjtiAhRYEQ6oK545wjgALJvy4dP2NQhdvW+qLEa+J7OUIqgoThZ7nORBpsr
Z/44tp1ewFdrZfK4uGwX6CaCGzh+O++oXEz+hUTXSYo6htdw0Up6B+r56otmZ2ye
0ceVLGeKBdRNJoBNGnHaVHPgWy1cxq2ZN8uqR5hEeJ7eQawXIpkUVRoRnpQz9/W9
3bntuCYX3ZzWCCa6brT+0UdblYEHyX/7QKmsFbOLZ0IUXEekxKvXz/rVKDzUR+HH
UwOrHwEW0KPEqfY+9zWMQvf9ywA4P/upXPAwHBuY3ympbm83gN+bsB0xWjAFbvRo
fJxtl5FVK6hlZiLsHBjAKdTWaEyqoC6TLibCs7fnI0DnhkqzwEH0bUAAUpLjYOjh
FQn1/2xRkHMRSTedmif/WmJBDdxpQCDd2iz9YSVBhp8t6wTTOxKHMWhnnS9orKGr
/4J/Kkc+J8iGvoaTmvArdr21m/t9jElxc0OwQIFygzRLfRzcjiqUFZP1yCrCL6pQ
WzTLy137HdEntQz9YKMh9kvi7APCXJuTIJDFK8bfnXpPYooUnacgv/+X34gHe5o6
yjNkWDh7ozBHy51gIS7fAWqMSAqMTpZLrK6yNohDPlzOmVR/SKW8GHiAa5qpxCqO
pNi7cbTKqePjvubffb/2fO3RNJ9TMy+uCFs1DWI4NAcMmElZ2wcXYyjxj30Tl54b
winnkjooyidO/Ert6twVytjGh7gzF9YSRWvyXYEmKSUxm4+WMjL5IIJzkFfU3+fd
D0zmLGs6n4dAu6aYwwPEaZcG+onsbf4zsy9tUKDGtEgeMeWbdLzjmzEq301vjpHA
5aGyrQdJFqe97cSxzp81YdUVFhukx2Kc1zxON9KgN8rZEXMg/tc3zQ9mUlt3XCNO
p7KwMMXwzcoQFhPgkWLOLdzFilMgAQ6yio2O3zAhC5MPXeCSYZkBhPfPBqy6oS2p
TVJtFW0XqfVGzkBEMX5t5g20tJEWN63F2SMNGMmlIJZv9nslvW1tJk7QygaWQBDU
okH3gijxE1/RETRqaUNBpxqmx6sK1j0DG2RVs4jRqMaa1JJin6xlgMBpzc7vayF9
FJjtrD6i06FJbMWns3sgNfxqp7AIsej+5coFwynOIImeWNbGWn7kEzvK6CUG/grk
rEl6qevKTY936yujr2KHbRrHW34ydkeX9kAeFPLNE0EqgJFevNTx9ipksn2bdM4m
09CUmOBXbWo40mzXXjBsGqZMKiZXeFGNcgJXCMcIWIRZrVj/IkNBkZ2H1aCaxE4l
bT6ydZ7qDek4fEMecG2gFaca3FS/U0fqsz9lhr64AVhlhdCelAJbfd1dbRg2PjZn
7SB45MysmlVhxkSqNTOy4h+EBqGJPNksJr7BPn7hLP6HadecCSQBJy2NSC88zMhf
NB48TsD9SOblb084LTgFGY9iHArSrftkOWwhh8qZXXO5mns1AtWbDJ6uuPDHpoJH
6t0EOfhBOA4N7czSbonqbwrZIMFOIUyXlojyHSuU4JToE4Xzcg6CYwWqJ5Lz2CD+
Vw4uQ5KxJjrnYkJqOE+x0vdwa1ITyL0CMLS3/9lBVhYvLp/2aq7XH+1i95/UWCon
XoUdt1h0IW15yTVoSVc2xy+Ez4Dn1lQN3J8f9fzDWCR5ioEYRJ4SbTGatuK6u8kh
aNwE0oqPjcNBZZ8ojTR2Qrl+2HaoorEA4vD25wtcfkOPf8EDPuMmHu+eWkin554X
fOP47oXInuc3WSRPmaDrFmT/emqf6pA51FQtPCikQdG+pOT8tSVeEEk39xjHJJfP
FVX1sD2Z1MKGOSHD89BVn92OQr9+tBMZgUCqaZq23WQRJgUc3OSdlhx8C9tgC2pj
QAp8ot7cU27p1IyMT8J77lpA40t9bAzAylizY6bzhRqjuuuNPczSCkTpF8a5+u50
fQXQdy0kyKCxk/qeUmMl6SXgTGQCsQZ+zK4eQ6gm1LlUXtlY5l1mIZxwW6nEkmqd
jvIAeGb0DckFr+Av6pwd06DdqsvQ/nbZu156O28FzE8nbMsfOeQRVcfvQKZHoR6p
g+VttvXFyR3inCfwxfkpqzfKt15/muHV3XI6xXU75RAT/n2pNOqhcxq3hCtmrgQr
DnkF2b3K9UQ5X2Dam4XIzWzd1Vb/G4fIFpkmeZ29yf+D/RI67XcUMHuMoc43W3Nz
LpL82qT97no5dxAHs1xX9ffqSE3GsGUicRkkcpu4/6yfXDyBtit7Y74N1DLY3aNv
9wsSFRp89NfiZ6hxi/KuXb6e84MA8kCf2V6w1eBXlH9tDMOXhwW2EQJwK54n4gl7
10acbtsfErPfWpLn4EauZxqMSf+aAzKgrowInbWxklEl6PzQvPaPcHWo87WWri2Z
VMqAgyqkxK9GyhD7xFYm604w1QtvXeDKOPfyQknKp0eBk10r8d1z5VP2Pl8/0gwV
Og2hlBppReOB/cedr7XnpfQCddRLfx7KvcoluSn1pHqFJFucj6tzibdf8Hg3zojg
CA4uuMwScQltHbPh1Oqq/XCVAGMen6rOFAnSYCkCMNBb7y+U7DmnAORUvkQ+hRc1
t6+GhrcGueSSG7t/X904VuywXHGQlEiBxOseGmTkhk37bsDjjNSynbPWX9miNzVv
GTdBwZhpspCb11+S7t8JFAowG60TbA41V19AGgQgyaxwkFLjWeWQdUAc2wxJUZaE
mU6Joyr0yVmusF4OHIUiANYiurfopNq6OyWUsmZm/JU1ceur1dqLEsug/sm/brK6
bbxz95BS0bUv4/1V0RS1WTf2LPpC1GRQIh+OhQAQZl8zfEH9PwmQNgzKsEeSLiec
sLqy9n7QKoZwr6K/fugiNTUiJYdra3Xn7yY94pyWHC0DBPGVLCUl2qbWWufkIMk2
APu7Xaq4iRSrM29vRgRwNSnB6ZrGX1abVfvgnsOzp36eJwfdnu60AhoP/X+ywlaG
/fo3uaiPOMIzWCv5/eyFMaX7gJr3+rQRE4kHDczb1IwOvckkTqfTtIlykaGq9ilk
KxRnXh+8ttzRczU+b1djPQbyDYlkS/yG9+2uOuGOuS2Hbbp0Q+EDtq3r316QhaUY
+e7Sr/DfLkhOWFiwmvraoQt17dxGHQWw5toWswA2hs3g1uecJCWS8IWEIaEaMdan
HO0T4nAm5+FV+R/Rg0SLMBiJspyN33mmRHxiH6npC5KpuSCRy9qr0VIPfyvsj0FA
tLNldwjg1hHflzg7Arip/9NxHWqPYMNEd6BhsowSxXu9c48gwcE+B/aF1ZWsF8dL
zeP614twSw4U060A+OtIELeNeupF1Q2AioMMOx9nAEX9u1XAvXwHO9K5Bx1ulIKR
RnGRNWLq13EiO74HAs6NcbnHNq0t8l1WQyJsyeP62LKT1QxgeEUbOKCEQnJTDxPt
aeMoLXbHLTNJDDioxn8WNxsWf1Jxn2vDoiDusF3LTbHSdBhStiWzKH9ZaNgtXlb0
Da0RVFMJ4Bzkm3IQTYfVuzw/X8mGo3dSidHdcHN0/WfwQQO1gaW/EbStwPsOwRno
NNvA38TFKViFxTmcVG++ov3wfPzSVXkzwEJ5oDwgUWHxT7ISW9WeIK7YX3RNNCHb
3H4cLnIzFuTY4ImlNXDTGyOQei4f+28kDB+vDjSQpOSBJ3yo82yCbgSNHOlDT6CW
cb4sZhSgerVTm6xJXhIsbFM5ReqrF4yM1XpoJc9wapAvcys5+etxnNjgf8ypAsy+
i3OUownfvQlFQD5i16zCPp7mfSIdi5elw8LqxqiBQSq/INxYkeTNxqHsuh2nF9kE
tRZncAT3OwEfX1083W58IKrg/J2zl9QrsaIWH4VqRIiNAlCDksbvHVDOF6incgY4
QrEGEQ/rHCHpeDqNDhUeUGwl275nhDalF8AS55+XscWplsTzc65F55X2vhCa42le
HPwlF7gFkLvpgr99kVd6840GHIT06bpS4zhi/uCltTqFTnAIqkBN9XlzxLdeScmV
GeZhJxoEcMazF1C+QEnvbEcg7m6lX6/FzcpNiTMaZ0AKkUflIn2cvX1PthIH8SyZ
xCMHJ6xOWNchHlWsgNFrk7asfuXMTOi1CfycqmBQpBSX3yMWRbZRoNHkAaB75Ywg
OqkUdJM4qyqx9M70Z0win10BoRd6z6ANlnFzz8fjfMmizhx/vGT+AbFkPRomFF4r
wbHChKScUckSl5lNhMmp5prWTK+z0xXCEMvH1hZMX/A22iA+G0s8VS3ZPAFVsgOu
F6k8e9+u+BTjI4KvBEqHm3H1mA7q6jeYCOa0FMj+LzRrQ5UM7VnQ6LLevccd7ePm
tHpXid49HfbCsuVfoK2IpUJ52/ZHiDxiNprI713oNZtOj/A7nMrKMkTyoDWKP642
alxW4gAi1jbJhMXbct8Kn614gl7BNCgisyzpMTYcYMOY2xmBnhjjH0GUhukf9AWi
B5Owu3gdB9w+wETIUv884Xuujz30RiOUSahbWCLS8L7uXRHl+YYMdc6IlHcaHLxz
rkTs7UDfau+NT+4Bll3dTigbUhycLS+zVvS0Tol1yXPcyJ7Y40PxUvK302uLnYRJ
JalAoFWxMwtcXfe0UD6hLkx7hwkVJt1jAcczik8EDovYYL9FGqRfZMo2V6ZCoLJ8
1RhLc6XkJpTprFnM6onFJONOmd92N5Eh9c6irvGttC2Qv9h+9xDGTmP1fsTm/Djr
8BWekeKq/Ow1T21febyU50n20D9pZSJWQGXXZVXgS38a/kw+mhe87OjQUB/x76+c
nuUZGcFfFhhvqPD0xBmuajuEgcfoqBgQn/S1yuL6tG5szzJAt70lKwi6oJCHp4kW
P/BIYUfneKbpdaR13jTVLMSXeToAyYVAcm+v/sOgzDlOea5VWqv11Y3/L4PXL7So
ayk10ARgsjmRUb6KV4uTH7C60+aJpo2gwYMqNRzw17EqO20SqUcNipl5efYZm4t1
OTvwlCLG82iMz3M0/yBKU0P7HifZ8RmQrRoKHfWNLQjRDMYH/9VgK6hvsmU1tKDs
MKoYJ/DOsExh8KiW5qSLON9GHl9zjvkRTP7FPaxzjwnU27FrigDHpCpU2FhT34Ji
5fpBfqBTVPjiFFPxZBLP8aw3I2c8LpMy/ZlZHO2+sIicKoZ1MREdiWZvERjLZOal
cZNA9BSPYkW4+MRmtYsHooD7sJWO87/6ks2/YGY5vXMWGVUc9oesnhd9egLhLfr7
LTDKuiW5ZCBl5xWlmzL+L/I7E4iSm4YP4qdtM8a2j8w3ATKuEwCCMvJPvI8Zz5Ba
ppw1vksF/RvCOF3uR1hO9Y7BsHM6aIalLrh0NeN+0YPU6nBU3YJt0KOpeUlZ/xKk
OQy/L9oNqG07uWYT6fiEufJVXLtOtPbb19SFRMZ33KMX3sjmjN4nOtAYVWsf6o2b
a8rLGYj5ojy0gHXD70XK5i5VTJhbLI9Z1rb2CUY/56PEM4wuKFFa8DR1aIX28Kvg
Lbn3E1yPpMEfRQHfyogBtEke8YzZl/aVySgdpuYphXBN7zgP69/4d6WONAipA+rt
heGnGHflq35jc4mrCbsUOv1beJDSDzOghkF9ifQSlX5bK0DGGfDGj5heEH9euxoS
AVrfaUPkton49qjiHhIP4V3rYczEeAA2VWd/Jz91ft52LOdZTHbk/5a92nN98iiy
Qcqzskhlu5XTPxq5xYWINVTdU0OFzcqok8NfqXuo7V9z5SkElQVulIce96b8dXQA
9EwSmBXcNH5rgpYnWdMEOjbzGQNIs3VfJDBJS3T7cESkWpTFXoAOxrdPDdaZgq8z
hnGJssHC3FLeatGBgU3JAINkbxMjMjZmfOLmS9w+fn42vcGno6VgPi46xmf6qG6y
39S9jCJpfbjDs9AG0hTcdXdDihRLcpfuw5ccOo/nLwUoPkfJqh8py5DPiGOP3rwV
AIh08iu1MNhy4MAr3tDeeMLawjNMY+yMl7A8Dw9DdjTxakUG/bbEGcUVv/rLu1tO
6sfy+k692OoqzqtmhYMdxNsdlF4sDOL9APrOzCajhyZGcppp+oh1PU2Uj6tJ/+Qv
Y5TEPu29Aow0LXx+f8xGOkccF6ILdm7NutDCB/c915fQxxQmj8jEMwpZt1QihlI9
6dujqMdRvcfbePD5zZ1BgiyNxaTqEbQsstip9LIvENkUCNtlYkqymmqTEULSsgeU
nLG7rgEpvGDLtFFfZG5f4yKEwBropNHKVBo8jikgjFFPWKdeI8AJP0FGSya3jMfB
KeYLJh2cuV/d9jaYsnaOsRB72y4bTGnxR4bo1ubYFvlvl35q2gLiWJWJzdIwjn6K
owdAinUunV+K+l79Y4bkGB5kBZJNtBPpQfOLHVQk/3kXOPVJwll+ry7pAdU2QJ6o
rDww5tS4yaHv8nA56lMSa58Oaw3Z4bvRyrzfc5XJR6xJvmIm6Zcck75j08Bdd1TS
i3dylpi4hwJksEOshE8ePWGTAgmOepAeF+etu18lVMHwIfywHoh3C0y1+yMLQMJU
laHO3NWQQkApcsk3TkxhrJtzxDKqDxtH7Lf1jr8DQXrNRWKPn8Z2H9CejtSKbsda
RBGbg/Q+FdLUGDgK/TAyY6TsJNLs3dobAtvtHITo1N/Poql9uEJ4uUmFgtw439Iz
kkvXy8noQ+8tPlkoxN38mTsXrQBRnzr6+f/LuJxv8sDN3ulwmZoq1S/3luaBdn19
qetc9p0xkyeZ/cHJ5NzCRzcojXWOiLYr+ZLdLZT+OiTSlIvRNt9/GEZBUImkgx4C
g2CWhegqWlqNnS5MRYIU7Wyx1lenUUZsGlTSsG8zTBo4nWF8Rb9r1rmPox0bJhxw
hQQ8nq/0a62XlnRWobztA14K4Wp0rzGVjojjBEBUken9g2VuLP2HuERJOQQ+4BBh
DUyeZaXqNeHCBrguG3NlSCOPyi6XhSU7W+8YqJY4+G2kiayHlQ2WK5nASbqNWAqW
mU5N+urL9t47D6lkErr1i82qgvy6OvqLjFCIoIOwTei+In2q03HezllDcsImis92
Lkmx45QSeLYsqCfkugEq3INSfCj4o8dBLKnEImnR4maKyWiDF3KEMkNum4bjarLg
ROtjUD8kFcmhsw9MSA7AcD8hwuk6Mc3y8FExA5p1VmRuMbA0VMu/kyYolfmeBLjL
KKF+6cyUUGrQXnAwGBJigOiWWTiVYaG1pqIDa3sQC5tPLKO9wnPgdIycjbflUK54
xJiMk1R4D002uBJNsl9b1Q7phCUcjjGDnTLY9BSZQjPPC48DkGGib5Ai4lxwdeJP
CgR5yXDh+jEDNBp/c948Naxy4V2P2Gd6jIErgIJe2EksP39UsgAST4jlxs7T6Jqm
+j3otkjA/VkZ6UVlj86FtRRvk8oFfKDRdkY7yMpTcOHb8GSdNW7+6phgm5X+aKyR
/y3rFIcR5PXuvWbYu53B08MOZCFTUYJXHUEMs9rwZeXGQNHFYkaFRhTUD2w72Bdr
Md8gLJTnH01GfuWt41Zm6BEfbCzObW2l67v3gk5EVVTyNZrI4dCaQUn1fQ2ntnEg
q++l7pIc3s2fofBUhU9LKcueoFFnfccYKc+Ut3BCDQHWRD+UCp9u0PEeX1Vx4F9Z
hWhQ/0qsYyHvYBtHVXywNrKpXW9goxy+d5JPZfT7mX75pMwWUVt7lf8gHM+JNH35
9NST/9PkqAhJw456ubSc4HKHBhccdlG78sCFNMEO0tltFyhxWZ19iJz/OLYQJMf2
NBOkQ7Bzi+N0g3hW47Lnix1EwbNU5bE7SYupoReeGhce5Uu919QdGKIpiqFdMlf3
iAtKmr+JHUY0cNp23mQ872tGN8r1ZuiDFFRCjqhsVp2MUDlYa0OxKPV+83YiCk3B
moDm8asDkr4UGZruL0r06tx8SVsXPKhjC/WaOVXd4FLRw1YZZWNuNDqzOaqyot4j
vP8HqPlB4j6cwr6xCynZh5fuVBgQ9+l8ZlcYMmIX48NTjTld7aCbKyLvbYl7XaDI
QSZw9dqTGLvJNlYJUy73DLJSmaoSS7U2diREH2WE9TOhPEtuCy+J30KHBfccM7bH
jsSC2m6qc+N0Xs/1cGbn4WLsCg68/nS9QFWPW2+39ZbUXcJx4qgJxJo7M7XxbmCK
kG+ijIkalWKN377VBGVlVsg5pBVW1yK+aUHzjY5LMtGCz1RT7OVnrB5l0WcitcMm
UUhH67xvoWecrhdfAGabWV6y8adoViq8Atyx1lRO2afCwyrJSYCmErI5ddJaXsNy
A4g+ZWz/JiEMCTP7uQ0EiIngkaSXamEee3+m75OhpXXuiVJ94t2BdRh5A9FedPXg
GvrVRJBvppsu5x6iz9ZCNpMLSrdqMbg1qFSDrONgtNZNXByOj7+XqICOataaKtBk
ByTV+spB4MWruMDDtK/oO0Hdyq28pmQ+V9zOcK4iFc3x6tOY/r4ZWT4b+8E+U0bV
vHTUtjiQDPU76tUcXANLhg7ILpO9Bhtmgq2miaB2d2euEvBhgc0IpUYR1WnpzL/1
aleE1edR7xJRgaWPKne+mwusz4FzCCCTeUuDIFsoY2TsXQTfuVDTp1zSlRrVDwxs
yfKaL2W+YTEbUyBFhejt7xfwrchMxxsydeaZyig7wSbg9UWRcbNka3YXgKRnQL0J
pYmDgMpsxLczrhCSE/CyrJDp/0/+gsuktWbelj8M/GvyEe0J0HJD5Vl6zcOoas/3
vnnxWe03fzXJVSCFQ3D5iELZ5aPU2G49+u7KUKZNpPMc9dVHdltC3VimBOMGYhXg
5WXllIUCdfSNMgVDUZKrpl/077aCo6rUsZyrmDgENJIoom41ahbw8gaqn/8o8YL2
KYh2MTrOdDSLeE8BWOnyFvyYJ9sBliGq4g4gDSouIb5bv2ZSEAac6d1e6fGZzO6Q
BaAhxXYMw3COMhYoKMcjFcgBZtDhJ2nCG02bUdTqBtbJ+QSelzgEa6hdXH4VLfW8
FYOxEk7aBFLXjKwuzc4QycyUU0FZQdHAkHXlv2Ej5x2l3vehnnkmNvrrGMINpwwU
8dX9hsQYiB0WAuzrwglYGnVTZ5/8dT1sqKYMvjh8Rhojgn7TowOKXNcs6RPUfZH+
QfcZmpyhohct+5BxpZgBK6svSzZMBXdyq3cSCF3qWqGESAuiacAY9mu6v4rIkSi7
/JZ6lUM+G+j6uYgXSgrAJLPzSqRnDSQaUyf1QouZ+XjGWT4ZV+FxFVabSGp44y6N
w+siXlhxpOEDmSZQT8QVxjISRzJuMJW0Z7AHD+MVUX5AoebCumFhPL8pCCCaNdCa
LJmw06Yfc58+Bl7TmYNOR3NsaWORtqG/CCsukrN8izByhkQTv8taOV2fiYGJB8kt
DncECr2LqcrnU5lgTR23m7dpHBH7nw0jocspdI1wELU46qT/JVdveMyUiwMFMcoq
H3atvIh5kboKGHHz4gi4JBDNVVhvJUEp93wtSb7lVb6rgVExKKeR+LVIvsYIO9To
yoJn35BrlDxUF5/di4kQy0wa6Z8d1CclW0qYlkMdwiszwPPNC/PV/P3MfZp6th2I
MLOC52LjJosem7VAwgnanKCGwIhRfOSK5dYIHXgjDRAJh6yLDVHh9Kye37p9DOfu
wKk34jVVW/UAmzssLxxJsw/d7IHi3PgsDOUZE8Z26bgo49mkoHfBr5baC94RJwIc
mtCxfWQVUOIY94erh1QfgkrngDU+Oiz6pQYCH88pVbo4azU2RUwHpYCIcALaKO3b
1j9o9ogXsjzR8GW4hkqGDoGKFGrrPslQl6kfTt9CgCvwEc+1ziQuwxnv3DGJ7YBa
zfLWuSKfKzrcCwadYwTkzSwfOOczxeV4iPwi2ec4khC4956akMn4Gqrf3+8pPQJg
eX6hLb5b9DaN5870gwg3mnHEsS59RzKa3I4FmJkoxSj5pUWs9QXT4lbinNTomvMi
1Om3AdClRtvjA3ZiLy9JRkDZ/prCkx3u8L+fpIWNFLMNtfPLi1Vr93FnQglbrxcG
53yEiKbwEGSI8uLNeEWEc2zUeESBZvjLABNccqbMzBUkM6Nl0gS9wnhJytlhkwK1
V4CR2qG+p/YFN80VEP+QMnJQTtQLdjcTVchVbXXyS1RkfsmVKbvKh6efxbgmrX5L
OERC4BF1A1tXiGS2oHub+CaW9cWjXcm9C2DeoVudiEbNhmN3XWX3s63UFTT8rV9T
gsFBOi5oQ9rgirSzoutHB/AYBykIelC0medbsZB33e91QfFmFn+aeHCXEt7bE+9c
XzkTRNTeLzE6MtfNayCc4z/q0V9kUqTwp8Ol0z4CTjH3Aa9GtkgnzGRc61RtO6XN
knEJap5NmAByLNh+2wResgwIX290Ejq+4dnYlnFEIncy9v1hPxj4JmEiTaOJfMz+
IDWS5RhV8P0c3rduBCZjZUH4vIQ7RyPIEO4/uz/XiPQ32xhBUGBLdy4cXsTxbA7j
k1OvxPB6TahsRG3W4BIBLkxu9TWH7DXqbxaxT5lzGXowECtOG875J+FSkQsiocpL
Z7v/QsEAmtUnd6TPe+wtOAd2nmi79iYfkbncai7o5hjz4uYhe11qLRmFyspM/esA
Wn/fsrujVqP4FcSGMtmbWQFtQ3cSXRuEe6RQgnX3pFXca5Zd64wCVUxu6uBR7MV3
B1GFOXz22+g+yWyuxw187CWMyvEM49X87E5kYlMNKNVr7QS5NvQl7+fhlgvcVO/u
O/rBxr5CTRp9rNn0NE0E4jnegCm/aVMPUHsTZQP/kJ2/gHBn6tlxzyozOzIoPD8M
z8tKdR28DmdL9rKG48Po08sxY6tdIyIZCGqUX6OZ+G6eS95wQadlZ5U/ZMzKIS8Q
RXDnuetCG2/hphY1WfjlTgVMRNobd7AQFfMSKL7Ckcfk5I4s+2C4olNZ6FqwcnWS
g3EcmV8BhEF8/TpM6jnhN6uSEwganPdIX2VXsCbFHmu1/bl1dAhEHcn2vUJQ4OF+
qwQkYKi6OgVIU8YRtXoEcCNMrWRI8he1kC/gC1qQpSNnd/ZEDs7gelCF5gm5nPlI
MbB7tw2QaNwCQFewAPVL1us6WucHwxChk6gIVLmP6Xw1cNVVSkNgFEBdhb/pxIit
I83AbZM8kbAI7uuXay3FEW0IWgH1/bu3PsO9Ticy/KUHUXsr0jz33ORRUZ6sVzPv
F/JqnRhT9kYjfqkSciAHrBseDKZIVMMaeX5kCOiyfuZQ7UQk1RFzWj9aPo9Jbl4t
CEDZf3zeCBJJWxnTD5NvruT8qxePZ8QkxeK90ivMLMPkCyo16OIV6+c3zbOYSGeP
qJzRrDXLMMa6aD8nvv6KJ1ugl1q+DQuP/Bbb67Hd+x4mbMRXA0DJ28Fodg2jurxH
J/c+FpmK7MoJHwm2TkNwXOfao0iQYiY2eTRZeAdY6d0VyvN6sle5WJsneSdwWt/I
8muMxiXX+K5odDHcOV9SNEMBlihcC40BgoaxsYmkKsLnEz/R/dFKYYKMAIPRkv2X
qCFfatHuYcTFmWc5AwDntIWx6arlvDYLvMUqjtGncM0VXAND3x6xs9+d83rAUi+Y
Vj2j2LKbvV7a8azb9XrO1XH/c8eFFoGsTXjCEN066uwMCg+UAL26xBydBDhtqWai
71P0JJHjxb0Rk7gtAlD5l85AI+IVlasm7HB7zF0KHagTQYdMK73Jq0ErWwm54vW5
hLINKCLh+W5ZC1Ia9kqdqUuv5gRGW9kZS7V1Z0uf3VBzsSiny//rk9EMSNpL8UAU
wcq78mGTDKBay5hE7zaxaYpNL14tSNoojr3sh1O+aGwQqUAGQx2G5llYKYHOp6/A
LnwZHhDy8CHPQbEkeM8K7l5fQZr15EqyUZ3FCue9tZ8QVFBjkD7qdjA1qVN8A1x3
lPw7ji0rle9oU1nC53+X9zBsbkY6ig66/isMx39PNFOefiXz5pDX7qnmOncLR0Y3
z5+OsjtR3iojRUhqlq1R+vyYDBJGEyHBU6QLi7v2eobY/WVEImvLCU0fwRd4Fw4I
AY4VeQF3XUoakML+xvEfRPEVI7IywnfOiuMCvw5+Hd4Yfq2i1q46Nc9eI5M/vyj/
XneREfdiEtzyBXiPQlQizKIpObNPpJLo5fq4LGvDRgY0avJk+nMvoDG/Y7Fk7S3j
gzUem5Y219I1XdQQy/F2Lbcd4OcKUnVPspvn6+tLUW6Xu2Ovh/afPrn/b1pCu7T5
CDVqPpAg+1IRVa5ySkguZjVt2YJobT/fQ1YfdLwFjQ6ThK0+WS/csqDfJ+sb3T8e
Vz9bdeUoLTp/VOzWpwD6H3EzhSIHzASGf/cW8cCGR8vPbQyGJpT3fzP/5nf+Tvvr
IEDHyMV0KPwElkDRsF7v+7Inu8hspAPqjSWbsAsy0aEWd66JV1jO1jcyUljSDjw9
KkazBmHRPJeS6eBoaQAfIOnDO8J5VF26OWabQTPnUnVtoziz1Y6ExHbeh95EMya7
CLEt/TmPFM3zpDW16ORATmqecB/JPHrP1zzMdVodYdhJZgMpqiQc8GUFK+eJhwBP
e98gfVZ/uNBarGVIZrL2eymjrHzPtSISjz4cvxcII+moByYiaxhzS56SQr7xEzN9
BqT7O/YD0/fI0ENQueo++ud1f00JZiDIvhF3B8t/X4RTB8Nj9iJTnL5l8tjNGepo
NlV+tD8lec4y4Vx7daPB7gCITOMz9UTPdNr+XsHFY7RrWS/bDPLNCNKlwaiNYElM
WF1XI9nXQPiemiFRebJf2XkJBFFIAx0RICBGVuHp/kt7m3DYtDYD7UM/DB08Hhyx
zZ3C27Yin0IYqFMEQpL2sWc0CoLNcFwZWlSvhH+2A1o/KOm0Lo6scxBQfj5YbVa6
eCvveghNRSHjXn4tKnEhuxpym/W19/YuII5dp4giv8RqXckbnRbdzVmvR1kV9Hn+
ZhtfQFdAn5EtvEy6e4wKg9XpNZ71qUlRSPBcaF0RyD4mRvajf2iDjQ/FRI+OCp4D
Iyr/gfqRF3C1i0TwDhrvuqxKggOq4o3vEmAPRa6aTaDkGeDug0kHyZJXn8vP/Gn9
CIRt1FBTRgsqAuNsQLaGZEWwvRzCTZguPYdpY8s/iFLCQUepPqUaWp4Gzqx8uKZu
jumIscD0Np4EE1HTtcKA7DWDfr6coi9aC95u4SMeDc8wicVnN4O0hEFImdjJ3jyy
Rt/5fkTagCa3BhOYQamJJDOG9jHaFUoNPTy3OyIE1x3ob45cX4s8rgqyL7Zyb3Sk
o09GiO0svA1PH87utx6zdAjIyMI6mwt2MhrmRTKtXoYuaPgNVyIB3kZmG4eARn9y
nXhwoJ+GS9bifCtNuxCgmsHfI1+3ceN4OKV6bY6YD1MHGzNu6kHqBn9onAco9VWR
RO/pjTWmXXjHRr4TUgDbsCFdUPgRCeeTDUwB/ztbr80SgcYIeXcXPlQbAEZHCYtq
fEXlbprIsTOgdEc4cisK2x17rxXug1gXAWZp0zXvFvUvTs1tpbe6wAn2cTTCRP0L
uxwyvzs2QKiCot9WSdNmzdCl8RRYPgqC6IawGaidAaaG+DgsXk9Bfpxh5NhB49Mq
NGpYd7/7RGOI3VtjE363J5Wof4FrmvIpJ6GkXuHfCTaXpWVQwBr9SwiuSe0+dlM8
tmNqYNwnqvsDufbvffTGVdp0ex4+FVx9foik3zM7hhKxsam+9GaEWRWSFB2iN/et
BRvfrfZY27wgnpQYgXF0TC9Noofu3FqJ/5kbZF6AuAoRCGb9elb/wRTS67DDJgrl
UgN15y6Wo5RRmIPIH9mzl/1H44vkiWe2xpNBr3ivP9S/VOAFkPvaeonspTY+iJxR
ZwioshDy/QB4XuT8dN0z0GcOM4aQuBf192LeX3An3OmnEhqG+WSSKkIu1f2km+eN
mhdX2ZobpEAiEcfh9RauFglhmkW8GxMj+JQjXIUQC915GZD8Sh9x5SxM+NS+LlNg
kMnqLrVWbQlOQ45O4SDA4qiKLM9pPXFfzoYxx9uzETx9wqCKhPJbQmWXo9DypI+Q
yyfQQKrGYwZP0rqj2mOvjMAygeUVBD27UPlX3DGqxsXTHCF8kf9jf4SSBuSdC0yU
jeP+BISGJmQPXlaMPfA4J1Dh4kz6EQwrd0mmsOucpta8tAEwo/sXjpyxQTOb45uC
VErcl49B7E65vfUddv4zIOoMp6Y08jqszXVcdV+Dl7ZM/DKzNS1MDDmJUg+S6KIz
ft3251TjrAHENn0+u4ZgAtx6WozriC6qLPaxOVOja3s15fmiv8PdnGClT/xdTeD9
PhYgAVqW3kXoCYM5bgE65t2zfiyPOoUFJ6tQvN0fXZZyva+emyWJDlE+qtD/n/Vz
8pY63xU7Df+bc33ooefWWHRZzCz/eHcsSlOOwzdFKKgzRAcnhcvOh+bB/iCQudb+
eEcCxGqrXu2ftLe5D7rc3OUK4fBrc5mD5/WcqC8W+LaXrgekv/+3oz7ep6EaJjZL
hn1MVS8HQoGwBnyTXCXqBv3WfaU7KUmaiDWlHZs+3jBHLFRNoBi64SgU2AfTG6oT
At8I4p4qBvezU4aPFRubAjfh4AYUCoY9ht63sykvu+HDLMEsaeJ1b/sFDzn9UJCr
BdMol9+rAbUBZ4f70L7eOZQ+vgEFZHthT27ZXkNJ15+GeBuvchw+ZTtFkWMdCaPj
B8tpoPwlZ9awAatcDeIi9Ykgd7KWnjYgkrD13yirwjd2mEOu/+JhTE1foxZ9f6hW
CoMz1bFXeaeqLK/hcxJeV7OWJrQ+oW/YQUNW9gYdVJ+63is1ziJrpfFhu6ZCovVn
bNUCml+ZleJoiDOfasUX4mhbtn2ln2tcJpFptErB7ysazhMHWcyJwUBXfQX0GRiY
FQZbD/XZsXU2dlB6L6f2XH+61BCF/7GcJ3bGOyrTkXzNYwWBmJZQYWDaw8OyHpD2
VEgzKYTlIMOXedoCdetjEYVDwV8VpTY/e1wLhE5oH7z1DbFqJZiQ9+f43BqZedbo
uJBwqWzq4Tyz/ctECMCpNO2h5xna/HB7GJneDojpYqQgNIRHTMrSvOrl4OmTGF5k
72xp1iK2vnNFei3mJl9MkcMm/8D7oPnrrGX/LSZT8HokaFXOsjHWl0/UzLsvFkT/
xYsbvwadlvUwB4CNi/7C2BrNKmWDUJbwtMX6wIffHv6gz8LsRaSdfutCuPADMC1A
Oo9fqU67DHZD6qGUzLkk6L7yGhSn6nc42HDUoEFCBGBtdn7JEEwz1z3FDm1gvY1v
u813AVKuDcTPmJBOTrqC9s5Gdz4qQi6ujmbnCM26WjKACUnmef2XAUyYxES6clZr
BK4YLVEN9Tuz2ZUUQEk+f35XpSF4rD4eUmmj86/dUyi2Z9bTlQpOPZNqakHQOqia
AvrGuP+cRe5Q8jCySK8nOiDZ5axEU8QWHE9QWpaodvEpct0GsAmzZgp7BuC/ev5W
57OiJ9T5h27oKbijkob7zQJXBLBLuNUuhzPDlCeUo0IfKwAEQnl0u6iOssix17Il
5lx9fuAzDgs4lNuMawm1IIKqjJIyg9xkb1+PrFcRaZcviUTrKhZWva5z5TEV+AVA
sf2mjzLJQIgN8ATPp4g3Gv0IqPekSTqPVAy5L/Z83FedM5XclkYU7h3UI5MLzoHe
mf16iWfCWAlkS9e0mnxjmIL63XNus/tm+ice/OX+NEoywAyVNK5xRJ6cEWTPSLcD
hxT7XyXBnKVGvU350rHA+DqIBlB0hDaHZLOSD6vxH85cDKjiMoenVVNfobiDHxfU
aMnqC3N+BjOI442eQUZTcE2OPsgW3qWbZGa4Nc/s6VSlFI5w1R+6qp2G31HP1C0L
2VerzrV+nGALt5H9HmRO3/KhG5c0L1S9XVv6drvyuWCrLozeOh+qQASmEAvrkcNy
N88p32qFwryLtyQ591yd5t0BudHfwFZ/TetYcANyangLGpbJTxJpDL6n8hb0Q8IF
0lxWrvfowKaGl0cGey0cN3o86zQK+KUDG8Q/yxG27+k83Pigg9iw5lwVc70rDx8h
btpfNQrHxipMey99yFGCSUNLA3y4wbr+UNH8aihyk7YwYQfrPR4HDH58QgCJ7a37
oSQxWoKGq8O/9VsVGK5jvKhzFis9vLUgzzhGYaS6lacQMRv+cg6YnPsC8RoowFGZ
iyciAFTcZc1pJDEz7Z/Im8CNtnbncAJxjLVJObF6jOB8HH2jJ5ivg8XF2U7jR1I6
x2BQ0P1N3iY6MGo3MWJApnnlPJT5WBTWt1WFmexPounQjEHZQd4gDafij6tZARP5
YGc5D5SKwHdz5XMuTqlWOQNiyiQPTALJMO26VHgJa0o66gJTz2g/T+84rS+GPJmO
UJoVX7C6mm+FRuPiIC77T9qfiFY0z9SeM0SGh2iKO4qotZtVrA9EQOLUuv3Qfvxp
VEnMkDIfoQZ9d3OrH1a7zMJ/nIoPc5egT6DPnrlZb80B8KA/cV8OOLsxHasUPRPw
CqsGAA4SJNl1DUISP1/s6m/NtIPVmemGpCE0o85wJku7R+UDrvq6TOKdDfV/x+hw
DRquXSjbQ1hPZMGnoquC7d3X8eFYqF6NTh+n3koJMPe4Ubz81ZfR0WRPtamrWtxN
FDodJaqMBG+HBnWWYszjMe4SkJfgeGGilbNeUJ4x3kdbWW5vjqjOvZgg59L5NFtv
+DxITWrk9ceNU3LvSVGsCfs5Yg0y0YNhWZm0comUjxhfu7+wpKU424esfpWVBpI5
RC3XzMrBi4GHq8VZsStE+MmNWWTbddGFzGYgpYJ4lL3dmpyUL42ZUYEcF5GvswjB
VDF3l6veAE9WWtLyovAUBAyLhPbdRm+rAn7nycbego7BmP1CXzLV9Sq1igPdtMGJ
ji+NC05vhyUy6+kXRu07kwyparKSwlB275WWSZ8/KkX5etwo9AR253OAmrhaT9Jk
64l8Sv/MZ2UA+LuLNl8dqpvT/5GzGqi3X47VJcy+jM4z6pf1wB9mwawIfsQsOMfP
mvTeKZeZDe5HHwpysp5a3swJrmRk3AYPn930Bw7duAB9/4mWPWuUW3giuTW7fzup
D89K1vNCEm1/sAWxDrmbCK0OVwSSu/55rVc/da64Kbv6VtVcxnS2QIq3MfZONQky
0pG07q8FUyBPN3KeOPl1KJ2EgJr4ROlB0wKZ0ERuCVDOOsCYa5+Lq9RijICcnI28
mbvryqPeHZt7qORfWM8MMK3Rn2vckQ3yH0DxHgSDxU9CI9b4POeoQK8T4KZPBnxC
UvJOfxfLLDeygFlQG7VAhW610KWQQ2tKn28OD4J28p9r2+lshB2Nzn84uMOiPcmO
w0Jl7SxfGhWhA3NvCY/3L6I5eKBpEAvzpPZP2kMCbk4zzBFNF6J+HyGGsW/SQqh+
P1/TIHiq8F3v/Np6SMPiIsrat0iWriic2upErWOjNfcypYz3tCXChw8q7t/lZHF3
mtcRfDQdweHqOOaUX/k7b2/iW7nYC6iAj/4G+3GugSejZl4XzeMu9seV/f/twf7Z
rQDWxhhWil5QezTuC+sdyWPV/pYf7mAVpXIbRgLNCrws5GxJRxZuIyYNPXb9wCFl
UJxZkdnIKMU6YqcOg7gl6r/mVC3KtkRI+kwVs1QceZgFTTHWUeRcfdC7VEqCP5mJ
bYXVT4vmSnEoG3u0TBIgs0Dsf31oJHqesuPmClpu3NMlSompvfFPx4rzwqLFIT6r
JoPClCJiG8m5lVx3KFi5UztXa4VyMuDsghJa3yiPdiCHRY5U0xVVXrkLdr9QWSNk
Xqo/XTgMbReT5U2VMBNFg25woBkJWUHmup+Jo6mHxhM7W/VtdqvxCcNO6bHqqIxR
OfAx7Lq7Rt86ycdV+7BHJC7MHAt0abZkDpuH68BdX1hkGq6TzdPULTCZLfWaMoap
TQnpYCd9trXeMNnqP8CdEs8mG/0d2xG9+Av4ldAi8yfUjxClMnHdTNI/guxARLLr
0LhyBToCaJmmqB/itii0wZDcgMYgYRez1J4Xh97n2/j+KYinp6J1jolwLSJT6HX/
SYFEhjWb6qeqFDe56w/cNO2LYyZOV6YHS4poXGFTzshxx5elWDWoB6tXzZ8f2WrA
vq6pjiOqjzZu45+1uut46z5Suq18bHi5IeicRV3tIpDaE28hNoPy6NG9jwCVA8NH
o22gAvHPjc1C8m0Ve1q0qADm3QuLwHEqJBqf5Eg/z9R8oDAFcJIPEdpuAhp+I3ey
EypXMBKkx7afTnUzLcVlHgjLVl4YywHHmMDO3zLhz0KLsn1tbKqtnPFz9+rCg0Zq
LamJ13JAlIKxsGrvCleM8bytd7KFVQQqLaZCi5FMJOTpc0NnKRx2jivpcjGko97y
BkWaTGkBEdsLP3Wa3xBK8qEcZ3Ostk2McTbtKaWPMtUp9PnD2Ld/0TTAKX/yiN/7
5wiX287SXeJKbaCiJkkHy3lrUz58j1Prn5Ohm3qTTD9ORap9fWYpJOUwpc9RAAtH
ycl8igKlA4nxJxULXHBRt+4AhkJkbXXwQa5I4DhAGaVpAznABZNGmO1Dy9woycSg
VRCyQPh2KLDkDy48BWq9nKIEnZRqmAGRox7jh394n6wNOM4UzWJRK9WgOvkoklGL
D5SBQlUEh0ld98K8QnRibkX+Vo3hOBssTgBM9E9mI2zwngzn5WBJo1BbVnvMsxXu
VlD1/jH471eUczMp+R90GGyat1LfGDrsMz+5Qsiyz07Qqrjp/cEOsYhOs7DPbGs4
Ileg6uBTM88r1/GKGFNifoRdbWICXwbrwXvFySI1OorPcVxIWNi2A1QZU62CgPXv
fRcbYvXG669+WUIPgFo3R9LGLZOroWyukqUjUkUfW6CyCAkVTMfwRXzgWB6rAm6W
OzLvFTOP9lbyo6d8jlPCtPtLGOkie//Yx2fBcTzlOIkWn8iTzDodnJhzbRc2lm2h
KJRwrqPXNd/1iqcA9CkSHaaULnWcGHHZDCFBHVJnbrCh/3gRNnpkZa28sGqxDNOb
+0mdmPWPedUTojNhKsp5s0pAW3ljYpL/9bfnDCK7l1ki5M5nVyJl2jJBQ9mRfgNk
TFJ38zH0oiOSrUZ/vgiO0PnnzAAgHZRIMTfrhIbxjktbG2vLP6yfK/nanvowdg20
gtdrUUpZniRuoPyg+w8rgvWXb9SM6MQKU+ycVfy827xa3Sxl2S5zgI4NhFTpyHFE
BIoKm95MsdMbKjZS4CyCvYOPl/W5+NhtLorJBYOHmcMXuqrGQdMnFOv7eWFa99tH
ufG6kcoB6t7JqJj8wXIsYXmsZK0avsIn+7jZqATwydOEVBOiyV4p1H3OjQKdxMue
vgWwQH/ZPDR+dXjzf5kHXJnRDLPfEgqUV0DdyItxviYvMKk2goAQYvrXKjyJP9aA
3M2dEz0lLOMRiFyeR5OP95t7ChliOk3S4SoSTFdnMax5bKb+nJGM/jpG7wvcPoFk
bORkllfrxDUusWv2A7Ih9zVpLI0z/wMN7Go0CvoVLOIkRBFRFvsjl95lIjrzNDX1
+gxRyseY533cJvV0p/1rSQQnN45669weLzOrbwOBdYcYBzXkuxzrHj1wd6ZsnHtZ
QaYV0o61ZMDcKsQLMAnxtHiCjll3n5gKdbDKVqnb1F4nojz6xqAPnhxAx6J1irW/
yIZ395Tyhm2juP+EisiwKU+wSCwLmRbxOqyW2Qr3qHTJis0xFQN5MsWEicqZIMr7
/ty1/fNg2x+ZyORDvV3gg3fjeerPbcJT91PQ4xjTwVsRFUJU9o2NnuBHWcyKlkvC
0NiJmwJ5SOLt1xLz1GUvDaGsfwcWvj1LdvGRei6AHOCkaw7zy4OuZf/9r/tWgJdf
zzJZGkGghtAsJu8uhyy7MvoSSyt6KIimXurVfT2jJCxQeZt983LnLo3cJpSPbVMO
ngx2NMLoH8FimizyoEhJvliXmdkYhRLyIetinN99W1DcuCrT5ynhjhEItHXr613O
RL39NUyyzenTQCJsZb6cGKTigNc341+HDEew064CpNtaN9mwk8AFfFQtXwYOAuUE
ajjjRU/M79w8U3Gzy6VMKKYUtv7qTE0i+CdBoKomtQv/lo9lMlT6Va6sQvR5ImYC
SSsMZ0/2EV/gUYm8jZZXfT4++Rk1fTJMzfzZaLt2It0AaNzvnbvH9sSgbwsPH2dc
eRLmPWm537mzC98eyMc0zkjNm58nUh5kTZ0fZ6w/wVEOSOTeXMROLEj3jUFLwKv9
Anoqy5TNyZtF55wDuNsp/cgMWl5NXYiY6TaJTOcb1Uch8XIkb77SzOQi3zRpdb4r
yYmBeq7yuYI2x1RWNQBfrbZgWlWB+1+dpFxV61HbLxNy9rt9rKUJG8fovkdbmTRx
P5mpwpyUXGziPsxiPeH86TaD2crFrPNHHmxGCOpLTFPNTr/7wU+WptMgA0CZ0Hj5
g9pEhmCkJh9q9sEw0BKl0EpkE8/G8JOgdHvjNxbfQfcFELu27oRmbJboC79jgKCr
di99mRs8Dggp6vW+68H0D/9NuD0Cwx6WBKBqsDb+r1tj0EqfrfPD7NEog9fzfj4F
d4gaNSk4uZ8TpQ77rRTuI22aMeiAhEbMQq6xdrELWJqGmcBSuktgVIUoOwld1Fgy
vOhX/SCCEAE9Bx11eDqV3vsQ+bAXmjMwTZBT1hQWO5uJligtiu16gF9Ha2ns+qmu
GbGJytQWCGa3HEXKpvLgCxpbeCL/3nVOgmBZTzFPEDSXo6js3KCquBuxQzZpGRM2
K7+ZbcnXoCw/lGcMDejwzkSe9oEvlr+JZqVTHh1Bs5tm5tVU6LgY6dp6Ti5mhwiv
bnHxFLc9ZKHPKWd7LRiY9KYwoxW707jaJVAu/WJtVW2zGQHqBb6WU2psw1aY1x4B
LEXuoHlJRmBP6xoq8akjgpxo1hbKgYep1RBx6tnv4X/NiFyYwb2qKnuDA514gny0
Czibyxz4up5lW6fRvoulHw0fuAB+T53Q2/CMQnlZ5SQMntiUx44i1LJlRHUqKckB
ovRU3ClnhHc24b4rphaogArkEP5MERjvArJkvoyZZl+a85V4Xn5JvrOLkCIfaesQ
HT5+FOtAXni147jD7Elnnt+ShwKtj/wB2ebXTZw2jwhNxlDdlT1MVEC/RQ7WokXZ
TDPQjLS5OkMUtFI7H6Ehvo1zVE6xPB00d720J1JjVhFdNsKGoipftE0CSncbckEL
mFIrvNURg5rAbKEGatk7ad71NxNWvXbBSF5XhcGOgCZLG0n8lx1fOYIXpcn85pQm
tSvxJfSPy5dXZsLHE0zNGvNv160Hyn35DIWPj9MzJKY+AAB/Z9ybyDO/x+lGfAGG
LwKwWC+0oYovsZT6V7P/iZUAkX2HxMp6QOK2vlP810+TyPh752L7KzQ9UucSJYoR
vTaNSauwUpOkNhJFa4p/1Z26VPbMu2Oucc6UiE9FTcTW5w0v9KniU9WnbVllnDG6
qL8eBNpqbwA2mO1cq3IJGLnXNRvOYg1IvmMWKRCMy7iDh4tHpCA3ol8suKQcb44f
QXkND2HUzEPWLAKIlOa4LrC32giPCNKyGxiSuDQmH0pcsXMhBCA8EEkOZ31Ya+Qt
GSQuMevSNXNOFy/Cvr4Wr14AWqOFrwzHaNAYI0LB/Acy5gz8gOVxBoKgUkZK1NHl
kCFqeTJq+6d91Onvj6nW8EnSIwVtn0GXiELRHNKRsP0o8p7dEW3cnkYW3cJwUnCM
g8f7AZHG3zLI1Ld6+3JBSKZCNvGyF3nplFsLPtq5Nn4FpL31sHdlLooOtl/Vxsok
adHp1em4aR21ZUxmy2X488vMuFynRYcKtS6hCerUgyD+vrK5TmReYR3OM+YWnzEJ
aKVt8aYexdNW03Hc4gr1HZS1q9t7zlc5atMO70uZl7caZ/udC6OZkKqsB7Dqhkm5
X4KSYJvp3x4G6O5ygri9aC3fix8A/GP9l9BG+jidNWC6mVRQKgvNUK9KVlYOtsZO
Z+N8/SUKgITkGMZ6M6NVjDxzaKqsI1ouFoF2uPbpue6jsZIvWopWuoRjza2Www70
Xjr1TLsCTM0qooXclbCMe44vHil+/xWX1mivF3WaJG/KGlnggVUSG6vbXbPReIXY
YAMNC/6/lO6Zp373aC+1fgBp6hCNmymJ/7Vrjy6oQP7EKcJQCvhxCrmOy5qpN+pV
6RFRPYdbHhwjAiYNRcc9DCKk0BNEYFBIxpRPjxR6VxsW4cmqVFMmHnIeK7gar0Pi
islFepCeo7RLS7i+N4YlyYUMA0Lp/vfNZIe7dGGpEka3W4NTeRGGoUWy9DzG86CQ
SReXFzXPOesZEBGpwpb8OKl+w7OmPpz7EgYRpW/4z0S1TPRwN9xe8VI4Kz843FRb
B58wwehFhf972KqdIQx0ueO8roWA1p+vBz+CqfEkWLZ5SfFoo0vj/tY4ATdx6s5k
nkSVdVVlP1ejphr/ckiwtCm3Qo6G2aLZxgpgq9FMkBP6uGF6wDQXeModEAEzyzfE
IQs3q7/Lb+f+v+PIMgeBWYx379fs58TIp6pvLtdg9LEjjI1VBrb+BS5q7cHeqAxO
oB4Pjq00T6Bh4LQb6EL+X/yL9euFapy95JXAkfvtROYTDo9Nv00aOjCd+2rhUO2b
H9IVO4YgSIi4Cr2LjERH9c5Lw4PU9eyNpGBUCgXobGs56xr5tpmzq5W+Io51iHRz
XcvjVJ6e9DzhYn+WM+nnPLGH7tRSxMpWw11+CR3Bnhxi0l64wZgq+6zJExct0XYV
WBdY4YruvcevXtwcDeL67sPC/AcWQjfHX7il+CvgnNag+z9k/65hdfMH5WOwTeBy
1KhfhBvnnftAC3yk8w9j8zjFo+Cv8pu83ZkbEVDbJ71ZNpComm09GF6RG5+xqxhK
SmBf3ksforbt0Uio2tcIH16h2kNvhXH30MtSHOxdKAYkTnNlo2YE+XjZQfD4zl2n
VPybeHMv8U/3m+BmwsMQmo2lwRn82PewEakE/xECropc/KAZ9JRxchKz/U/4gVGa
JaCAeB9dAfpTM9IzK5Fw+TBMfyMGB248S5ztfewsr2KeYfve148lrLrfnS6a+vRH
oEOZyrivJjNpqHj+G/LI3ISQu/f6Yf/enToXGf1bDHFE1zzABjw+mxwnv3YtE393
8toA2vqvcS2aNRLzeBguqxxn8NNoDYuH/dmTHX14mkJoY6vAsUXX83B5Sdqfg1au
1aBOS4o9meMC//DgULy7VvjNKrk4GuCk+S684av54ozG+Hyqc1hNR7bpRg8U6b4m
cyy90LhCc1ja+4XZoF8jG0yBLcublOQd3M2/DxzhjitRCGkCzbXSxFv770t6ZiZj
/8Ou2QPh3wO/9DjP4Hc5V7jBqwXNQegvlCIdYxBkgmZwpHvFY3PXU+M+M7w40KYa
Wn7UI7n9oWpOsMLxdwJoQOky4Ufr8V8biaLuPFyplFYgFjVlbgj1hEZsBkqPejMw
D6GePLvXua6abrrn3JX++sMRA05VzNJxptB71ABy/CiYq5I1LbBPln1PqtWfYrEd
g7eZ+iTdjUyvq55tWL3iRvCVZHLgQSEx61mSyXIsD4wJV1zvi0fQ8nasWCnifTgt
NoHbq6WM7pBv65GuZY32V4WTjknFjZg/waMoAT9mnVi5/g1Cz6WSQrEN9hg4Ziqi
/STF8jmtGsBTRLljLIVe/2ikKJtmo1zTReMdaCNZfEUU3t4+opzLxGOyazso8XQh
WsGRTvfbuxn3VSn0lC8jgQuU7IirF1DqfXtgjSq7ww4AsO5UM02obEnL+4HJCLmf
7TsL41pDXn6LVvAgtYLPokrchYGY0TfPZPPJp4U8Gg/ReVI0buvr7Fo37C9LR47Y
ppPaXYBHfZbxOFV/ZrPvlRszRZhhg4WOWjtw6pbLOHIfqNTgHCIz7GXp/Zwe3Y8L
Wr578bLrTV/xuVOT0rcPXGvj5HnG/z9OHRsWxAd9Hh4n2J8r8ymtRjhwIpkmi7L0
Kmt0ougmoKeRpGkYXN2pPbvO5lcsQ1eCfLjRgxBpqPzjDcUBC6un1TQs1WHboHXY
uDH2V5SEYjVdjXc4rHzC2O7gLOvpgkMP80bUcrAiT9kEhlp1dzhLTLkPG633QODU
OH/rOHI+fd3C5MRW7ttbZNqpLlzKVPDe38+BHEE9IdEg2ojja6PDyapyb3jm+QFO
KmO+PJhyuqukSHGlzSyFUuGRxuItPfmkLE9ufpZWZsS4BSlx+bayH2tR5zwflmWa
xQ8TJXWZKnG0/RsvrKzOQJoSXCj+ZgvrpnZ6tBqWWKAQMOIoQAcs/lChyGI6gyTo
E2rVGBqh4kS/5NyNWQpK84UrTToy+rNNwvzFgSoNEjOmwMPPphyeldY3egwkvKIE
g7F1FIegdr99sUXCFo/N8xRdGyrmDVc76T1c8RDeUxr+Crjmsz3V9S30oEpBozgT
2oOb7/auHKrZFpgN2RIuQASyhB46pPynp17NniKLV3QNdsYR8AH/fAtviCZFmj7d
pWeCrwLzehnJv95g7a3xpyllGXPKP53RWLkBSXCxNgSOdy0Hqo8S2St9Ysaf/K6p
tTiSCC6Hon3JWlXpMbVC3gVGaqEcYjrjF+PLf9nGN2xh2i1EyB4yJaJUvicsoH1u
aA4FEKWKHS+rX+OTbyG3Y4xzCVqjaFRmU/1dliVkEoOkde/uehm89gDkrYnrRZiB
bQtgGCVA3N+rtkn/6IAo3e6neVBqvUVZR/VEftKgHCu4a4XSymY2SlErO74zr2LX
9s2Tu6+D6xWQIMex5dKhXuCEY2/XxyVL7DwaoIxp8zgmns8Z6NZUKNO+9IZCPZTC
SZmIG+hHuNOH64Bm/OKG30opcAgKTFo90dzxbLVGXNh0cFtHNraSECHd2rBm8nSY
yP3Pxq75IM2QXzIGKQcq+g1P1Ej25e7RpquM2UD0EEHuugVSJkxpHrRcrke//JUl
GZnSX+XooNYa2/sdKWGYSX30RdvATyC1yWGiBaYvxDzbx/rCJ0LpZuoE+sc4o4uc
XiUY52KnXlN7w+ES+lBIgCfFNmNWszQVouqItRQTJ8zji5yG4Agv1R6DhLLGL5V3
Au9czpKvMxpfZMxZ5hMivrr073hfmCszW8EoKV2fSGiCkG+7umQ8PC5feb7e3ols
b2pWGOyAdrogmS9cNBkhAA==
`protect END_PROTECTED
