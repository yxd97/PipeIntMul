`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZwGGDlL8hqyHQeU/PoK9RdFgw1RvC3+gelOtSrHM0CUacgfZnFS4/3iZHkaepdQ/
S5rZm3xibnFisCSpRfzx2ZvmTWfbGvAynMKF3M4e6vJ+qZ60bqJQtMLtACNPyhDl
3rNDUONBN2Wibtv4Y132aBrmO2Y/OSP+wKpMeekfcOCVitLZDY/xdhUIEjsl4Ks2
wzVJkFkjEWjIW9EXVIgBpLT4z5cW4ebYAeJn7ZnJHD/SnQj77QXb4+6vx1yqSRjc
Y1+fnptc1N3BRX1crOdZBy4NAVNXMYcDVsZAk5d6EVxe3OqyfeXmXaLjE2Fu5zp7
BordT4LXNJXhKRV+VTdm2KLisxRauI/1UK4t1OCDOGFzwo5fyAeXo6D1dIeSHIIJ
IO4nlFMBoTF/6KnFwVhHDA==
`protect END_PROTECTED
