`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EPJseuTNs/5FoCyFHKJHCepAf6by3rmdKXay0oAHYTat/EwXkBpPEdeTLERSvul8
w4J3QfHSAkbmancFqUE2FAoZAAKN5bO9Vf+WH0LRj4barrtkykkc5MP0cBZHW4nU
e9nKn/VdnqgCrljrGxjbsihonxH4GWl0jQ3wHKmQW1goZ4VN55zvWhZi9I76OsMo
yTinREjaqE0jXbnM/+jEVlNma725tz8QJ4f4FwB8/BfV3o+EKyiwuf1ekaIxRUVd
HpUL60HiX/CRrGTn39jhkrDOK0khSKLWzRZSTwOSp0z4/ypVxjuB10Migcg5vuZx
G+vL8kSA7Bt/gfyJTv4gvPXwOEfkuH6Udu9dcgPQ85OucfNQ1acvr6iwPqscTmcy
KRBsQZsGjW9jwE8md2JtiOfXJYxU5thY4NS2atHPdrnTxZxMBTei2IRY61IVGQZt
10IeoegShv/TPj7Bm6FA8SMHDfdzWi/ZV9BHwp9kAaOsPpKRxk1aLraRHPM1i9tz
WhrsC9uwrqZZq+hXVucVR0WFo7+ASnODlK1azJKm1Yocb1rBfBjSyvvbDHWHQEEl
LQhcZHHOiLAVmrcSe32dAS1zPBjqHZNLXUuy5CyrnlL18uZTRiHsTsdhEED9Ebhi
pBNsC4W9Q0M2S4UshiWqAw==
`protect END_PROTECTED
