`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wWO7dwJdpXE3sj9/Ad6rVRjnvFSqQfh/q/Gry3fYdZaK5M9RA08zhc9E5Zab1Rti
VV1A+eblHtMuF3tVKiaB6snvl0sz0jw8flgjejzqzV1xYr8saPttasddQlJLPGKn
DVQBLIY7MBJ2Sw3JUUKRBCbKt97o+dp6/Gxd7l9X+GcviXJmk7iXVTZRs/2VuyaX
hq6SzPYasYkim9cACSxFuBhzcNpGStAYk8sQkaKFnOLqHBXCBcAzKhUOihDF7Gj2
LRFrV3qw5Iqsq1mpU+YNtKaJpkoNxhO5tofwh+L9QgEYpm0bkEdqgKU9EP9YPd+v
4ovGuOMpwPyB6M1rNUfsPEc4Oy07TKkTdBFS0S4dGkKSWyeCdachkvkLNGKaD+9j
4hhvkzIhUafXh/OpVmuK+wgJeliYadLlU4TJTCqEwiughG1l4Czh2ucUePaZ5Fr1
QPRiOlhPT8j8uMVVO30VDv1+55eP9tSAtFEePDfS7PdB4L4nslZDFEEDsqwXKar/
1BypxM99gDlCkO5aOwV6EMAinJmcDjNo0xbap7hF04zq29GJkfd5V3fIrIRoO4OM
H6iA59GeCfe+eFMnuZNuQLzoA1lFcSyJmUj0HHxlJMjnKubM3kWRMzHdxq9VaN2u
hv09B4AIO9yivQ6ZVpcM01DbjEEt8HvuXe8QuSbHwxHAZwLpw+Fx91But/bEVuFi
5HHggFcnysa2gQH1plNRK27IT6cK6G+/+Tfs7lMs9BSHBDJIsqUqMkAQZbzJPsQN
GiTe4VJIbhaU+wEw0iFQAtC/PIj8IYpRCOmv40wiMkgK6MUG7UkdSo/qYRx8vIfY
J16jWRoCSRtE93Tafdm+AwVilD0n6qgorGWmCelQHSXL7DCwzlNksnqW6m0vwVvY
rjyjeGn/LdDvMXHDgjWhDai5PFqDAdlS0CIYtx8OA0IWYYTGb/V1C/y/Xc1Attb+
ohTfglzJ+KmhfC9OCwFw9AuiM2D8pv9RetPVYb87Xoihubj35W2Vyfq5FQwvVZ1e
Y2OvK/mKNLwhWUEbZN8d2S2lxymU0YAWhLtmCfseqO2APV0IU+L7bZqiL0IIq0dL
DfxSSWQE1gzyV4oO3AiwAgjJ+oE8oOK2IapuqATsnwqU6+weKhzce4uxZVhCAsp6
esYYJN4sA9OTey1WiMWw6nJnd4K6Ejarma7XqjNGuCKEaEME8GwINLVpp607Z7qI
cd9IaHd9ClqNy3GtYghZjEaLSeb5DUoK2GdVTekYeQ6gJfJ3LMVVR4W3XajjwFtu
kp7Jc1ljpEwpl9QxxBKeoYFZNBOXGRgtmtF24o7EYUe4H1PsWn0mFdo7ETQrgCi4
3JBFsxBOoepGTQsM4eUtMgUwAwEs8Ev/+iG4KuTrlWvsnZf6hogNGjWJ3TGUSd8q
B/rMf/7UJtbYrsWS/0Ym4izXSX+Jru1fiq6YI3R48xLT9Bzqp9VTNYu3pR0t9Tnz
8deaRv3+wT8Ue5NWn6UrdpOLzDQdYrPtv+tqq8lW+LENXq/mojhGLb5m+NRp+XcM
VTEqWX8HLFK6YDsgPYl4p4NK5qzL0Mf5Bl/xrWPlqLarM/tYxZDXoAv179ql/nZp
XpJnK1r7J8N4+R7TCcTCxn4AkUOUt1VlFh/hZ/ZCHteQ+gK0BDWTS/LMbzVCmXkD
6aQj6GA9NtfZraZNQzLZvimEPKwczaSD8zzgi4aXvheqNZ1UBbrKkZZpm2KQI286
6EFPAgj2wVHbiI8aBM4WnWAFYmDBio2AoB98QHNi3l0e1hcvu9nFE5mbACXFZeSi
b2nKqYdmcjS9o+j2/Idtb94TS4cQ7pcrxYP097a90MPnJv0QeFuCy+kDducjG2jO
bmCui5G7fqMPxhkjFf6iYrBy937u6cX9xdirsdz5MBe1bqA8IciCD9t99vhOD8pl
grPQ6SRFuqSVwRy8ECmMVIQXMy4NaJwt/5kYKhhojVkDEiNOA0RZhqQEUfuAU5vz
0XAZVMQAKqHIH8xLKwKkI0dUOL/oIOjDgkHDA7K34PdYVYmxYmx9moJdmkA/UOaV
TGnowrQ8VTjeZJK4W9WfMEyPWoKUinG/pLsLX6M6rUyIHxFhwKKs6NIDiGOoOn2U
y3PX+C6nVIuvNx8rDw+So9RuO+jHpIwO8TLmMBJ+owkVsFRxRR4aedgN23OXFfhm
hUTgqJN5b91+hhkpzF4cXyYZpAGzEu5Jy1Q0B02GGHdQtj/5zEsnbyj/JNCqTqVq
WB+/iffE1v68RQk4TbRRF/MgfOT2fGaSmFaYrmu8YZz1bG8O2QVa7/fyPW34cl6r
CDBT8gTjP7Y2MwrRR9S/uUHgWiMFfpoziEOk1gGgu2qP2rBWjvyd1XgtjRvTKxJK
GCCjvvKy7sip0MFZSyn/Xu+8VlT98iAF6PCxcgIlxEeBqZ+esCxlWEe5PNoSqYUe
d5NPbqPKVi20SXYgpWUZwMg/his4Jv4pwTJVhZj98LIC9EP5/0UzmDiQFysxt+/B
J0HvpL59UNuW5VpbW4sVVxYWop8znY6MYIX6p/504aCYsmz07dldyNkJRVdDepkz
Brt2bkmfI4LIxes9SqMsGPzMHTVToYoeCs4QhiJdDURYhKpHdNqdMXfFbIyQlhIg
dMrhoaS6ebDDo8IucCb7Vg4MMoAJFNk0VKpmdDLZ91kK1KUOuueGl0dW7oUVB2mc
FDiC8QKWpdWuAgy4ZhAD74wOrCAmUWaeuHWfNVupEaAbCPWhI106dSPE5b3qxV7g
kV3KzBEqugv9Ry/y7JuREsH6zjSFPEYUwkLYqgWJP9ZGR2UN73Xxuv0YBd6HC5oN
zAtjR7rSgJ9VfRoQJRz2FvVe3jfN2tr6YWR410SDWt4StSEA3wwjR30AEnzK2WCE
M0Cy2u/O3yB5X8LXh5wXmyTWirSM+Uw/ra3kUkD2MhdApkdll4I9QpLp9t/+Z+dS
ab7Ia4O+Nk7/u2antsQzpomU9TAeyEL4gwXeVyZQt4JbnJrH040/aC3fkHl58nuP
nC6/a8ks5ALB9GsFXi6a7XyZAjn7wZJFWtXRHz5xFqKwUcQdLZFnYGFDlngx0jZH
q398ZPvTMCKGxI+Ico4qpcuPGOUwIps4O+hO6uqbOlzEOOFZJq5/H4f4DWhgXWtc
KWPQrE1fUX1ONl94RD7fs3xsJgb5j/ZCcIdjpnylw7MTX4BYq43Icon29RU039Nj
6BjR8AZd1Cwh0d0bfK4xDfqlzeAkoF7jTc5dxb4NLJW379eUMki/fKnyXyyRWHsu
q9+RAeuEEpqUuuQA7aT/QjNBasEjrTVQ46u9xxg3b+TXGHMbJGZfYM9pgS+yYdFd
5AxmnZGyLELzm1j68CTZpsw90IAF8R7fFlcvmd0+0i26Q8hXciMgSEcdKm2w2EPr
vYpIv0ViiAUDUiDyggfdt244NWmxKAVhv/CpuMXwGKSFitOLxP3h7crKcj9ueAnb
/TZXPFUJ1gDshHcrrBlPR0w2efPzgCI9CFtBlE0iOhUDDZ+1Fa2j8yhUBOuU6mPD
AeKQLHpD7fLboz6TO11QlC205t51GD15erLoL4d8C5ZHML1jDBkVHT6TFv9oUqaC
gOu5gDpYIrlncp0A/91zl3GeAx5mljxI0a4bdUN+LLz3JT4Z2wBFW5Y52oRYz6ZB
DURFXHjsr3kW/rcViK5ALyxAr5muZ6ZaZP14/CfOWOMLso1K4li4VZ+rNaawsTZd
K7xZbIozQLYK7vQEYIpmc6xW0WGY4iv+26C7pMkyzMKQb4Rgbgzg8m8ZPvTaZj62
8DtopSiaVJk/ZO6S5eYEB0GZQmRg6NunzfwUpjYKVv3wLkMuiVUFkbMipfQH2N9e
IgR1MGKt9PlfSNvoQkSdgO1JUX0fjVoVsGgGJ6mQ0BRBwuUIsEEKjrn90TbT45i6
wbquTqso7xxT/pnLrlvo4bZkkO3QdKu9HAk/5VcRS691tVUziwdKbY1T6IVgcVc1
GSq4WkzCZwlnOrotCx8CiObe03cbg4ec97a+IrQ0V/FWmgnh+JXQXRPNkoq6qAG7
CClUB6bh/0kUbhcVJ7EllJfVTN+us6j/ckfZCt33laQhM2kpSu1InzST/udPz1lA
lg2CAkhLMj0KzO9F+Xg/98Yg3gFP2X90eiadPG5uABiTwk3/7UxjMf7P4DG2byvh
eob13IXipZq1KLRtdBliRy4o4Es7+YWsysKCO7IqHdw3TmEmaJxdch/i5YsxV5CZ
2Oj1NcQMZaDqpfsC6olTSMcsaObwfF4bRtWO/3mAX9O9/xToaxRUYhgAgToZWOUc
YOwElRApEISWTAeUfviXA3N5Fe2dhnjX+8hgTiSq60iaQip6fIx4XaIG4EuQGEBN
g3ZWN1G8iDTmuC5lIR6XWTmsM81GpB/tI2LWl4YQPSRcHZrIaQUGGvOkjFAlvXyh
YBMoXY9skwULiyFkm3m00MZlzooLXqQpbdpGLI8eTbwpYACG3srVUCSl+aLIT4DH
hSMgUISAjrM3uQlESTycKWxcCyFCcZbPUCWTFGi3Q/BmxG2wAmtqoiFW5sD0EmD1
ptEvYzlyb4eoNbrqIUDVvmSL8vYN9cmcs+yAzh/WFpsbet5pOnqshfKcD5Uw89Xu
FBN7RQkt9d9QTiW+HuREZd/sar0hgUN+o35bBB+0rtk6xCZo+GEBrUg3/IK/mA5N
5J7VnDqq2ECEYm46Xf5iO7AK0Pc6dwiF/hB+4mqktMu2Eh+bcvs+fKws3QAP6I7H
r92/g2WZ/qEcj6BSZ3iNANK7H47d674Ndqf6fcpGI5xS+Wxklny0/InR5jkXMmgS
ez3VAEILKStb66x+kg8anDb5wjlrgMZS9FlrgpF+0XPyXjK1+M17UZHIXyP4DGiY
N7grlsCnV6Z8Trgkr1yFrdtnVQhQM8nNfVsa+lzq0mIeX+AIxxXWhvQkwdN3KoLB
wGbKLuOCatLii5H4kliGlKnjzCha+og8MlmwgjDotoSpNZvK/dpdDv5wFxozMt4u
Ymp+fub41OChfQjZ6jDHuc0/7CIdy+VJipPslofaI/Fz6DF7t98+wUhFMoZFcOfw
I9/p8pBIUelNih1CDGWuOQ==
`protect END_PROTECTED
