`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cEbFHi0msdov4QoJiuhpIpSBjAysK3tlVY+SaNSTRpRqKoAvWFQcoqLUqHDsEAZ6
zJ0AiIlsZn5dz3zR3uf6VeOjJWzVw4im30LcaNGWtdJVa5oX238i3mKS3uh2196c
7eIrup0zljbsT8G+DQgSVfMG0SOHoft5ONO30ENGvyCjQxkJiZYlbdfTM0Txmxzy
IFDOGnDQyybH9Nm/5gfgtWFNQEJr2zBnevRSSJB3LJk/UHVTAqbkwvZIjrGKKYyK
0iFNVc5tsDYeh/ZPB8W+MxZmwQYTsi0k7OpOhxoicPwkNRYwZfqq0csD+3EyEQI+
ySbaFGrhzS5CiAV7+MnvYkgw2DPsQVF1RguMcs9UxOZZGHJ1U+skj5khMt08303N
g/icFL7JjCoGQbvYHy8QQhJBE6Ad0holRVeNk2+YMhINFYBAgXT9SJwKAjaHq455
1IMQUy9Q9noLzcGbSHQnHAQUR6pVDIAC5zIyY/4/p1nsY6qIjkJoxTeEHzxuF+XU
SyhJQZtj4vY2BzOFD18v+Kgs4EgF+6/R8+3oSeldAf5smncVcg2iCxDbjiGCIeXw
B/z1pxuxyk9+vWbVUKyQIB2M/93fXja9XiCGUZR6sn5DRs4tpNSTFTXKrQ6Hj2I7
DCQWIxkyx168fL3s8/iJct6ydXdQiT+mrbEoGAg70EEFG0HT4Es2qxXkyyY9w74x
8eLDgtQaJZetyNZyjOOuQh0XFTsKsZEGlvHmy4q2qNKw8mhj7Z4bfHkfffIN7naY
NW1PuPDsUcF8GlGeFBmd8A==
`protect END_PROTECTED
