`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rE/Se1foWOMscuJxDRDEdRfW5RVxARlsDDyzAT9W5QF1b9gW94GaLbyt+0zBkmbh
druh5dLDvDZWePFukYVL5d3as512ARs604qseKO2u5s5F9mH8e9xOyhMzVa5RNDD
KsA59xVCRoh5FwWL9xRoHDHZ1ACimAW+k5On6vOY+Un+doXzX6tr2y4Tqnl3JTqq
IzL3jbguAF9QJziqH3+iCB208ma7xXsG4Mn5HheqeDyXLOOevHE4+e1KTM4IuizD
wgzaqbFm/lFXibBmh16Tre60jn3gQLxGyPM/tDI+s/sna55gum/pIvogctIii1BL
nZkczS81EbkrMF5B+6KZDHF62HzZeohJy50Aos77oaxUkBdx3iQMmKAE4ULXK6uD
r0psV2lk8YXtPg7i9feaMYuAe2bwSOEZOnX6cMGmydNaBVzjhfsst7sq7OBlTrOp
Qfo7Me3LDVbao/GECqjPRrQJGpfEeGpozNhZUOuzSjcwrUCQgAEKKVLv3R8T2YYl
F0aWLI+bX0h+eeOAT9C3ufCXsi5NSbSSakZQAdCvHa4dy3tRtIHugPTElvF1Mko4
G+aqYbW1ZaqWVnjYiaaimpr2JCDxUM9jKeDEQU/D5N8hdbMb76R4Kj1HEWgVCzQY
qIUP8o0qYVNhLpdWexlNxIqgCi+ba4Q2Klaj1K9tCwN7ro93HQBrTfniaqOLtnpa
pzbBJEWUBcKPqas+rVTN9FnaF2eh1if78QLDv152ncRNNi3QVU3g6cTyoAo4SO7U
D85C3aFVTKAtfOgF73vUkfTR614j+dorsg9Jjn3nKXkovA/ZxK7juxsfkzCCC4Ue
D5QhNbFL77ON475vAB41ve8TSGb7HE64gAUPkw52edNrpbpYSLLoGXpfrbUrhmCw
BoXef7AxHqWmcZECXSItiOjaLcPdJF/lr7Nay52LxRE96wopSW7GLr8j5eCBzyVJ
WYJnr9UnJBkr0fCQ6XszfuNnXS3HRWLC5+utVnWig+ipuSLWoc0VYN7CpLIe5Ff3
ZyYutsoFbT036NSU3N0IjF4pKYgfN9ekow9Qt3PfpWN4uYA5Qs7LexX6moR7t5DM
lNUx1PTldR+B2mQcRT1Zt+nle/WAfixjKRlEGWHrE26SgMerSHJBe4qywsoxNMJQ
KFqTA8xWPGtxhe3v5PhSCn/u6HOAVSsnjG4DxFD20AEtX3PS4ldAO/VgCcvr26Gc
JHDa9bIeDX9shtj6lld6wuF3k68tiuTJIOL8os6uUVQ+GvRTduy8bYgyAQyId98X
P+jYLt6O3H6Z4vaxs8PqCEIxgGA1DP+6d19jQQcoFr1bQ2Bkm1w2vFFGINxX55FI
C6RHEuvxwDHHZ4l1IMDJr4dD0/cUTsDGct1iBH2lKeH188q6Bm1MHSfx2u65XIYm
kmlxoZw9lvSX+cfQrC6Pq2aRQaVI8qaJ4R+BdpUTgiZFcxiOrpKhH1GTQMG77hL1
9GtI6XcdJWGp1FdXamaIwXTIJSC9kI8PaOT2wT9DigsOz2k2AWXGuKnWS0ysauCh
zisGfWmcL+AW0h4QTPnJXBLTVD8tXPdgDVl9lXJLpMFJqxiAuT34kxECLgh97rPr
AJoBUPx/UsuVSXVltoz4RrUS5BpMKUuxtT3+57Bs/+VK9rlA+iSl8kMzkJxqUZWB
tQIcW8v/+793j4v834Dw7Z0NQnai5J/kn8O+8qkS+zp9Oxwf85U3BtcForBT9w+h
FDiw4y2ozSo77wrD9A7G6RC4CCDS4T2EgIpmpSboWwHoedWogYPYJmlLsFBuXp50
UlYDXReqAVlt8megHNNopiTG9fu0b5f4I2PbEtgUDQ7AnpCdnSi0HLBgGThd4oxq
GdVIHML4xh/uuKkO20E/g8+8CECxW7aIMFJOs+zvpOV2hjNT2V+Oy4eX5c1UCrVY
aaGJNeDbkS07uT6lehojqbvh+ljp2xoGBNVKpCqtEpwCEwa/n1bRfqyIRBlRzuaX
NTjpJyx0/JG1IiFSfhMFASLrTU8M3zx05fGtgXmFX768L63dALh3MFj2dw5YnZCC
pkgt6g4vW2igs32rxBWEb+q7L+E4h0o74fG67NVnEQcY9BXwxTGxl+pqIoMZlMbq
7m3pXj0wLAR483uhl7SigSL5dvw0NiX4sGBqN+yBR0N94tL5lX9ySFdGQh+ObNCs
WbQdAUrLXV9NSyM7tKAcsFJJGikr/auOLFyAOEO9+71HAjaAMnkFoyVbCb0XJYbh
yRwFtAjHMt+s2ILE3AUu/ewq3jBvHWzkupbuEGmVH6BeAPAEmIRADXohM16Ryj4z
KO/H+OpAGay34u7v/05kXHgW+YVC/q4n6UsyqbfDHD+hJU/sBhupGFxOxRY3QuHW
aCyJGn3pypNkzO7a27jQyzUs3vfvvBM6C4VqSYOt936txNWQwoMohSnO3cPW7/p9
z2RIORAQVACQMlb2QjIIEGJQeivDwau4s/O2FZs3Utb2uuf8MwL+pCaOfOrr3Wa/
w7UvEw61uZkbTFOzT3xZmK8sK2QkgylRkPolmWY5q3nnYJHmy2szZzHZQLcJ/K1v
JSaquTuXSj3k6Xtd77RXOZ1WyUdkXRHYrGHj/QWzFIKUIYGopmO+pUepif+hCs+Z
C7TsH2ixFrzP89cOUyxesOVZiWl2889B2Vdgfqpv+5/dmyFKJ+i83cpkJPUT9dU8
6oTe9q/91F2zcUcA9svexxlYcbQMuvjX2fs7sCxw4wYzPN8STljdP4YhXHUhZa/i
eHCZTy/5N+84Cao8BW7wTw4jjCrRYqL5kVD61tlvRgVeFBPtsC6Bk50O6ArreWGt
PYRHkCysdkPzy2OSzzbIGbB4xwIybwBcD/EBQL26Wfk6E5w94KnD720D/3fJVMuz
3IuPuMCB6FmrgW+s3BTePmDqe1k7bRYTpXvcB8zkizRUkL91E+quOqC/TRlF4MjR
kmWHPojnOXS3NoFJj4EG47sVjtRowoH61JREQwthM24MlORevlY3ZE4FCcQ6cBeM
0YDmLI4woHw3MPatvTIPGkVLb98kBNWE0r/AZOzb6Tv6fmK0a08rojA+KaT/2feI
FIcKDRrop8Tc+0/i8bq/GW8/D2L9Ro5d9EXmC7AjTZWd1oMIROnYtHV0DwdpYi0j
3oK/ZmQ0uCjnAJ+HdyK2kdt7FD356d+xqvcH0ALQicq+c/9edEHBQ3tDs1U+Q6d/
yYi9bOGi4LyF1/2WNj2kDfkrrK2atTGtbsjEdlgokVFhYoatmsmzLt3BbcWunaLT
5Ka35bdyYSqjHblMyCv6LONia9wKI5pqdfML5hl6jbu9e2/oXToY9PjIEURfsAVV
ShfyHBcNNKCQbRYjV/dt3b3APeiHjvIL3wA7yyrYVnr0/m56ni3+tqNvsIlkFTLG
+qpn9C2TrF4EnGoSZw+zuyloDOWzD/M3Y1hcoaxCD2NfTH5OZFQi/CX4/9lbsBrU
NgTpadpBEEIGCyMqGndauKRuKDYopewGAXBTthLoXSu42XmPLzITkb7nSqNeCMZV
a7cwciouqG5k2UxPQXpRp/FJK7gkPNKY8n/q2Sy1N1+JLmYqCcALNQRq2zQTbJaa
5XdWt3Di8XCRz26wFUbv6TPcIXN6oHWu347QvSgPCBLWja81sh9DtjtOcpjg9njS
nOpR1+SZFhmspH7szUKutHrDvD26Nxn3xGxd9w4YSI7foCBzvKIbo33Gb4S+KSm+
OBGnpzfNg6doOQD+T/5F5UvDCxgnFXGgBrcuKcatLdkgSzmv/wsiUJvhnFYD9x3O
XdAyF/tygfSfB/5wMasKvwMn2fzmbQHZZcB53MifN30ObiKg3tGnsiqkRntL5VkY
glADzp+NOcGyCVx9VJ2s+lcw3RIEAZiYVhEo7o8jcROwFUn/YQvHQD7bnKcmFOsY
PgAnhCdIaProjUVZZgb21omr/QOgIWY4D+xUhx2WGaADFjxR8g1NycVu0iPVxIBM
tLXQEs+MeRoawz5K38/qQVc1eES1psOd61eJq+fw1Ux61AvEr0rbehaw/i+6wUHu
Slfi3cN67dAHl97CgUtnJEw57VUP200cepzDNm8dcekW0E0A5lhWMtLlkK/4IRQ4
HsNaA8v+Xvx1dO4GuiXOLs7PsT2WNwZLp06XyOojH01og4zD7bov12B6SElKFbW2
0s6GbPZL5DZizaEpSfC2MzK2HCYBb2NM1caVp7/Uv91bplfA4rAN3VqHQ7NX6Jk3
3DmnTrxUXgdBvkaqOz/6ER2M8h1H7oBHy7JJsJZTD33J14G8Gk+LbE/IaZGvgKme
EapxTcZtXsCaA5NF9Sd6sYPwIog9FODUnBgbu9tQicERMKxereXxS9A+UWEq+coE
N51iKkMo1qy3Y4vL4cl2gY3AIMBkPEWClLL3DKb5+mAnIttfss6cLNR5CK9koKYg
DA/woAb4guBHuQ7BQ2hzEs0DkrX8FTKIkk3eRwJ+60JzGmy4dnJmpLNgg+BGau5q
bViZgi8R9XaDdZ4EMaUi1QwLUNDGsA4bVE9t2KFxGoX2CEyLqCQXopd5TtStND7N
YpveKvFeLlmca1aN0kbu5sV99ffzHYyF5K12QtqmljozoxmwUL+OoLiWcPR75z43
Qhv+yeAovpZObg3vX0kh1OopDR7yEmsx0nyRfQ5XkUSPGfB0Kn3SrdzzmQt3XNqx
NCkdnBTscqTK4ZCPVvMVYFkHVa4HjRaBT5+sYAxWwzDPyQB6rgAvRbeaHd9L5tWz
y/STFV//ceYtQpq1i2uR5g9TYFOhSkh3I+qLoQviNje/ht+kfrZNRgfJuo1jLWS0
8sDvVgfANhWQpsZy7eAVwg==
`protect END_PROTECTED
