`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7O8J339tE0Rvk0taKZi3pblyey9PgOoE+cQIp1bsQRSVXkACtiZZbWQD9CSAUa6H
60AcrbGwmHOnYE2bK8+/liTSnp1QBSB98anoCRWcw/Jd4Q2r/mzvqlZtA7VwEjcf
aUumoLfrxnDbd7QnoKpzHLwU7nWKSDyztPzfY/OBLVFw1StPdHO4byWN3+OJx8ts
ZvO+S1p+QPDvvvLJmgkSd6RxTRKP9bYLfgI4ncRQ1p7YZQHABQoW8AtVNmYMoNTZ
PBoxe9+9AejEvydz6b3LjuclmlhRdEvNYZQLcT+I8RHGwR6RIV4Lj87eiQqRIIkX
t81sYGVPvbi0g+OLuqA0ABKGcyzWFxXZPNKu9GuOzbvpUZzzVNA1nRS60GbHFzWZ
jb4GdGNOV8nRj4xYadXqPQCgl+o2inyAPrFz57p8Tt5L4VEVL6ZD/QzmPQIQHcU+
vL+tLJQoUIG3qyExyJo327n1Joc8N3+iUWjrmW6B+WKXiL7JGGdFrB2fQkr8HUJp
D/y6Xw4E8+kcwq/WVE9vX7UTNwjXwlp818urIFCOareywLrOcprCtEafj12Y9uYV
E4UlYtpsuEYlk+DHMUVquk4M0FIPVpHdWamzMLceBXxXRabY/UIphNy5qGjdrBwZ
FEj9wQLvp51z2ApemCdFQIfKPhHiyUXnP0RPYdwatK7vnKbMwZwz/DKWay8IOAPE
nZcYPl8LifoaeWP485xYa2nKXEZNweSuwLznfH8Oe1g=
`protect END_PROTECTED
