`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aXZ1ihsCxJnjOnhgYbONNLMwzRsAcho3rifSD7GehI7Kt6EhDV9+eN5BtJ6E8q4/
i3CefHS5GkRsdGo/SombTLuZ+MhtnRCs4cGq/IoasES5IcaftPrH8JNjAXiGPeVy
AS90xs/PYHyQQg5TOdSfGD/ov5mt3ZN706PhG+6o8m/RZ5RyP9dXgWQ180dHVIUc
mVaTSpbsPZ94T0GlsumDidN3LcNcTGwTwWDCqK3P/IcLPDZz06YovPZYMyi5I6+i
3Cgj+CyTrmMPaMK9/IOp5o4Z/p5mQcxGruiIfMimhSWiuhRsG3qHWEZFXqj8j6Nc
ENxLNnafTVOFYPOA4IXl8NOxc8jKuK31SkzYuZEnTmZzLTozhZxMxdctJo9uiO6u
lUU3zmVx8waFjqGMNc4bL2hO74CxR54qEpzH1Y8cRE8D45eOrmvY8soaTj9wYf47
FrZq4IIl+/c+1MxgDMMTXTdYYazD3lSKbJQrTpRfuuiDLq4Abve+u+xxW27X/+Hg
kUWWHyfmztIJdp1QS6RHtSISyHyQyFLFxTK2pNYYEeNqlvrpyrBkeCkZx+Hf2LSm
nnheWWiyPKWwtuixQEnWkvi0tVZ1loGbKLUrTip2xrnS1fwXS0dhBMikDVl4iq3+
XDo4b5G6d2ibBLjwf81YgsvAa/R6DZQrkbilCFxjsHqz5LkUlA3+e+Gdk63G/U3+
2PpHVMHVe8sygZZur5Q+HYdZLg2hbauPjbx3jJbHoHgWNSCb527PyPblWmGz9wsx
vBk7MEI6nBEOY3ibh9Czg+MBP9uB9ZlP0WetX2CLkSMBeVZ/SZ/tpDCA/3Yx7On0
QHWC5HCB7e/fe9BAgkqYrbRYWpkl7pYVWkZ5PVTxtzssWo0Oh7KztzBlaBcZ0a/e
LgOPoqoo35fb3ABywUgAIEJ9hlZOz5OtKguQ6WtdnSnbXMDalL4yRnjbCMvUrBAg
yujgcH21h5P5vaVTF333IOJmpOb6eyxm7koA/EZ2Wd1Rr7C5t1VqRO6+KqeZj+5r
egbPMAJglDgkXH5impk8yqltVBIEBeuOuc73MW1e8Hqii/y5hb2vGysNyqMIahAo
H+0KzwwU+gd1LEklhHQMiIq7xZcGGDkM7GIBWQV3CCbiI6iFI0bhgew034C1z3NB
VHqmwVA+bBK2ZGZEi3eMWzllSAjvNGvFmsIGozALAHZff1XbivUAUE/lB36RoAB3
xMcrvfVJseQ1A+4gwoVNDwaHr86RYr8zWiPmOphK43p5hktZib5E7zDIPzG+aujS
oR0qs5mHVcFo8DcBtoXqPbDUt6p7j/B4rJVpvfYTdi4=
`protect END_PROTECTED
