`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+w9Mb/MpyGlYT85AocFkNa+saml3/ysTsYYEXnj1wUnivMFYaCqUN98QLlRcpRl
JyUIIPUp5xH8BCtFwu1YVccpxBnw0Pxo9I9SHTfnXpwgZ9EZEeTtkfCvpl3ulGDG
PKSOKE8OFdIIWTnBnajATSHHRhbHhPeYZa3Syl/WWkUjIY0YO1iT83HYnMCedI4R
DOXXKVTVxMssaQDg/1LVM/PHR4FJ/i29wTwBo2+xf7gtE+Hzik63rpDuT5KSWCi5
xND0wFli6qEQUVgArTWTcLmSOdoN2VhoMRXLeEFK+nFdaU5a/O+pWuvhqRfTTFp3
oqPU5BCVNJYQYW5q+QVNe2SvQkneBdSbT0SlEq/rIMaBpxomPVBZItOrOJTxbcho
ECO5Zny+I5WCRTdKI3sBum3M1KbwXHdgmXCzaIgQn760tU+s4KAuYLqHOeNTdxJE
rm3KStOdB1Z29nhmWduRW7egnYtdd1dKGGIx2XV7OtqV55v3RuGk244Y034YY2JV
TJje9hXAZ3DrGGFPuKXnXx+oApYtoZKQ6uMD5Gz0QNL3gpnXbEyqlVWHMFvZlpjG
7UbU+zjJAJcquvJ11yr6r/2NiFP5ENOT6hngJDz+yF3qrqHBVeL8F0TEZi8ntxJU
tWz2bKTiLCZNfVTOme9orKufjxJoZNkl+aqnDO7tWf5VE1vKTGKhd0dZEsvmexnu
tzglUALSSSTER7FKryQnLIVio6/r9ij15KSIYmsKNxSyE30QRGHLGauigMYQ0N4j
l++9KmI2khVZCzdYKOrmphAte7XrgdfWJ4VHrL84qOnIKUJgwm7BCeumXOD4iBQ3
Quzyr25QgNj6rVjAPU05qNeROLUlFnHRFz8w7nyeyo9r9uLnUfXu3jyZyueM9d3B
AvbcLRklxBZ1cy2mB6ZRwUT1PdNUVhwR18cfV6/1niStDuMmJJCF4AaB+RiGSwKv
yFLlpnPiGX6AK2edQ0xwyYEo/ISNwdyBgyLJM1AOZX4dqVDssrAnfc7DuKQNJLh1
VNUuif+RRMiapcbDRYh9gQ==
`protect END_PROTECTED
