`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJT3PHgsla4pcfayMSdW1EfQUXTOiuNWwCMdJdKLWreEwg3kXlR23CLaTpUWA9q5
vwQzEFDsetFLybAGlUjRafCYPVSC0ay3EuvQscFoHQi5Eig9k/FWEt5Z+keU2xm4
cXDelaljXBqa6JrS8RHIsxCnvN/Eg5RZpWSp7p/worDBPGqtj3p7IKqDT2NztALo
cG8LMLu5v38clKstmWBNJjbYlA6f7PE3BRQjYlzvJ5E8FMnBnoNXIwTVVbT9TXes
d/mamRDw5N1AvbV466Wd7cP1Kr4ynbWh+V4M5hcoVty27OrdXSHKUZrE5vL8Y0GP
b/X6Pur9+UXlBhyTIX3qc4L1nY+oAS4m47Ly8dTxRCqfdJVF6jn2api/1iJYjZDs
D/lopYNcv7TADZmBz8GKzlfM+Pz7wYn/wUrtyIrzmomNmWhm6dVy3FdyobIAQvwm
fVaLMny/wrr8R5+fUpC3oQqVLeM+aK5rz0ns91WVR/kPcSjpovq2c3PpBxTOzHdC
Sx8tPyvSq3c+iseLgAtpQMs+2B5wqM7XVOF+lJt+y1P7C11SNS2eU7qJv4UsxKnJ
Awd0zo6WHliSUfzxDPG3oH5lnvyhppDFIa1UABldU5Y=
`protect END_PROTECTED
