`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NiDGjOVLxPtX79wSsGEQZ3CccaZEOO540MEEACR69JHZHSs9RDoBuP4w1g5zbYBV
neiGnlEOhHFkVJiqNroMdYJOB98/3tdpKWe3dEhaCc2oLMcljcThGrLq2gF037zG
6fyje2pDh6FWa4ich9TXWCQ3Pd1cp0GeS0rSyuSS6d9o3Y3Q5LxhRrrjw+SdIr7O
Ry6ph+hyc9ZtFzG+qTx5TnUSl2FpHKTZw1CxXWIxpuFtY9MapiXUfukbxjE4gvoX
GGVN3CKOEuDu24JKPwq1GcOtNeyYnSoVhTJaBKvZD6fMn2oA0A028p1uhGmSHYSv
L+QAA84jTSCodQHfsv0/ypn8rNaYlufo+nXmqNYAbQfxHV48CmWSLiGKSzBTVLHV
6IqX5HFqPbSisvsO/Jz8Sw==
`protect END_PROTECTED
