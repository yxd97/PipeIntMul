`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0ukwjMvari+9yTjdqOsJFbC7Jw2dWu3ozqK2G/0qAL9odivDMhGdZuQkuLnhn4x
c0g4Dulo+M+lwwrh8aEvhersrM/ZyDPSgqlm6LyABplkTSacCNTHj/OrFuDvw3f8
tAem3q8zqj05NITLHRxeLPjGfYyGpGjHIobqes1ZlWTlxwAkZPs3At539uFjADB9
4ATfa7/sS6oP5HP1zSUo0IR0sR/gZzcHTYFBPx9GNQJ9V3I5HpJhO8xI5xWsR9MG
KC9YjG4L6vYFtBJ3Ic0gMYS3f9DzBRBKEM3MozLBvfasUNddre28O9oL4g5IDq2Y
rJ1SJ4p0BOEwKcarsqc3psps+De+irKjf1433c71/DO3HssuGUv1j2oF1h46GJsB
9co4UUPEs3oCeUejrFIfTnj05d/WMS6Q5seeGLaA1L8=
`protect END_PROTECTED
