`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YpG2LljiYvkg1oVUspQqKyztPWVzuI/YFixab9CIGV6HEvvEAHc41o6qG4vK2Esb
xilVXTYGkTpMmQ8FVVD0uBeeeE3/x8+G8dhq8FQQcnzhaC2m0pVhmJJfaM4drQuV
9ZxhR+Ed/Y6Sl4SAgH5NGEUg8ixTcje1rOfFCV+0QUa4fdOj/UOWNEeFGzJQON2R
oRBcDng14IjhK2A4zbU02+p22aipksGenCymjo5zeXSr4T8+1+m71jODUo1UAPG2
NmCXV/tFJ59gw2lTRBBRBtVpqznN/tholrgmN7NLCbY=
`protect END_PROTECTED
