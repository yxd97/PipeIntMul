`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V2W0jKdn0puwVn9ajuRjSz0UBXxNj1nkTJT7Enbd44EPgEvq+xbZmGTqxRQKZZh/
L8PCgWu27LkkJcaEvxjpQjdKBDhOroPANJVLwDdtzQt1j/I8m+498whmAioGcaAp
u+Q6CONnwRUo2l/qB3/T5EKRHlO+RwWa7D/3jLeDwNgSexCb4RcmzjPJQd8wRIEg
ByIxUz5fU4IQ4dRYjv1uF3dMpjLXoavhiJf/IPCO92/dzLbuAuKRbhVMmBBPBZXt
pJXZFXQxosiPIvUplQRpt/mtU3g+IigEVcq3WQfASCCXpK8lWNJIu05TonFJhvAp
GbcTYBB0oz9aeWWg7EpwvgMxQ9suPcXhyK0FlU/8fg8L606JX2569EldA924st0A
jwbZkhJgmt4ve0sssDRFAKZnNH+59fYktxYFICkXscknRk5PIOJXzNZWMD0sQiEJ
pqNkWWnyR2/CITraSjv/oJWDQAF+3NXRdqMoq67p9Xuz+k+nUYYwkjS0h1SMk2/Z
2rIrbNUUqGJTOMQklOvdROH8Zra5t0Vk2D26JNDxu04ZYoXlkT1G3p58A+7UDU2r
`protect END_PROTECTED
