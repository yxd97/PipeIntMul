`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5sgl2V9e1IRLWn/d+wn+13m22urCKqifHBew+Vvdrs4HTJpH1VhkDF64Y+/rAyG+
3Qj7mTuuyfZTKCyMK3Id6MtM0uiXNfpAQ7BK7SSsgWZ4/9Cf/3MUmpCPSzcFr5q1
U+cppIz4gyIB8FtaNUDFdl8U7BvUohh+JPmRuM6v5fCskuAtjbMkJPYibVEKZyog
tOPugFhwGiLkMFEpDNW9NMzDFTlhEaiy/xNHjhZoxlQh5VKLCrPC3ZiOYuH2+re7
7O0bDFllOLKhHYM+dTB1GVlTtSZ5SxHgpEmJI/ANT1n5mVlbiMHRIsS1HZ50MZYP
SllT4UXPHQOo92igiVmc6DNWkXt0X75VEzgGr+cGr/7OWVdjGtxKCLSptg3ClMQJ
V7q6lA0abAof5+Mgl7YwM+649Ln4oZNCORHN4o7U5wC5GalZraN25QjpDJljlzNk
`protect END_PROTECTED
