`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1M7xiHOlWD+Q93ORD/pigQAhENTqZ0Nf1A5EkA4GPD+5viuth3y0cZY6BKSDfP8
0Edx9XVEhIgPh4QfQIZSTTFTHEappTbuJKDjBgjYWShreXapQ2yNFHnrRXBKugAX
ink5V6cmacD5Vp2fotpdcIBiliGlaBW5COJX7Hp5+SiLnKkvNXZTBqkv9d9kQeWy
JoONsa+cZy11B5xpygqsmOD7KD2qMX2yaTc3rQN3L9yA4z8foB81JU5UP3Ra6bpT
uBA+luvZxo0f8JQgtkZQ/boMxg240Z127m+j5OklzUyvmk7YoU7x7TPWx7d3xUxL
Oh3VQVeIBH1jLYkfyEk5ZyWAYZHO+L9luvIpZiCWLvl31Z743FLDlHHS4jzSpKLk
3Y3JI8hwvaBGdw/sd5a/ie6zEiGonnjLaqZwqjwCUu/UMl92JNNhSsxc0pSoVJwl
A0GVXHZoBLTgh+OLOvLHgs0d+H1ZMYS2V+eau5dNM94WZEk+bsLbCKxHRu75AGDF
/mnddyUPwBDYRNSbC9zSWHzxGOpdyUEMcpCIdfq3V5vEi4D14UuWvVyUqyAbGIk+
PM7kIEBQ/UqJDpBd/ijsIIOvxbDEOM9GXnkVOqcK+NFT5V/2Z2Ca58UxXu7R+Lii
LLY5IChHOSKqsEnximpTTu8eaR31JcUHZIirVjfWNP/ui3xUYkRQK0ygt4lxYP3b
bQsRGbu2eNZfb8BxlLOEjpSNOkWRWp4Vxiy8eI3RzQqzlAPTOT8KagW7JoNrXc2i
O+zh0eVyhCZxgI95K+8Uee6ve30T4aWgh5FfSt7sCMvnpg2GKlqbuYVT9fOTjGTD
88KTRI6g2jLavv3AZoeeNA0RhU8sOo7p59SEfrgA35Qou/2ZOPEBAER0gUU477eu
E9LQGjqQxk6WLApxy1on4W5OUZCHCweSG1VnsjspcYf5T8iByMlbrEF9cxNj6/8/
HzimgSUo5kP7TiLf2j8d42oIcCPfDNqH8PSyjTe+8dRr0eCx1Ot3mJEK4c2ZO1F6
6qHF/jmBKGMyN6PdPBapauimn18Ft8POduYS5Q7d9IrV9mL2qA4KEKPKKBvNbmCL
9apeqBpPvR/eFBkPEgbx+eal2rtzHmdrNGk+GZzHMsAUVYujfZlWxT9f8xNiKATI
wm+pN/3EzqKZ+XH92pJ87vWUQbjyIh7RZipp6weTqCxNDM8kOWL7D09mOFqu7Rwz
HoDnFWBLB28YX1NqVIGWplayb+aVsad/t8uA13V0mH/zY7C1vThV3OfcOuqwFmt1
TwGYMgum6ttVtcLM9sc4DXpsGVDQHUiYRTc7wzDsKSOgYoUyoIq39mEIKweXR+Fk
DG1lKlhIwtEFbarsnt/50thFdA1VXhpZTipRYC7IvFUoruOVA3SjqSPRzkQipDRU
qqDY/KsklgqRfrXgfwi/NWaunJvTUEMgKgG0zzx89LmuK0TdArFcfCsxsQr5+U9V
98hW2nS0sSvD4TjlJTJWkvvyUWaWrt19UTsDC0+Jz+9NjjiwHv7HwBXz/Iyqv4+Z
kCaK79pFZvOYOPmVLZivrKPlJHIYpH8/odABFbgtrIrFH9qaLd7P3nfYxQ6Ya883
RZgaSVjsTkntjii2QOx5e6vNey3Ls5tCavtOobjiMZ60UWWFU0xOv9BkQdtGU3ir
ur9CQ9rgj8mBhyRY40KXPc/P/CoH1S54D1Sn2QQ8ukHuhRuCzNbJFonDZVnl7Gtr
auQCgJ2WV4ys4vps0Hmbky6RWRljamPcjoABHlsiXbKPL3kW9QjRCNYlvCfLjIuj
drd8NkjruPVP57xtwSJGrXP8QtKVUqG3yVetvR/tkSSfSR2EqQj2pP3uDgjLokH2
PFOHkZL6f4ShaFR4Ipjw4zXdHBYJkWmB2JCXZb6krXYPxbtQezJMG9iN2QtzwgdS
MkSF3eOuaH1bje7u9Eg2jpnp+FuhdiTQc7NCDIJnguav3Yy5R14nPU43KkzEXb90
6PwmAkT0rgDu7ZqSu7+cHivCmi9//6LmOBKGAJ8hxkYEgKoXq4XP+NRR9TGsipuk
2l0TZkZeYO8gtNLIShNLU3TiPj5dDUlMNCrRKsvpwrC8hAztLK/hnfbBOeA9J6+n
9ZSZbY8/N+HaoMkvwtVdYNE0yHNg9rE6DY0F/00hxrxTGpC/RRaemEE4Cv7LBT+s
e09jECX556bPge3q9RtAIRyFAKBEaFxdzt9urgS0xVJ65QrehjBjaBe2BaeYMfzU
JIjXWzBcPw3KALA0ZGbIXe1sLwalewQ4w6VqT0dhHMsbh65NwqJ7oC4DCVJiDp7q
h3j/BTIlFNBY3EfZVli9Mm0vIwGEh4apANpJAqwpipUWzI0RkSdOgc2s+1h4/g2F
5JqPs7dMBiDd2TdxmvYydYHBjMBE4A6hwKQYrYpnbbPCbGTQpIwQESbpEXI8q38s
xkSX1NqAe40GFl+vtfBngFkRdl3v+7boDr9woIwRMJTCQWzvvcBwC5CKenP0eD8T
CI1/GchlBEJe8o88QuLeJSZxla7nOkzuDOBji90I022iqsDpWnO2bS2oFny8pq2U
M0VE/O7Z2SF92wbgABpETmp3UZJPj3IOKUyILOn6kbubV953Ss/x5Mq28wlN/t8c
NoxPXl+P0wCv9ec+dJNj5Fztk9PDk25RSDGM5qFLGZwm75daAHf0eGm1uvFpHMdo
6BimigsvJhQ+72/blIflZqeCNBEw14cjOCMN16ddexGhH3wvhXwkSAMdX10D5ZWk
/HWG21eB3BNY0lpIem/NYVWi2PmsEW2/9DhvTvF/0BvpuATJDi2p2B3kmhl0OjSf
dz6CaTldvFLx6mv+QYTNtq9m11cazpIurb7J17K2mtR+Wzu7g2yy6fNE1pmaADhp
O6bv3UFsmfR97JNl4+N5Ii3Ux7rIV0/EE5zGRHdiA1dYVbDSMvrMUNy53WDVgL0g
BrCJ/g56b0GtANoWYTkeXQwXhP+cqTugLhii6uugGnBAjBn9CwvwePItHP2L6X9P
xIr93rRatpoWKtsTVAyn6m8g5wd3ScPZ2d37jpXSj9TKqYkx7kZLGJGv2HWI5rlm
92RHvePydTGpl3yUJvwcvpSXtpIR6ECANiZsKGnoJ3QD4xkclm1eFkf/ZCyk2W0h
iVR6do0uLxM43VbgGiLJvErRpE5PFmH4maXT28n/N+bim6dLJgAdZ58RjeKy0olj
Aw4LhpGudEcYYDVac4C1v7LHmeqG8eKzqHOCu0YjbWux2yTUrqHOk9lPzTV61c82
PuDSnQKJPQsYNoTiMk1/KfeBex6cOD3rr0hwPQXE41Cu6ricC2VWW0U/IWUnEqr/
Ojn8SAHOAUnxVoKwZ8ewn4h0rVy8jdpzW3j9FT2lp7k7tKkRzwNyj/kaeaD94o4a
TO4MckH/Ocn2BVIl7Bt1mwRasgEvDuaAO8WYStBoBB+fQMa+ro4nyxFfiVWRLKhw
CDtqdYROz6h+pH8s/HzLYQJCwP2RW5FARKiDRzg/1p0Mk4aARN+D8Eu9GCq7/b9R
4eOEXEgFhcRWWpQ6BVwPlL1gYx2cmJq9pmfAOvnmnHZNwvohLQjosDbyl9AMniPZ
mWjp8tucstHCcRQIr5a+RbJnxos1RRMf0T7qm6ytxDkfop2C0Ee0ipdgGOrdSfkR
rnlEL6mPEgas+fSLmlYM9KEKUjoiCYDdNECJe0ZsN2fGgR32XNSBjGJ4sWCEprrE
e04wXlYsNDDPQzacD5Dts4RSvGBiQG3/SRYyN2/iQBt+5m2Y9110RboXgGpbbrWi
t1+aOGGF6vnAKXIDuXdSbEF3xacibJeaZFktnO7OsZT9AbIx1Z0ysl7PIYYTimDi
ZShVGLMYWCfJLBJIjXNVxl5UJfQ1X03ZNH+fYO16QkeitjvVbU91j69rRdmsb5r/
NpCzOJsJojx0R9H2mAI7lCAfYeud+nNh5LXwpRBTNQBd6h4cf3fm546Yuz/J/gd3
cLuv1nTe61M4U9lALi0WZogT9c6O6PFX0pLgL1E/nj2o38+U5oWzqui1iLH2i17r
1R8Pnuf1vt5jH4+B/ig2aoauUZYqd7uKO/dJz6cAtQfyOHl9xCKBgG6cdNsAL9IM
1Bxf4hkBX+Zi4v0IrOyYwliiHAAOEMClqzQYRahXx0UJ1E+SNYyenZb+xB0QHefu
XKVQtrl63zeTn6g1BONVdHLemh0OMzWBdfwiA+2b5qMBHv3+/HJovGIipmhWqCRY
qfxXZpwbD9A0EeGAUNSfQ3bZ0cs7V+PcSiO3R8CLnia9YVzH/vmuyzLh+mfrXykq
XxXi07jRiYxANeK5JQpv+dMZWwVgpyxtafOlp59EA7Zh2BQRqLthJRgNp3Y7yD1f
fKtAX+zYRVhpsYAqqXabtH8M5usgflpdNEDZxm3aHZ1G38AYsN0FjyzUtiMhKQQy
bRx/3F3U3CKWNwp7UmtTYcOdq8zF6wbaYcNEFzaczCHpCBbhoOnJgiEsrvzD75DH
9w+aafvqdTZBhh57P9D7JnhTUawHuNf2rw/bxzq3ejVQL6MiF1hXz6mJnJPDNqiy
qBfMwGlnw2Hc9BW9rH6t90ks4+OEMz92EOu2qh21AFnyuU+5gGGd3Q75KKyYTE0G
9MSpKS1V6cRmPYuCZY8OpPgn7PM/+jxwY9jq75D/vJc4ep96bgPNFhx9uJcF+fW0
pmEz/fd/ys1gTKlJ+s02AiBMNGSzMBdgazklTJXvgrzeF5SRhgazLCq/F2fL02aV
JHOYFWhjlz4MVbA79iJzLHg9IggUzp0oBmlu8JKnqo5qg/8zp4/CZVSuVHV3JbBS
Zz99seW6/WNVy0wfcObK/7PFRGaLvRkaAGTfF1Ey5jn+UDTkF4iZKSni9g6Y2Ka3
h/TaB1eaMpMcbS6jI4319UDF8dERxTljsb8wetKSlaGB7vkP8co5At1DCugDOx/u
pqIBIoMtV3uMKee6DQPSzzG1TNvlYL/bl/uAAZlkpa7j1NUfS6qW1BEtlcTVLWi6
j0MYENnJLZL7GRKsUQ8doFl0tYN1UhjTypV8zxxoDL86e0guF5+SHXitvEXe/gEp
iyjEvLX+A9KBnN8ArGbx76z5s+3zK28LLAGH7NZKYu+2L8TIPrnQYov8OJesU0pg
SgS8IPGVHsKyt21SNzjIBcGSznfACbRcw5sqRxd5O3519nCmGQHZe+3CK1PZjnGp
9ogQ/trK4zfjTEAny4dOWFmsMq+d9n3i6oBSMGhtA/XTzlHEe/B3ZDV7hFuZB5sF
uMXpQH5aoPQKiSfQ9h6tG2ypzNOW0mhLx7NZ98ENKY6tkIfi/Mfn7jkhPODiJy7o
4ype80TnqLbrBUaLt2srND2lN6k48peAzb50PdIdlH4Zy+WcW2gqPogtwahjLuLj
DivSXgxjiMJD8QB7BcReOtfiiOS2Ay2lvczDX7588YKJ0NtXrbCd4O1Kbi6rRopI
IfCanVUdjuFOZWATzm4OoMnaxM+pA9jWmIKFsbHjKCphoZ0cQt4i+AjkI0GJZJtF
ejFlEws1GXbCKVoArCmnTJ3YgW679xDurdw56Ph5h4likSYL9r+Qcxd2QYWUnC1p
3vitxsCjqkuNrVv3UZ5aRtfp9n13Oz4chKcD5nisp7UiNCfxxzJO8XvwsTV2H986
eBgXIy0JbpXsji7CCp5/lNUqa2rZg7Q0zRPIaL10cpmF4+PsoVcJUr7muLbezGvZ
eJK14ku1uIDYbV3ojt0JiwshVoxpOHcR0xpQ8h4KHVGxcG0bLMNFHo/U+iX4wFwW
wvIGd0M3Yc6v/Rqj4DyjILb+dI9KxEU8j4o/tGddv5fHoZyr23kUwdiKmOgpit3f
rfoCA0wARLMPOZB1V++4vfvalxfln1qFSpAOA2WuRXF3ctBGEu6ebwxOIFc5ezQ3
mfkSAaEoO0MARo0dFfesvV/fdkYJt/FWbyQIL2pYREYWPVA5fkPM1gCwHcYVM5o9
SUxUsBDBLSmauuSdvisFXv61BIn+YbLjoP8C90n0jr7DXM+9EDHMzUPwdRXziSE2
hLwx6LJRjUmXFd5c4nhmWM12fb7SHJa0R398tk4JlmMT4zXp+QIT33gn/EAfmU2W
XilJ3XKCQIPyOD1C7PoTDIj1Z7nl5FxoLnrAt93SrizHzHGq1KSZuRuyCQTUNrFd
LX1yXuJgHMWtErbYqFMagvHkIsx47mrhJ6c+DJGoPiXWPIa+wwOgSS3unPWQ1Bce
6Mo7tJv9YtzKfWnBmuEuCxzeh2Pr+IC53xUvJdB0l84Cfb+QkUWAwwoO65m7Ta7m
VTGtQKnE4HNCQ1d4qqK37YkVPKXguzQvcyJLj/HyQnHg0dW3Vwky29+/rcxDjcwC
6umD+L4hr2Ydvd+RHm6tW6w2/tioE4PnnlIYvy0ST/3jPKGiOoUhtUqgQgrJ4ffR
fdsSZS/mvvXDwflAay0w0h/Px3wcq098RZjy3mLnA52MgnlqYRxRxgld0mYvuAII
gNwR/wZrRti+QYKMwfPwInGk45Kp86VeD2jQquwmlrD8NqPupchnZhlcG5RSWJUL
7gaFvoIxTvO88BfsVLvcP3nHh1sVbJOawWdijOb8EI2hrguhHE4XhYln9ia2hy7c
ImzD++ysV0yWmdFfu1zvYifxCwoal0Wys4sdsUKSsZ2oW2Tbk58e+4B3hhC0aTHf
N6pbv+Yr50UTXlXZ0KKMo3fVhq9cKFRLEEYQ6Cm5HygMFkPiVjVWWmyhZ3A+TEX3
4pALmtx21rwPZMv+l/0S5gllP1PauigN1rLHej9saOYSdFFphXH8weRiuUr139DP
Nz4EAt+vXxhC49oECxPmG1VW4OmceXI1PTZsYolsVcrZNdUZ90XV4X4ph55CwIg/
2HOcwu6g+C5c0Q1R6p99PLy8IbP7X6v7R+Vxxllh5gWw7Qvv23IGlhyXDVbratYE
bPl0+agDWmNSJeqoIgHtosdUS167hWluiJk9/r+42wbr4w1E4Um/lH7UZvT1Lgw4
5otTu1DSplJz3nO7ITo77mKF4DBj1Q6eu5D2Q2k2CuFZ9m2sO/ZsYKc1q4KSEQ5y
XppQ8lYtFeyRNwOkcpiRuFqV7DJW1erKTJHBPm9Mm8MX4gaMBokblnYWRUkWHE+K
kO1mjGEBJsFh20KOMmSmao92LlSaWGDe+RwK8i2oTGS21NV/yZ7YD5A7xR67qZZm
2rx6HJdo+r3/7oJaEL5lFQaImj4mA9oGE7fIthOxlGa0QAaMx9HmzALc2b+ke9Jd
isRJxzRbnsBt+Ybs6BykT/AFzyzTQIfD/4/3M8NKo2HxBpp15GDtiAUz/EcoJPjp
56S56glIkudjn9HWp/bg5NzyaZUyh7mmViqXKXvcAPBO3eswN4SXZR1DEbcVCwKa
5QR5kl6sUMGmYZ7VRaqV4iSoiYhqL8vicWzIAcNA/f1dVdliEI6d5E6GkWpg5AJ3
jKOmWIlLmjfH5Ac+Fb8VeJKRyLaBdERTBF/xDnmh/RfL+fucg0yrN/vqWFKEz473
KrqJH0gl8A4cEO0zewJElq/A4PPuhJLCeJqbBep0Vwoa8NnZ5SVAMkUl96/ji5yp
zjYChqNyULmQh8kQuqZA8rqnXdpLXWR3IkLSItnMNcmlmQiaX0lyifNGSqUXKtzO
F69RUL4wFfuUFgxt+SKkmnbKb9kmaBCoUMZxKb7G3fnlJpKlvaU/DH15tcXwyTgq
jcAHdH+VznANfP0F9kBW+Crlw15BD3j0cpMw3vcrbHyZKnzbCcoWcfv3dubDOWef
GbBawCqE8h4UaMYOIZbTMp+rtZ0eypEnMP/kChQGVEVrtPnZgdn8KTnhuLWL6TC8
GkAR5QQoh1UdNX8rcy9ReE1MEPZDgOQ66ciGlauErA4GBFdE1Kq469wIpnt4WPma
UbzNHDWWArIOYsiqh+eERGXq20twMhTFexHhOrIJoK9tipO2hZwcIZZ7zeCjs5Xv
vxWHZD879UXI2zaMSrKdN9ZsdHfXI/23I2vTT5+bYVdEBcJDwR4m43ni62yTqMXr
3pf+Q6zkWdzZ4tJjM30xb/GDU9qhSBTIroJU8AaPi4vdddahKD25ORIDcj5WB6A7
fxsDLx4iScmSEIi9xYzlOoSWt4QRcfJ1Ge+l5NHyNF+HMs/nN42duK9r9WvS0aat
9OrV56zEsqfp6jRkFbhi1qPQio9pd6yIM9yKs72Es6BNHTQJFl/pAR5g/jA1wwfP
+I4T3bWC885OMd8XuZWbPAxSU23s6JTFaKcBcgUOIvwAK9dlbL7bab/8YZmLAheU
HhfRd9gZEXGcG+RzGb5chFb3Gs6ztB0EgHnH0gmI9gG74cRiGgwpflCQHfSzOjRj
gbSMN0yDfbaP6lq6m63twCNW9vkh+9zQK6eUthsbwddbesUg5MwdS+MUsY2ymi9g
a1PIa6tps1HwHgbuKRAP+N6X+zP4+mCC+IubagnVcaxYjcBM6KhmBKTyHCaxb3J9
FClRZ+M7Q9BbGPCFOKVzeiUPpszF+zayLNhjyYMF+XESNseakQ4tVRDG17LVDYAu
6ABHrX7XMKcWgeNx33ibEd6EHbQAOuzE9Tou5WKCQ99bdp6wbGOEnamX5RYzZNfa
/5b1y5fIXNeVi7Z+bhSB0IxiKKd8SNg1iMUcKqWrkZnfvQWgjvfvA2xDFMLrL0V1
GQLc//y4axvAsHN4UhGtW4W8cEKnkDFK+MfHRW9YWKNTPSM7FEwqHOrw4dPMcNXV
/5UDZYWpO2QE9CXrCp0Z4M/4h50hOANIyyGuahoTf9yEpm9QI9dckRaf5KuBfmCt
yigkG0QiE9ptRkR6noeDnRtxq/G8CbqXTU0tyIZQFMUsPv+NthvuD6fFEU4oNs1F
aAJCMBHppFNOVC3QQWivRN9LA+kzbrPHoucFAYawynre+a39wBW7U2dIsljs4LnK
+U8SCweT1FzB8F0djDC8I3Mkl9woOmnx26lPaw9V7mmmvFL1++O5ZKFBeIg8hvD8
2ZWZSZ7JP6P0YVvJEJERm1D1YM4hbQTMXRUGC9B6HmcgF5+Agm7yKm3ZDwS5N+lU
gO/Dq/H56wIRydvZ2Q7Q+bBEztMDWW2mbBty1d30hRH4D6OjfHRBNQTKtbh+ZVZ9
i1XdLtNsPZOI1Ly2I8O3477or+Jbn0FBK4KjSp4sZbXdox378/wikgKQOn4OU8v4
Mgc8ZmNlMV/lO7nOuSehbSoQCocgtxczL/ZAN9rd04sRi8K39msUVLm6Of/Jvpo1
c+BRVHtXGwuzigTpPgqk/QEHXSUvMPBN2YMw6Pwri0Px2MKa76JZByGNR5Mn0ce7
IDGgNpHL6PToZw34LI/CpfrInK5FtdBLRTskD/HLRGDM5is18hm9cATZFACWxqO7
qMAris0u0dhQqUlJZBegVAU03955jdDv2CZ+O0TgB79YPVT1MSMf11/dWkZm/TyT
pWAarpQyd9zBe2FL497+NAS8ojQj+CnhJiE9XfqKCD6SDvyMKQv7T2Q/vKGg6JGK
gkbjIUYGAFHD33Nkl0y1LJxd9G4p/yunp9r0FyzWayDd8alKrEDrBhdG0xrq1j5Z
PYJr1DZC1+TLSiuG/owspyo8iX9B9AN5+uEXAvrSP6k3dmt0vCw8kZQVlMWv1no+
mtOx+rsSjTImMRrNjiWZTr8DtHbWqXpQE++HbFBTxfLs6aupFS4EHd1IveRSZkhJ
nve8dRk2fyhFapgk2NJ6Gfg5hgMisXwgV04RFoXGfrav8x5V/BOGJlYsQAw1/G0m
2HrBJ0nx1DiOckYhpIK7EOe817bqyBIpCk1SxU+lwqUUw9xWyYWKEsckRBPjsQ0e
z9fgR/OEdg25YJIhKcI+rr0oC2RQOUR+a3beiKXT7q9FWP8kXpqS4Lb+WRhb9Jsq
Oisb3soqg1yoOXCIhp/I9HlI2BRbY6sYacRp78H2T5q+JTCXVb6Vrvsv1i1cFH32
/QNEovzZnJ3aXBpxN8CSptSrZHPHQLT3+nPEDag7nmbP7NXuINQikBDrWOF2xA9z
zQ6QM74+6ULSvIhJ21/wvo8OyvFJArtBZO+momr+wFNAm0rw6NOKACmwZhMvQOK9
gddPNHqhq1g3w9gDNd4fBlypJkkAzIFvKGzoqSS6KPPoOqbKHP5ukqcs9fBCXnoG
MR4hu9gOb8oo43AiSl1Dz4QSoly2H/+h/cp0+DsPcaE3io0sFjWBvCEY6eckXKJQ
g8WLt3Nz2Y2YiMShDVP7ryYJk2rSvKoZw2TMgxVijL28dDguSuAFDlo8H9N5VH3p
azW0w1dnRI+oYMN/22PcOtj6dYcjQcGUSIvtjRMSfoxLqs9nB40nZCxld43yUOx0
++JqfP65kqHrSq6qimfce98CilRi7/0g5KPcv9fRG4xivvkqL9eI1z6ZqdZoB3uE
PzgYPr9PzKs9iBaTMtz0J/9qkj76HNDc8o15BsDY3Iwef3403LB9MnVCuVOoKpOK
yM0nmDSTqPB7t6P+N5HhjK4EKt87Qn6iLrNYCybo0pqgxqh0QothYmNSEtVGF55h
4UKMtFyx6PtM3AJEfWm0T0YYCK83ZBRjJQZdCWW8zpvih+Hfil+mP8Wqp8cPZOcj
spNmmm4H7f9X+Kal6rfMVYF/pd1wlxXuqWnAE1wcSn0=
`protect END_PROTECTED
