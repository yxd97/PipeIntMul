`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpynsiYQtMR+2fjbEWFL2EXvmRkt3ktJWXn9Pgt8tmW78z6RAVFY46UxdAQrrP4m
vCtdd9fUCMgFtVekGT43wAam6xux5MHdrjINfHjRvLPrDevqplsiNHBCFhYZtLjF
v5EoPPqwvo7vvcJNtz5c9n9f9Y8RryYqD/pLFFKmgrImwrvQEOPlxSSTrX5wxqK+
XjlASf/aXs+mViaP4wjpQ/LOzfWEfXj9RnA6eXvvH4HEVJJSatZKRO9IFXcqSgKb
enfBxq2BkIibPArlzBHfj2tGUhzwZbHy6DHFJtlQYgakhufzNVqQ9ApLX40GYLsq
GvH1cv4YA85tR73AK9mTX7g21PfZZ4k90rb77vKdyLziTYZuB0ZSo/NJUyBtW2j8
Kzgl+hxy1rmZsiVKpRcXDS8yPELDPl5EwlUsSfIs9NJae9H0mpkMiSNeLxSP4RpF
StcF4BxNjtlK5voYZra6bwDm2OBVEglUlugbsk6hBEL6YAjWJtSb7SR2Fpw8siIH
VfkoiWf+Vs86rxejui6Mi1kwWODyk9pY6O2HrsXXOms3LLZJjcSZugHVWkv0FTXF
DL4cn5g1VbY2GMc8bt2NYVxH2oebfHnDPVPK2SGSsChrfxycGmcR97yWSbU6KTsD
Vp5FUET/SlailQktrcURT0aFcsC+GSxhv0OwisRf/jG8He+jyW4uJ+sD/wxTet+3
joYV6z3POYy4afV09skf8T34ulCJEtHc+FAN3ZCFUF4=
`protect END_PROTECTED
