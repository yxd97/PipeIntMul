`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RkMBsmxufLYda6l6Au0e2nAggqLNF8BU0E5rWNdwNKz+flFzCHKhekBUVHWNHZ1s
clLzwQJTqYxv2X/+2EljSHApPQqTAm35XF7jLYfR5xs08UD2hLAF5gAGzPxAUXHq
kXJWtrmZQW7nUfcLavGBNATbQn/5lac642Qnj5GV1VNp2eT1sF/RMDmQd6ZcuZEy
vYNLL9eiMAU7icbYO0e1vtmR+6tZ7Y0nl2Zcvv0Q/afLUEQoY9eihacPOVvIzdew
v2sAeXaqdgBv/mVhcFOz2qaXNjdvO9NaGgjTrWdIPowjLomuLJ6E+Zmv5ZbYKAp6
jst7Qe2MB+U7ervkKi3oPpUMqt7DFD2eLYXwZ+nT/BIOE3vlOpm2GIXwMcqNAfEP
ihPZq+UN1kizgd+nEfiodtXgCnCvXqsIlhhXT2ZKZtmt3BU4TxZcXfMd7xUnJvu5
qf2bOe553IsIaMQpY2FUH82+LDxH4CY5PBmEtoGKVtwKopJKhjs9E48I/NTa6I+a
ltR/mcGHSz7WB5ss+NxDOjecPykTjdUzSWhrfGdclrTy7kwx9An7MVtNnKGsJnjl
v3NM127+RBOirOSfD5b+xPDygQkwiJQpi9mGDq3cXpO/bRMOcGQxVSSCLdH6ilXq
PqJeQOoSgZUG7vNZpJ9cYTbT/xm81DE9WPQ+YRhINNgTsyo0ihc0baeebyUhwDen
+ZeOHoScri3fp2pVuju5apqzJTQHREjXQxsa5pBU0usUQaYA8HbCdROpb9Tt/W1u
ny5B5nBlZE3Wlrfjqpktg2k2fEsSr1LoeDwye2fGfawGyc3cJ6AiGC9qrXmEw2tK
ZWQSznnpTW+V6t0jBNbeq7CArJj6mchU/9OdmSVgbty0WD1Am1VJ/5zQaQRxkkvI
0IwCqNxy2gUDZxDI4AQFvxM1YT0NAfImGTIOVdEWUAnftkyGBHido1E1X3LeukwF
fK7xOrC4JNO+yxLDMm2NscUW7ylop8s0MP4NdtppcxNvNfP07e4V5cx4h7qNgwcZ
pKgPj3Y7gPO+8PcvNEyv4FqNV7y9f5o1IUod3Jdg8j9jF1RX2uvLWq1FXSk263p9
ohgCLDQURrgMPO6Lfgi0RN6B3Gd6Z7ivsTXnnLWgXBY=
`protect END_PROTECTED
