`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9UP0B6BUBQhJrKFvz+gi9Hn/GjHDOuZ5zQqXPDM2YLYHRYmZn+BzCJnsPc2kxeqP
wfT2mlIk6KcNTZ6LHYBCbe+/hXUX+py40VsavNhLlEYZoqr3jv+kSByYjOjM6+36
IwLhU1dd/h7CyAbchgdspkbVgFeNzQrsFBblVMd4wtBeun34NMlBQrCf7dMtvTgX
uGDdthn1V0wspnxCMUxlCAG6XRBr/OobPrh1rU/SQVmmXzNHTlNkBivkZRoD+ai2
xAoyhbfIAOMI+9Oe+CXkAed5MHRukd3/4u59nDJDAauL6feiZlyvgDpqZzgJ/u5Y
WxnzQgAO3Bkku+5+aB+wJRJ4PZwtDeDy3B3q0TXrSh0LnSqWbhqlVrTbs8UISqIc
/Wkp35ySCy3Mf4fS/hSLMg==
`protect END_PROTECTED
