`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wAiyRxewSvllRulqWF72BXcPwuRB0HlVPrG+7tFSVqrPyrQ+4bk3gp8XjL9Rkekh
yFztObXT5bbmi8PiAZxMmoVjaSpVAeRrOGhyLC8HkHjLhIPzdf+qRMtaKh0xD2ll
45XTU8Lu0gxs1UzpdxVGVUleCoQuvL9NwTLVturNeZGpkaNGenFfnwOWCusxA1zj
ZEgIsJx/hfdZamVDihb43X52JGQ1RzFAbNyn8wxsunCp5ntUMZtHh3zyA1O4iObE
LMYpQsqCMZKQsErTZzK+Qko5g45K4e+mSlDBVdOFqij81k+5OYkt8EHpqa+T9RVv
nVEIxWePJISXxrkvyCPa89PAs+HOF/O5qLaJsgR4sS9nbCu7uxM5fpqY9EB9Bik9
wsR0efR2/xxF1moxHKLaUh403VD/lYZQsvMUy82oOjqGoG9rEksbxQvKLrOSGazr
hMCD0lTldXPU9kgzP34+SZa1D1R2bE+A52xFqG8BXJiV+tdgUksmYvj8g/Ki3yog
2i1925N4o/xzgKdKWLNSGSF+EC74KThqyVTyYwNkUxTVAr5wy9/XdJDaaH2usvDb
bnXodV2zAsm+PNFqcRuPMGhTl0zZW10IIaYFAhE3xBg7y4NX2OJkGXnpe+LyqiEg
LtPxu9Ux4xJ8AFKqmoV9VP+TU/8LiW1VvJRkMYcIkEaeIRPH69jo+w3faiTfWpIJ
979joZTCSXObUf1wMf5QF2/9zf30wZ7Zi48CMJ4w2dW4I+mYelogfWhPn7u972a8
au7ljSZGzYL3Q7WFoP9gl/HEtMmlWZ6jhGRa/dLTNmuvkUFZtjcBsecZeWgJM6IH
NP5thO3Xc4xBkQHftLmyjBR1LbsTJUHTB4+unt2Q+6bzvhLxKJOXIPy46pFAmOhu
MAJ/+63wDaDPeceGZrtfUotaatMtpsngi+LjdDv9ZzhDCxqXndre4Fan8Og2hnwX
ZMFNlEitVeLgqixRCkT3I2qoplpw0pfVv0BMnlkZCb8Y4ARWK+ljGn45GjHHx8QJ
WcRrxiPB+qpJ18j7CEFETbDo7GjbaGkAVo0HkxHdjSGelmTEHGiQoWB60mK9/9nU
2ezaqQu5k4GKl+qx8WV+kk3EF941UlZFDGrDM/NWqA5vMQu7goEXMiIQYrWoTpwZ
34cRlfcfCO0hjZeiEA+nHw+8674dW0TklG/GAfZ0MosxX3JqkXMFdA2VnlUpkaBv
Wmix/gI2sNVp7B9yE/wXdF6BPViqiJaHiVU0fg7y2ZEABU+LPYmXQrJaxzEZny3C
c7l6m1lfHwp6VJptc3mkIZI9/PzvaaWveEEF/n2X/iIjpSwzOeSDrELRvjtI6tff
hssJlmsRCP4I9nzWpqEldItpWJ0nLgYcIFu1KfueOaSmfLN4ksQBTuvv+47ZImOu
GLeja/BtmfePrFwCt5HeFLybrdtO3CZ97Xxwt/rBGiDS3orNNOiSXazPVxcVgyQ0
j+wbInX0ut7E9fc5Y6+js+/WAgQ2/TyOrbgw8cF+ZQ7aH816tt2UuRS6z7G/P+OY
82GvOj3RKM0rwoOacuP/+wHbwvoBD/qBzpvpt5S86xD85W05Kr8N1YfhY9pno1W0
dD6eEMlq+g6WufkeUzdqBdwytXHqBIlJuHr/ZrkSxofpqAH2O0xmtxbtoC3zuT/k
jQwaOuhuZEs2e8uYvz0mdlMQm+8d3gpDCpdA9NhaBktRVnZVhMksAYnfkr99esES
MN3+OMkl61TS+iyXGBGXL0MwawtyCHGckloWLHkKgYVhc07fXXl6WC2DCJWv0aWr
9AzGWAF9IzAtdNQRRQLuxX43sf2bD8QB2xwk4YR+eXQ3hojbUiYxP5qmkRsvj/1d
S/t+Ul0viCQQzqjOsrwTMGMl0oeBI2IvXgjKfSCxWUXft3YJR/pIxhYr5ahnvuit
/9o+GH/5IzQH1n/fAdbnRsZDSjJK3gaQbBihcFn8iTJzK50DxH8uPnZnJQizkBFD
7MHmaIbcSGKoklWmQyEDfkL++7aLuygN9WfYh8ZyaeVsQGOtzNy5iOFVeNwaiLDa
Sry36tfdLTfVxbjcnr/Mg1XZ8Kw/KB28bAkxAwcJzTqUO298sV2OkEUVyTPq6Hc8
hELJU+1yPert+ADVFzPd6vn+Lw3RORWqbvkZM8WIbpiQKR1q8+0q1ZdpCorQQ9aE
tL19jG+mo6qfeZn04Uv0raEW7foPpuI/klAuGucWtwPg3ZsEedQ4/YfHNwoxhx0h
TArO/NAD27YtFFLfLOYOA2qtbnNaCZx6HRA0OSmwQ8VDrbSXEQDe3AUnMh0vbcGs
wQBdN6rE73mGtlPVJMj2tiyEqvxmos1vBCXqGVrGyZ+WzMcGRkfIvnDdt/yINClB
SKS2PE8Mg8Bt4SQ4U9SB4qZr+pbOg5hexM4wkQSmuMwWkBwkP6E7JOhdzzjDAOa2
OMDT87FQL7rtS40vb3BwjfY+uu8j2XniXr2g177lIMwtO1HfiBwx1srjjYfhFVwG
K5HEUj3gNCoxQwSjTpkMoRjnIwI/EAwWDNsuf6VeSpDz81TX0ZytxfrIaq/El7Ti
eFhLILf3FYFP3cdX8NwAvM10kLLNRnwhdnB4AjAv1amaAboJStDEIFOMF7fDo8Lu
fxdQv/PVl+fpo3qvv1d8Vv9CzktDNNxWTMBhGih87kAKFfjmOFjCB+qEi5LRGzHh
+6w/+yMqGO7NMIfTxibygJDvFE5hxnEbEx4KoJXk/CXVfMi1Xf1RiuK/5f3yVVOf
lLui/8IcbH+WJSg7BUA4yHM9hQItt0ktQ74Jv0tTUyOnWZBg5p6igdBD2vWUsk4X
vH/nWNHixrE7pyu7R5P3xdk040B1cbGMZTjoGs+GAwW2CSR7qnUu3p2cJckrM6GJ
AENDI0PXA9pAaGrqh5100WpEoDyQmp50wPKJuKSSU2Nxz79OLEMD//h6uvCGRWa0
skg4CVxMwly2YD3cf9xXVMTH3Wz89rIkCy584Zuuj+NBtF99OCsYhY/kp/mZl9yY
/FZXVovpxjYm32is5GOyvZLvPVN7dGaaSh9RWbLrmhM2I0GW+xfkdSWh0CKOULdi
yw/VEiFnP5d1B59y0PxAp5BMEWWgpa9/MrUFXZL/EYqkdJQPFRQwJd6uiQ54b3Dt
yXw7UEdUI3sY3AQRvd2GAfAeQhKNkLWudhO7sWSZqwQwT7ZNpD8iaSw7OaQzwolV
dceK/J93sfz45/VNDbPLEBBVyhG4SmafKAAQBCvjs51Rs2C9AXGsDOYN3R5Hijkz
TD/zwRjMjLbm9D58aiesUGZ3fpiA8hBZu7y6NDSWKLbwj+utj0uBnuzB5i+hSZ3g
61dRL2nnaINmDYTJagoJXpfuliDcpVDTPWKTNsIv3IlV96jQOENtHrA8Yn36aGxA
E1x9c84c7WyYiUrwdii6J3/UV+YsWsQYLpUlRfKceLoyRQwgLaH1ENvscdV6KNzE
Ie5Ipv34uybtW0nV62oI6tJzMZzkXsvrnq/ww99TaTbWxZozzTEjGl7dpOt8/s3Z
l4yZDMaFcala6vAk3MMzlL5so/A8wTOI0iWWbvA0GtQg9XudRrHAMJp3ibicecg8
dg1Y3ADUSb//ZcC5AFQU+DtujffL2P9fQKRAGsctkctjLr1MwGU9sB7hZnxy7vOf
30dd0yKTEc/7SoIqZ3+JZbPJ8GHkvJ4HiAWwxH5ZpdrCHUJRktiA3dNU/0he+BGE
ZtXwWt/CHXkGCAonFBsSA0Oo9kqFwvk6t43FPH5qSZLk47hv8IhcCHXsTWmLeR/k
NSRzOlytLyqZd5ltaD9YV2A+o7xciN7oFUwXpmNdZHttD6yHudRcseWHEPm7rnR+
RZ+wZbseMiUEdAE2W9XZP9KUXhxNZD46mJxUmwgtS8O/K5j6GTBMdtlpz9OT8lRz
vLobJPfcWuPwV5MdQ36NXlbYW9IcLo9zvXL8LB2gpbVuu9T6U66XJHgSHyir/3G/
Z/rLlvQCK2g/WZ6oaz9xsFH/OGRLkRlc2W259Ia/w0yc2XnglpL8yxJzohkcGEC8
DSlNgEZ9drk0LegWuVw4WE2SWkAVwSydxlaa3gawHknn6NARbn8u6Ed80R104pdL
rnfH6qaYWFx19hXjLl29v3a9U4WDeZwswo6nmV4D4rkuvokB91N9OQMT9now+oFi
BdcPvOYKErAMBQERjRjmxwBNzXrXJLZuGfVq9rp+92pgn3+8W8LY6DEjcO0Si0tK
wHgSNsKA6+D7mmm2dLut1YgAw6GGZw/r9Jk/g3UKLlovHqw4EGMApMJmv26bRPe9
DK6dA0q7+J0IZMdMEGZygdZf2AKpSBsRlJMTeVIfjj58pUOgMyrATehACJBfUSEU
nBYJiVGJ5PckjwZzBOduriBs7gcYADDEnovlXGu1BHv5gyD4P981ZFBFAcayCT0n
SyAZPewmfE9v1L69SxZExkswRqqe3rX3f/i5nsz1TRP2LMOQSvG6rCmiSOB37XUX
9Xyv2WmdLvi1xwbTUlMQBSTlPBAMbgqOhdvD3WnMiMFPhpdsTSgWyJTRcKaE58Qr
5JI7v2xM2/MBUsgBw5ENdj0VjZzGNUKCML2Md8jaRdKg2fDBFJUjCO4noBYj8Er7
j/Vq0TGVzH5RPPxvrc4MeVl3FteR907fEVOWOnXcMYjgF1jv1AZJzSIpeSJulqql
JyH6YBRvV3+7EYuUpvu0wSXv5gApSx/60ru8xOLBzKYN46AOY1owJJLbOwrU22ut
sdeArmQwcdgUZqXUdlmQxJJYUOPSljK91O4hmsgNS9QNSNCW282rBaJj1mFHNxP4
WwfjlrCTiaby4JMbpzJnWHo03HbNSWHzCeDDF4AlZE6fX2OP7C+hapoC2ksDaO90
dIKBIcAmuSteV49I2I4bug6eY2c4LwbpIDozQchP6Td0nXp/XdY4iWOYUlZDOxkO
aFLdxtb7ktxe9BQD43lElihtVENpApqOmEV7dELJLW5A0BJDK3vbV6JxjrFZx3In
hSHXfzoY+ExHDczYlJBg83cyZ3l7QaqvKH3IKIh4RczU75r5qRNzIcgcSlFWcGhU
4HQZqYV2nDxR+iZ9QEP97OwUd3ukQuicKUskAyOlubsPmMWKzi1aoJ9AtnhIekgE
2w4KPx5hEOcBe5T2kUSxi9+1U2DgiK2+IKjVmCe2Nv3fbvlUkOqmnQBCXzTBc4vO
RxKPz99zCdKYRJ6EVnNHgwitBLe1cuDgYyj6QeRyyKc+f84PiKw3jhTt7dxNkH2D
vv1viJ3eBP8k8o4QN4jhxGjozQbZ8F3uxym36tdrO3ydcNRJiDs+FS5s/sXAYe4f
0tVIa38k3ewWLHwPSlMYjzublYR+AYYJJ+kq1nCLuwi3Lzx8BvwehPtwrqEU9k9F
ycXbf3+7zlqixfWnwkiSJrrwu0KHqZZlURw6uIcmia6ejQuYGqWCSfpRI9q9ildB
WMCpy9q1sbwvYBoYi0JN5HDzeXMOlTBm5HEm2gdxJzB1vqkB51QhA1rhi5+DNOkY
WQM+teVohAQgkrEjf+mRYRb8TRXxUALSK/TjIcXPDCGXNW9yV/zS1Q8JUPlAicEt
1lHl19BgiChG2GIwXUrjhz+2gF8f7+SWNtzq0kokUYIVdvx8dGNPWPBmkogEkZnL
5FWZiijJikm13C8vOEpf6Qod1CRaxkaiwOQ4TqTVb+25z4PGe+KzcdYjTyp12yI6
r7f85rbVtpjjkWNECQs1b6hMyzw23scAb06qxJxgxQ9kveQ8sa4LhWi7Y6jYmb0Y
hrnOURk1LDz+tkOWARXrpTxN+xi5rfm+LrP7NeQWaTl3NWZh8cwNOvXlwhEcFodN
HiGZvhv4OAkIXqgexllXcWWE7YU6hl3Oo9znq/YE4w0pEH9jNPwFsbEciWNcigZ0
Sej2o48+IgWxZJk1asW3z7KyDF3f5CnmJIgsIVaTMOC7bjzwLe5i1yuEEctx8xV6
B90pgIQNj2JTJbaIhE0NY/bhYZZjWy8QSzuBYTpPOioIHY/mWtFEx4/m1aiIZkfr
yzztqRtD6dtyB7nVe6Z9WAUz5rg1zXv7jRMetYzPDU2hImG0nzhcKzx7xO5Oqud0
tUAJLwb9I8gl00A/8I7DDEdEO2E90saOkrvejFI3lQhWcWsWgXdqrD2szgxDodYe
srsFxo2ACGwa7Uve52NNlEoJv4lY6Q7jh//JPCAuSBrI5jY1OTjZW5fME9iFuIqq
uMg4YNmxLh/CCpFEDvbaOWNCzsudgLFFx+Ka9HNcsK6EAh+2C5niijYFT9a/cuv6
Z91VI26N6lby25EEZ8dyDdVSumylNuf4gYHgE/uSVN9rasHceNqpK3tpMnqSXFC0
UAQL4i6PKK+Y2kuByddu+zKVH99yNm19dwFG8HnfKGJtDDMNcqgsrWv838N3CLAx
EePHwLV2/OV38E3EdsLpvfH4/3P07+DSsM7f+ls/ncV31VWehKfVbiQxJzaU1T1W
ztfMmd4XB6xUiU+RSS2anpaWq1H1anBHzI7y9E6T+gK6bUbm3Vvrgj/6VdfYyOKh
/M7ty3kEPSGAoiKZDwL5sXlzjiOUXH9shsJTqwub854=
`protect END_PROTECTED
