`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vl4hDtClLuqkQkj3nBX9HVhGq7v2s9u1EJBoSjDDgekKT3isTEyxOIHO5eUI51PK
Quw3Ryn40Bn9fidheSIdE1J+0obESYNuHCNEf8a55N2I73/vjFFiskszwb3eMU1F
u41cqwIDk7Vpf8jYsWGPzYHhLOOFyGM4VWGIpUiEsxYkqDkhcIe+EGzt+JZx1ScG
UMOpn7eSZrd+UnTghBAS6BSX4JQLOjKTAGxFJRYT/WQICQlzr/mJnhpvCEEer83S
CNv7aiu0pVxqM7u/30TymXaC1rESXZ2zYS0Bafq3Dj7kZvBf6Nvz9qJ620TMemZ3
I3CMA19XPunE/70I/oPqPmoxpI0Iiq2l4zDVtROfakrJMvLki7Cv7hgpv15FrYVr
zVKfrshHe1XnfXkeJ32vjQpAgBQ+gazcW4gPqGUmt+AWRWtJXt5ajvaJxbVhWztm
svbw/oZ3stgkyndOU3Mk58juNWJAFFT5NVU3runruRfs00Opde+/uuvcH2frXHE2
6088fqzE0Qt6Wc9YTfZHRY6kco319iMzmEksZ9jYKICaQa+NmoWyA4rNQhqkz5Wq
ZAIwCLyorQIeIs0ZN9XD6gt53Gtpi7CDOU/R+QJ0DrY3Gp0oJtFjP6jFBJ/Vwcx3
T3wlj6dP+IAV5Uj79G2DI1M5AcRmWSUZUceYRxO50qF3ApR36m1MLVLlWzi8Sco6
e7FulX3KDut458UVjp8n2WAuN/X9Owtmmk6cQe5IhurZH/BEO2SJ8GCp1mCkb81i
EXG9UmIdgaFjPkSDQs1S6TIGOfjxHWdqmbLFqGdYbdVZTK1cDltatXNeBXTS28rj
V17grwHxWU3u20WzROQaHMTomYZDyXMQ3fEI+/L0RY+qanlo3ZWm2+L+TJa7LwLm
Svf7BLaxsPcXvSsS1aX6AwgMwe7Na0mISl89UCQUWheRwkwneQgvAj8yzQEGAZcw
hE/x04RhnU6oF+W4lN+KHAS7DgApxdniEZdLUtyhSBFxe1OusAkN6Oupx4bB9HIq
FwW0Z6mPVA5zcgODGzw+eIU5xNacVTeCWfB3Hjlh3xOJCavwY1MhzJ/XU3AkrtnM
WzMpJs26g9Ele97VlvZRolVL20v7apK9tzY+7yTuSqkIS6H4WT4BYL6xH0oqstXB
NQLGgVOKpT4yamOixWfgKrll753+1q8GbgLr4U9GMFn07nNNEd49kjuq5G7ZR0yo
dNe9VQam4cM2y/5qJcPj8BKvWFYaGaMtc9Vtxi1j05D9J/vzRin30zmHBxKeoYiF
VIkZ6nXk6vXbS7Z6bMMzPg2iaUYVJ2CFaXAG1aI73U4aSGnBQlSu7vRhXCOf4Uuo
96SLFBAupsIh+UxsKto4v/esBns3ERC+cQLiTVw9gg7yW/uw+RWnc2CXKa3ehGzm
QfdjOHYlkJxxpqYzuEfTZaVF7pfO9Sd3blXjGRpTirTTGOj49wtrXrWYCKN91L4N
jJ8RSRyhlpUqRDkSz1nfUx8fD2CbGCYOLWr7WBPDO1484N4Zj6+vn23lH8P/ETne
Rxc3EUxy7IGE/YtzOVF+T/MkNSEWrzv+MehQ1nYRP3sdF8GHKXS1eBUgrzGu00i+
uURVcfuXypzy9Mi+gbhmXx0HQeWCWypIA0dzwV01lD6aZmlcJwJheqjYFS4F6qc2
7JHwUOjCtELDmA4dX3ZUOjuF5SVgRMkz0fObDEyXRTTZImLBf4GdVSpUnejTXpuY
53qiBkRhpCjqnLIgP2n/yVuERFDAlJA3tfc80mwtpKK/Qy7wwbgqDuIJ8lizmz6g
ra1e3dHn6TgOIHtbBZWGfuT5F88tC/MYnGgijqbzEuF8DVJLXvHIx2P+hlLPJ6B3
kP90r7kPmEr+/LQBeXZtCezKpmnwCxUpRUWA8C0j7A0Bt97xUQHXDCKZhST1pxz2
wqPRpkPZ/N3+sXSjsvYfBdkwm6d/4SHb/R8w3Cqg5I0iolS9AzBhENP1mTn5bvp7
fgl22XAk/TAiG46lD9uqQMKdLeJQugJmU2UIhb7rTNvUNn+Hvh1tHgc/HoUmbvk4
Mj76ilhvv9rnmv0C7pA7MKi8FuicYdXBOfyyHu0M+hZP9JQeb4JM9so32xLTedAB
0Cq1tnOUYb60N0oTae8g6LvngdT9/LnmxSLjYQ69jrPIMncm0/gC47A5EDWQpubu
ttFJxywhZMi5z7MSus5+uhX90vfgVNeINQB7gU9GKLYlmPNY8IO2AUsgucdqWW00
0xUGGBW6agDynZh1BEQMaso907SUA37rRm2VjD4LxDWVxdpJI0OnzYTIw16+L1sY
4FeDfOMZIHckLxvlUAiDVU6P6SsWcsYrSvLeggQc1+WOq8flNaGC42W0irZxZtcG
FmVNUQzv2Q6E1BlxuMuof5h0+slOBc5vNq8HDKxjaOv18uM62Np/4cpRKmHUnRqM
qYWYQ1LlmNLwvY8sYZVkTET7D4fv9w7jnI8iI6jOkutGKqGHIZyoml7UNIzhqF4t
lJknXJc21G3/vavBooPRT+wB4yq962OhwTeGNZDcN5tl5ArLwZXuE5ipaIQpvpW3
MbEo4qXwxYaD9pxpVvRX30iz2cFTK2zBVHtHBpdv2xZJNkHT7JdHuDhqMQxVGIua
PQ9zMxi93jmARf7qBKwjAI2TSIqQVZzfB3EBV6E57+gkvOe66Fyq+2jVHd5y4Gq8
TLInVKBqctjMaEofWu9VT/SQYxrLZ34wIeWFsjG4dAS21JetwvgMyDq0pjFADDrX
d1hC5XA5YPPQjg90ku2Kfyf3JZchopMgXbeQevPmFC4=
`protect END_PROTECTED
