`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hSs0eq+9S9ptyLSzBKlOlab1K566PFSkBUaaadBbUqYeYQ6bZTWwHPUEhP1JQqXl
+8DpzEGJAy6kncww1Bj/tMoZ0jSuq/3TWuyXpnbZD9zgdlRDjpNLT++ZuTW/hrBn
KmKX7qTjYnI8LqeVUNBZkDlzL0gxSSHVWPFR0YXCCAg7aJJgYaiCc/orOtiDciYa
WT7rbTG7Dewb7MSVqeURkPa7nH8OOaYfd7HFuUrYh4uyNsBqEphQJXLta1fdtwTp
5X1Uw6W3T/or8oeVtn6wDfn8mqpGOh3K7jTe1fLa6Xummbe2Hql24x69ShT9JeyT
YqN8voWnt9ZU60UBx2B3jMEp5e2ADkPqc17ZmhBb2ojTR9JrAbOnYbAKQ9WaAQbR
146+hOZgWpDPahrLNImeLKqu/SG5pY+f9EIjetkYuamMVLD6YzyMqq0YJS1WNQo9
EdgiJ2m42aaRzBkXf7FgGKhos6JP0BLNdTlXHyZnzA/2ZMtx9cPy22snccJDGOXI
Z3i/Yppa8qFF0g20sdKst2JbQb3R4OwRXBMUQNvERHDxO1XWxEuQam4t5S03kMPp
ENvvGMapo4kt919jlsB5zxSjtvmv/Scr15xdt2Q7jznQeYr5v2sQ6aDZg2baQWIp
XCKvoKdS+SjWdtiG4awnMYkccWqLSEpNyUYpEKzptbbFIZBxgpnJtG75O5bMyKLS
da5VRmrQOZxMJMQ3EhvG+KQLcuq4sTFCtjfG32yRvD/kGTqwPBc7y7Ah4sbmN7id
ApmKtZ4EvEkpOcj3IvGVjwae3F2dEL/RPEyaupTKS3iFaXYjquNiwwyHGiEl3jgA
Dp4ORrr4Aud07jh9d8ioyPLTT135USv73moRDtk495Tvqdp0dkHDfOohcD/pNQcU
2y0mBtOMI92bi6hF5+fN3DNRBIAZmpAssQEF+RAaKl1bc5zNw/UoTfhk11gc5nmE
zGw/o0LwyAuqvEP4pDb2T7Iu9hreatkYooH0GmkPtg+98IYnKYqrGlbiD28eIvBG
rJX2HX2YI+VDecXf8g0RSI2tzyeOTrkW2sToCCJaO2lVEg5oDWhFoA3kpTUoV+01
ZpjdiljE8n0yhhm/MNq5F+THN82YgVu9/pQpFZuqrygfW+YTDZE+RDvWyCiZsb6c
VliYDXId5upHM8pEUmOmxDeQK2lx1PXna7q8iPdE1nSnRJ/skkyHym5JaeN3N63S
/VV3CgcFxRB6aS1YpGzy4zU5eIcdNuOJhaVHewdBV+aFv/6FNuWN11PfiugH9O8N
ri9KG/8YFgZzDfttP8UVTtYAT8dUp5a+OELm7D1mPXwZSnRtBopR2+7q0W2jqdSB
S2J86RmZOrrqQSntaJIqB/qkOAIPNkD3DZZKemIABNI5sppP8dapDExIb1tQ/XF2
icd29IlgwQeJHO94hXpzLG+j2HzTaU/x+IJBlwJZ31Y++emMwkcYZ6h96zK/Vab2
NT91JSX+RkBv3TFU/S9TSv+bCSHnfwIbI2ZvL4EpmWAfmY2asT4a8HXUWKSkbPFU
Oy6MLOLxGnvA8Wt6elJLEGwo6tfO1bertJ1ffpWDqCanA+H9LEMwUQxJgZjNg2ZQ
grOdvfEqn039eLQ9uGTSBDCchngcOoI63fxkmpKepa76IaAExyH1fJ9uDVfOBMH8
9auf0XT3GRQYExGaeANvLDrp5JxWcbs/MO9kvqtUoqpFq4Bcv2XS07iOL4gQ4KC0
A77xVMIfRQdYs+dbcigg9xBMub07Kd3bYRzB1WUKAdzho1vjqbsEqfsKDNvWZq5B
nYjwxbTFcmVWMy2bJuRqQMqL4j0tXOB7QhFvQ/xkcSofRBS8HlbDhH9ic7BfzGyn
SMzqKHdO8PHmO7sg7UMj3Fu2hykn90urfucSQVBMCsRnVvxeV/NfQdk0BgAl45Qe
Rp3twbkATQxpW0KgHYP2K91XflaDKVNTfgMSQ/tHtjxOAPLDZX/iC5rZQKTf7WdA
0e5AFbyVtRGRtVzqMmrFiJ4dwp+azVmkhE7dSStVOE8YTMXwL62k5iWrMp4MAfHD
z7TK3bfm2gP7yV0X1p1Z46N/DvxP5vAI3F4h9buK1nx02kOJjdHSvBIGDylV/BGg
j8YkyjCJKs5Glp2a30bY0RCkiObwTO75HeoLnl54gwB3rBdRwYOOjltHpk1GAmUG
8xcNM2BzeNkoxTOtcZHh2ySC6M9AZj6dINgZpBTwxU3M7svxxYUhj5CmcCUHX4hQ
dl56E0y5QSSFd+Sfr7IHh+hK6msAmEQBGU0q+gq/howU/8x0EbIV69FskyzkAi4f
A3lgXMIQiFf8lzxnBS0csB79qX/4CNNa87GIIIs9lIfCy61HH/CP6PBpqLEfeAJe
6vvwNtcSs+Z7LS01MvsVB0pGcsT6hQOkDysptIefJkeCwOg719e6GSFIdwQjotU7
29V3jiZ8/gwimUeigZdEYjTVvLp+M2Y2rLKsJy/rT0+HEQ0HHI2ldv+O+rgNLHWD
ZHUGbPeQ5CpMlgW81e8u07XwzBok9hxwA0tdO9FImgT0VaRotC0z0HHOBMyEg3dS
CKLwcoSz+lRHhHYhz9WZaYiW4HK+Yo22KrrWfsmpQ8VbT28JIgV0awIsd68WFZve
DDUhL1cE84hXiW4vknMie4/1wjC1o6PrDjWl4M7gw4g+vbkMx05dcHEabW/GNpGe
dhv0LxHkB32k9tiwTPnyHckTnEFrh05J3L9oJ5hFdtNl6yZxBSyjVGM/h+Tq6iS+
O1A7acj3kuIrG0KqAfA0Rpv/IRHXlF9g8fyeWGv7Q7fprnzMCjbzfpJRSYesDDys
ekQF9TROimlg/gtpNkbe6+HDdIPEXidZp+Fsaz6JiTpLzzqN37X5CljG10DWNlu7
0MhPPkyYo6+OqWXh5uPnzrwbVm9I6ilIAYLhZzuxkGzni11e1oYp+iwLA7NeClLI
dwybbpXN1uPCOW/V7srUeF3krbCa7CNXlpYdXiYESTMWuFx9tx8CzZWabN10OhIZ
4cmxyObCEwX+bunWfVqTCVULJxCq7wy/iuBbL3BajwSlyl5IIEjo3f+DRJhVs6F5
+9Rb39GZa/upEpLaLYxtBzpue1xpSLvpWICKSiQFsh9G8M3hDH6hISOMBJKcHtsI
KXVFuv2kqzPuA8BaJe5tmJnzC0jMWrdX/HesXDsc0JeRCzI3XHMsEnC3UmVHPIl9
ZmK+Ys43E0XTIeoFJNHdo1GiTdbqhksDt23V7Is+5uZsmkiPEiCuct3tRTK/SkLt
el31zVdHYWAVI3xZdfcKVsowZHZo3/4fq+QjcWCIwgcWEiqtmU+OwJVufF9FLO5d
pmh6oXe+uyrjqCfJE0bLOT3PYy82jyQkBdpcK89FN94ebl50Vfz9SO2jPtWFSlHO
9TE1Qk56BikMYQsBChZN2xAGZJC3UJX/fh/odCmwmSsM8tfNIgHJSvc7JU4FU7w0
an6e52wjaglBYnYF6bZnCZUVM7o372FrZ7KTqpTAcJ90DbaAS87omFoZqOXckTXQ
5kvQyYZOBrO2oKDT5Viw20NHdUgS/SaHUHKJPIJGDP67YsgJPRVvoMcJr+neU/Bw
Ncu4n8kyXinm8qU5HugnjJRaRXJhwoJxlvZ6lfwBKFdFtPsmnl7zu7B+TxYJQsSJ
fHB8NwAJkXSrDEgmSswEpg==
`protect END_PROTECTED
