`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D2DXLeDwkslJGU9nga4CqXS33Z6Q1cCtoH96NUIF9t/jYMZWGLBNPxITKaAT+KJ5
4dzyPoFOEVILfyagZ0FuRkZqrF6JRNUunWZy6nG3X5v80hiOhWm+NRSZcJiV6rHk
PlsJOvjllJOrTExR68UiTlmiw4zRSg5BRDECADmYKxSCRQ91oD6AwtLGxt8erUeQ
xjA1Nz2e9/0JEoDKX4gxIiV3cXrrM3K5Nv0sdOlbJGfe3Gw7B2+vm489gcdKsDjP
S4G/e8qI0pB0X5hU4RQfd9xTlmBT00Ou79AOOLlJbXMQA6R5jI5axDQTlelcwwRl
bJDi2/hMmafJWLXI16LNBcOgcJKxMcFxOMkdPlVKTPISqE38TDDNf87F1tgw6ruD
CDr7/cmX6eb3Qrg5Xraucw==
`protect END_PROTECTED
