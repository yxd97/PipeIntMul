`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jM4ivXTv2d26Wrttq4he9Y+AdLrCQQPC9q5SDjpRFBa5ndrnZQ5cVPDxJmwmP1Fv
be840scK11tBfRf3IoqMQPaIl1pd2Cl4hkBJWlzD/fCOxt+sEwwA71jAQB0LjkjI
kGk7UB5atuQqMK7R+AwLPTIhuQnzdfsAJKYYNcxL+UWIm6WP9/uSJwBE0Mg2LqSx
4S91zYoV8zZW4TpPbWThrwOMK5XeJUXIcj3VdSNJLRn8xcWyD7p8cX9DnCA87WSp
BW34hzZeyfp257SDSX0uc2262mpbK8hq0INZveUackA=
`protect END_PROTECTED
