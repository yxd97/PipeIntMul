`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fc9w+hJatb5HUYGgZfSqeBOj1pIU4h+Ua14na7sRJJL2RB3qwaWnYEi4+ujHdFke
YeyYN8IKW8VuYr1qCIvRmAq+DE4M3xAMZxJT3mJOuM3fjyVGoRMtpD/NJJPEwbeX
0Spoc7snWjV4IG9cP/V5hwM4iN4uz++3aCLj8QNul/4hlTXHQr8IDdtsGg8hGq6E
tEH2+gtC4OYofy0v/RtQwdCb4/L7Dei8hlODWqmCNn/lYyt6NTk0LBPrLUUacLe1
82JYehAX5AMMflDKZ7Rf2Gh3B12WMaVkJNPlQjRf7iJWUD7N+UWRIm8aYVazm+TL
DjrnMQn6CudZKr0vSoMAd6PGX1ZG9rqJ86CfSb3CfilTcl7HsTHmtS9yHirH11tZ
zOYH2kr0P5T9WYnN96eep49HxTHzSvGTuCRGhBOy+0HdBfov4xF2BrKPxGIjdhRJ
`protect END_PROTECTED
