`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t57f8EWu2OrQDbfkJHjIrLrT4I/SnOHW/JYInAU5gsuds9/+yhdMxSN42OJSxY/M
Rtt92//OVpUXk5xOd6vdnPCre7v6UV3qZelMzjvijVBAxYzd3YNqDCOzPsOpPR1k
hO63RUcLvxv6wqApxE0lW8rT38Bho5ZEq2dkZevP2+bHVxX8KF7KbRMNNiV8Qz69
TNmjXW/u8jGWk2SPH0eSXZy2jp+WK/Smoxx+KobXMOKOpFYUEi2AzuifrqXh+Jrl
f+t1WVmrWSPHH+ShuTxd3U90uYZ3vKDEvXfBbwPglFnsx4LZ3y+jkTYvUL+lHaDL
V+uCTy/SXMTD6oirNUTuimb2LVibsGNLpqQuTW7OfDFw6sBwBGad/Su2fx1RwTIX
fp/SmiDqcc088FnsnMcC7X/W5bf7D4h8uWtWw7zn06s=
`protect END_PROTECTED
