`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y0qpAYH6qjBGRdSHxMIeIsqfVUea2gtEJLD1x/yftpZgS3oLzaUIJKiXLUUCIm9G
A2wJP/TBvW9sWHvQsfZ/qal2qrPLOITW3R2gfCztZsPGRTEuyeKYkInAone4qXRe
JdAzkN5nQzkHS2JYppMFzLUKkdv3Mn8hqZ0oLpE5R3fbT63DQNK29ZJg5IVt/FZu
1p5aHJd7YUwHwUFqb+AYU+PT1BTK3mGNBhvdTmTMonzT7T01BZ+QfO04fXj2NgOM
tpbLrhLl6RebaQsGtlIhLCSSBbWKZRbJLvRsDV8hLXeNcuDEmow5d0LflKljaE30
fd8wvLoF3krGdZJha8oSQ8IvEhkILrvxORTGnZY7+iEke1XYtCy3EE/tyBYSVag8
bKCqauGt2Kb0zu46av8I2UsH9ahkx7liMEoWyloxR/U=
`protect END_PROTECTED
