`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zCtPBaG7KOBiMimNVwNj2su1BIdv5w8zq5Ck7fbhDMOYzs6/qSkI5U1yQ7SgUTF3
PCAQ1smHnibNk4x7fwTASbff9NQUa1obGklGudoMv3Cn7M3gEPeVKa0vFeY82qpx
s1OZ6ERMXIvgQXD66BR63ldwzdMpwKX3T+czH6IzZkPehzW6CmK5C+WGJust/tCF
qgPzMmFzSi4cOkTLGc5c8xEkLN5WRKYNMkcSH9rn5M44EoZRSl+VpOEeZaY62aTk
GL3xj8lEJ6yY1uFkLFpehs5vpXyAPb4fy+ix0rYWWREaVmBTiL/sebli5nR0tog0
puiMzSJ9i/VDHHfaSixp1ZOLqRqqRTUiUXbe+NsGIRBzaCa5o2DkJAkSPYn9nvyL
`protect END_PROTECTED
