`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1HqWfLxGYwICgqeI//C387PevzO8i3mXISEg/PigLp6tk/tOtBuG5SIRyF2Gu/9
KmjFoZPlRpXAK/uaH9QQKDWfm9ujmjjOPbHhyZneBZH12uU1AnElimCoQNFP3NK/
g9Z6S67UdtHGMxXuSOJQhbnIoP3MakJOOyk3cylNFcFOYscKMAChcCq0D327bzZG
PJMwUY4riv9+DGHkvN1wn4Pew5viLLoVXU13oz/t/LUaIHjgO3fnLtiheleevpg4
9WreJvRwIrSmbGONMWEheLaDRkzwQ93mq1yshEm4onxWRjTZc6+s9hD1zl7+c/pQ
fgKYPyiwmdXqVa2ml92EdSaGqLSKQF+ln7FO+yJBPmwzIwosoX1a29jbVPu/DvBc
aOAmVIavkGvvplqioGns+A==
`protect END_PROTECTED
