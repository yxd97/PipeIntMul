`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRa2Z8FsTNrCnMtOBupu7N2xzlzfLVfTEOZpLoI3Lk+orwYtaJSHVZWdUMetJ3zS
Qdr/Bspko1rji1uyByGzEQ21/ZL4SjjB4yvhC6/Okh+81z19stEGnQLHt9A7RXVC
sDBmBHQYTBHJUWF6+uwsWKcX/PL3op78Zd7LAQrnvlRxbBlAfFLIvaRGAd2SlIEh
x9QjMNqVWULkxK46rSMvlkqE24vfWnyDxIrMT+V4onOYi9IElFjDrVZHhQbYWD/A
YZlBiK9rUCAP01Fbj7BTig==
`protect END_PROTECTED
