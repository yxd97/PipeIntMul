`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1eAsOwQHhYKh/U94FqKcEIrqD1iAb6r9d9LxMqrc/Nk++Uxl7PipyGOhLlJG7XM
kfbJQvoEiN2KPk46SwRUYyBBck5w6avdrTjHgXRZOvy/INS8RRFzFg31jwP5GogI
TYHBxNMgoY6JeW6RWwUQI5kfXP/p9fRLn2xwTGnHh7Pj6Up4Yp9D1MHR7X02dARp
KerKGjuxxe24s6khXZF/I6EHXwtXGNLH/XmUzjC/O2Z/6Hg+WaoIqmbX2Ah/PLDt
5ze/YXwh8UhcaQWywHBRYKTCLKTddb87uYtAaCGEbBzdj1Adj/aOM/HQnMRc2XOq
JrHar6RQVn7Rk26By8xLUmhxQNmEtD+/99N7hKE6zoFcDPCuS8+ZO02/RSZI1o5k
0GFunMAG7B1xhG84Oi4L3Yt+0sajvLnaKHEyBQZHawDUZJub2PTT111ESubeMJWd
LU+EBpDvLDBPhE2eQhf0aRtLjuBwSW+dpPfJ3XAEsfKKRJggqXfMasyDIRZUMc9c
CcVZCWCtgL7zp1uqDRl1uSFfR6es9PK1KzsHxJCPafFeUUhbm/EIj6Q9JcWPV72E
wlZNUKTsKmot2ZQsNUSj7G7IM/HYTSO/1Cfy9p9PHxCtwpWso/EWAQjb8GDP4B3y
MhLZT0ygXS78R55trR9LEPy9BIRFKZtw9uq8DaCJKC3bY7EvYKjOABU8ZPmkBegV
uSbdQoK4T5fvxpf/Tgq1ZQ==
`protect END_PROTECTED
