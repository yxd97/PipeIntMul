`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
phYZcwR6bvC5kvVfkZk1DnSc8x3qXvp+LsvF6aG1qdc/aCOZ8KMV7d5Xnn6/ieiu
Jr1LLaKr0S3+BeynsheVHnlvL6W5kWTosYW1z+bq5Od8o39lQgTepDgu2B+TjOGc
UJrfFN9v4kJXaNTqL/ssPYGqwbyyUDYWoVFr/6rEp31oM38MyuNaE6cVhhHo3oih
zs83hUvljhFebowOheE/UqMaQmRBYevbPHaPM5CKoF0mXSCN+EhWYcmTIQbCnBjq
AGZWSfctOad+4+Jai2MxvLOc2uYkDZEVaVmDpWilhRHt7vqMl5RruR0ei990/2hs
7hiA5gkIXFYDlrMvPWDpl2Xo1x1DVS4TqdSmBV7ZrBNSmpvSw1AUwuqWhpSvlLa4
g67QnyJ5M0aDe52SkuSzXg==
`protect END_PROTECTED
