`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mnw117UZP2bt9wnf+cRJJZtJi67zhRrHfLxqLFZbUS2WjXXcS9kppMmPhPj4tbDJ
P+G7/w8n9Bkwp9U+YhAmBKthvqubZucGtMfRZn3tC5JrBEhnwho4V4A1HNRSP1Tf
4kPTNi/Wfj2jDkXJQaf5ikTjl8FganoekD38E5v81MI6H0Jh1oQlJ6inTEQNtsAN
TOhWgLToxWJ4UMobJyH3WyLb5tpA70khqwSc91EFlKntLQ/MMTLvp+v8BGLf8MRU
ZeO5gVCornMh6MQ/MJ2B+TkFk1JPMberqTY4TKxux+7D6JyQa2OSNI6UjQeCSZbf
Q7j1aiEcOx6biySd7bkjIhOr2o/+zp8Jh4fSUJ48C+foVQ1HxxmtMTGOcKk61c4j
FE8SyqUlprgOIjgWI3+VoU6bkhc4kvMjRTlwUtIcqjxipZt6cl6auyz4Y/1zyXPW
xFpkymCf4sBBTGgJ9KRxTSFvtTmhWHCBD6t9gzF8LDy73Y5j/gdhxkyG73mMk5nq
IrQj5QJV80UIyhwaK8mmeVtOYD+iinTRICcEccxXEWv4JAqWodbRnJACj7K2suvV
vagImiGxwTG/jWqxI1nwW4qexonL0mkcD4F0XsmRRGtXSRlIm2FW3cLZ8i95XBMs
uwSXsBW9RbtfMAVcNSDEJRD3mLOrpIFUud4+WeO7sBrijnHXeZ5XHNMw3jiI27DG
nJH8cMe/SV2MKVQFkQ8qoemAG7aQZhh35M4J6RmGER6P49L5wZxI5XWZMmIEHs4Z
VDmEXlEVvUH8eG4c14UUVA==
`protect END_PROTECTED
