`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LzstrvSuAfWZW3mNg4jOW2XHWzD8Y+/bqWztb9qI0ig9G39yA9VVl1cIdrPf8TBS
7C1zOpXlamqncEo3T+OMWKYPkVkirKJLrGstpIPiSNX1cq+S68+n+o/p7oCOTxpd
MfMulfNrOpd9rlV9/EDBeSc/CDnBaeqbfwNyPyaMNGKUG4WsXrqCZomOK6g+TRUj
mqWwt66Jv6Ekqkj8vplA41sofFofHS08XBWFdAb/E8dOehxZEEnmMlbHIo7l407u
lsmuWWVjAUdeY0TxB6S6adH6a/qoGI+XfiRSibRSRxl/kw1ithDP3RoDRddKh44x
iil7kReTjVpP8bhZYjrfdhcD6x/1HDj48wPSQ+vz+S/U/YYRRu5gDhSywUHYtz3Z
K1MCzVJGQXTYmbuFdiR4ns27S2tpASVJmVqTpsTjZZjMJVYa2XmxT/MQgybWwJCy
kq0KOT0voOJx1Fshj4F/Bxt6M2r+UAdDfGVV5yOrwwDLm+w1QzTaJPdFSag6g3I1
NVYF+3BenEqaviPfuQfN7SfEYf++2oNVah15lxYC17/0Bju0j1Zj34qDzZHpalNz
ExATFjdhvohkiqjgpRwsChMpyRViBambCM+YNrZRlktp3JaN2zwADPLnPLOpODAW
H64dvseBLI0eFoy1fyAjUpSgtH9achTM+5g7IHnVurS6vFqTDWmYnYVNd/wLtxll
6lfMg3uQC0OYqgiQtQ/9uwTOabFYzoyLXlzVVzlEQ3IHkCxpCZhKjsmQ9um8wL+0
AnYd1ImjnvnTNJFYgPoZolKWZwPHs25T4EcKKO9fwul4q6X7fsvVksLDGZwjsr2+
2sWVXcu5495U1jJhkfTdNvkdIyDMfi1mpnHOqZo4zHfa9j4MYtQGxViMoXA2NkUx
uacvV6zfjTRWCsiDo5A5D2HvqYxm47OnUr+j1VgY3itzlpn4bCzln3n0ExZxSe1R
5d6Z7B1RlscLboe/6pvu/swzyRFaiPJ6Gm0ldJK6mlWdCLdkxzFKKZKkhrZQryWt
Hjfark09FToRi/2OHduny7ajJFA5sRKzLaE+v3zEreVRZzsqnln0J+NGotFhGLbF
fltyDas1SDpPRvY63ZNc4J2MknoO29bpt3tOOV/exWUyOnU8utHzwkEWWDLKI1wI
7GOA8wP8o07k/5mxr/C2PYB2gHaY94GT+BqcSnRwcS2jPUADymbEdQJBuVSv7abU
AFVTGRdGa2pv1uu9AhaIVVsWt9OT/BccUTy0rs+o8Bv7UOVH6iF56bHUrqvLg7MS
N3XRvHTa1FNXIOV3gLLujoGvLEsV3LaZeERB7A1jyJwl1Y/8H/q5PMj5/9E/Y/aM
mIp6P6qPUBpatmA0ciSd+nvU+COySGHLup0yf3iiE8no0zJqU3jbLp27Cg2mJ5SS
inWxffl8xSgri0T620G/1Kf5b+B8rZf8Bwo+oPJdavwgA8WL2d6aAGQtGTjwk6Zp
JdEOrCH4lZaA60LL2VQgMXHWemnA2s8agb0d0uyjXeRX1whndQAsbF6QVsmE6/BV
Zw8WIwvzSFqWrKQwikERlt/EWvVQjoESPq0ffWzQPkDS5SNVviNL10h75SGocR8T
ovkFAN0YF2jhCNoIor9UTKUqsS6NXlNljrqVtVTDFHDEt++cEY5BsjS5fMwOI2b/
fnHLYnNEvtZdtB7g87ef3LIE9n5bxJhl84RWPLNFoP/65xcUBiAVDVILmWwZOE9s
Wv6jh01p4usVLtRx4LGm+PcPoonMxGfYA5I7EpHeGogAyLaeOf9gowXe6kNQ7eqJ
VrRBEIGHXGF1NnOzkO3tlZnc54MW0YJNb0VHkusvlidMjH/5Sh6PLhbYZX08l8yk
yjX0Jys6wpXMoI67sBKNyMwtoShTXYoPPtgMs2rDGNY/ssx9s+hbTCm6GshapwyU
CjVZy0WXsC3OIxTtat6KzHuwoHKhbN1rwhoBJQgObuybqtPukPRWDp9bxK4iUqdf
rUnzRzWqcSPg4lXSWYrumfHYpFUJs/lW2YfT3PRG8NE=
`protect END_PROTECTED
