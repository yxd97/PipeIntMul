`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uSE73FW0C27yMWJXRpKKnLdujkElRhaupo2HU2ayy/NUZabPIxU0MHOSd86E2R34
h9/2Ja8cFTOSjGpfYCiHetv81Qb7dL/1XNbp6Ynb1sX17lEYG9z/A++C1DzklnWa
6NnmE8JmBA12fnfsUH5trk3ykDQeWOzqFdWO4W5lqphAQHCmhpRRFibNbt5lPVEP
6k2UXSL6OOas3HM+V1AIdlughlZJLzai3ht8m3Li448czZu2V/Ig4DR2i6hMAtWK
X+LRcum7eeD6tNq/fFfxaQQvd6KKSpOi0AJz8GMzt2+RsaicEu35oR1fnNT94gk9
8l+/V3hqsk8mKvVF/2P+r2JKurtICPiuwi0VJnxgVyw09EM8cOvmke85LyTw5D9f
6UmvRZuNYmEvJSUWcbe9rasFl7Qx2zioU5pWHa29/IGOAgsf+V4eH1iCEgoPZ6/X
WBa5PwNVWKz+dP3bXungDgmuM/2gRZZpKS8qn4fT0rCrdSQFRvdLThIRbslVOdhY
dW8+P0VjPffmkN6eSxJ7pGXQ/Mr2V0HHm33l3gQ4utOEEi7JOnuzPGQCawBl6rCw
BUKlyg7lBKhVkpqfKles3WC0o/TlP8ufdMih7DJmSjDiESkXN0vS+kwp6ASH26Lm
fCW058iP7+6hBTfdf0WaDjaiplo1stF0HLvrV00P5Ujf0atqNsYo7DA9ffRDXZgG
z49E+xFcM43pQRXmACiUQpPMbUxMbRvXMDo9dRMj1LQShqYxl3fBB8nmjAvcRQey
QB6+2On188AHXtvIY2un3GokzCbd+PymiufgXBU/tUghqhsiZvg6MbNFKX4gfYVO
ZXBrsUeYjZtnQ8eBNCVej95eXU+PvIChsOjyBML8D4Y4LU+wxdF4y08ggH4lsuuM
umeN93iJkUbyOXQYS7O7+2Fkvm+kZNWiAiXznXA77ZN50CwtUlLyOwFKuujOb4PX
LdJ4F5YZ2ffNFaTGHMkRpdii8UxC5oyhi8dz4WguCca829T453E5BBFQX/eZ1of1
ofSIhMRrc4synU7BjysvASPaKPnhy7fPChRPRLeQ/yXWf7UnYY/KN1KsIMh19LY1
sz4xF+ucbbNnwAWVaHVLwoAzm4sU7mwYixs3/4HBo8WldV052lScVmN9sI+HUDpx
T2uqgSEW3OjQcr9jDLv4nPeuqwgmKq/nsPbHX8fRVg2Epbs4kDg6gD5o4w92UG81
6kypig7QMlXDH3ur9n2GxLwZr7da3DbsiNQYydm/dR8VVBnxV1T+krnLArsxNzOB
eWmCjzxvdLrvsHDRDZ2dMHnKLj26JkpVd9JOccsDlgD5bMPheiDkELvKcYLnJxgo
+Sv3lsyOus7oIaz+S6JlcsA6GL5k6T7YtzidiVacdotkNsVOGkqhJ1KIBninUr9A
VdkHhFu9hjbFAoFCCVHNk55bzkaNvUKxhboeyTSI1cY+qTKMUc0ii0zSA3pTNld4
dT3N0a1s+PZ3mm4cb9phdhNv466onXjN91E4WoK6uP0gKRELkrTbqzWOyo8eANIq
Eo0d/mPrUrj5r7L/9uH4Q3wiTRzycZQ/cEugSt1PZ/OI1k/TFjSYJXjhgIeBGNac
aobAt3voNBMXgXm027T16EpI+Kak0agNJwvOHnM6+pDuu98wp/lM03Cbj1iUwHgH
xTA+SUUrGK71vPgs7NiYk93SqsWaBl/cp37Vz+K/JGMfKxspXTvbsv5U3kDvdEQk
uwheKvjEpO2eWnWKNWJQbdT6S/xUU0L4871bARX5RWXGHl3pHnTnPaUmHGM96N0t
8Nl/1e66sFtLlGxHIO7I2FrwnHwByAAUoMW2maQWcqR3G5+iCm3HT4IAS6Lpn+Y7
h6dzR/ha8Nk4wR4/kQmPKXDR6Jg9vsXKN7nDavXYIDVFakaLokl8TlF3HahhW24o
3fOqY7FOexxAkSnCcGo1pRAukUyVZaPx+p/Ipgit9xHGQM0uYNfMgTMzTciGGY+D
8NDyCbCk03+OuQw9iJniqnQd31hPA2BWXtZNYTXAilaa8fkiSvQ+a6biX9VXmR7R
o3oYMlL/CGGHAq8yhcCPIl+DJ4njcblZbtapQ4gsGdNsjXh13q7+dHTW57YrCvop
SVn1rtggZly1k5ORC09QJlXyQxCsNIENFl+cuU3jI6ucGXODkmqGRLCF58Y7m/kU
QCaQqyA7DR1Ar9lKtZMNs0kUPHr9Ebs1VCBQ9OaXMdr7TFmF705H92ln159dAzR2
qAETD6Pqxsl4fKGFZKkjfqYPJsVWB94yh0lzDBrsX0PX2fESIj4MAhQRKuFLbdFT
2Lz6D7aXYSh3/HFVK5ZlvjaY0NWJ1BCNQ3FThaDlxSW9lAvTsiu80EG65XPZ0YXs
179aRupuAqTZC3MzG3xa6V6j0aoSJmK5tUoCQrx8+LVF9MprZrbECCqmZ6vohDhi
Q4YC3cWWlxAQguMKC0kmkbjvR9t+SLrXqL2D+sxIwJpD6EXOeb2WV4HYTQir6x3M
SCv5RO9FBDYUA8qtZyeAj85YsHqG2lFylaZ4JjfRaU6WoWoQZTKgAAPd/C4s+k7q
4Rgx/7NA2yd5Tru4Pp/UmBQu0d4qdZXyNYJNJ6XBKcAuLCbz9hFLkKrcUb5kmsOE
qmDfF+Uldnp+/Hycm/N6isLPJ6BaBFI5HnKMyy02RHVtnWrHwvOVobqrRdFy42fB
Fg5s4pkUrbVGDPRnRViAOxl24vgYNZt4bZRVcUhqNs/7Ax0FNV2DVOEE1MUZtlkg
uE+VsINanuYALRXfCLmrW3ok6GeMhRga8UWo5MoZWL251yr//C0JSE6zVuedptBP
ylgRyT3hNVtYW/y65zrOKqc4YZBWr2O72Nqm06eg7nSQ6bVSjuKyZb+UoCHcvYcp
oiklWXDEyo8LG2Ltdc/SBqCJkFVGC/EHVqxo/B3xjO60uLqK1xUEHa3l9Vtts7AT
ilHlR9OtqpR4Nx458iMvrdq2YbdFn/VHxX66Wr+eNBv2sabJ4zgoEBF86h26FGFu
w6MJOVEKBdzPPj5sk3XiDOkxARBYjcAQnZO+XXkHsY/nopgqsy7OHsdV7Ogec5kg
iK5X9Sk7qkDBfbeW7pveoFQ4+SGVWqTDcRLzka44UPXUTlf0GUId7rBw2nysKqSt
7q32CVUd3+lnM6Gsxbp7JEuBRrHdVsIe+97ky+N5OqgJD6pJMmfnozZR0k1Dh8Uz
37rs4e8DT+lhVfaAXsH36DESA6PN0OnXIoYkui+5ltuRN6Ty0zJKCBaoce5MUcIa
JgPdyVYfK/AFqFdgXA84UEuH7DAFqYi7YY0wR6fzBEOdJ2cwpK6M+odCVFqPfUZm
UJ0XPMYL/R69oPwHNlyDKbV52bxGGEEurPV6ntIhiDMlP/PY1gjm0tZkyMji+nsY
VhIZCHi1DsEAYKFy83oynatjsJJgijXZP2ofC4dczUMPtY3oUgxiP7v5xkB9n8JD
oMOUNEWN3L6IulVuqHh4FfjwaGt6zE88V9WPnIF5K/vrG/3KEejqe8GeePWiUlgR
mOLG/7MVul7vbLaW34wnETIbS1xiD1r05YXqktZunr0lsya1mud3oZnIDMCT/zRR
hDSr1l2gefHNEoututMu623MjQucOv7ySILF1eWmbyaAim3BFe/W6rBdoW4V8xlQ
BpFYqmg31d3W8jOs2eKSS3BRv8UuQoib5bM+Ipq4aIe8kPoAJNDsWHGa76lL3ZTB
rzcFc76e2OEK8RzDj/4U5FL16WnmpdSGkVG9/xLY+TxBSC0x/WmBXm6VdGl0s+bI
agZm+TLHE1X8ku7RIlhlbRcYqcZmv9HIxKB5Et06t/yisisf7h3bTK3LCWXiUg3R
aRZjG5DFGnhDNzq9LaaUOFFztbAe1FQXRird4T15U8XE3ZwdU6SoB1HggZP9h4CZ
3ifxWpDBbQa2EaPGJlfE0yRgJ29eECw7ZkpHkZzmkmRB4IViac5uy2jI7pKGJTwh
z3YS7xPUq4DYqCgpg65XjZdwgBIwLN+8saEjAHz8BvOpuhYkzh46hwjJy84ypAFx
Lq8NSYzcKN+EG9RfQ6Y3BN4odwbrGTiC6B+V1j4sXS9zXe0sPXWpFr+G4C9Wo/6p
wZTZjmPD68WfMxfCvhOf4hqhQy1lbrd1JG4ZeWjdKCZvI8763u8q2PcsxzdiiyxL
XR+qpI1859PTgMLJ0aJSo55CsUBUKHoGmsC99BAUvTWqYaowOlaqXn8wx7GxEbre
m6OWhzV6N1dfuLHq92KFKayOAlE0CdUghFtQp0Uvb9YQ1fsqCUYhH227prdvjN/L
Ef+w581EyLmsH8Bfy7HCHj9qN+h9tuSPgm39nlfH1zmXRcqfjjunXF7vG6A3ko5E
w+as/Yp9b6SIevUBJGiKt0K/+FyQEZS8M3plRWnkOE5xDyuEgLGPyQG+NRN18A++
BeroCOrULwmprIJWTExQfhHl4Bm7iUSe0RXPVSp9tREXkwlNez5dUbcNy3gXCaFg
ZR7PUmTbW97Sq6IbnSYOMxfgJTwX+0vWboqJ+5Cvccv3Dli3lcioHuEI2vw0m7uI
7db+7su4bUFbbi48PaV1U3CnDf3uSqzdNdK6KSU7HJAj5Ti78BiZHYkcWcyrnR4G
K+h9BfkndnKyDi3IqOfgpMGV1soLRc8S9JG0Z1fTdc4fE76+BfonJPfsVY5XM52z
4aMYLXklpgOhxBA30nfa6ZCih4X0p3Phss2YkEB3SGTYjodr/ai9/bpZqV5GXs7Y
FSEmccZM8wOkDtmWPyhrkrudGFXwCyNJWW10R0xY2q2Bspmjm3plKcW4NpM/kKD8
KVRPGqZQEXbOOM4+Ce8YxVOHjjTk0TP95BCvYEMLy+1t/HfyWbZQNOZvK/mo69UA
7rIXxN2y9THs22Ld7xph2GxihK3hh5YtwvDLhL4gqIZo+FBO1Gb6twGCv3rm+kBJ
3aj82LpfIltnhkBrW3sEZDhv+uerucwPxtI8Pj5qHLXzgCfPz6Zse7mPF7itHcdw
dG6DUzyE82mhcRTYOaPQmh1RCPufHbVCbiootSi4iT3S914o7IktFf7J8Ce2VIDH
QcxepShvLY6rOxICqKsu+trGVe55cE+QhnDXzGYxQV4F8wxHz80BPi/gpaCrEx6y
wUavHXYxt3l5BK9H0JRT1SdIZEgOaHG522sp6ynMlO6Pix8HeNTwBMQhAr+MReKb
ltg5VUQ986rCMzXPAe2XMwqC3ohqdnjeNvDEk5ir5Kv9713EV3AjNr9babcF6GLA
z7+yNP1mv7/NoGrA1tYrwjz2ukisbIN4paPZTLWlxocY52ncbV8r93Tz5sz+0q5X
cyHZPHWgzVXw5Yfs9srGJrq94aZp9osjfMtctY0Wmv2XbkyoTH5DToOQnBmgyOtj
x1GjLqVfxOs3XJIlwvJQAxFkH0JdAcb1vabVtBwKuiGLShGjAI3FkASh3m68Gjbi
DXU7VnjvcrbKe488AY6YzCf39b466k9S2E5vhJLG4iHBvVwjaMzyx/l6mzkueJsz
FLDpIEF/qBRuBoP8cx+/ctgWKZ5u0HO+SrTdFbHKRnRZbRG3f8lhw0ke32Y35jnL
lC+Lb8z4/Sn6pDnivY3r/FT8QKQGZ2Y4LUp91w+k2bc5V/1e0vty7bxWdNSF0jtK
gi192mwHFL9SOzZzcHudC2J/QntT4I/UjowzVM6t8FxxVT8+T/OWnFCC5QDz/Hs2
pc6acPd8NvCbcIg/q77c25Btk0hsJlU12GaPaY45AqbQ+NHU9dKK8YgtSe/a74ML
lKPNwUsXRZfg+bZ8QZMJFrWX/2j953myOkYFzkqworD1pSM2PwpVv9EsBMHw5Ds8
ADBkeRo1MWVCCezOSjai9eA03O0FcE6Rtyo0bbe2Oan7XSZ0y+OoLjueFN6XkODM
Jyb5R8UGd9ydTYm/5fPa0OjYYXoscGesXeA3yD61FaBJwMUDop66QFO7x6ASLQ3g
NBYjdkNvSAMqJhFTFLKBW9fco/V5OcNljb/zyxC+emQybRyVllYO3Jet/vmxwaG+
F0uiskys8lWrlnOY00k1aiI5YK1fd0AYS6y3AD2ZaeZ7lD2u0h7mEoLt2YT855fg
fZRMyd7oLf1OqfKrD3TVR1d+BiNRadszUTAGl2fMF8omKoWSW3IMzAXRK1fFAVkq
duio9IsTDRLhSoFMRlrBPzjgXksS/8RNxVNUqYE/rFAzyteNDk6LC/hVG75PN06T
0PbSeETLgZSlV82xW6DriQ9stAu7YTP6djjZtVR2ngRnYvBJ8rHJYAAWAiyCMfkM
a0hKvDkyyXSm20Svd6F7CmxknFFNArqhYQRzu06ZsVpnJxbgFWYQcPmnNepXQy06
DULAzg/0fP8L72mwZheJttEkRmguh73YckIX4o+g8alREPX7LAQDQU2sU/E6MM2L
FOonC7hEMBLR1pzcjGTFDz2WN5emUUQ7AhCl05z3HKlpzdFgtDh9VttopmHDrhat
xbcsj0E+8RUECdcKwRJusAvzvhJiMBCNYr4ShSMBuN1mD2IkhBM8+5Dho05qYZ+S
V4pZhDMJVROYITNutN+BR6cvsyMvTXbWTbbPFZiEKWOKtU4P0jESatN98dcFLzYH
h0VaQHW+pE8vy3ubd6B5Ka7t+n1bUo410lbksQme46+Tv/dhywdI8k/F6S4bKJe4
JvZc/d+F5DhVCbpASi6sedN7GWjd3sNcTZ//6VseR8i63XyME6rNaiRvWbXt/sKw
DAWBwgzJmo01Dbvx7DLu0zOgo0m3bt91HkNUrKu9hivVmHm3fJ+2J9XvtTajJUM2
oCd2MDVunXgDphtkHtwa/7Rv62Vf/FQIRTSVDdba8tnpi8ITXYaTXrWZZE0spCic
DuGHjCIesbA37o6KlUzt0Xkt/tjxY6RnGhXibFacnOwzzBk9c2/yZUkQikLNJmt2
lKtVPzh1U7MugIl+8dAG2+O8IPhhWKgzuFjHAPInPXmyGn/zfWZH8x+cSEMp4Otw
05eaV+mM2u37/1HJrfYvgLO9NZWLcM48J5KnnA6OtV0Lpdy6K/vqxOg/0s6/P1Gd
sVY5YU6CrET42IKBsrnbZavsiazrbaNpoVUL3MmDVxl0Ef/MRXYxrkg27CtacYcN
C7ATq/sUmpld32g9xQcnO5Lm+6C6XoMQTIPBmwQPaJXWUuRi786oNZv3oY4T8uVD
ftxxKOM7bJlG7+PMU3Otz8QwAifZWqecqArzH6y8VRbl5sSYCCo01aEMy4nuVnTy
vgg+Ci35CWQwmf3IjnfiDk2gHy6f89/hoMB5pF+zG3M3m+357VmB+CoiB7lPtIFW
qv9Yci3z25HvjESYJSNLoS4RW3Ipq+BS974JvzIlfrDKGbZZ07nDGI45WYAN8xtV
GXhj5nIr5vbYbxAEzqhULVDluumZGByLJefRU4M7mesaqNTGEKAcjxTnc01+Hnmk
2Hh3ABabSdBd0+l7gZgfCMc9yJVdR08NbeN9n8Zx2TiS+/ZskBtAvFG58bW/89to
SFS8Oe1Je++rcJc/INupO1towFkbJ0G/RghMHzxgjPLuViNDkE3j0RQDu6tfXAaW
q0iBdWRz1fQsJ701wkYUaCMWXk+fNNConUkk7c1kdJGQGz2cgja9jcjDBB/GPX7u
Tv6pvmtpnsSGlK4FuqLNEkP+sJnXp0uQaou7u2ufmoGCENx21B/FNz0DVrzKvJfx
KgP53PtPx87xRd9ijDzq+3cr1+DgFYqYWLmEXepYgVah4Wrkpm15SWxCL+C5eHl5
AOcexz2nIFIjQbTjwX70tjJyLsETYNvRS1v1icyMRQs0hHEnTbOZua9df8n+CQw3
ZFe3kypHlpPpB1Ly8jJxCjiOoSeHInYpZ3Mc5ci8Sbt1L8GSdba9uwRyW6FPiF9k
vYw1kzllznDinvFDRyGnst7FMKJs2w5fTzOVDTt4i0sHiTde2HW+Dz5n2V5otVAh
mYmn7WkjiIDhU+orjs9kHEYQIDgmklvZ7Rl1f5f8gHo0l65mAX1NukcD2+NR7wSj
gCmu5SyBzkq/noMmfqFk461sK+WIq/XESOi/402T5nIuntxkh8oOdKyU+GeQQnt1
Ju1sOUsrjDpmznon2+PzlReBqItb5SlrOGxMp6QNp+wPh01kajpzHEvFewd9zjid
U2HkfBexaglMgEmplvdCPouhd9JuHLm53Nd1WIaUFMdS1uzSgQAcoB/vDBnRY0Xw
itocouo14ksXivIPwXiaMKeO/mtoP07o0wNt9EMMDHqRTF58nyNj+7l4baoV/WyC
ex7IOzLDFLp1EFPmocrg1QJ3XDFDNbGAbJcs3/RDJAT0fWAwLbniqwpEzhGdatUu
nMLs+jvezFyFJgi/ikV4TQwFxGlMjsUSxstOLVTEwMscvZQMm9D59tBCGr7tRJ3J
yQAYNqfiV/HpgzJiIzDF/ywi81LoHVm7UPjfzY3rGZAZnqTxrm9toG8QxZjGR0iY
RGoeqYfr2DOCpYviVxyRpSDEcsPIyHBCfLQuupPoyUJ0qbi6S+Zu0nVzCZeZilsw
wkhD2mTNq6XFxK8TaSyA0FhCi4aI7V0Bxeg9nYUiQPiMSUnVT5m25EVD2A+YX8CU
a2Rj7ZyhOqIqJKRP882xBpYyXWlUWwsjZMRJq0s6rLuSaaGd/jgM4lgmc/wrGbsk
w38naH9+mqsUY36VgFp3QhrE83lyPGZEGacwkEqXj6oyrFVA/LhliVstxEegjyyW
dB1LQzQ6IjEXoHxR1fA4BTwoRQjc8aY91ihWrYUwuvpjCS/KpykuxZSC4IJmRFJw
UYHrGSEFUitlEvyqlrHabhCRXfpHmUfm6Uuj0RThm9hwgFEpmTJFcHXR7Dcn6Vgm
5Oq8kZRAKGKWIQDzVYdICmbqRaWDlPvpw+tKFGMQgqsTV+JtS9xjVph1UrqkU4nt
F48i7fnylt134dDaxQOR6bLJ3+umck0eT1HPbq8IabSSIuBvShZns24Mv9ox2R5m
uj4DNteMO04gMyHFteK/HiW7ePy39LXbbbd1hoEXLMn6ieHiMbaSiQJvSiHw13GW
pl/2yuzJPxKu3Sp4XyETlqaA375bjOHOzIwLn3j/mTR0UEowyqtqNjwfKZUY50KY
tUPwohCZPoqYqWHLWwqJppEOf2UEgTn2t/O2X+4pICMqLN8Y7di0bB/tzNRbasAS
MMkNAjU8oDimKurxa6S/zjHUjVBCxHbOqRPAAgAMHC7YnYJj0PmXozrMS1EWzyUp
zFpD3DqZHkjAS1I6PdjMVY3JvjMshaxOB9md4+qxy3I5iM5EHf5sEY1egVQqUj+Z
gPZswNdZkGZ6eCJYXz8O1VAMwPvYgoWSE/x8LAvBEXpT31ny1+kq/67xqPoNbY9y
mjWZZ148tZooj3ApYtzIujkFLSFlY504KAcLEo/52eYIdfAD/gVWd3aFqFLVC1m8
8Ss5RYyYjSo04CsbyqrtBtTaYnENhkVksR1YepGIafydVRKyiRpsn+2JQBQhSJUn
eW46slnCIMA5bFpYtopdU39Qx2gQ/KO4PBIZ890yy1eWcY+gcLYZKfsFl2vAVeZc
0gogd0q81JIAgKXQwsuJt8O20zJ2osnfQ2I5YLkF0hzSPXdyyHf/Nje4BmaZllln
Tc0Jz4YU93cN+LSPHgb9uj/UCoW4SmK2eAsgSAQPq5MybzKtyqTUeyWO+5yM5b8n
agDBtiNpttcPa3Q8E/+WFEq2uVuSX8NuKkgN3yqHTgjoeEfZEF/aAq9+kK/PBWO+
ceDeQGH+nfTtLZ0KSmTIenPGrMsodlKFULX2EV1/V396GuGk07TTy66irVfgXZWK
K8G93Us0GglHZDoOo1mAiopLsiuj5OkoVlAhCRXiENMO1DsSnrCxGw0VWuQYQ21o
EfEzRQqHmlUHcTne9yKW/rFDr2zaftPYXKTaqTEoibRCmSxVZ0OnkltSN8ArFCyX
TWIh8+s1mFIjZWiLVMJSI/e7y1aUk/xTk9PF+VWfh+L2xdxh4ycKIRZXWpe3sZXH
Fb3y2iG0ylH8l/es3NEq41olaqGDunEPrk4z236JrZPOTksF3VGqc9C75o1+rWP+
HA24/sD8x3d/1nec/6M5Xcu1xwfPJghvtEGl/HF4AQuIO/5qAZzzKgKIxkslaTbf
1er+V5sM6RA7gsL0kNkNNoYs5RGTvh2WtvDWVo06e8s3U84eVBKvbhpj5Xm0qB7D
GWsAt55kkuTjtmKas+xC+nDxYhrt9TivSKu4oX/P9NwKi4hS1IBSOXFF25RmKmo0
cklAUQ40ZaIr7RCxTGP0WRxryaiIsCJJRjIAZvCOpmFObz/U0e6TkYhO6USI+/08
Kcvpy2JiDzrXSuDWYXZyy5SG4FqCOCjYcnjot1IOZvYO0lR2tLR1RtXKuXIu4bkJ
O//QeyUBId14TSkC/xW+7M6TzXEz9tFq6d3xYPZ9ASrE5UbONIVeOgHDNoYaOdQ7
e4MT5EEkUo17JMO1c+VoVZo8uFU6qGCp+vHiqL2PWeSo6WPdf0bP5wHSBURKqfLd
m8cdngQt4YNGo3I2MZgl0fUUBBRARtc7g/EMyynnPqvNRfOOlctY5133fPTx/6vj
EHGqTtDTIow27vxFZzDaQMQgR9/IvFeBYsMk3UIeqssG6WyY3nhehS/IJ3f6Yk0i
Xy3mOAri4w4IbZQCetu+kJbCOtTxR0twxRIZaoDTlgpMEf3L66b5uSN3FTzGSpDK
oHY4dvdFPGPfH919byFywnGYzhL4IDFQOjGnDuFoklUk1t7Q/L93ObzJlW08tXJR
qE2dFqpJevk9qWht4aQXhA2zYN1sZRY3jY0bGpshf3zmLZ3olyRDKEeAfV0T5O0X
jke4ljWbSzU9zI248VUISneMXVF/jgNOqZu1+2q5RRa+93D82so31SXLedKIng8w
Ve14E2T56sQ8/WGzqO1hJU+2CW6n7QguFrP5ZnoKF8I/PwbH9JxHSzYSAexQQB9X
uQl7hdaLIKzeHx/R6MoR16aIH2FIQ5piTSvZ4cdVNuDxfHi8XtMPnVWcpJnRD5fZ
ycsaP/K1vL9b39MXOXWetvhD/je5po6uMhmLITkTut841QAevhFGy3JviuxRapPi
9J15l+0TBftBfRw1z91gC2QxUJuer5i9/8uJS5/rb8vVSltwsRTmK8jaWDQbCzE9
qlQ0vHIh1/Ouku6uQkIpjQ==
`protect END_PROTECTED
