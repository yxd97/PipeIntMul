`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0getqQHshv9qDz32neOGJckFgsc/GGJPjhivhnJUFNWB5NBfM7020pebvYVxBKH8
9usg+50ryg0PJNpPY3R1QwNcE29OD/bWhrPOU7v8FqE7kdXAXoZrFZNHa8eys3WI
+e7AP8qgWH9iu0+5RfxXIGcETmqtpfMNzQGMoqJbBWkytCWZ1GzrN8PO1AZpLv8R
4qu3jczsoC36MWFOjclldJt437ePXQ+dlXEx2T1NnexwDQDz/tqBia+M59LgSdVw
K0fdz7raxW298BNPCWuo6+2mar/3/abqcuxHoBD3XhcahTqwyuMfpXx+V8c9hREQ
Twk5LHMcUy/3ycbNHNnapg==
`protect END_PROTECTED
