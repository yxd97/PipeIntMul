`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rTS31vBXep+mjA/+xjYVxTO2QZmJU6ej+JIvBwkwVHgkxmJj0hDflCG7HpTC/O7E
uPQO+s6XQ18TSVW9fbiONeqCtA97g9N7+JkqBCcdJyF0PzHzah3oqWa67qcSZghx
fyqQL3nkfPI36dxP7KDJfMoG8/praD+zFT1KyNi34rRdixM+BD0w6zQuSBIQEayV
xFK0v0F6X24iTiYnWYrtGaW7UUZC2dVVTvrTpMmw7DjSmy0HSQ4u5I0+uRr8hWQr
OebHskfw+IsIpnyFGE4rfa4DzdheX5WR+ur83AFhjidzueHh6TuL/TVjsT43pGj8
23rO9QdjQiSn1PM1zcy9twMfYKOuq4kPAfh6uPyLFz38pA+0JGKFvT6oHN4KF+Mc
24ppGPK7Fw7ZG0XrGiqqNnm2sHxaV6slXVYnBMW0LPuCjKP/oO+Z9uY4SW/LNtGi
MFABhRNGwVvyim/dBx4s8EFPtoQJR7nLxbXxfIyfXPHLjPX95Wa+BbMSRs2fb9jQ
mIdTmA4wfVJtHk2/JUuC3uv6R+2MTkCbPCIqKys+t80r6HUHJuQ5L8rCzWqyDrg0
5TADsH4r9GNNvi2H/HjBpEwqIjC0IZ/6bqKqNC4IH2VU/g8KnTo2FC/5N19v5xVt
zxN1FVskNKhbELkDXCfxsLhd9DUWQrUPQVpuyY6wa2onBj9RT0fXaSf+7Oqoqu3w
193IDqw/zKPn6uDqUQMnPQ/h/GDUFOHsIDC7VzG++5AS07n+yMy1L/NhSgLIuTbF
KPqKMbl2PbOvCT++R5bpMDldNUsDyLm1XYQk5wFK/bDimW45NROaErNMJN2QOHWc
ewAn65extlsZf+ef/xHFazDNDphEdPF3Zxo4ZVL/zhdmfano0R1hzuh9aaibStbB
dUDZEkZUtFdPi6grgzp74she5AoDSNoAa48n1RPOajdDWg3LJC1lNTqxS1ttQ8Sy
sjadaER1TGCBS80DR2qdX5ycQrmUTC/A1H2fxWfeX2LV1AZ9f+YACI4OnlupRU+2
Y1Ip7R0jYe9COPxjCuxgHTqzRNUurgnwHP2V65H3EmmP2RcMEL3vRroxf6AVDvil
VhkS3lyDWofF0psXfqAN/Y0pbsPo6aXVapKAPBjM8oD5Pi0YANkNcyMxWN7Dp41K
6CiwmzXRyWoNi1a+vvNuUsZuEfD4vJ9E/sb8pWW7udmGlK1DBrHgz996d/O3M/Wq
0zNdNLgeFRPQGwL3bRGF32fxWkceVmc++0CNAkqKqnmYmJFFUadhinm1yJ6kPtGd
I8eOqUuq1zaAJ62XhpD76zUtA3yJVkXyMX0dwykI6OmPH8+biifCrcf5er1tcem9
KiOQl+PRElWPZGlyF+q0n2T8AtIXmGmQynhVEj1o/wc7sVnME/lfOzD4nfPmj/xY
FCTuBcOB6lIsevilsrFdeFARDkw0L6cOdTRArJPw8qK8dY4qfz8eqxShivzDfw0x
dF2nL3R/KDkXSTeG6xod0oU2E32XsXqmbghUk9hXfOm7+1Kc3BB7/YzUaw1T5DWE
Mpz4+DJzl1vPlwlc93OeG4eXpDeUKossRYiWZbQ3qObjXgoekVfGot1T1sBl8Bm9
RZ7s9UuILdQwke5owZ81N0TqVNZdJJC5nMvpf4g/vDh0Ktfe7NXBRN31UO/8wcb9
mcO60JO96cFzwDyzctOeudT6u98BBgoqOI+dPzs7HVIich/ryxFrjZcdUPn+VBgz
gN0vG0go4I+Ul96AEHl8sOzlKQNqTfC1+LPrAwey1FE=
`protect END_PROTECTED
