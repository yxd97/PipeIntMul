`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZv+gtyguSTxaxQ2ApCR1r5Lp6kmGbp8K9GM/4+QfeTQVlAMCSjpb45EAa0Vwk6s
5jXm9tCGbpzxBWqNCgAjQDUE4unh16AWbYuei1+dLFgZC3s3/+DO9XSvw8/GApSp
a1QiBoXHyjXlx1nTxFB2KpSZDhH0CSjcXxH9XMHcFYjuZLEwYFqETjjYV9YRXxhP
9/snENswUKxlGv3KFBi2jBQnCzZR9Iz2Rv6GQSACkErFhAz9v8uEYvTiw4OfhBbP
NMln+SLvUZ5o4ZMmyxuSh2yV0u1uIn2fAgR8dRvWzgk52Q3gGnC3jmeGxxpyQTBF
OYErZZFGtMDpgpGazVKnM2HlvcTzKoujpxlrUQqAbZHs8+YwSyiMlZDhHqZQABhg
pVmFAaW1G14CYzACAeOvT3lqlC7nlW6HPXjcSIME+nXcVVTNsX78jBJSVcKaev2S
x+z2O7Y0mcfNcEz3fJ2hrc5a1mP6sEr6vcloP3W+auYqsB+IhbAjO0DBiO7B9xeD
m8eiMNcP01dmMEu3Lqr7Qer2w0Tx5YPuIh71rNPjcHGZhvs3rL4IkiDQb/yvWSQ+
0jsEYWYh8orMqUICOdO90uiXIH2VA8ho3diB5ctsX656Mnz42/o9Xz713e0YdiQh
fno5AxWB3Re05NdT38aA/Th52Gm5U6it5jMv40+zuFT06T6++CgZkW+z+zwaVxlB
3CC40+Hw1AwAVfI28oqSDsRs/g17uF6gIc9iqpAwKXRjIQtJZJ0CGeEEmSef/qcR
I8fEu9pAatJ9zlmjDuxHbOxblCnqv378eHlBTOLTlF/0Gf7m/jrY1X/FcmgDTHJG
mXInAlF+HMRtylZLmgIJGw==
`protect END_PROTECTED
