`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXnqC4nP/JtB1IhD9F0PHUEfOkwCbER1NukcliGtPygEOrqwP7lDPAPUgkpuNRXG
Dcm9jHjXvmb/5Kqcy97LLndKF+GdgTj7aGHihipK2O1Mya1uMGm8B96tz8dfLlUX
s3f7+ykXShQ2p+juvzmnS3C6uhU3KGBAHgaSqYfmMmvWyebss9AtWox/iVZFOA3S
dTGtSew1SyJbywoW3zLuZZDJFc7PaNaXD8bFgiQeaeSruPbXPNrbDiqpWiLDMohK
+6M8VPKpJq1F6uGjQgjBMltpBIJFTdyF8YO7NiHkjpm/LVEikHBCS9JPUv/nvCbS
LLQ7NlHr3900d494cRw/1NbWZJFMde68vlQgNva93ObQ9PWvFEShFdpOKinJ9KAs
4ZAQBUQtijKH0QNUzjY6+YgsMojP+S4kGp+IchLTkjj8jb9lwcDOMCn5uvooqbFZ
K3n4A7wYuE0hDTFKIsa50zPcP1AyYqxDL4uB/w1AlisUy47Ys3ihuTxOOEgriFIO
IckaL8jYoa9NxpM74Yi4Qc/8dTxObG2KYmNwUpImqDsOqMAH/PXwsfSAcvrRoSjv
JfA/miXEp45MRTjQ3eIBGZ2xl6oACGobEmpoB78gWYIoNKE1HsJdYRSdEmScu5p1
E5ZVHTMAhB3feB4ndPIexJfEGFNV41/LMr0ztzxybNrSecu9oSvJokXA1BaN1vfE
I6BAlquMnp6g7U+GkC78/LI6cNROYs/bLxeCGjrK/gb6rPBU0VqBkNXa9q8MnJwi
Ograx8vGWcz3egTI/CmHs8W7K+kfMtJFpBHH8hHJmowOOFA4ZdNzyam/T3B6othK
DNmnicC+LiRWUnvDaBACVa6jioynUR1QVXIMJDdhZU+uAGkeZiPGYHqzhRfyYEEU
Sh57pl/BWauBVxk7bv//Z6/O5Gw5+2e4yDuGS4e0JZNFXnUNBXplhzNfY5COIWbc
IX0yFf742hxqKUpPaoKo2HfC8xVQ+5HpKevAgljRIMhn+JxvZRhGXnk6cmGoMtxu
qGe3sZGKF8Dy0QrV30IQ3cWNIfZ1IFW2gxEKLOvZI9t9SwWC57CLQ42RFqtpInH8
DoORffuMl7fQd8yfl3dEZKmHoTTMA1eEBiDXnRB+Cn0g5os9j1+qWCDB0QBb7j55
Ez/mpKzV6tDe2eO0iGXnBUI04L2yyjH1C24qFxZYhkayOh5grI7I0bY5zhvDgAjU
CaU4MVn3qZX5t4S7LdSBrBalHsABxek+hqi9ArvyiFn0WATBvcVpfyaFbGVjRVVo
zZJ+d3w2OLxhiezfMu4ul++OffN8f0EKyhm0sB0cnvteAzBaNPj+/SbWwNp4Rtne
4iP7QuRJAhLsms3ggpzkZk8fpKvhuFn22JfbJyS003S+5manvv9Tqz04Rea1chn6
I8iSrrnhdNBX1g7UjQks2tHQbHgKyGD6/PJiS1WTUic=
`protect END_PROTECTED
