`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zJGL/9j/HLaRBjgeJSsOTQ62y7DP/ON9jKesyChYzkVOvhgdIyzhelZDuz1IpqP6
ka0ARaUh+3onn2y5QXXA2xKq6tV8XFy/Cbx48HVkgtqhIYseZvK+EuLTHcGsW32/
/mBO6bNSvGPF5Gqb5QdO/posJGRfAuImoksqx8XbTvsh5WXTAfILbKzo1qll3ike
2MZSjfM/k36R0rqkyWKUv5V3k9dsaf4Gn773UDJ7ysX1NRxJqHaFgWQcouaZ0ue/
2h2530UyqH1eHg/Je5qn+Bjg8oXFwZrBdf2eBv3WR7/p9WsJNtNRjwr3/WmmwBgu
pxnN3YCrXEtI8JYVJcZYstLyE4sH9x9QTATlbemLGAwAJGAGWW/hHZgvUMQkX4Xz
iuPyiSwvm5ZnwCy+JXmMBfLegBRwvgoMGzyeE3cFvbbs2hlF5hKeLkJEcmDKwCkG
QdkQ9RnPyhFTJqRLP+4DSqU2Kr0f8y6RT46kqPNo0dIp4NRrHXFIoSCHa/E0M3Vg
lACpyHTjRAi8b8LATgWQCtyU2Nyk5g5wF9VhsxG0DrXmjRts8xra08CPTpKLLa+E
qalN2okHj+3bClczixwU1wbP1o9sdFtT+sSO4BwC0gEkkDWcZinFX17ZsjBrylcI
geITD46vRoJf+BQvUojvf3zGXEV1cGgX1KVRuRsFNLiMCSHL2TE9E9EKcZffh9ut
KRa61JejT74onw+zIua8mco3takeyoR6ig1e2dZ5Z6xLuHCgHI12kWE55x215B7y
JuMstp6hiIsBsmlYrwSa3U7oWNzrKb5nESzo2hw4exLGvDc5Sz8oMiAtUITpTo8D
+x56XDXOSFKbcWoH3tey8aLnIGptQ8oylHNc5mAxVa/F9zr6JMVMBeGFMelAbteH
ZIulpYagaXuixZnaS74PMPCJFW9mvUsJUwUIZtpVBD9QkRoo5mGdwPlIIhhi6pY4
8HbWlneOF8ngzsf0yRNjbJ5uiBg9qBkZkKm4sgzD1ADA+WNh4ur74uCzYkQNRkAw
cFF19kO56rCkF6UsaWQ3dZfUy9J9b5QloZWyz4T9LRhO+G5VI5ke6WEY7/c2HGQm
iewP7DoPXGBKF80jGpFbaEcIYZRCGrD5dJK/W9Wd+rlMJDuuGjT+C5GLTJuI1Zsx
FDY3B5XEv1ZMxkW6bifO5JVipW9sk0nnVKJu+cg4rpPZEnVYiZ/VJbomDwiH/219
AbIDd6JBwgj5Qg2Qk/4CNXsCzd1QI5kKJOSv2gtSbKa5g0EkjcWH6rxYSnd0BDOq
Vs4fsC6t3v+zglQgsvEockzqpNpWvzuvCNEarwp4mMXegnfCQ5+JNsx9frjjvfS3
sUOEv7YHx+k49jbhZ7r6Ra+ghh99Ar31dDT/XwqROg013v/zZLiF0uAYWS/KsU7x
w4fRsFIvnbUZXwD8k70njCfWpnbsz6z0a2Nf/7tfbu5NlEYB36KiGrs/ZgpP5SVh
RYy2VO2abcfC14KjeNwf/2OnPEAEobLKQC1wRRzm9XtIF4UJkF3WDWq4m6/Sbf1m
QF9ba9sf87Py9oWxdCzeTjXHsy71CSlpa/JCFa4n90ylQOBQZ8KGUCf5G7HeoOgY
XNX58UNSutq+P70uEtqgluhV7h8EVBjfFZ6QwEKwF3UItKMxAjB2LJvb6hleMxdk
tSka1DCJh9Cp9SW9r1nNaUO/2JU5QtPEsNzAgixjwy5/dGCrGZ71EQyPaoBNxqD6
go5zKRPiWbwF4CM2o4Q1SQDoj1ds/EIFYVOZVixQeGrbT9OxXlJDfL3oQeIcFOge
EEpmbDZEUiuJiBaNVp4c/07w+yNOKRbqLql/F0cqxviyxGn43eSuOw7/+bIF5xVY
IV2V+7ygULry5uAY6BkFolVVshsWsX4DWKzqKHRLdM1wGHnMhVhOoZ9NQ5alms7Y
R+mksd3BNty4e+87z6FMFCxUI4Fo+J/45VBwuEytCCpLbYo+buC4KyfQzWbGLZy5
66h03jlssz20KIz/muPXCSIBHMgJsPgGuSl4lbK96EAKCBWn5oFS+a39XEMUnAN/
xigw7RrUotJlaNLBlvKiBd/LamzWd7cyFGaaWJYS99BQPFqcTwupwNw1uyIma5tN
SzvFeTpu6i7Hbc56D7iNplAgJBR24yjA5bbMV9ZJxuF+kkdhJyz6nKkErQWOPa/H
fKkJ58puZjTFq2ke825CaMUfvaWzhV7UoUGds1DpEe6zs/YHrZa9C8EaTJFEYiSV
sZzF2bDMA12zKNwnFRSZ42Ek0x2Wuo/Iu+d/v/hKf1O9Nd2eZFNJb2/7U+yoXtHJ
SVi1M6duj5VhU7WhB0ydyJrcWXXGHSDYlH9rjf+K1WwT04f5wsFk6Gj5pNnG2OWo
`protect END_PROTECTED
