`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XD5xGmJ43wo9qmt65w+JVo7uKGr2E9YLOvo+pyMtMll5KYupO0QL2iMaPLXhQ1bA
gbMirXYSVMsZAtvA+EU87vqYEyLkkbIc4vdGJhIWrdp85iuEGtQZwByT8V66gOs7
aAskBLhTarmKdVj8t96wj7bOBdQGbUaw1j8b97Tux3xDFHYMfm7Vn9m8AfSZ1SrJ
YvewhOZtD+Gc2ik04hpk8MWsmFcxeN+Ubvc7TdF+umWZtlTq4g34qrTNTtvTQ5ln
5cn4yyPuNK4L7uH8mGh64zwAwbRjqDPvZZw2PjmfPMT/zt0ZyyQXDhFLdI2s5pCI
+8AsmrJxH9kBOeiRGRzzNrNvaaCsLl6XU1OR1OjOj5QSooMb9ftehyTLoZqT1AWo
F4ExLXunh6iMY5mN4ojqOoyODrsp5uHkE63jQUV6kwJZVqcCxL7uk0O68m/IfZzW
iPKRMV2vUVul5JM0UteOKvUkRxm5ZYjNrDS+ux1XZZc=
`protect END_PROTECTED
