`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GLrpYLLZhMZ31DRIlGrsYcvUpQ9wvnD6AS9xSzAW7arGEZxppuanPX/nu0lofYJ
zDxrljg73EV8K96TqVlM5pZou7JpllvpEwuCJyI2xDn6bv1J4yMw1u/PwCEJTkwe
vj93RZBI7v4bYejNPUBqd1UrNsFzv9pBtZM9yFIVYhp7vYDi0/WlbOFmQQ90U9ut
JwQqNPDAHxpiR4IH3EgulfaBQOJQXHqGCqDwUfOXUyMk+ylXY7IG56/evXJ6adGr
Sn2cMvusb4VP9FM7L3oz+gLuItiAj/6yTwpVHymoNt6CZ2jzCSxtKke2AM4oJ1/8
Q1uvcPrSPL64qeohZ1u10relkeva4jATvCx3gHw1edsmtnx3sWDCGCT8ZGP60/Mh
TzNXmc29gPpqykCTtjAzyVFgNZGPEM9/M8Jh7RfiSNQ=
`protect END_PROTECTED
