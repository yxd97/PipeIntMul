library verilog;
use verilog.vl_types.all;
entity KEEPER is
    port(
        O               : inout  vl_logic
    );
end KEEPER;
