`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1yDuVsf09KnVe/xLWsCvH5eCIL8XSdJn80fi5Ii8Ewm78C83B1E6CNO0YY1ljpy
j3a8gO9c3hWWCs6z95pS5STBQHSRxORlS1A5D0s+LrETTb1qNNI6R8nf1hwDLCQH
uQf9yf2URBJaGOY4PdjNORXGzdlAYd4w2VR/6+pl8o5QRK18DrhtmRwoJCsuBGno
I2HgmPujXkL+lGx8n9ustvqQsomNfCSNlm7Y4Gh8rqAke2rfVYMDwNSOCHdLmuDG
+GvbcZKwv1PNpfojNkwQTIQLX5YEOSLDd9pjRcAwzaM1xwEkFFGXqspBoJsC1nbN
l5jXR+iQQN/bigXSHk7eo8lVEKm+MZRTB+u+5OjcFg8Y9P2b89LeF6ijVX/hVODV
JLLacja/62TbXUKPJ+7wUqBNBqYolFmLcU8CLG3K8/IjbrRrSSCjK+mkO2TgHXQQ
r/EUt5yAwB37N66ylc46wPd9Qo3D6e4i07AhsOuH9pIdObh95ZkJawX+mfB8NvQT
k/VFyRoHxwKa4jG13255fltXzoZvWpgVEM0aYYn5TGVFk9eTQJRc84AGBYaLnvvc
Yhkjhhsb7mYuDlEvgXHFGQiPrZ5szECXOEa9+rIWREDpuwH6ZWHhZteJhHDZ7M8F
nKcamHRJcYvrLexsKoUhCISXxh4YTrWUH8gqrIvo2XQ3DbUOmnRZ41wmZwfm7h2U
YZIHA2seE4xgNZvk1oAg9vqB1zyJEskvDBm6KD+UNmD8KC7aHPmgSpHJHjbN0VSs
n1LIV+bCQBNF1NUFdG0bGQB0xlaAe4iyrG5YKBmnuI074MNNZT+CEwm61rzSpwzt
U8Isdt/rGGLS0GJIk3EoRZvnJ2ihrjhjdr9oWwcAqzQlf+uGCQ38mybjbqV/bOjR
Y5BUfJwp40Cp5ibM87Z55P6KeYUqBFWsTlM75wAI0YNivK7+eyPYiaSZKz15qJez
CBkkKmQL7N8LXvDzCdZs08IPtuvjdAvB0dFZ8B5st1rxAPmLAjU7ZZmiOC9P8dyB
5ui/w2w13OyL0D/pC2MetukeanYmncBp0gGZ+/Jmg7BEPPmJhMyoufWSSMo+PprL
1H/nCZZA91zQQsmb3caydZ9y1T7WyVp1rmy9mvkk5PP15LPwTRPVLFTq031uBx1A
OcRojg/J0o7jQCtS1aM1ygCNuzMWKTq+7UrIXcpqTJP86ni++w0vrnL0v4I/F+Ek
AdyeOzPJ//77tSTMJGMBIMQgqlL22xGqrP3u+0KuGiQElYndLil+8m8mDwoFjlQw
DivBRKlrs1SuORJKATVUPXD/WQ3yOsGimF6FIGRZhIHVbu0BFcu85RJlnvTadex8
Rs2Ytu0pnYDLdCnxd+VK6opLBGYv+g4AB5eH1xVmzXnN9eGnDemuXMTA7jW8vuej
BX7HCRtzOyt9j8JOIBH9xPd5ooxs70eRydl2CvSHsoy4mZ6X1JlUqqSK2V032LCh
UoAiavpOGEfbBNKMnX5CMAR5M46G9vDX3IaiH5ZwgNz96ldT0diHAb1dOqnW92Du
T4UruCl7UuUBbvmBQ2MDPctq2Ra+xnsT0A6mObKL1atUrpsarHCnu3Yc7aL0Gaz7
BntRd8II3QYYLz/VA76Wo4eRJ01l6vkAqC/82Cp7oTeDZJ9fPR4UpipnFwWiNJja
9uSMfK5VBklbJFXvds0EZUorZGk+NojfggOQ1yMZrroQpqDzS/RHAfqbmAmt9jX2
nwZVI3LP/VrC5oaOc/Aa5ZwYMUJzi/le5fEXNkunPS89JAMc3T6O7SUB7VaNcbmC
OyuIEp1OfCBWxq22higHWZ3C2N47b6Hz3FAng9Vn3NU/Z4N9zPU+eWznDFDuDl0U
2VqmKTI2dCbPfIbqoMEAt1ph+IzRQI7NgpWNAoe0wzuRh3AN9/p9zvNn2hEsgULl
8Jam4ENsbVW2NayG83u3l0iUuT1EkkT3xg/FuJZDi/c52utstjcZZx93zTCqnkWH
xES3FZNt9OfgXSnlCRC7THm5jSkQGa5hTzlGZPZk2ymd5Q4ufP1REMMoy7EaHhSb
GbJPb/DMbiBbFnlQ7Jk+P/9yOGWIGVZtTZT2Lu1MALrP/Kk2DR3oDGd5CRJvYeVl
Li0PcMWaGx3FZOx40bwhdEO+RyyNGeX6RCesN2f4T/u8ZaM6aF81JSO2mlLT+QCl
g0rphOQEq04NWIuQH6eFPY5QVann/TS/YlPCKzA6XrN4o+rwC9oQ/+GDkvvFNKYt
EAFpKR5okIswTSdrl32fxNXbjoDZuLLG9hrl7KSQzdZMs1IHQLgSelfKm9Y7FBsL
f4fWu85UEqtbpUH2U0yAf4/M4eZSCF/raWfapnMe0c1HFfX6+lg4MD1FvHB9JeZr
ZgTB+L+FYR36Z4S9dzrRXHD0UKc3EnekyxYO+hW/JC08R4etmMTrFqev5yRLFbKD
4WDejFrN7YCUJEetfIbUfSmYY0YXFlU5xuN1qWveTld23FWOC5GK7BxWjkWutzIK
d03mFIVAhucUVKA9mDjPzWWU5uReRtmYmOQ/yk3KbvAgWl9GRXyqXsfg/7uwmf9M
RhtWy+RZYtTHFiUQD02Tqyfh2l8vGvTFIMVXxaNzaqtQqYVePA6kEZsnmg5bw/Lj
HRo52aDtvKmJ8O1Auonhnvpvqt7QL5PPA/8AV7h6H5mT6+2+zrx8HNi4WgV0Zw10
hnDsRAdj2j3rLdwuBvqG5/YAYV77AXzCwswWu5P3rsNCsfGWhqGdc9EhNOKfjrqD
LIPWHlDFiBqG7fBm4lzPEkCeVqYs0TIV3kcI0QZm7M7YE04nHzjM/307zza46e7n
2NnRgC589q3VoQ2oAyf1+EK4Yo9XgZ5W78O9d9kIBN7p0jpE2ZN50W7tOND7d5E4
dsOFJTu3Rf7YF6e/nYhro9ur4hCKwzu5TrNNM0v7TUZbWV5dBhC7tLZbLAxPGcPl
t4J2vnSoC8/gnXa/HsvK8EAoIIHmu86RPylRUAWdWuybUL61aTeX0uDBBMNiVzBm
yVsFdpxO7exqVQCDyxchl8SBMaEAjv6AvlQX+iTz2h6ogZRL7HiYQIhQn96R3Pv+
0srAkPCdA6mhdKeXSusdoBKWvfM5ppmpCZi9Zg431LaqUvXwAiD/7VCMfnWlMArg
YApOFj5H4u/wBo4IRL5P6A3tAJSS5+ub/lch4tNn3hL8fQRE1tqZkT8Uu068DF/k
Fly8etGx+dynpCvzDS/Jd+lCBL9j6MnP7cBzGXqkmUgrfWCyO4Gsc3Y24CRIrzir
ZYIZVvwLBFD9Wu1IGkZCFRFN5DnIxNY3rF7ZSmZnsfq/eq1pXTRse/BH6S7wBK9v
ra35UF0buF7cYiXbhknGVkmnyIK/LElC+JnBW+R86U1YZWVLOz5oZ2EQlrXma+gR
GUHqcqGK/xedlqb2HowEZnEnb6jIn+BkjbOlvnwcxzYRHonALvpTO0nQvs3le50N
UKsVfdJuHNk/VxjsNKkSY4pTXthcnTNGOfZs+I7k3T+uKlmDX22Z/sKU59Hpz3TM
Rj7NY+bJkzkHC8FTcRzkT5epKJlMj7sT416VzsmlSTaN5ojzpNdkKTQegtb4xbiM
mJuBDCuPf86T43Y7zIAh66HRpwq6v8leLw8nxqxShn/yXzeyzN+idEcWjYp6i0fz
0npEi05ro0YETIXa6870KQ==
`protect END_PROTECTED
