`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMt3v6umH7Si4ddI458qK2Cg8pk+OMkSBOS1YIpMlmaCaO2Hi5nLmkie4TT5ROuQ
lgIBtXDXnC3o30WuvmgTDSqATquyk0cbNBTkpc9r2vSNx3nvK6PZ2Om4BAT5FR6P
kI8P15/FxobAOUkbHUdCsWspf0MVIkkMPgjqo4UYB7jJvkQM5DmGkSottYWJaJOq
HjLEObEXC+gzIP6K3EamF37QVcIZ6pME9tIqD3S1UbQjLudSVUiXcyyW0aOOPvIM
tEzE/87begtgV4Kzp4XoNA==
`protect END_PROTECTED
