`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJJpq0XRwPobfwuupT7Ux3YKhPLLt/p+BgYefcwTY/biBoy16SZpcRSHC/r4QJDA
ZyKw3TaAgrHoRFcfFaDv8V1YEMUgKznAQhBCopv2GZedXhZKE6ThZTr4NalNiuit
G4K7yYWktyfZ2rDOt538BZtC64DF9ec/OLoGNIH7aR5jxE2Oj9evXzTUDNAc5NtU
6cqYytoNlEOydgxCo6bJ1pU2xBUeRS3WAsnmjguHCwbh3/tOShEPqh8+C+3afWVL
AmU5Ufz+juRwgNExAKvyORvBS00SrP3ylRUyW67Fwbs80EIpPcu8BIn7LOj/8mQE
s1CsNgHDX7iqULJfdaXNEqwyVSV0IhHDmbEQ8s99pGpH3KogjK0VsjtA0IiQ3nw9
xMGFlFlTNKdD6LB+OjSkSUFZzLQglHObM06pra0Jl64XwlWMaTLIRCI67RmPop41
vHQab24yEkwxs94kJelgW03oA1zvV5lgZSS8zAyqQUIlBD53KYggctexltPyOSiS
SHpUd5LiIQvTROqL/C5tnnSbQODG131IoRWqgkhZU2csmRtI6/uSOqDMQn1mwVKk
9npzLYN0gqntpT3NuoPQqwl/pTBwHiqJGK52tKclxQVZRu488dUDSGGbWgi7MCrd
jLmqZfI0OKZeXI+f9qPdX+HWgh3+Boqo1qC/JDVuQhKTWEfxY5+6hp02mVDv6qoD
rIFM88WhIXwmlZkpItrI+h/UPkSHJTAuFpaFJF34mOX7XBnDBckeKMmoNAD7RzAH
VdtDu2gHpN0oUwdwZzoI9Q==
`protect END_PROTECTED
