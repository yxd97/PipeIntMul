`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gYG4k4DROHgcipchnueKNV1fNSEKw1EzjAt3JpB+naFY96RdEEbtQDmRQxOxUdtb
1P/LF4zzgGiy1lmW+gwToKdDgtHoSb21T8jH0u5f6+oN5eYVbnKUVkyw2wJANqYC
W6o42hilvMhJkaD76urbGZ5BfhrBIGxsLQwvyShglUXM6fL/9MTiBdl4ReL8CZ7N
vuaesoNQSqWvv8GaOviSLx4278vaUD9e6SujfexfpCJUnzGHN+jlfOs19kocgc2J
hiCf5IIxN9EOUsfY+n4e0Ys/zjrT4dWnJsiH4ihBKqZ/V0JXBAL0T2Q4z0Q3APOy
3aMfGVR+pJpRhww9Px6zDVHj1nL0bi/IE4Tgz6TqDXjtZuUs7lBlps1/lrS0ieD7
DFgdLrL169L7cpzznlVoVekwVCoHwntPTFiREQPUtCphWIMyrDvg5QnYgcAtZfSp
hjQNoX4wVbcQd10x/BvyQSVihw1CjWsJeei0oz0lclGVx59dYmd5jfMKQXFrDQQ6
KpcMzkm4IRAih5gQLmEv8xAD4BN8Jm4L4uAL3KZxB17dT37qSrAI6NhBnURdRwzv
smd0lfEuEwEamUYYvxjDGh3Qk9bc+uiZsyUsRQhFHd4gOdrQAcxm1oB6ESEHQnfG
Dcm3A+YDJ/kHAQMWb8E8fORCaQyX6ZRz6U/UFUXJ7/gpVbPiuaBkjwixbFGC+lEG
TmjTsoUevAniG2BkOwSkPunf1xFpNdB27yy8ajKDkodxv2xBmLYfKAlpuxqGJetq
Ko3xwvGBdAQ5aGG3PPZOmUmEM+Vm1Fn4reM1kJKTR63MEksmC1vdvveS7C4by3v0
htEjygkVlLNHsp9tnfbYepC5bewQ0pXfN9RlULnIzMGRsquUABxTw492Yi03V3Bx
mftfkw+9PYE+u2I41gxjBRzxh+OE7qx6aVvMclDavhtpM6Vx+bISyTWu2oCcVPcK
CMMyEiwz/9dxBgokf+FqIdPTkHUyk+SEea1D6raXnSamgkh3sKmDCBon4pkIafaT
+ZY8wWz/UdptY7RQy87zMhxkoiR0S8R9c7n84UZ03ebgauBBRHjEh1tkmCa9o8a0
JI0wnPmnWNw339r103fx23RXEL3wdJH0G2ggcfnw9yyu3HTc9/c6YQ/edFXBbZIA
1nCUuUQpJiyA6j2CNaY4ffWthnwAZJCX9OyDkR7+pRho7Oo+zmVd/mF6gmjusHJ3
MNEmJWIoMjZ5y7WF7x+yql2j3ySjr40QQR3HylEHgXB5aIpDekHoJJF9tt1Xdxi4
g27lMXCtlHZP49WSTnsZPhzRO+YE6yao0zWxO7tiN36Kruu9zQ4EsjEkP7o5SktA
qJ31lr6lSfnj/moRP+r9TPQq3z3ItWdKzLMlOaUbqikg4HDVJM2wDxVQukAlHIyf
AHQcs2FAwSXzRJyHX8tulbCCrndLHTMnwW729nSg+jRITudADNyHOvFW9YpBx+Dx
wvcKfYmNbKCdxIsi7CpkJLen300mVBl59Oei9yVz4fnyIdW53ImU697Saa7pYxq7
OYY1ETZ/W5tHGh5+fRnhiolns7g1UjR5eVcb3Of4S/aheNudzNtNfDZKzWuMP9KV
djYw8VAyttQYVClSfEFw7KyrfSN5ZA0sEyV6zb4Q/3jV6qqVpiwfbJ8GLhqZWuMY
mDaBmEJa5ubQXiSGZKfupo+nze68igGSHRgI7IRMRsL2lMIf+XcoLa73O1hkfEZ/
NNKZEnh42i7i5E0if75BdhaVJjIk4EprFmqAvaf4mCCLt7vrWiEkSw6gOSTUBN5e
hvWQ5CMavkPP01JjKbDI4miBI8sFmLL1rd9/ewtbG2JGo0oE+EjiDpfICftGg1qF
9aKiag3r2UfBvqG56NiX7dj3DHnniD+ulGEqbNidr/50Yy4bxrLm57rFptT5Ig6x
8jFKMyhjq/IhcAKneIhEySFl5OE34GSwVdqQ2ylqIv4BPIocd+Rch6SJo1EXdphS
FVZ1HxCrkdEncFOpJXvskUNTeNZH6pdlWMsjTRKZ7wZDW81A7OCOSSzVfOlFnX2Y
RhZI5MdV7tMj5zxu+ey0R8rZ4ByVHdUwwk3L3dYGTIJLvDH80vOPgsawiLEA7f7M
Tc3LjK0y6OAmtNC+JLKywPiX1UU6D332fXPq2mzdDjY8RkvPt6kCfRe4/DtJdegD
f3aXtMEPwrWfDPAz5zBzJwY4xCB0tzUaTlsQD1Ty+yUhS95s+MrlGJxtdGei1RPF
kecuSLPmqWDmv/OfMTVEOYOv++2EZBgxpPcfklR/lPe8tM+M4EqTixg96MLUZHB1
e/osmri2otXueLVdBy5Q4m8KKftKTHvdphCo4Kyi77ziVXxx4iPTMiVCFnpTsTsx
lwgcHWo4nPi/G9aRnTEtPWxDLrtdeAlgnYjtrJeYC44ahZHdigF0Xt/BOdKyCvAf
TaLAnbhhCuUgXzTqjKgc/U9xop+0VylndsMLjUTOD7eqY4dV9OIiRByBYsnA3oFt
JscO8nSEvPP3sziiJpW1PVcf64/QpOz1uVDrEOZC0ENZCAuHoIiKNed4gZbpjsoD
oeyWiK/FJTCaaY13xNMkxAMy+2CoHyaXLk0NjVx1goWoncavVMN4VKmKBApYN53W
QQgUAAkWRH08t+3BK2jZGGoV9J/tOQjWZ3ffUX4c1A0MEzfeq6mgqniZWIK/+0vD
LwmiMV2pHrAPkZcxKh2dTsVqhBdsirjVvmEmMGAlYzToyilI243liwOVKLKuVEH6
0lIrkTKKTvJ3E8RxinLIBj2zmAePW7k+5ce1prLmU0WeGsexui3uD20HEpBKluUw
DAOoTeJCO5bif3n8QZ60lc9i918iXbwCEniq+vOPUEI=
`protect END_PROTECTED
