`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQtqW2XIXJ5fGJH35yEjvGl63anRAJgIaKGi3swxnQ7pOPTvXPWYyQVw+HvhlmGG
fTcUp4Pu8kluRFFcErELXJkE9w27lOP3nwVAh9dwWINI+S+IxBgEHo27Lnyo4mHc
/wSfruGHlwlYfxklJHvIjwBj1A+bZUOG8NgQQVC0BZhWIZa+RcqQJnCom4AX4x6v
hMfMFJXiCXRjCPj3OaWKVl2m20Mn7MLau740Lt9vfz9iHOUIPKm8MWrEsWBe4ZzV
5r+0WOfbk0R8tTVfCzywmVcKm9iTyB49QzV5Ef6Pqu/BNpBC+wZlE+mbqNH2ufxk
MizWbrf/Du8+p9wy+H8izeIftwhSZkCDS03+cV4AnrMlXwSHwIU++2v1i2Vj/T7j
yiHBxs+nClNCRxOqfMILjPuLbExf2IakRjcTBuWWW76xQSX8iUPk9CzOJkSEKAvn
BMlm8U4oTpqrfy/U+BU0gROJnviLL6kbhacKFW12G0lfeCCwyJlSq4jZEoebh2pg
HLgBgYzYwZId6xt3xVNYj7Ffd96qav1m40T4J6A1AaPQrGXzdFupqM7LAqW1GKlo
Yw33H7AbtfStPaNedGqSJpOg8Eta6k1aRHz+26NEG2LPz8r3MwxmBdTuCQXPJ9QI
YiA23zjGBUkKuVBc19kZxCkqskWH5bFANhugbOxMw8Lv/zBfeJ2kDnnSD0I7gjNT
OAmQjW0MVgQF1VOzf/9ZIh3aVV/HSFG5qebfZRXK734oG1Ous2HVVMkQl7eaYiHp
TnOWqO86rAV1tSkFu54PqWn9cJ8VAQbAz04I2C3FK7RGS3k0jXEDVlr4+FLifEPn
48hOhWblj8OBLlqT1FzW5bQpLCXtCfmDowbJGWAR/0RFo46g1scH9o3Ww+FIfPne
Jvs7Yk9//Mccm1pN0LKFkflrPFVCzf1BufocU5nfdCkL162Z8Oa/agbcJ9iHXWyW
nrpC1AxwzeG4gFfp2UVV7k+BCNw7m6SZmxt8MoCvJOjDTKqs1I+EuDbxwX9S6Z6H
4gB+2L6lKPS+ccUSWcTNqQdrP/oYKCTXSk2wG3dJRN4=
`protect END_PROTECTED
