`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/kGnEUm+/mRIPw+VB/7I+2SBZ1wNVaIlwQhteQBEbr9c55CyxKcBpNVfyuBMQe9B
eAKGFuUFHy3VrfJncdxRGJNhk1Kq6jHeRH9syOn1474wJ9PyaWQrN58dQ3DtwSbs
mcyqKDf9KmL+/SnB1J6buRdIZMrgmV64GxAGnn2HFt/WcEhX9k8c4YXaI6/O+Whh
6xEPO/CNP7mtbt4p3NcXf+zcG7n5j/h2ZecDKx9SpVW5mD6HeEmAKo5We5CiCESH
YgyhIEz9XuG54HNKEo+nyRJaY2us0UqvPB/VB3Yb3zGPezlNqPV73y+7YL5CjaYF
SNJUzjUJezrPZhBuUHwGlP5xgPJBXyWA9GgG7/BC9r6uY51ZpIUbhwkRRNSQdsjq
XyVNLtR6o8jQjDMDxOagoOv+/jm3csBLzR4Wsm6hWWJTaRtHm/KFbUht9KeU9Q2s
b5nyAOElE4JBELuX3PReImsha/q/QcfjGOkZ0/dgH+Op2Lp+meSX08/cQdTR0TYd
FSiMC+gKo/1TcaA9eCYPoFHMWILnJiG2soss6B1LqyDBe/nFjjjj6orseDdbN/h+
K/qlolr1JGKGlNOiYQa853MtWkGP5D13z6mpKgiWRBxhyJWukNIojwgvE3xFkYLr
MmGSLgWoMHWdItd7Ry+Ceg==
`protect END_PROTECTED
