`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EUx9A9gf8tR/UNOlJji6k+kFpHN/pkoUSrmDZTkWUsIPnHAKbidjj5/FwaslYdOZ
sniUKBPeuW23p26AkzJIstg/jH6rISWCDMPoi1WohU2hg3oymC85EPme4qMqZ1Ix
WDmct9IUWbP8+/wS0kMfA1/Vwf57mPzKlvPirxOQg2ygQ5OtkUtgVhKkyWu8qI/h
RslSIr14ASg+js5pH3hIKbPxzX/f6qA72koSPXku80haGPCiyldOF8neEa3WwO+I
uY2bbKcPzmZQXyE+Hc9kR1SI3nEhbBCRFPx2DyDW0h98i0BAHvT9BC1sNQ/ZvWMm
4Agu/b/jvwjKID2wFiQukn8pDu9bKGCRIcdBn9+AJqO/fOqmgqZeSWCGa0CZ8tud
pev3fTkfAaihEe/7w8x1sTlidHSjUQokMkGlo2oXAphUI4hPzzwseODs1HkbLl8U
E1hkWV2LZrS8h/L5ul96ThdTHASD2VamBgmA8kTkxw8o76ZaV39iOr0uMeMSZ43x
IRrewpp5LN1GzqLswrPjVCwZlBOYpsMgA4h30koL4JsLkY+FZRnNN0X0rboVR451
ONdla+Ob5kUGEtxi/TWGPWYvxNz0CyXWG5pXJ8aMZU+seZi2OM9WRgoDzrX4ZYv7
CpNwB9qa1kXffghXbMrJ9gazhKGtv3oedFqZfWe0SU+GWuX0dWLVfzdxlXpsu5ef
iFq7dQb0hVwZ+Ymh0bhGtDCHKC2Tgng75sn5bDBJorxAPP+smRfDdMVTH+xK72EO
vHVfS6UHOtEZq93ecxBohjiOChUvDz4R+pFXj91133HUhTZJfYF6fmSJEVBxlo/m
YgKZFbja56Uw1R+kXaxyTjDz4oY15kMms+zlNb9ZfdPdSoadkOjnqN8BZW66rwvP
x8nt1doJVP3fKqUxHHnd8swDxd4jg/KnIoOapQpIwdIFLJM31ErOV9VdqJYyMl0p
T4qhDs4VobanLbJbo3xGfSf2vQYFCuruI8fn8v/qYqaXhJ1j3BjgJFWR+DZy34uk
orC/gdZ1uyw8IjzZW6gVlX+aiH/DyHB29V16WMkDv3T9fQouWox9JR6c3Qe36Xuu
`protect END_PROTECTED
