`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
imSCZ52UKzMnaHJRr9A3PikMVhkuzlXcivhFpvsb4n7/ypXm52/uraHB3M/YLa8w
a/Sk4o/Okx1F4je8W0QrROQjbKHMLLHfHxLs9n0UgyWnSzB648kFD+7wC2nQ/pFV
YORjyGTXpWBqRhS9k69JfuZLhvBT3QJJXqMfCWI9ZYSvGtHAnp7QWMMfiReQ95w7
+f8uJ5AkE5ZTUE6nF5svogF718tHq2MhBjih6FRHlL+49pLc3XkDW5Im/9hfIJfD
ONoWo1reP4v8L1OMiYz+BtMh6hYNu1gagNtvGW6ExxgP2aqC4Xi4iajoebfplEib
CRI71z9wzZPV8sQNY+U6eZunfEpXOBQMmt89Lj5+SnOPwq+iyD27vmO55t7G1VYW
7UKNoFgNDImADUqcMNfWu+OVQq4zcqft96Q89klTSW+SYGnShzWmjzxZpHaEmBl/
/snvwrAVKY1UZBkmTqcseR2Irna0ls2i/h29Klqs0x4D0amF1m4JyOdzNthZqYFE
JietXDKkP0s9I3sj3frv4hTrZc69YWCdQnVT8P+Ltks8lFP2oXrqZ6CkvqDSeOAz
4/MPixVMlMMcFTKPCg7Xx3icQ+DdJKsbyDl6a/De9ITQ6vFzXqt9M0rZOEDFpVPc
DEwAjaoWVskan5k/oBnvlAheVeP6YpBAgrCaRsjL4BH8JT0ogWdyw/t2lY3mvEjT
FcqYyGxff+Aatyl03cV6JLeNvWtPlk1iP8lz9bsy5mc6R29gKA/VKDatalJlFvet
NSvGJ54pMyDlzxahTCdMf2PByQaNAgtr0R/SGQ1+Lb2PNtOeVVRIV9XrRA1CWWaN
3zY6t/SaXxPMtyF60QgBiel0atGtes66enY6RKBRXu1joBkoITS71sxgftVKklk7
/0UyUca+ZSPaWhlUdEHrxEgUH96Xg7D+AxaFr2pH85c8EYTD7fdZDU7PwYdxG5NQ
MdR3PLwcO1VtlLqmiU69S7Bzcc2nQZPvqdWNxTBo1vvfhJ73bn/24ntPoVXv5SCs
A0rYQoE4A5TeCPJYAVQW73/ar926ur0Ownjl0cctFrrlPICWqP5HUp8oItuU6KWx
1X4hXMnKDsqypw/Y4x5zYAAr8Zg55hTp5zd8WJshAvKORP2NJ+JfBLC9PAGNzlwW
531VoiuaFpVw5kyjnRJ3XVdflYW9uxztJoeHc3JAWsxPbxQ6xTjDJGpBJpIkH6Uz
kysqnmOlfMxGRx1lNzPXp/l06RfTBKRjHrf2Gv38yyZHLQMyCVdTyHsbR4HNm3EC
Glrv7PjqaWVfAWbZjFfUa71qn5NT1ZS0W7ydkEp4bdBDuXhYgL5+7paZj1YJn2ia
d2J5tbIe10TqbNyNWAzbeUAauAZ4NI4p94z0hduGq7DhGmOkWkGhsDrk0NY7upr1
o5eMafoC6LT8IBaRoaq5XTyyvffdANcBkXiaVqAFogXINrCJqs+gDI+gYwCv3t2J
R7hW72VcKygrNq46mm/qp9dA11mIKab/sIsU/+FD64idYzceFAeGvpysVvTbLfRn
c5OsdeRHqiV1Ij/nibGWLzhRsiYIuTUR5pkCP5bUQuuzzjfEAvZH1ghpmJIJRDXm
yuZQoXv1bPlkZbxkgBpsYC8qxU9S7576aPmIjqs0SUAFxu52mKB8TpFTgihRmhwZ
9Gy7wogROR++bAJqMing8xWv98sJhhIaiCPbfvQltzvV9JL/Erri0kilhttXO+x+
PROQAwm2WHdGqlSWZpgB2geRoeds2lMmcNX6XuLfqsXu8PQzaKdIiL0taPComyBJ
21vaahpCDEH+KPyeDcfInbk+lDAl1tf3QN4G2f6mJrXaNZQbIpF4UW92GtXDYmdF
02R1BV2YoLriMb6rPt7snYqyz53jNRszxmni/0k2GHGC/N2M3/yhY535HiiYLGlT
lscTbu6ECnrfo3IyPIVp840oXQLmE7KC1jgDbffCH4EGn+z5Gb0bvlcW6yx1U4ol
0r9p1N65TWnD0fiMOyw9Rsz15jLJ1MbZAGhTPaVoK/Je553QhQAn4dH14h5ZCvWn
BNNCrAYtrK+8+WWW8+auh4vuBG0UCaLSMiisukfTcZiANXDRxbLocPXZz4jiKgLw
MQAY7143P36ArxgYeM9ZQxvk8WYKmxQO5jiwtnsmzVEBUCBDTQliZ1gEjmnoVCAd
kMZeptkY0Hd3s5KY0ayWKvlT23Pzx79ftCjLmSs38tGBUAITLF/2yJhrWykfjGHN
DGDVmZDalOEQBl/2SQdzlSKKNPeRcduppq+hzTj1k3/SCyX7lM5EOVtRKhrTAQvO
CqHEB3MCJSI5vBmrvVDZo0tDYeT6D0Ifh4dCh3+UUgFc8OhB/am6vR/73q4TkwCh
nLb5YMzeA3dgfrYGB9WMEXrAFc9RJMwYn9NnlEb5MBXX+92sQjpf3kkzKBOMeGw0
uIzz1A5tu4TrQZKzr61p4koLstFlQKIbTYOyHSwuDEJgCdMIhHRb/bKSgzUfpAWg
cwnGTzb+npT8KGCBcRMPkuipej6Q53nUoxQS5xqwVQFhf2j8HpO9YYvl60c8+hvB
bOAksWNs7i19u2cXLCSORFzGDByD8F0vO3J5ylfWoJDYy67rlWPTqIJM0DqbFuNn
XllWQwVyQaupB6bj/a2GX9Xs2XPhnFEa6G39PU0PVTIvjtp8f9LC+r8WB1Iljj1m
JKIm06Vtbg2DCJHPshZovzMJ/+aq6QHsXz0f1hayzkPwU3MCUJygNbjSjwBZxwm5
pEmQyht0Y83KXta33XT7reaqO9plAK4xJ0aM/4B/neZXZOQvKjTN+MbPowfjiTWw
/018mGsOkdJskPD9Fl5C78nATLNs88x0oqYtSNpZhFFwnAX6vOm40LhzG3wN7WAM
G4Eara4RGuygb5PaD08lNz8oeD45ajG7+zvQSIpmlXelKNPhMdqzstSx8MM4QH9S
mO1A4MFeNrTcWqCdeXzGrRKVrS7ksn+axWhzUkr+qi6ABpPy5s0O8W31soV8s53j
sf9+Wss1pVZmmAM4Wi5JiFc7JGrFMfa9TBr+dJ4oL5J/iYEm6P0RZ6QIwbEEbrUy
4nNzwc3343OOvQ9QCWL3TMJS3NbKbcy13jr01QVJIHj5JdqYIRDoirbTF8wjLlKS
nY8tIByqQXytQX6eWPuy0LoM4bViZQQyeQcR7zAwsE6JGf4YDuAX4zwl4oyCoNAf
yaptNdh6hmnz26BQ4PwLlWdV/twbdnAkS+XYByJkje5sYDuDo2YW7vfyBNCeX6iN
P/MzaTpb4p3s2qYyogxMzb/GoTnjRnDudEOi7oRSSTiPOdWQ/Na0WvjQKS6lG9VG
c289mY9yLjJQ+mdE2lK+T0Vl2Fd26LlT0tEf2N5X6P7ztC8uBJtb0oqAYVfKMBW7
1QvGjrTnoEvSgpj+RV8jyyIjPlVHKnXuKDxeCht7s1+ZaQho0lj56bETY/mEzgMU
cdJPN2iuZoHHPBXBWxuYQVWdjkYwyPMZUm+ErJpL0lbDuolyNfHMoMnJOtDbTJep
wXpjyJojRTad4aH86SU0Io9dm0PEDRkXIJM/PDKG244FHm8lWYJxrQZbeDHwD1AL
puLE1RYGT2zYQWJh2w6oKIVPq7RzUvQ59xgpUXJPUcWJuLB4MXhbjqv+5s+VLXj0
j3s8zQm0EeSjkzjSxWEWdFduZ2OazoUDQNlTcU5TV45+dxs2OxYNvp2XFtiwaM5Z
PeoXhfcWAoEsP7h5beXqgS14gl4FvKyoEnKhUbPAObHtZhhk2cSr8pQdSwLFsWqQ
YVw/rjMOi62bwZoV4rlGIHiKs77qbYYeSTEchExVoFAxvUXyV1QvSH3Oudpd+2Qd
B7x7BBcx+yUTABY8fAPExbAClbMSaCgml3RXDLGwibNKARJGMGpccfOcQcW1/Uly
XKEQ4hkssoP+oTU9f1F/17syZnlbrGc2MN66p5OQkyzai6b8lZzpSY0FuiI5h+LK
X6OGbkliwhjVe5dPWoOSeZtsebIp2nHb1e/9aMwjXj2Tm/PdqUEGpgPC9T5hqetw
gxev3JgAy9pwvHKnn/R4XLJ7fkfY8PZFzvcXsgo2Ym+Fljx3r78XbUK4vx3E5kgR
qfrKTR4rJ0h6b9uAzwzY5pjkjRHFVahPTkOatIM882Env35NKVczta2mV8kLdxwF
8MBVDux6dJ7+BAVM1i/THr4xLraaN1UGIdJKtqQ0tE2S+DMyXYezV2+j9s8b5hqg
ff2RRL9WacnPZcWgECS5RLPDRkO5nXaRK+D/xH1AIV5koPeY3QjX39paT1/ue42g
NxnHJ7ZLEpdejLuQeVn3/lPsHJgGtrU80rX23QDgCLmEW3YMqaYpZnWLne427vMi
8DWmPBltzeBdBd6cEZMLnf7nQ2bbg9L1w8l4WJwfGTDs6L5CIZ0nCUlL7LZNgkLz
kopVdqId1bkl4pLeUMRa9NLVKucS5oZuA7UeQjFpIynR3SwPAHs6SPHb+Wyhe1kg
n06bVA5dI+e0ISUmHQxbkwXiioo5YybYtrHCPwhVm8LaiRq7wXpI0DwBzD3S4VxH
FXH8iFRZD7/BuVk2O2dNEvZayP522/L9nR5zr2UANWQ69IFvGS0g0J8bdc1iDAwl
71GNDhlA114N8hG25rj52/QrsuCvv6ouUNY2fZ9GRf/TaaEO9rZnZgFa/m6ly2iP
zNgl/GsH3b1DUnGlDP3XYYgA4NqDxorkldKKGtECR2EAj+h/EadXku6CtusPz+6B
pRP6rDu7qoA/CpFA5a87uGZdczxEkhmkGiKVFamZaAEIsASB93R1JX6j3a9XhVoP
OpVX20fSGmy6ihGyaueNcSMf+hrJXlnJznNsYV4fdMJ1k1vFTGGKuRCCoFu/9Cp+
HvUTMUy4TBZD6ohc5nD+NkAEFKIkZWNzNxzSOJh5D37ZD5nL83a0ZRxtuTbKaeME
XXV8DISTB6q4akWZB4/BV1Otxmq1ZyT9U0WGi+Jsb5H8uVAsHSagTtDP7SglUYoS
JFMOlIoLbmghxnesrJZymWQPcwTj6LxR38lgjOF11JyVxgGK/PkJ28ec7QVQJpFr
d9rSO8C8E4keRaLSINvg0kMa0QSTLqiRdLqkW5Dn3HRE62Ebm4owitvKAt5JpLzT
dG1ogU3Ax/gF6Uv/lrno7lGQbtSX3buWIA3CpwhwuJy8TLqcyEkOFPKDbeqzAFyw
+wVZBsbHxR6d0ZnK5BUnT+NS878BKBRiiRZqUc6cxymjLZJo2zh4Zqo+uMF1jom1
6O5JELcRQ9gMtCWrnxx5s5B3WX79cNYJG4QkN/ekYedviU/jablfJB/2aMd+snXg
cZxUTUt/aqhbg5E0Rk4QVJoCrCmtEhgGkFGm2umq6AwjL7pBpxdCeV5I7w/l+meR
4t3bP9VPdTEAe+p048XPeXz0A74a7IbtT8Zl57xbESJYcMmVGqyDCQcQEYBTLLhv
P3bH9SsXmjZOdN3/j02pu/P0lFd8vO6fCGwN6j0rOI1R+4U+bEmB4W+Ul6BES8xe
8vj+yGjyls5Lp5JFY7FULhC/u40Tg0eN7dwSaXoG3FpwFrk7+rS+l4Dhewt5c7vn
+HsZ+4pqoe7c7W9A/Q1WbFAOKsUd/ZDvh2vyt9D+CF+/AgdgkFeBN8Fak0DTV1vz
uFxYy190h0WOHzvFJ3+iQTtSK3Kfh4/4X3DqcjA4wsWvLEuGA0xbyE1TcLT+b2Jv
mjHNJvzCX3P+OeHOzz0dFWUzaSYaC4JP289NeYwAz9AacB6+r1WBCzklOITO0olh
psVTLymNdLhRQyru8pm6X31FQyYnAc0WJ97cwDNjYi8qbVQVIS/i/dcj14o9TPhM
4Bfly3Prq+NhzI6KuyWdhseYvuSu4iVjbkzNFS3SupVWHFzOaG9Bogg3mpjrAbvR
Cl+jjxETVa+Ii7551yzLSFXZECdm76dQFgh0TBFwybHd0x0WJx6ZfsOlD6M/4M6D
ZL4ZzzUTfY06p1Gs8poUbtAKwh4ZnueUCqEu3sd+12ORs5j5Eba1t1BxMx/mQnZZ
KULYBslxVHXkr4+fgmfcVwivwS+v7/busZ6hCaMHndJ1A+G42LYhF3nwDy5EjLOJ
DFrfY/tiRQXfC7VuVIPgC46AMqO949vzScW8uqXFOFjhEtloUCg8nqLKWS2HlSm/
RA7i8eRQ0qLZ+ummkWOpsFqgR2R09WqvRMgNEIGUG6ObIXq7LW9sIcdjoi7srhrs
vBTRzQPVzccaSuMzTyvF9y9mUo6ZJEhNVY4dHl3DlZJhfIzvgR0ALgp9QcXBT3Gs
AdhtXCvpJRZ3wD1zG3KpY7Gvx8vtRvJJZoMgRdFrBXQpBsRgCYCkQWg0Xvs0SIvh
wU3kEsV8G/COCKPqxnTITYqx8UURuN9jlpe53E9FttdRrkCkpEvfPgV7wT92cq5Z
ikvIk+oLm+vjNdbYzZhw4q4gwIsb5UvfWEvUnipIHWnUHsxwJL0SAZYyJ6RBqJpo
P8SOa/bk0MY6XTKaGaU1leqdPznW91j7REIOTBAVEjsm6XmIMd77YcJt2QuShBoL
7oyjDk6xRW2ifHT0hsM7eyUwRpC9EBZ9VV9GnF6eDLOZo+ja3Usw9I72MqYUGzHk
WCGktDXhXqynZtwklkGk1LH6XWIqupiv8HnSihn0O50ieKzvvfWQ8ZkOMR19HVO3
bBDgtWXPkPpYnalTuZTurNa85KXC0HTkjr9rohbCUblZ9xx8+bpyzXAwOxQ2eIyQ
l28vywohT3zyTh1oJldCDDFswRRYCrZyFbhhvY8U2H6y5RHp1o9IOPNUXsftJGGO
L2N/SAvwapdcA8su6wVEhKpxwwJW7haZPoJ5yWHOrxDUiALLGrT6IY4KfxHIQBVD
Fprp1vD/b1dJ1LKTKofOTV/DiBy4d0VU4SnKSLA6GtYWvTFBikDT5QPFmOK6YRMP
rAcdKZcsppIG35cmVhYkC71LvV1oU5acVkngbGrsFRiQuvTQdq96U09CqOwcI+yW
xBqp8IydItrdhOAAliRRfPjwgk3Rmks/tO9dcuIjtmAA/4vF0ez0KVGdEx4M+9Qq
QUU/uXROpY+juwqfLt5x5qneoXgo57F8PbzTDyJOokvxJmMNK3uQmq674jGLrNf3
kyvneMispOv5vQi5dEeZhTHQ6qA0NkQgRsjfm/yh0E/hfZWeJKFwLR8r4J36cQCo
IIvaseXjHS4HFkOyYsH/SbBJbs+whuOcvZU2Yg+GmZEDpj2xlLZTKImvjeIzF2bs
6PgZpTpju8FajzLRY6CtZoXf3JigIEy9RLi4HI9mVuNUB9IPtnIWfRVo8xOd8PSc
cdVPDM4eNbwaF4vxZx+ujl1XT5y9AVd6EmfUlht0JO8XUQ+aoq2Uu6ZiA+T9e5u/
pkd+ocQ7S9HIlXp7sjHdBpQ3QmX4c8NA8wJ1KKrFRzIx9OQJ2xIa0MeaYVKq6tBh
zngiNfs/iyOJ5WiFhUwBIOED5mFwYFYiV7EMKDyPjAsRAB8TOg6cSuif+aMooB6z
Bfm0S9gjcL0i8IrVROnwcRw6GMRuCGjc55vHCVF31YkhXGXt/leutNpmLNflrqwo
ePiYUKyxmv9m1rk4D1nkxkINd2ThN5OkT/nNE++hQVrGCRStSAWdvhZY78EsJF/C
xNJxpRh4miCKBel9GMJ1OZ/CZDvvBOUFgc4o6S1Sn0mxnrUc/o0cVtCljGyNVTOc
rlt25CsVUKDwr7gqojed9L1CQ73uAyDEqaUJjduKATY+Q/pNmoeUrCeiaQRBw8lQ
QqKwL6oFxwrhLOT0z6Pn4Nt3uo1Sb0sM4mM7xNcriVMdatYIUsrzZDBqugghHpTE
r1fT6qEDViQmKeAM13uohT22Hx9J8gznpaykf/82W74JUQepZQbFl0UswUvM+G4T
Dr8ORL7IotPOiY0REse2gf1UkiBloALbXtOT4M/kGzMBX0jNfD24yjPWkoc3W5KC
T62DXeSZJxC7Xs17V/VJ/6AAy/TCh7kf5Wov5UgGRV+ukANpp1JCoWMug++Ljbhm
mHbPQ/GOZu8sTBm+FYNC5YvKJto7Fgrta+E8O0Dkm0FtL0yrf8S7OjAEHaJXZipd
5FcPDyTnAoarl/48tLjzmPK1V+mwqTYY4EJDiouQOSa1KYaUe5wRPQVQc1Zqgrpk
MbI1DnseWLQYauUIVWThTFGK0pzAMnjyDpYBz5phi/E697SCCJ8kxGSSE7vmUOOF
JRp7Rd8uUd36V2eWehFJ7VDJN+SW1Aq99bgP6lPSY9NaqcBDZzfu0qsa+Cwxmthn
+m8yicDBFBf5shtthKznshRNUuERZSfO6vSzbUa1pfbCWz1Pidn/ANu2mcN64mjV
2EU8hnb6FsaUidnbeXsHfXW48I9lXShrHuhNuG7TomOFm8sHXMkZOK53Y16QmFHR
EBSwDOd+FVJ3asXj0D5MeDCGL7/BJpIsgkjdRS0jPRQOHNHc7Sq3U8e6/1PY+WmK
OsO9alvYLufJdXT5kq/kakoxbh7oZ8Zcrn7bDqazKT+fhDDy8Fu/ZKgXuW25gfTP
uzfNGyUCm0XOYgtvN0V2qmAQy5AJ4UNQArNTeJVqoFncJH3eWBTmIUJbi9DNIlpn
THaInB4OtLH9ZnfJm7laIP5/0u6qkPdelgbeycgPpYdi0oZiIWPKayBxHXp8/+RW
YuMN2Oh+7vFpm12fvl+eU8Nn+/pMWLld8mUTceWVlIJriTP9sFpg8vvkK7qJIqaq
kb4/8Zyhc9QKtGH/o91auNheQ6bFlj9vkyOy+a1NA8Fq1TUi2WvRoQ8f+fd8ud87
yStmjGWuXtBd3Qhm1FQVW/z7NNPfukCu13mOmbu0/LZp70xY9aNz5ZiUvW2vN5Db
CxxxyYG0IoYpeiO+eX3IUEIENiTRfMtBR6RZ50JWPxGcgoUtNIIN7x7akYAwBioI
/Mg0G1FnmOhbZF+hW9XlygCl/7PDCOv2Tyfh/duJbgPt+JxhKoDy8VeXuuPmnF8Z
j3lCtU2m5mLm2Pza0hX5LstaZUiPhxF0ZWc6JAx0inhbM34U95YWMGqgdBXnUjh2
JQZA3hxPw2TCqaZrHyh+Sk7cZcQrzjpORbBWixxPJ93X/N3FSGzaPCWgkNSHAWz5
i985a2lSChh4j3DdrideMPtiSaZ5ICbxNEVJhyuABo9HZeG3NkVNC3XfScaNBG0Q
L6mu0/c+g/BtxgWeTx0T9+PVS8ufViPSREwYNFULfqZgxsT4J43zOfa2dCwuYbel
L3sV7EMO6n08dCWwSimwE7VsZ3biQkxwNmg0iGdD17ZpClZBcKLnWgVv9Udt1i5J
xB0c9vQWXjQdaKWwC+XKgwPtICuF2Z37jpWFIXiyImkufghLw65RM/Ri5NFjW0kv
fC3s7ZwfO5ogjpSoaPcoK15VNCGYQSwdtMdgIFl5B6aSyTAJy3GLUXOAnQPPsR7P
xO1cRI4c13O1GqMGAuvj+XOOqxrUsjYL2qxGhySBJvMNiV8zHmIx3jfveeFKgsP7
E42kxrpp3wI0XnYJ/NbQw2BeFVwP4o4+2LbQOmsa0POdaFYZUfvwDeIIyb9YFZQn
hhFb4u2TgoKUsEG04ZycFCAEXUXDupztij7oQd1Ab3sfYjBqWLn2o0lfSWcWV3xu
G7+P8n4eC9NWj9aisf5Si7CXkc9teD8tB0zqzbQRtSEjBmIQtthlD4yM2IXMgGgi
DCLdOl4v+NxMt0db7LDG5Q2DS13cxmGZjDP4dJ0rgbLegaqc1alESbW+9LX2bnPV
EfKyvuGrKt1fu0T+DvDczCk1BHQjvat4qv+p544mzNdzZOy98OAP4KpeiKqTQ2od
x0Sq/GS3yLeQuoqR/cdWiySnREh19ulI4eE8CM5oloFJ75q0kuSG4KNHSGqCbcBu
rG9AtIflTttGkdQGfEwr9qYKX1Absb1/Y1BfguPk+3XzS9ycf7gP9OBgktb24ZbK
gYqfXoGJBFOKBExNGQRJStiJbf7l1GWnWu1x/N6tDtMTWZ9+z1Db2bIF/nz7iVXF
yPreYOEJxdqu7DMy1ynBnmgPZYj9CyaygkvzaEyOXn9+Zwu9XAzN0Lwi0ptywiP2
Dyx202nbqWI5NokZm0ns0WEzR7Zw0FSHg5lCB1tS49YV5gSCMKhiOHKr8iduEOnx
/Wu2Aui5MH4z4Xf2xjBUcDHpl0Q1KAg/T+KOGf4YVDuT4Othn6Ox/V0J93A983uq
JX1TKfm6DAS7hppuo875x9UQ9CKrJ3HwrZ4wPTprp79t9PyxxvUxMIWlah9KnB33
Z9zxUPqLmQv3PlcAk9wEp3FPMOMBcJltIuHuU8+ySu/ITlek+mKN8LhhOTOy76s5
jyIZ2QhV2DIk/Vn8XpC3K9zy1coE4QC+FOMtT8mAHk+CTy2L9IfVxAST3gW+4l7/
7PY8uQhgNUfCWbIplphqgmxmR+0y/RO6ihqjMmdx9G+fw5D5H0WYzDvGzi8/LGEf
xeAscXHmnN7bgrQnrHhFaEYU1VQ4C1j+2d/37g4T40nx6E3VSXGJqHhIpWven5P8
IKFZgurFZlwYVEdgV5OtRFeXYzcgrtD3Rwv6lpMmATdq8BQYztzIXIxIh5KRTREH
D5TBhOJceTz0Zr+owFaUKrbgJCWVCZm3NxM/Kmhu35x5h2LAdkQKwjToZowqEeq3
j84cBeFMZJXpzNhpdR5kzAU19CQSeRuA5DID8vf1FQrbPEWQzL3hHTmI6FdbSUYW
SkRjqOzPBCAcu2e3DqULqnVPeS1yun+orm70KlAh6/RqBoTRaByj1X2oroMct49k
cirwkNN7X3jGdETG/DZC/ENggUvKujEdcanPfO5EIHgxPUaAmHN0u/jFhvCT5q+k
tp08DgUjy0zJpuvdoD2v6pXZmXcbuEHXoK6Q8K+HvdMxoGyr6QmPKObfpX+FWPSO
nx6ycTBND8kO60P/ofIyrpuc5qe9c1wvqiVkwruH8LmpgchIWnNFE94dwj94HlqO
6kdtnuUQNCI27M8S0Jv63ERaYi89sD+A+W4earFVfDTB6LwoFEYxeReRXMFG+59v
E+F7cPLwHMjaXrMJkykTFeEMEtnS3yefj8Z0FmYzDApseWuv2SDQDDoeYitFMMHM
C5t9SJNVtVjZekHjjHPONe/8xm3glLHHV7Vo02thHh7fZyjSxPZoWdvqS4RtfnSf
iJ/MbbXDY9nb1zQhrmtJgTj2NjAmtJYh0Hw3LYOdig3+gsgz6Xh4v/elNVv0D69D
4YiNeV8QI90qj8elPhUP9Y8rUTqtuVcsnAgpSTHs/XXfduJdcsq7qOl8ugufoWnu
T6A7Jh5uIhY+jDnAit2nZzX66F+EWbSn1PM1nWk8st1QhNenX/T7gQgrzScxSiaF
R5q+WnFaWAz+qK3fmhSKJ3sN1I2sPEmyF7lAuxlczU0IbMSuwAB8NTn805bYs286
lW7VEk77URvExm8yTBngQ7mAQw7lGziewpU/7z/PUK5BxnsyctKcIaCVyUqzR0hF
+/TfZPqWtKU32miFU3w/kppXlHeq1W8e7KrrVBAvhG94i989WaYNa53UVFCk5KA5
dli2bqSzbAxPy3gO8/Gz6EuYxYaXWbNhQ4EGhnON7hAz0YtAAf6MdvmMw6N4NIxW
EtQxJ9ibBDvE0PG9GfSozDFZyy5IGpGtyIxjIaJlPfY8u8yZboBJW77al8aLkK9P
AgpMv24iHU50g0pdluVZd7BxJSK0E17daKXMJtKNMh1GmSH4YkK0EG/5hGtReSIU
2s5ydEfGCOhaPwPAYtPZDRfxegVqk9A0wPome7YmUBCaiywvh35BpkQxOPI+Kf4z
tZ0UAn9mxtMR21xbaBcuip0FlQVfGY4ns9JfyEVgTfmzREPUPyAuSR2/l4Ru6vIN
Sba1oWm9Tjayfmo3GjEdwkvfpO8aYIw22xWSdBLBmgHRhr4wO/8Fb3aKaOASu2Lf
8dsIFVWsPAn2siYm79U0+gR8IMvKxtyZs/o8te3ujm/1ANsW1wwWchkExyF2mDeq
AXqM3INQ2yZ83zwymL6xVJQfJTyEOFbJde0fiF6To3sXD2EpcgjyRnRKqRpqxjYF
MDScGID8dfMiHVSZbhnc3f9abajVFzg0gcDGQgRH2jIckN9kSirL9ECrLeZk8Xd2
S6agmTyfOqoGncB07wLZ7xsx+k7h6curM7jHMQGxP01BEP2Z2gBwqOjwPl/HIwoP
nda7ulf5GM9voxTbS/T7Wng7mSkeh44o5tL3j302xbe88OnNqj+TIdM4iBf4IhpM
YzXi9JnqE2YNyAwiKoGmLXkysxAOZdyRPmhIAs8rlF1Gvt/X+O4akIfr/EwoRqQd
cKFkNTk9JWH/9fIGUNBpiZKfQ7jZY1SIDsq+pzITvoqHGexYa4ZzBk9KQFUVfjWA
JHbWHM+dDS0LfULanooe06rGvZclDzCS1hPiVW4l65DJurGuEXXCnJybyzlDMk1g
zv7zotBCi74aaI8D+eoNktWg2hjVwx6ln8upTCUacAqTMD2LHs0TjfLiRpXv60gG
WHnsb1194NfC7/xngmanRiQO6XTPY4FTfEPwdh6OyOE4NNeymKD/N+EjYXoI7xbc
gwKsYrghZOwRL1SxjBaHGQYfq4/DeqsknGwgr8hzkIR6VNtut8PyuhD1m+zFEwVP
WdHQ5xlVndOtVkVf49UuY0ONiEqIbqglMa/E0HO0C/jowPhYumBCVtEMcLv9qBCX
fRUD8/HPULrEwVKOCgdwR1jtj5GEOaxE9SyBJZT3rNqyd17M8RLU3UO8Xf39bqTK
x0Bux1ZJAtgWz8A9rrLuC3m1zq2jsfdaolHz+8qMnNZBuiwNSmUm/KLM7tF9Eehm
rYwg3/3CX3HuRqITROiOA5TMqndEOs6SUkZq0i5RaWoaZA1Pi0XS/j+xgOJgkmjT
NLqSeY5ksyuZluaDf5rMlCycK6UWZiV6oaX0yPb0UyinjQHQSdYQYBsyULohS2db
p52bUSGhx5Mlm3qm0gXSpVLSuswxTfE+VqJKHJs+dVLiL3Npgs6VkfTMxjySB7k0
6d/f5lQdX6s0ow0JGGOLO4D58fRMkXMwZ/vuYfCTbOxaxCQC71EaiTdTNMYjWn0Y
a9NSBjN0lF09iFXFnQe5nTImqOTYJUHReDZcWpV0YvaB7jj6fdH1ADEpmICBT0I+
kexFkLd4EFTv5aHd+OCnYcS9COnyH6Mi4/XYbMHqDxbrj21ozGhDLbO1ejNeQWP8
C+49KoShofUmGa+J9eyWsaGnI5wjisAbT1oNDY7XV7sXVsxx/2eltp8aQ3sq/kfq
ZhN8oxJi67vlYPoA0vBfPxjSdjUuahrc2bQJcdnyaePJFSJ0aL53Yw5q0zB84i7O
0CkIf0U+SjhwHw1wUvlP2i/zjVt0vtQbuds5tmmKhp+EgMZ/SIomBUizFwakwOed
k1BVSNjcVvMeaKT6IfR0ZZzE4h8voMkfgPqPIX8qRwYP61FB9c2ySRIh8sdWnt+K
TdPT08dfj+xOw0dwqXNZXGrIBEs4+MPOD46RRPAJBVUbJz4ZfRESoKFmksFRALRC
u2elc+a4aq16CFoPKNDKgWqkZusyMLydIHGReElXTl/ft+TcU8LkfjCdLZNH3Cda
KbrRBVMWP7tiBMQXFWBAb7tCWIPs3QvyL+uabwGqQFStXisPZzWp9pch1dLWr/hN
KWGQuwWBHFuJBVRcsHUT1dvOk5yq7+p/BiHtVjBn/3F8kODto5upRuzIvAtt90tr
nFoGf0uyYAcgfgBaFP8tIpp1xTiWXQL9gqATrGQkA6R6KQ0PwM5bDLuHaBY888Ex
b50RpsF7/hecmtLOTqm3cI8SRo60nTfI30uOoYdk9a0TSWbs+ib+gySC3hAwZRb4
qLBvxoTENdjsHGN2nS7spaWtRF6peXO7pcvse2MmT5A1kg7Gq9y8PyTQ9HvFgtfy
ICoTm4jMiHq5KblKCiq/D/PpEYq5mEGQLEJNJdhgYgVTtf23plLFtw5RHJ339RuL
uVV7jZcwEoXIkHzWTK66OC3JE+M6NQ7ROCj4V638HJ/Ys7eT7ocmt3SWj0CMK5zy
tyN6/1/4DG5uBE5xJc+bktOly1il95R9HjcsVImkal2FcazFSBm8Xttl8ZetA1dF
tXBhuZODXYY5pugQOorn1reQFccwqckpWanq4J7ei/QyBp3A1/Ldzd/LF+9AO9F4
96Df9dcByPyyxlQ5EerdpwMrFmZgiN2Crs3mPjQ6EcZ2LcEQnaHxXKrKQu7eeXJo
2eITwyIJ3q//rFgsZGt9Q+CYdwhv1oIssfYDp3+QIjEpMQMqkfOsGXY2GF1cDS6S
CVbTfizz/aTloxs05Q5T2IsGE99Z2FoBZ1g1E0hrRTayK6d5aCyb9KetRVvaMllO
8JPxNmxEcVE8roYUdcyeDBWHLZNaqGkSHIzcRJuTP/Z+y62J4KyHf92zUD1QMAsC
1UAgUghvMWtfrOk48fmbZvi2EeAZlmcEC23atafdwwEr32KUJCa9wmzazG5VAq9c
1Mb8K39YkEBb1O0yf/9E5iGBbEgOKB9+A56LU03/mmIFt3JbbgZeIPLA7EyLCiR9
JdCcZMadz3ue6e8kON/DRsTmBu/slIT5KQzCM+HhgefYk24/qzt8Vo88eaoEsZIu
myzuYwKZK30iKUFKqXzX3rhoVe2sGA3C9z42q3dmLWq6seu9iK2XG77AUupUNYfr
giuyDSdCMlmq/8rdY6iY5YTqBBgUy4+VzqugZfdaBZXhtjEjKy6Sz2woY3cYkl2d
4UZW0aXYd0AG78OAbQEhBwhDyIK9QBzE1FmJZkE/gsWI3VnagY96qv0EyBxp28mV
cEvufJfcl12AHY+zyuoqMkSba8YcYU9p7NV9gfWUBIOhoX/Tz28wpE2fSxiX9sMP
vqtXGvnNm+Wnl+GuF9TYSAU7rRLBsaEQcRR4Wvld6WqxvnQFQTws2OMadpD2mHKj
gqs4NLfFjdaXvNB9WG1LlrdCidJuC+I8Uk7M2dj5a4vvOUj3kSFouSLhmU+RHciX
0aTtXL6fs7taktBNl5gsZn9H2jRrkvPo3+WzMWD0oNnAPeevlCgg4//TglYb4ndv
liIibtUMgGZUtrNKFQW0tP8FCHDRrKgjGCnkcMQ9s1e0Bjj+viP2mCeUvaL/yYSp
Z8eNdmElkB2vONVmJmgrEKg4mWaE2P1OLPt7pc0Gyr+CefSNzf0SedlCrYKdu5Wd
B5kkCpGFaA6eTdjMI0e5qQqqdcKDznH+7tkS1uLSbX8MVvr7Ur8XNMgDTrEG3DGD
SaZ6bCB/97waDGN/iR8xSBZB+W/nxcJBN+ZCUrDhttLQxxTeDxWhxJRXZfH6SHsl
YL3QSzKRs6kh1ATvytWCE7fKzsi+xgvWq0/Z5RsGNeIEAkV4hd69dHp2bjUsw49m
mDY0Xtuduicl+/x51tz0yddR5ooMP0CDW5HVo3EGwA5mDo+dJaxXl2Ept6F9ijhR
6Tf6QN7mA8iUNLO1E+KqUMduh/2RrnvAESurCvFiTayQ1ujEdsgKXZpK+nMu4TBa
DeWJ234hdFYTF2+bGvhKyXtsf0FPpG1xxiJ8jWXkUS/ABZj4NFxhnFTt/wCUqUkv
rJu9wlpN243q/X+DZW3RYNbIpPSDh4u2YOOi78SNQb+7dW2Ig7zOR179Dxm/66mD
8mQu7oVEnNGk/bEuPFxqf/+YCelbmnWnIS9aHt/v183mQRsaE5A9IWq7HOolN3Bd
nfrc7nZWA5vLEeZvZLhA0kP9iktU5i685aq1/hw3Y+xUnRD9ES0QkWQX9EYUAVyw
hvc9raETpetXRWwxuc1s93K5ybYSN+wlzx/yy4zHy0/ZXt17qWHgplpb0gfgubpa
t77loHLm83cMTQXyhf1t1KezmnxMjyX1aCiL8S+ZsVw7PeNPrrnacV1jqtuIIhrf
JR01eLqncHfA4dWOgSNFHY7cXivD7bRT1XT142sngMMpz4XlZOjzK3sHG7P4RUWx
nxHYk1uXUSfppAUG/islhGGQ+2YoVd3rc8munh3v5+usUhmhKXKKbgOjvleetBio
ec4rHJnm5mX1ZiXaPHh+OrrbLMGYjFQh04sa7dN2THR7wvLS/EKbOWg1lMScOkQC
0vaxjey2lkmrv5oYbbZzfXTEq3GRpLqKPpykuRAtCNMQLrkvR0XdqwOcF9lKFmh6
ST41fXc4NaIKqnJWZknKPNGNGgJBdzPNnqYpjtiEpfPLPfKjlNJD1X4czl/R5BJo
qBpc/9KCzaYDqoP8Vw4KbvMD2QPrzY4+D7iBGxZU4A3LQbHHwYuE+IgxXmPYkNl/
QmS3ooiiwOkFIpaoWcospFnTxffotptOZ1cJLIgRxEQWPdGXcJXyA3cmcdHaP6aA
F1vEHv0B+ttoplpBc5KfC/2HOtlIqCMjA7BAb7pH37/HYr0K5V6cVyinOb2K/QfP
Uf3py0kTTEAC+iZHlMLkDBN66y6V8q86VoTqxzk91eCtuOulCVeEmST8BfmRDNd6
ICDHQZBFG8FsphnxRAFnGnTJxVM+Ut+yiG/lP3/LK2tO6DjQOxA72i+cAeBrcHS+
pouavw/OEHonFK3iq4C2ENh/p7WL7Sj8mywjVmxtgTK9TAtKOzBBxwAIzgrJCtJz
oBd2KliBKAcOcK7Uv2AALSX/ytflbwjK0VF5Kn3+tz6cjkJP5rT/73++vUkpghUs
UbFMv5tUGpAJ8gXKPTB3aHK6lj8BjpgToejKNwVSNFdzLVg355R0URiGnBM9CGpM
68HFXCPWXOiGq0gXcKq4mphAJ8VGN1UPz7/RIvj8QFzBrGDTG+5ImBdMjxc8/p2H
noPasY0TfKsN/Y52KrLTw2hFktZI9xP4RXnwtsRMANXkofvISXbVa1aEg6fKYl4P
JBmAEsBjcISErNow0Q7f5IS9E5lCitPotAtsv3Z/t36ls1zQRvVexW3de+FZksEZ
d6KF5ZCI2Ic0kCPzT1wm1Dmy43Kfr9QAf268j19IJobjIiBzHDmcdp+qoqi/9nT4
VJG9/xshU+VneHpSwExcC10bdKvTzEoq47NW08v2lWUG+HiRJZxxDruH2mISIGJp
NQ2NdIJvxg/D9kzkRdbOLQFKNiVjU0dCVJf65b8RcIy4MrYbkkCW0mJM5xd5z2LF
nbfaoLD8oEDjbOKOURo5U3Wywkzyf6X2IeHZz6m+ZpslghBdKPV8eCw4IIzUwxIS
lWKZrWb4JCV1NhrGeWQpow9LuKk0FFLX/WZAKYVfZI50fIodnXWKxAdiKDxdwGpk
IeHwTH69VjILKq/xPrFtr8pNvv1NJ6174HIkhPzcpIdAvtlXbiQfYSBwpaeVhy6o
s6X+FVJQ2Z4ouyCTWsuZf2d91w+FENbHgVaL0rrOkxMBGpB06YtZR/kD0FhtJmTe
ntmelPBSe/9If5zh9Ecq1iF5aic4PXDcXwEawyAyOyJdhSDUeyKpKsn7oknoKPEY
Pb5mu9m8AdO86DKBtPMZlsV1CXrX0sOAg3YgkjlsmorIKKqa47A1uUKp7lmCNWzj
u3akLMEAVYr7SFOQiPqadfWXypc9UIgN7SlSQEetXbQizyElslWr0zVCorxodfef
QO2RZMi2sqFDCLZVfJlXGZcP9H8bck97E2lF0iheJt96RsAjSvkmE0MuzgEr8TQH
QFsValKZ0irCijuDUJraFYnpYGEbMtRZni4hsD2+NlAzaL36LbDlRGqnWDK+nu64
/fD9muyphfPOcqslcLRjXAm2K5eQNEULSzlnyYzOuJC2puRx2dxCfaDk5BSLZU8P
cAyTOPyK3nX9rY9QSFxdykuOj4h2gp1eEYHo+oB64/JrfXM3RgEoDtiaDhrAKLyq
12eXG2eUp647KKz1Bytrrk9J63eoxGtleTJnzViH3bdc1z5ArFHe3Ct5hoKc9MB0
hkoEq6UJW6+CfAyLx/s87Z2rI/LCr+5OApWC4x52BiYdRxa8aXaSrs57L/1n7gn8
uN9JGF0G8bkxs1stgs8Z4cq2e2+jAlR+/5yoHqkAT32Rylk23eJMuGavfZKVVaI/
rpCYiJcgsZ9ctIJpvrG6fHZ6UHj87SoOyPABcf5AzRYCXLbF+vpukNGt+PMij0B8
EfL462eq/oKfh0fZjum/dWyOVS6aO+DB7HQCys5zXmm2aSIuZN/41FRD9q60hMaZ
81aeQq9VdBgpxqmB7BfSZxMl7jkHPeto8aRUS/en5XUNszBVvHPz94xac86q3k5i
wyR739n00ddes5+oLnKeOtrw4JTiQ0pGQOi1mSbnMNHuPYDeIjLnZNHzAxQVwbOC
ZZ0v6rMnd3YSxlRZs4kR3zuItxPoohK3V5XOafpKIKms9NvbLb9GQe8eM4yWsKe6
BhgZV8I47h1qsW8VhFYak7z17A+HRcttF/WpcArbi+eSppCIdwzxzsqREQZeWOin
GKIAZGkr0puLwhZdfDu4S0hjosZyQZmQ9+Dmra42BhHHhUc3tfPM7sc3BNOT1MjU
q044t8+L92OI2EZAB8gcqbn1XnQ89v5bxZZ4v2xVE0M6fiXdPjBrPCvnBggMQsYh
44KflhQ4Qt1LnEEH9SA5vSapUuG1dNFugyeOq8A5nyxyLJZg/GstEgwTpd8HwkDy
gurMKco/mFTO5B5PcdcLM4jYOFK15c8SLKy9nLI9au9LBamieVB98CYZx8mswAkm
SvHTqoOLbk6zuBTNnwT9RY/7KWAZFWiP3ate5PTaBj4r/6RJzZGEvDInj3lYv1DW
RxCCTAOoRbuhIlkvMefGzUJRyHdYylJMmFDHrX+3M4SYtJEKdHsrmO+e5JiaWKLd
iBcORW/DddMpSNSBosD2JdqnQcpNjyz4+q1amL17XOFLizWmJJ7Tv3KKZAhdGm7O
JGjJ3HsnMUoJINRRHWg4hxovkh7vgAvm429c4PDfh0uJoqSqZsTi5M4R9HevmKmT
qwqjPp2mEyhDTY3fcpDBDEtmVEHMITz9T7V+2BxhOD2e/4hGbCLGrlpq64ZjuFEV
y5uY52A/rjXq6+s85yU2nm+qLgf5+rYINvZZNdyq9U/I/T/L+u0D8fkyIzN2SJyj
4IjoGO+g1Py+LMJ7Rdt9ml9wYC4Nd8hatICb13t6mAihGlI1ubAs5it1BYssVHj6
yCRqGGymPB3HsE5abS5pFMLrvQhDQtb4XvZDgDy118/IkEc7K/B++XEhhBep6I1J
G2XOj25Yfv1x4PzpZKXwymPsh3waEFW/Lt0F8vQgIKBVHzkXgWDj/lbQYQin5cO8
MbsBmIa1LBXa633ajgqm896okx+3o31EAHsta4FQ4hElG4/gV743jQwtD0zhf3lp
U1ADvkns5ecoA8e8mCK8AR2KrDpNET18WDkuWZLAi1sfWjfsAgaYuQI1YQf5rjLO
HMv5JzWSUNrpNLEDJzvMjDmtZZIwzbVsut7N/v8DW2YLQYccgNOnv0w1UR+5WXdM
ksQ346WINmse4yOxoHzUWLSeCvkMPto48nK+7q29pRlv+m3LwuSQxOumaTQMdymd
U1cKoOZ9HSYFFQE8vkHaZByQYAe168786EPafaNdMH050AaTy1XCJ70d+gJTXtHM
8kpDBP3h2w8W0xpZkju0XJGopzpF5Wyb/0nANK4W9Td3DMSUVrXsbbsRRDLQMekp
l9d84sWbQ9/aC2AzYzEW4JIxmEs2Q+6OUxyLLMLTl5umeOJz1fgdm/VXunQF8jO3
k5+av5vB73cac/2b2/g1+4QAuE1laRdtwp+HPapQ9ShVxFYRlCAZh0FpAalBpyG7
9nJEPsEdXUjZB3dPIJRyAdCequAvGKhb5Of8BuLoSdQ2Wtv+Hy22SbBCwWNLjEQ/
Y2ssmzuhJOedl9MdGhmVbvMEerxqyd2iir8iUW2gc4OqPA7oB+63o3wuhfCbwrvo
57Pk4cq6lyT4NceZcOQnY+aaHT3mFVPwaM09GDt4Z1C/idSJcZ0EBfkd/mGBEWc+
YXPWXg3SlpULYUK4j7ZI4Pi10wwpujF4v8jlJKOAMQfF7+t+6zoGtGDrIR6bZVvd
UrBBWYHe/ajOY37o6X9g3JAA9FuyfwEnG+swXxH3i3zT3ntkvpXX9jOCP0DYgmlA
ySYOsNJAKAS2HTRwJyju//pgL2/x8ygQmty+tEbDjG1kFApft82Bb0oXdgESFrfH
nj4I3eCEs7IrUz4rTYnvWcBv+j2YwwTOWsko0hFXd8hbw0SikWuCbuTteoH9Shc0
12h5SZni3ncfDT9B4TiAHIE3vW8/9dFlCqUdjFE8Ox1VHL70zGavQ/L5XpVWzH2s
GRYmdHLyqiHYMrr3uTYl+TGpsFVeaWC3bxnLw972FqXByu5X4GPEMwCb4GMKK47D
BCfo+P9dIIyXwhZX+5mYvD9WfE6YsLCDt6VYxN2G5lf8EvPLrPeb0Av5/JQLy+/d
5XQ37pLGA6o+Ls3Eekj23hA0ZLvWTyFBIeNyMsPo5Fhgd3KwWaxReGG7/gCoHBWG
TKAuE5g7aeN3VI9caUIWGUG9t8+lg2hKgHRpOITBcCAQSU3pZhi2o67IO9nw3qDC
Nd1IRERQrV0OBNMd8h88Vhu/MMS7dMp2sVPb/lbMuOZ7ENiiXH1iZaZpkF7CFD6Q
mQUD22KrkaLvDu83t24nE6S08j+QfCoDS80Lwt5BoFCiy4RTvqlvRgxReWDXonkT
DyWLCZ4gW7BwWLwQxFOMFYjjRGVXFtiNnLnIGn83OU8Toh4/MZH5ByRqg10t7KMW
ky0AYrPDkE53mswqyqjd9RD1X54sy0Y9abuT1e0nbWTUUTK4FqjEtBhOvPWMlXVE
gVJQ4MZph+IaqbIZA8bGot9o4rKNXf0ZH1LcHLsaC1GnaFiLKx3+iwkBxISxgcin
2HVOZ/Fpc697agDSIljkVsWE5tOTvXsjEV3nIR4nSqUSsI+tDUCbqLnGIb+gk9FY
3SaQufIMVWc46h7XBJGspymgxP/sFKo7og1fGZjegfpqeSP10SxnolRunGYGq2Ba
+XujQxL+hes98+azaMtbrowvVNhsOBbyWaEeM82sNV/hvFaUXE4/qZgD/VVTyW7k
Na1jWvyEwl+AXM6jozh8CSHXVts+8bwl2nerMVfPHiLduKmVpDMALfW8oDdgfQVU
oqAOconw9tDAQdq3gQ0+WCkOESqlx9ac0pr2GbkgYoo/5vaI16OAXfx0Iej8DoSI
H6KqUKOGXWWmtHUJ5N7ewAYpSxzJGLq+CuEEGt/7F/XZA7Bx4h3a6Yq3vdV/A4cY
v3fZ72rrcYlqfYhBqHWIzGA5bxO01Lv+0ZtPYz0gIEsBLWYBMrWBcfXHWYzpW7G7
A9WpWvllIftjEQaU6uWY0rojx8UDwuL9MjZKX1czAv9g+52J8FYGDa0z42DDpB6F
fhrqZV1k/xX/IQ1Gsdp82iU7eWVSFmbOxuCz4JyBDhnp5+x3BFIFJJeZwU7AssFw
ek0Iu++xYAUoF9OUTd7UXY4LXvLu8uL07Bfzwp4MAev5xkDNg2F6BMC1AbkeogSu
zy55PVCjdJ1JjlNZ7TzJBOnfB0RUjbNxskHYrlDXLay6JQXTlNvXIeenR97HBNS2
OrDkIvau2iuOrNgxFPqXn8RhZ9Ttxi4OtOzv1WnIS3KSKGZV+A2dPc11IAQMkZjl
ybFa/PKHrc71SNNpIecjwrjzlCx6MADEJ6n1GCGwcmvCHpnrXjpu71daOFAjgwVl
0XvcKHo8iz3UP3u+se53Sp6tpwCieSEd+rcOImoJ4h8zMq5YTwKdAZhQMB9XZDz/
ymCwZOzLqPj32DV6DkswL0ESAmEqyaqPEBDmH/VFBNFTTGyDqSZS0UsixP1taVU5
9GURLuFtqYJJ6JURjy0x0xMCI6qYb1jF3uRfzz0KJaH/Wa0VitiSAEyQceMOmSrh
QvV/ZW3PTbxQLRp1wQIIhcCEr9ozA4vdUym0qZjIPymdz7+PtFAbrL3XW7mTUuQS
WDBXt+bk7jNJre8XAIeYgpWvfWcXSiBohBl8wG1ZgKYQ28C+peGROJivJxgIpZ85
/TuSAolEQYkRR1eYenBW8nzcqRgnnfq/S/GvJjGmIKAMlfJtXLAMC2mr1omwrhAd
f0Jh5a69mVDXZA7lh970kLWDR8LBeb9fqv3GXN6Oj/wKlgP34EBWLJ/Kleay3mXF
Vapne/woOqPYVtIMRkqm1nWzi6PMJVkKlDavpmCgormYttPrpLSD+ugKtT/2yTJB
JNpkseQl+dRqRpKPpH1E63EA+C/9yLaTBUa/zYH+4y27MV96BzN6KpPBTjnlyqft
mRnoRpH0hC65kDXwyC432eydGaTXpB0uBmbLPpjOe+nEzqLLam9i77KvNG2DLEnc
EH6epOpnEEVT1qO+J8nbaBdlZ3tpUbbk882i3vn6ZFwShhykXAbRJUbmYMfX/DKS
tvTMm5/qAq7GQd4sdvnir1NUfrdE2RH7rbMazsEGeS35T0znB1I/nIc8+WKpITKi
q19w4hauU2KUIYdPgynvFnXfxXIHYXQo0whLQFsLh943wo2e65lR4mgVtXwFimsm
VSIDHmDMa0JX9zZ1H/zb6wH0MFzBU8coq7zLrPnXS2tgA2tqmpsDCet1t7i4UtwM
6Wz5TFLUsWuXHlBFnueg5lA2EBL9O6oJwnHHQzWtKdU9NHeydmK7R8EFf5Q4q37R
xseSgTOCcv3jomlsW+PmdmykPEfiPksabk3/wusGeIweKN/CWF1YAZMXY5cmxygZ
3O8C5Tv8A6YnnFSrrpSEmiL5kqMoKEX/D1LhSZT5AvnQ4GaphdPqWczyH+KKiime
RuwC8ZU5Z3H9AYNQNwbS9wGT3TaKhtdU4bJWUvp82g/sSW24gf2dgiKm8Hn/Vj7b
0rfZjM5mp8XhEK+unNKeZQBrksnORJMEx+Zq31VTTl2l4wnfr0e9i0gXVPp3c3K2
KB7Bguy9R73LdREyFUhUv6CAw3J+zteXqp3onOj6Uw0AARkUGQekbmFTzJZM4AYi
U5c6KiK90Txc3iZNoQqxXhol67iWDBylmdZt2AmgxFOJ96NEWYvls9hs2gzmo1Hi
uijgzLv7wDzolE6u0RH6FiVMmCOxT1AcEP8rQrenQuiBfUNXBclNwCkj5n6v2LJ3
EiOq0WWf6krAQxs0bOfTbnJp0TQd5FRbMv7xM3b6+16OKX1h0BEPVlZ+gcVLBexR
yESdPfCjoia4fJDulTKmB5K0haCnf2DXQKjQeJmgHnSXvsqCZKeCL8puB7As5NnY
ykz432Otxlv3duFg17itdRd4ugYXUumgwPJmY+lAg1FrF9+xddI/dQN/qLFkRFoo
tczQN5CMiB0OPEBvQJLchrZuC8ABPswVRD3ueU3fhlKUdKq0c0/6bv6os2jAS07z
vyEInwSUUxle4+gX55ms5BrXESpiIYoC+nYIJR37H3ad+emkwq4B+4bKR94ySaZx
x5K7bsNydOfBliv5WIXXdS9HvIT8C08dKUrOaOXEzxkDCqwfiNuCylvyiOUS1GiG
+rWDKfR6WzGzMIiiASyC5Qnah8fymEuKsnxCVwt+s0OrFXOBI65SHsfV/op9cwo8
xMCfqX4HLVz5R1Sw5ybh7wPjNBXLsvyehRiCWxwAs9v6+4Diqo7139pBdTg9Ii19
xhBSKZ1FksL+t/unwV0+N2IkVfd/tX5jUxTM/7xci/olvaHHO0fAFCdIB0Pdhd8B
WQuEOZVQuV2fvvnEwl9rFuRBLNCA6q2fmj3n3uk0JD6uLo42WzvExxAqjzujDWf7
oyvayHwoagf+q/+dgKl7MCUgMyS+Ul8+OAGwwmAP3m8Lkijmv7bOueufmiz2TUBW
fSsqd1NwTeCdBR72PZA5awTS+lnmVNxlXwTbBwBhWoQ4hBKePCtwyfSu6cm4hY/g
Rk1jd7bd31k+a535m9DuPjTIRO+1PTUSaA3itB5NHSR8g3i2r3+LRjMLAbDEAlen
PeHT4pglQiIoUxLE2vBlb7FsFzYcms7xYEpGKm7kxuh5JFPQ/+lrJhdrtD3F5Njb
MTLXwVrU7m34uhhYh5lzH7uRXn32PmBdaCH2LMLkVMPOLIg/beXyhgeJjuBaOUx8
5mb/nhe9Aw0hyHDb8e7hVuzi1HB7qPqRgzMQiZS9ne0UqmvspsT/QLdkm2V8B5fY
rxUJFtPcJdyyPX7a3tPq6MObSJW0OMklfOV8zfgVHjuOd96Zpg5W3p59bP03lIWX
WecyWc9DKndAmXnC+SSp0VuJxsS+PTcGEWNz3iydNmY9FKRN2XWiwbkhhMB6woOg
jVNZQy5YwU+GD+gCI21T3aEQH50h5yJTXDnZ5WD7s00oupOJZfmDpDBeNwF8265z
XOmY/qajCbE5St8OpiVzm1MqxH6Fuq9V5/Upw6rXD8Mq7Y5RF4bI8WeTfEdQJ+vD
qpToXWOVfh5btFeug449Rzb89aBjIMmAo5SRqxf+1YWlG2KyzTGgaLLiOQiu6yih
Ep48GXWSRheKXaCCJJIll6RFX3JzbB7p9eWLpShSyiH757m6u13PR2nhGO5swABA
sLMznOy19AlVVOSLJXIW149Qr+2T878YUSRaeO1zcUEOSt9ExrDKg6bj3KGrtqL0
nwRWyBznwDGubAjgDhM7jNjgrL1JPndEb4ZHVKUoV56GFYpEMGZsLUfMWgpAbqcj
gGRRi2UvIK6c2lVLeqSykb2Ev1VYs8vSdbSEOqH8TfDYrJC/1XaB/uiAUVC/dQuk
ZLfjKVYyK5wXKe3STjO33Baidu4Jqy6y3o9bl+eUkJrHaVt5decHAZVCxBkiV9lW
LHDg8052hWO+S7KiQXslu03GY+b7bVokxcPXClEsCl6UONSyncBV3Qx17zrkLeXE
g7fUs/taeugjrfIr5f5kn0JaaJ0x88n1bUPZb8UWMdcSF09U5Mnnx7OJ3P8zer9S
0BEqgBGJqsuCKqZPmOOYongwHVVsSEjTdIDdrdOJ2tkKhcjigYSNb78sXv+A9LN+
w2LVEQqdH7RdCdpY6mq1GghbCe70u+0XGEPUQ8n3PpebhYpdYQSEL95WL+q05MX3
2Pa4eRICZv3gj5Zo6yEwg52S/KjYV7L09KoEjIBrlF+Tsd+bV3A6xDe7tAZu8QW2
ia26AdMMTN2hYbbMM673MIJl7lkPKfTi9pwm4a+8wfI6wRYlajFa13zCFAuWXSJD
l71CkFNqwd+PrSQW56buyZmTl89bj90xFGBZovnLm9KJw24spxbXrCiaJaKya4uj
2PrNzP4jfY30ziOZ1bxjUmfKELFw4dQYpHOaH1Wb9QN/xhZ/tpwJMHuLIZ/BdSDi
AC78LYL9na07IOX92AMYmgdukAyia2rtNosyQnyEsBk0O2wOAfqFv7VOLgMXlyGG
YDN/dFVFN6wdgc4oP0dIcGC1hpQlmwLgsLUWWqxIMLE1P8eQM1ti27O0mac7I7CQ
LDOkgwDzjv47JX25W4+al3ScE5wUzL/diPMv3PlbTrsN5Et9VWp14WXOsDxYrk8a
se/elu+XYMnG8Z74ysPyCBfgK2yJwuQmNipV6BzvAXfLsegmElsYiPSkoDPP6BZ2
sGkMGV31uuUHPIclnD89Vn2wF0XHFv/qX5sHghtem2yBb5IJH/PFlSuctSiOBa9k
HS3nhLF74sP0tqUjMWrmO8Nh+dAimDdpipzlTXFU8IpWRwEJ6GkAPo45Dgyqh6iz
jj3+wM4qluONXIHvFrAniqPkHdk7fpf6PDAvdROkDcaVVKfgVfGcVRgOy18+OzJY
w1tiI+Jj9vWf9zHxkGnw6q1gfHEmlbMRyP42k2bCcWnkxA02uJ4EPGHZN2Rqa0eH
a1++KmfuIELy3pGI57+fSqrw9+r3bW8cfzoFyvxt6uk4l1F7r58N6tlTPTedULmr
8CenfN8S/JmJ6V1p6P/ALNHTAuv6GGs88RP9hZcvUTddRtj2y/vNQqevfrFqXG+t
MZPDlBVJlAtThHSUQPvRem40WyChjjgsY6lM6J3MDFNpMbsrqC2nQaVkdBMRLfih
7tY4J3uDeE+mYbb1+y/cbhD8+HG9VsN+cutyPa9OyZcKJD6twgmd7om4xzdM5Lro
C0ChMP7GEdlVldTUJq/yfjyE4XUagnNsyMl15JrC0QeQdf+FP4Q/bbf6BsWgsqAC
JtipJo4usPqrHL91UwEVvibMyYCF6ghw4lUxJcKpHCxGOWM9NsTaaMGYx+NYTVwQ
z91v4hh2hN3hrXkHPTUyrKkCKGtqGpgRFJ+QSZ9bKC1BEmD1C2xlsQRxhv01gPsq
slhdVFdgeb6SBiiHN9lNB89hLvpyH6CrUG/54D4TIEvOx/MIw7o6/ttF7FfQwf5W
PcIqJphPvN6WIVPBciiGD99ASyKn3tk5YfUWkYjcAcY2M0U0idtZfs3TBZZTtNJ9
9abo0QdskSEb48U46s5b3ZmAXIp9yXJLm70i6dOGd8ajfA9zaseXuziwwdWT6BVW
JLe/QF3Hngppno+6VgjrFVMBlrlP3yKZGriAzgX0KMvYawtOfKiG3E36PmvQ9ZM9
acmLygb3bTrn7CNEDpH9pcfGe3I2JbuQ+847VnFq3cyZyxA5yU8IKcPj9ODb6ncX
ygGyymk5Nm5KrtE2JKRnowgZE/VsZ9fVjEGUubdOZl758n6lAZC0NNIbwvru3r4G
5+9oI2Zf/KDI6uUvkDjSN+R2iA6feXp7k4/DXPzleHQuYTxbBBV2nvyZ35NRlsOC
H+rCbax4x1JtHNcQ/QcXi0swZ0tXMjKvxqTAsCd2sagAWTJvNV7ety6obBq0Gohp
Ev9mPXjdd/JgqAvIJImZxgdeEqTFnFQ50CBIVLgKLzDwVd/52PFpaBUWPyiKA71l
GfAXoZkBJTcgRn15xRJPFnUBu4zjKyeTzNnCS0sVw8WgkdrjHWXLs9tfwYO/+zEr
bfH1hR0VSmjTMWSML+6u7O1Tb/XrLM6mhswqgnzR5Ia2Ycd4tXAQzy7Qf6IU6+bB
stzo/hVGh89LRdR1X2XAtm3yhY3PeTIbOGfzkxVNodM0dV0k2hZQJDW7SEpKQv39
F9J3pB56DsIMYH9GjfkMc45mnI9zAfIMk6hhTPK7mPlC7NORs+7dMSu/wL/vu15q
C2pu5YzlOlUau2DK2LmpssVyCm8pYSWsDeIfovZx7eUJfPQMKP+lgYqn05cjoHIP
GQc/GcmQeuPcCwAFlWLDVDFxk5g5JuA8ur3MZw4zuPeuCOy+fhEB36IwsNnx5Zf2
5HKPpAQFJikWyJ4i6GB8i1qM6Ra4gVPjG9o2f6u2ul14CMYfAiG29VohJ9wzLjJr
cE4E+h5FrhwaqOLcqVbWJatSy+8Z6Qfu0eIeOFNze8HANsWLu0Pq4d468mVo7sLD
t78BkD7Li6ixCaGB20uV2k723U+AWmeoVYxwPFLj6vJX63dRhNFl4G6u6rj7xznW
dvDo5OfBYqQ0gLhs489fW3Pz6Ed9lRzaXYplh4P/eYOKER8saFK3TAHwoHE2+28J
XvuTMO3y7EaWhcVv/uyyMKszK6tEXSTWGbsBfMXC+FAQQfMvk/G16zc4qwxz56z4
IHnodhbej4UMv5mr2QxYOvEoS1z8hcrC/6ymiJTjsPLwx+CN68PiXGTFnR3nwzw2
fPBR8Hsh5gkIK0a2bpqFu99FZbiKom5Yo4M2ppGGsaoBXqmwRJ+nWZgmpexIN/Ro
vnpcSWPvCHx4QHNxdWotpMTzvAawwPRkwwDQyWO20jItQjw2yy7p0j4CUNiTJPgA
p79zIw2Vr+E8fbWJK0AMa86E0n5h2mFNYYvR3Gtm5oBZFuAxE4L3uqhVaPru7X26
ndK/Rl0kSJssx/NDvTlx59g6gbDKJHkmy7L4M8EVHonxWeo0TSjxCMWuGbG3Eo5w
V0rszq0T7yDJXlfMapqAmVQVTKvz1WcxPnM1XX/g2RCtGWRwo2r6cyl2uLj7jjIC
RKgIWi63GfWzGSDyYXGq5IDmh93kQyzc/ia/2Tn3ZnAY873wgRBCQ6SIdwgkUmg2
N6TIKMnQ8wqfuOpacVb700z837072C/tIPfygiEgm03X3+UMWNjYIc3w/8E7eodL
Di9SF8PUKppp3lV2wQSahABFLm17KoReRAxXzwF2bmajD0h+Us2bhcrauLfPF0/H
2fIqbTqB/XzU9Aqx0fe2PXhlTczyC+8HBy+pv7QhZHvLtlKpzezvPXXyypAroYbn
ejSmxTr4jsQRX34nayS+dTQS/UhqKUx8SoMnZXzAnTp4GsQj9YXXJSag6ZA6hNf9
X0n8cJgCTOhFfD1mI1qUb+URw0uClwMmk9PWkAFeWmGz22dI7l32zrlIFXcFYtYE
qT/7pHbYlo8SB7li7q+/RbaTyMZumFXN0pV+ZRTyRxybAauyaG+02ZUb7pZYJXyi
7q/PQQ96QFGsFzSvV7MyFD1+wcJLoETMiqnY16k1ZHcYzX9zPPYZjMwW5Z1ucTix
VgMTlyOwO2wCsOc37T/rQhsVrX56SCcF6GKFYUKSFa4oYL/pA+ElExWpBaCc5HYL
sPLe7yHnFkI1xy7OqI+AawY/Y4USf9dhPZdA/otfb6t8PYJ0YD9djfgGsT6uKFvE
zD3bSzK37/4H6uatV/Wg+tRgWjx3QaAtIEi+rpZf0S+QQOK65yAALCdMLTFq+y4s
6/+n6OKZCs3a7ZsMUbmVTZAKYYhOVoIBWSqdzJxHxBoTCVv0Mek/VW9UNs6Bviib
RL8SnMg0qiWidmH1CHplHxH3DvlQHiiZgZZhgN0zYmRCc2H46lV6d2X6N4C9Bkz8
sYCJZz9YNQHUTtUtDsjgUZoPfYKHLhb20eFKgPpe+WJ0DQx78TUF8uuOdR4UqjjP
tK3z6LcDsYtxEeuyc0ytIBkfhfd41aFMp90qECeLZc3KLoyB1fPfzyDbIdUoW1Bs
7u2fnIxyvm8+2LzV7bmIbPgsswBFbFfPvmKGBdBI/wtauKlw9XYjCLYsCYNP6Nmm
cxbzoudFORq1uFfWSvfDRaWSKMLWY7uldVtIqMkd1zeczU98HAREuK/P3TUNNsD2
Yfxah9ottP2lZKisdnpJfWfj5aFbl3AyUeQhiCRWbAX42fnKfxUmcSV0oJ2rvXTN
s+/KEUkkrDIFv2L3EcwVW2YnE/JBWaHaO0z9Tr3mKS3UO4mFuQ8m9ytAbJCrPSnb
Al/GDoUhIPGJiVLFyaKfnx9Q4OffDJHjSCBlIAiJkyddt/EHoixwVXTMiwKHZQuo
wVPVribWqjv2l/8VnzHSt9PARYNsx7dqVI/O1ezsoIlLkb+iFnfFrBcTpJH89FFE
67AmxTVnmGm2FizhpLpVH2IcVWkp1HtrkmJl/q2DwxWRQyelWho0sHw0970vf3qj
D3S9kfnar5E49t1rlNhwq0nsuZ3983hV3LLHQ/B6dwG5cewmZUeGjpfGPamTU5o5
G//9tfdgvqFlHsrjTs/zZfaOMfass+C9MXBZL872kBEZ92rDVStkuKFTmPvoxsmD
P7s2HWIBCuVe4KNOfRQPRGH4RPk6qks0qiQ+B/Q6aXDjn6ZDwv6uSdBcO4JGhcGg
TsTjDRu0EJmZ/sdv7Aj2cKJ3+Dh3TcuL1AiIruGhF24TWYde0IFDaw7N+ndf7z3S
5z4a3z0sM6ndMvK4vHgcDeZ7yze4HsKvpUC4a+j1nL0eMhDSBErIIgJsE36cDuz5
hsOtEryXCgyIOYMWP6ply8HYucrNijClntw2GkTS+WfON9sktozfkQdsyao9L1G7
PmKF5ETElB8Dso3WpDwntrI3n6Kss/vKSvxPSmQGZHC12ZRxGIaQiBQhDFSPK4Ki
GWtqx2aF+jnzp1PanLOEY9nRQFR76HSpsLGOZCFMAEpgwR/2uY+YWmOZH7wBjf4p
YAKXe7vjUcaLogWGBItUA61OGZzJYzjQblZ/NZ1B6gD1Z/Mf6say5DwiRGzpGqVy
+IK4Ei/jOCeie2MJSP4e89UZyx8dAYwOvWftRBqzg6K5as2KUowNyxvEh9dVADEn
I9na7M83FSnVO+5zuoIqCpQyspovhtYo+L1/uLRyBbLXU3Yr/5Py8xOa66CcAorY
xZgv0LEcw8bZ7oAATHz73qqycxV4QfB5GH1nk2ZRWDs31YPuuEc/0NwVDjd4/WWX
u7aclhozkEtz8fwxk+4jY72VRubYwzc4m9C6myBk1ZFTYqRJLIXV5Qj0t9ygWK3x
BWeHV+YnT05O5iePP2xGrIErc2kqpfy15o4x9YnHKcDzhc/PK8XDn6QAZAKdIVWO
EaLXZNmn/tD4NA4T0Pf8UYKVa/8KA6g1QUjyA9UDE4zv+1I38/belH5eqnbmm9Id
eaUfBpHWX7HVCx5vJnvsuHp6n5SUnV1FlYB3YOzKSdN5gtw81D5ATiQfjDnN1xPl
WFE/tsVQ/GVwcpURYvvxBAqk/HrwUl2gBQF8W7Zdh+UWAFKrKaAop80p/oa97cJY
G60dEUsGAW/fWEeqPSnMXQEvJ5h5Jf+cP98LlQf7nnnxXy1SzOeryms54XeEy8mC
bcdlCRtGc7tFb1Tp14bfvHBKPUI93WoPlwU3VU2Ylw46JK07rBtMRhJIbowB5BJE
pVRgG+ihv3l/vmK0PFyIvpir4yPpdYFcdDw0rFWMw+k9h6Yeafk0jv4HrbKivioI
xIwIk1zRpJIgfodOUtDnyF7oz1Jf3Rpx07CTZGM8f+dKMRC9/z+uqdZ5LYNWXpn8
eipiPdcg/ZucW9yJHB55mMSpKs/+hoB8VdC+OcGUo+FdQOm7ZqP5rXOJ43+rrIs+
GdFzRuH0M1BdHLMwLkl1fVboHNEWS1HoKV8UakshB2h34laTTrARe7ytWy4N2JNq
IjAGNvZLhZlKfPX6QnzCa9Darp9/ZeSgXMW7TJ1aDDCDGeVPKGX45X51Shc3s0LQ
aLPmWI73hITV9XTVvthEKfIoRvrYZbgCPgP90WPykFfO6h4chvuSuzcuY6ELCTp5
qVE7EKueGCxMC8xaHJY97FnFEzcI8JKU2Re1Ljkok+AY25D5sR4rTtQsD8w8tk+V
zV8ANZ8ZVdel9yMoJVWGA6Ov1nxTxEQhKFctUj7kwyKylYVaztU1rYnhVQs6oZ1v
76sSowJizjdmq7ZLkqiMrWkgVj/P3BBpxPEhX0nyuq5fTCUPgxC9UuWulYmXaOwE
bTOFQuhFkRGvs5qC+KTBtt+NDYHpwKOHJAXJfe1uapEWczBNszFqsxy2/ZS8ubce
z0jvGIJEyQiR51wUhiA3bsFq0wsoFdORkrLUnIS0GNGPH0rwTHK2O0uF3O5yseRJ
gldKygNSmuchY+UJueLJtq44AtcmJsINKi7XguxwViW2a+xJjhAHa0Zn5CSv/b6R
kSxykgfpwTYCE6eOSc3f2dF/1WEoKqu5pjEriQ5pwGOLCumDBzkGkyOwvWuQojVY
KFa6pqLG4Kt7jw1JcYuVryamzU0Jp8l9fpLvrflg4DTqYdMRbA3IreY9et0r3FMM
WgNOO7cun3zyEBoZCgtB8HVpaYKVOTYipuGQgAlkAebo+8tH8ebKvPFUX0XD8gNB
k8zHMS3TIxOTaTIS8SrdKIdK5452HCt9A4F6FJiKouNqSUzHokD4AWvYKsn9P8Fj
C+MY00Ph/3JFEApz6r+JnB7RaC7Xu6+nF7S8Cz6BpVyj5HVukl9OD3Yseg56+/Sy
sCI2Y4n/J/s/qoTbEJYw3S7n96KRbH7JCQkwoNUrnNtHTKG0rygoJu5dxIZJpLjm
Ixi9W5ZmlzvCxjHXpeQA5LLVgtwv7WK1BDmTKhYxs6SxNNIn+wQtgPW4oOTxM6k+
MKyqnw+r9gvxKaCSiFrGrrORTKhjcYlXCYjMe2+Y9Z6EDZf2URWRu0E/zGhsoVnK
5IlLW2XFszut/RppoNT0fqe7z50Udv7n7K+t65liiWncm4oC44qN+rzGfUTa9S+C
FkdaMCIIn4t/5AD7cu5bHuIk/atU1P1dmWbR1S1wno+Uk/8PDSXP8SdEgPLXYVGr
tiTJyijc0dpQRbQe+r0F0FhGQAIErXEl5MX4DFP240bYk+w3wrC44+Tx3kD5KYPb
YGlfzkvxSwiE/ktucQRCEYgdSEvrR2k0dFAA+DuX6FryhIae4G/BSxFLMmPCKFmm
aJgWaAsxu/EyfIViiHVDva877WCjrz6Rsq3BORvpGxzGDuchbn/98pf2NUFRYCuk
pMvXfoSGXYWlARA18sy3ZntPByMQ2+dzCH6+7FBArZ06bywQSqSjXMZ+S/Mm8P3F
Hx8JuoEoYnaP+/nm8VJ4x3Tbdy0pnF4ogj8GQlWKMUTDnFJPaV4bQLaST/LEEMPR
aBPGyMH8t8xdVOXIqp+ch98J+evy7BCCbjM82Xr1MaYY4OUiQtp8ajBf56qxyFh3
SYeGlgKsyWcPk556gK+6kde0XH81RFmT/GqyzMyJn53yBlBV0v/X8YSjwrWcDkks
6dCRzKBDeIQO5lmlLbeKOSm9d0ZU19RVAA9mZ9YiomE0tlfyX6BsZNLbXLM4kLE3
ofs0cCtL2tFT5PMezzQjidMUuQIPrK84TFeevdOe+JqFbw8BiuBJgHaNrftGEq/L
BiClHhCMh06OilFvzxXah7pt800iWahZaJG8vkYwVllsxk7oXKUYJb7a3SC0zLAW
HmDqcaFudCl/8QB5h6E0BanMzy0ZVf7f9fetQpQ7FwExmxRfYEQd8shvNrrGYEZI
wHEoosIZPqyxn3L8esstwu2cFoB8qaHDIXX6N/dECk9q/uzGnrI2IhC2Z9USQdda
07e5L+LV8AAA9vyB75WdVWz4lvYOkw6lKQVQtuqhF3yEpKL3MFlCg2RZ2LjHQciI
cZ/9E9rq4jNRQpn5YT13jyXq6h1+SrnkZSW01xEt9MY9q7wjEGBUxGKFhFlM3veG
8BwMDToRmVQ/Qpxu0RDx3b7GT2TiH79wBWIVisc9aXtdquGl607CgjbGKYo9vdJy
oq3IpwWsSXmEri5jxhPdUWkvimMWCVmo0AJsT2nYdli6u77qLX+Ld+/27DsKCTr9
wUXmS08f/8yjBS4OSe3mGQ1HEFK0HF7aHG8TSLcbMWz6lZ2yjINfv6779G5lpPyP
DmbQ6gAExRDm4AsiQ8OjaUjVSimMDYkcc9Fif7aCtbXwsUU61McOMb4lQ6gj+bSp
d0wQ7ikZIjTgQm+fHkU+C05w8IuSLR946C156v7TSHgUOWpguAmlHmo8mvRZKopR
0zZTEL2OS/EaR0FdXpm38tu4w4PnltgxnmLWk1zfS06GhsXckgb1DFq+LbSogq+B
zVXgC/pQZdbhC49rG6dqmLBZUdeD9GO76GaekqLpFWIBmc/241MZ9LkNtNQ1zddO
H6HcHKAWenS0ufF2zcVAxFCjr4RdvXgudKuQb6A1+TpsSWiusH6q4whNGbwtP4N4
9ntgpWbDLvjth1iwGfT2u0Grl8pST7PKRGrSvZyfMlhjKtqJh+r5wnJEPLs/+TbO
pl418BQVAHwzLWLw/ds6bLFqTqI4HqkTZMhtrzIxM+cAl0ahBugiMSl6TfYHs7yl
ArxQGQ91weAWlu3j7vqSyv+tu/YIQrJGrdjVvJGlDmyodgSVxDIaZa+IwQF6ncCv
NaaBkPsE7LZRbFG0XGnD8/3VWH1MaKJd08c08hB5eFjEAKg/MEYDdJ2hkGNzWoU9
2l+09xPnReX6q84KLKpZzwEsNiPJWxEUzMuHpSVsCmcvEeKruF/ShHlJQIDP82Ys
mkqUJTOn6Vd0qd3qWVw/bxYRsIAM0nf2z4oQlX6xz4e4+4mfleXdzy651qtOHHIw
TAVocCzg9CZHRVu7DrU5F0L6kpPct/PtfAEILdUtUB6VsL4wh1ZOrAx40An6Dcq7
jcGQ4rn/3AwVXS92gxKtsZJXSNMCh26cK0QDF74lqgUGBqVmpmnsuSP13YL/mUpf
u4N3R181awRbUe/PuxyYN13DZYevVd+lq7Go6wK3TbchiE5C32oCxWHA3i0xQSBx
SUIM/kHCJFc5wrx7deD96kg6OgfU4ynzCQ6+RP3QdE31msAOZETGT2qPKG6NM+u+
FfBB7hWUsFntyBYvj6xN9G/Oq4Mbc66tP0kBs5PyjrXig5Irp4+Z4363ubNabOBJ
yNd7UxCJp5PHP+Z5QW4lyHmZqUtgBS1+xTZ/v2d6a5cdc/js97NnquQYGxIO/gwk
MoEfBodg4b0Nl5FFtrDWNAns94hDKHq96mqNHN4W7+6RLUTA6wEq1VNG8/R90OLV
JzmXtsyjVFxNYjaVpqxEsIdBtjOd88tf/pXQEBMPi3v/xKriRNC44QBn3WnLXHJ2
VU1DbSmwBa9S6GnBfTcsTpK4sGzB8TsexT5JqfSOjmTEI9irba2ZHhYrRePI7/tJ
FVA6oiNYH6uRxaxt5mwDuCbC0GpDDRcJWaOb7EteKPVWfpaA/0M1XWtzqZ/9/kin
u+c4msAjKxgshskaCrZmCtkQGEMwxaBCJkHZzGRKD/mmKW0XCxfYUqnXIkTc72N5
m1L6x08CxAPvKGWLJuxnrwHqfyo7HUWcaNOEG9IMsNvnz9u4p/4Y99BJ5kxxyfY3
ItvG9+EUQDDGpMUY9PbHv3MEG2CMpyWIh2bnbzKC0dluVJZs9eOMf8TTe0YAsziD
QDkYreUaHFJ3MX0sGKj4XlMdhNZSOsWHQKiJ4qqKSdIYJr0gar1t+YPSEp7Vwom5
bGGk9fZMSOwrs/c8q7CCcMrSYY5chs5PJ0i03TLXSXCtQPjN0ATooctwwaGB77EW
kQmpn9dEqeK3cXsalPfrGvx2Z73oSJNjHvNqbMvAw62LBEuRt/S85SWZQ9wVRRNA
151xuiAgU0oypNw2wtzXc/Y/ZIjGAOhUu1K0+MjuYAxV5cbju43sK9PTE2Sv0SjI
I9Iv6Za7gT/Fc7aKNTRaZsvyKK0Hr8f0SlcqR5rtfPYs8f9Y0fmL2+GgXtLvSIxP
5R2zrzpq0yhmAKeA4+1/Ml/1ewHa9x+s4mNQD0GV3yx9iNopkNs0uqLO51e6hl0/
Mo+O4KCWfhRLMEO7+tIyWy7VU/zt54fDTaE41gd8wWuI8r/aeHdFbGfM4B7HBWzr
UAMvD8TPmXMJqUC9KF1f5IbhwgdRICfrqrPvyXRvWUUTiUAsx5QduCd3zr2NpJWl
m6ixkFTRson1CH/QEMTgpMDf3BkBKuHc0s490NBGsu/SUyEm3pl5CRJk0R+xwvYZ
vQI5PZ0QL3VCRf0TCqsanWDUewyfo10WHp6qBanw7sHjC5SouJirpXK6tIWeI/Ky
yR2iQjTXqofexpLrOv1TZ+kVuURpYuGLjm0sBljJvGz/BlsW38ol4wrF25wUEtHZ
n+FfiT0swiU5alNiow1TuVAn/SmQf1T6aKmYCT+FegBb2J11O/q1V6VkvrnWDn5b
bQwzheVI+uRDiMzOYAlR/qBgOuFiPtdqCU6EmsRP1/1/MTgRBq5wQd6QqIQXoR7a
R6KZBoGOjGkw17MgMdoxEeovKF+12wDVKgCgSmTE0pEcA+BAF/AK5qWopITANma5
t6Nmc9rmnx+wIeUomOWHpiyvH7mI2a8N1ZlGL+jw6UAqHkXQKhR6PkRXTmg6fpRk
koXVIqm2E5zEUzt1f79iCSLNvrAY+VJe4eIIPl+VAk/vod83G4mg3TJRImNdSSPQ
8Gl4loG7vLW2HehjyLupyc5GOt43U6vRmLb/D4XwvjUGDRPwImTN9Bt50fvN5MUw
Xo9H+Hp1L5VPzbR5BlesW5AFoxDwYhDklvjpLxGjtcl5XXJMXbapcFT/BXXmcJTJ
RH4A8QHCNGYpwnSpcDgJyjevuMTJ5VPwq6HEuI9dE3eCpbYuviEBxD7BvvLaW+oa
e4WzMz3ubTQQhfvOZWLQ9kYveOK4zzUFY3OWZXHdVC37Gk6rEawQ96MjSBQyRdiQ
dSmUtxhknCatIRkd/dY4WYb6eL5+ydi9WoegIBt8g7ZOwRlgPwn25OqZy0K4nxXv
eSjTSuHUX+DQXsICQex/DGzaS1WnCWUX5nSoGqPEAQYU1YW4u5nFprj7XGvWAGY3
OVB3xiJXQu0E267m5DCVfRxGCXX4WRCkOUqEY1saPOgvE+ju/3F9O4lKNoYcFIgO
z6o2gB71A5ER2tNGX93/QjiNdt/KfPmMnQyjvtYivwFcs7TL/xkmSmHFy2AkWrIF
4bb2eHVJ+InpZOL5NBVgeTYkpEQzPQff8qUWs3lsoPzdZkUmZF5C81JaJQvw3hZp
CqQ0Uwexm8MYTNtWC8ue2RAKXEy4Gc2CEcp6tyZGDmm15Ku6shglIC5ZSiJcpElj
GBXfEaWuVVgw9FG+orhRcWUII0lIlTFoa9+e3z6S/D59AIy+UYF1QW5LWQ0C9vON
Zgzrim5YchYJfXu9EXVO0wn4OKMLGUGLB2JJsw3xvjg1xtgVVMp/ZM2tC1tHS1mr
N4BVDzxC2PtDZuLaAfhOpBULoUbO/A1ewv793IZ0E1xFxiqUn3TaqfMDH7kM8dKK
nruHpF27xzwUISS4jcESuZh3sw4++kbgmkWz4h2k8j6xyP9dV1B0j6dftOyKrFKG
DRaTrV833MSwbrMz++F7mfk6KNo8BI4Be7dFpFY84200bnCiYCuiKjg/Bnw0v9o1
lkvfZnRwGb7a5Cbt+sRoToGK6FPIvGO3JN4r0uwSKJM/srF+duCa6yPs69vIpWH1
ESOnPhXV3UdXxSUWjLpOjtl1MJeZQWt3VKvW1n94xrLYY2eznJvQ5DWOSW3eOqs0
QQTSZ3qBCnvZBC6BTT3rqD3JWfdQQBMg51qVWsxLsWQJ4Mpe4mKXGmttDjkzvb1r
DjSSMznnRQGKt1WXybHFdQ7niKfW9/xEiE3JYAges4TetNF2nkHztLM9bXSuFAXe
4ektltBErhvdADQHB4s7TNfcloIeIcXfkqNDd2maVchx0n1y4QLdGh50swatXpGo
V0PhPL9rr8RIoOPiqpLbDzOFT01YlPN7mxBxo2m4Qhpaaf4/U6R9J7JOT2WtFOPs
i09+q+Djv2e54Sz+VSPOns1Z1GIrCaoxLG89FqyyAoftAp1W1OIXziUW6gGoCyxx
4SRdeDqmSSTu+WXj8nuG13rc6VCXLcathQYTN+OTgXBu9Kcfsp891q9DNaa/MoHK
k4TP3+8xcforI22LUVesCcBlu2ibFHIO2YRlFVMFuPbHUJvE1eQD25O68hJQIFBE
s+S4XwATFugks1dp+3q1ur9/2iZvWrZo1Vh51x50vk/+FXE1t87L5jDrxov0OjY1
aVjUXGG55xlc1lB0Cu/LuVyIfYA7ZzOaxnaluEd7t21YW8Jsmz1XaodXcutN5++q
67/LKu3RnQ8BgfHffbdtFyNMmN8HMY56VH0gptw15srXX/+P4Cd0CbkVpt+loVus
/y/RjC7/H+Mge2uOdL9+sR9BnOxoFl8E0LN7t02e7pIz+VGcPuqWy5S8YLOFdUiB
6G6oH0AsmmThwb0MQfbMoSq7bBQR2nLLn4PqElBrXdjABAxWGM4SWyK6ENuTuH/j
Kyq/Grcl3swFdJiq9+KkE3RVEzinYBBJGw/qDTCJte2YbtQG9fyNbSLfTD3BCj8r
1VlO0dkduIuWtZRPyT4aYuhikUEnxsncjJCSGRkCXGN9D/TyQAogsMqNpds1fyr5
RVYSB9C7s2Kobptvmow2O/To1OaBiaiU3OssajJZC9EsiBSXd5NZxmPAOBKShqcs
DHX8tP0iU056L5n/zmH1vcXvmOJ8tZ/uljUDUQgWQsBF8wp4g3eS+WxIEssK/YmB
5WOwGA1MiNZFeto2fvWKUw70/wDtITjunSyCzdIy92K5efHhw1oLTOA0Y7HGhtNW
hwQCTTsA2FBE4uIVyJwwMPXTiIL3fqcTyRwoN4Ivq+GbWdY6GdOOdPgfghKXSksF
ioYgnilhTCQnR4mP2nqhXLWs756D1c3sEO7YPP/6vgq+Fhfs2aCRbvOkqjYuloPo
OQbXhpdZ60Wu+dsI/+u492MCl7PZgjomIvpSayawhdi2thCBcDzKrAQG08MSEApx
LqCVe+EEN9HzCFCCj7qNmbsq/JTP/Nljjgic9ZCthmLwUwTDvJWe5nD7BgFjwfkZ
3ThxfTKhEJMWy5j+SDRzfrdTLUxCnpenvvr9vLVwlvAP7o1rSRPovWKd5/vPrAOp
ah8Lk6w/tnOZtGIWZjmYLQCdVgPmpOeQKYt/VbxX0igCh+zUsd8bVVQSELYPwLi2
zxPIKKCHMg3vxs4STg2zjH9vb2Yrx9cBHFrv3haIW1k+a682xssp7BocKMGLFZen
ftQw641pXqkJ5/gaiChxyijqMSJqQmJqvANyrcdGcfslFgh8i8mrxEFRPwUAXAdQ
GJKv/UKLAlxHfEe8e6e8t1Q7DtrXEhKUUCHJoIQKngdVxn9qFbcnBIu1AIlTIGAE
K1LFN5CcSpIlqpF0s0eghm1BlXsHA9H0BFSVCzmz0ionINt27qSfPFeO5JEj1cKJ
xZBRp3Z3W66bXINK7t+uafRGFBu+6ivIUQRLSXrACVzkEWKNR4GzzVJUv6E8GSjQ
za3eaDHG4Oxal2Zh/ADUmhbbuHQCvB68xifztg/2+3hrBwdeMjNENt5bLJxCuYb+
34U25/RWZO4PTWHnOMYPg/ueJYc42bHH5qqc1p7WhiYrKuJxKG3WQ7rjYbhebhOD
SVVNR7craSdmFABWzGJ5Ij1tEO1kPp8rq9v+ZjjeZcNUenQo/oBdd5+ItqxclY+w
41YaqzDgs8YRNs05Q47SB2MRlLTZ5dCdK7lzXqEeYyQqKZTC6+ThfSHFy/Nlcv0J
mER61TN0J5nVNFgFEjeukOfoMbcEKhSSxA/kVKbyNEaZuBMTpyjQ2CK3BpINnkw0
ryM9gb/hDIbosKAJOuAktK/6a7dI6yVBQ9HxiR9D3U63OQ5lefiWd428kenjAC/g
evaughlMyzLBRJLGfmbdhRVYdWBYd2ocpWF+QatdA5RD+y9XIICjmTjb4ABfr25F
RbhnzwPZepOlFOG/OTjscAH++LFaTdjL7PlHPzRiJKUy2UMlTo9PY19cDPa0e5tu
GgLVp50GDU3Tr5ZThzc0iYmUtUuhDpoPE2YMOynsDbPYvknX9oD1O6ijwL6Z2eY/
caaX2uHxkmBazN/alEQVCG3TBrwBDoKWe8cZsGsk9JprhD6pM9Oz1fMS+sBc9xZk
7F9AOgLtMg1sy3JVTBep46/kMffKZVj9sFcVIZDhhZQL+8SWhQ0eNMgAYRLGlsWE
JrgaGRYZ+tR+XcelRo9PUG73o0wriwJ+oG/WnqtNVv1FlXyO+w0V9nqNN1hdXwZg
RrdMyQ0bL6oH0w8HU44b9b65gJPs4B+R4K3/ArAH4f07BC5OPzYYyBWFFBzPhNzU
vmZS7x+KRkBKBqIcGQArHAN2BEJXuEbcvQyba66mya2EPrtU/D7p2VK7cKG/M0ew
f08w6z8HqWjF9hmxTt6LZmkWrEuj/1K2+dd8tQp0uaFyBHyeoTeRqdekbDtUsqQr
G5q+qxy0fnt55qYBt7JAEbj/Eg+zYYr2XGOVpjwuv1PXk/2i7taqXM/PYl5sEsY7
cQzFPvrHZzxlUA9uIsnHT5adwi6r1cT6r02qaPoD6UKxQSuA0gGbKPMQS4YpGPH9
a899+KUj6tqiEEsC5OWlf4bRtOYsHNZOMTZwQvO3W3nSo1HdAp5AWQUse/bYQXXQ
+hEhRtj6GhGe3Vj2Et8ExjgjeBVbgkwqvck3FhCoHwVcZjaL6ahjVx6n4+aqPrdA
P0ouFW2T1iydXJXNrYhU3+gOt9zs1Vc1eEJ9YebOjwt2VbexIZu0N4l4xZSTC8fL
unl1Kd0qAjqkWRMZoHVlu98OGHFe5fm7hjBEXCgSNi0id+JmyAc4TW2i2JoM7gTX
fec+ZoY/5de5nYe1nqpQfMgv11gRdIYYzVTpqzeIQLYD7o2UiyvJFRnbsJUlFz3S
vWYURY5xts6UeVy+hGE7Vc2myhdmRQJ1kYrgJGzLiApa6JaB4IvLQmwripfDrT09
TosF5TTaxUXebp48KKTKLE8K33u8Fkrgsw8qqicVJK2G7eLLvhh3IkArgcZDm9ek
1tIWucy6YCnNfPL6CaCDayYeIUlgtz+qHHjI/yeaUpirElMErQiogFzyg6qzKBf/
gc0Oicn9Jb157uaJG9ELnngwFKS928ady8q/RilAu7h7qEe+KpJomuelejtpWKT9
+MF8tsDziKAzYSAGoKuuRL2n4VqXx50uomNx1FAtF0C554LNZAXed8FRlQTzLcXb
LDEZ0VReR0ZJyztP4rwQg4eSqA+1sGLxtZHnwbVl2bYuO5sD7xa7ZwfxxtC8eD61
z/dbjeKyEbAbP8mbxgTpRcrn4jeMA4T/WsbXieAyf9JlJq7EnTxmcS7RwAP+EbHG
ViB4GIZLO7p+Dv9+FQuQ099geM89UKWLDf3TXNfM37uZwu7fiRs/bXf8D4AUvWeg
WiNKdgtaXOwjSNcNgzUaSVH1EkJhA8DSN3eGuK0iY8cgtJsDB8YLIu6kpKqSL0E9
GxFL9uNkZmq69t+tarZKnZyVCvIvDh8+V+PMUt9OtU5Shtdndou0MXMoZST+z1V4
IZImMqGNyVcJpLMqOkFnQjYihsh9J6TFeUdEbg229DbBqmXyDjp4KcYiB8eRGHh4
dSdPZ70A/XmzEEXM6j8rHOjryzFzHJbG4aHHC95ka8POKgB72bL/1S81I9vGvj8w
RpZ93a7CpXCQTRmV/+Le5WqyIjLT26LjkcXMTaDaY7WeqFDvxkgGc7134vMCEhxc
AF7EQK7iSz3lopRKHR55of/YNdTMwe1N1OBvJMKhjwLf8HnbBTaPnqB0ewPWosw/
7Rjlp59yFdIzwZthIVZ5UIzEHcgyV89l6eb9FEU/fv9ZoXDfGn3CY5QZBTS1jx5/
Oce7WB6QF4DuM8x7GbGxGU3y5TuLTBEWCaLE5YBjngF//YFziL5T38oxxqTgG48e
WM/h9vxOfZzFFd6lFQc00LkZGHCc7/MKFxiqmJR6knsm6qRmEYkpJ91mUGZkfirz
bGGltx3lfria9FSPWlI0YCEym74+fJDn/c7aBho48xsNwavQGbCh6sKu3srfdIB8
6+GZq46jjaS+ttImoSFclZwnt/3S7AwU3gAaZfHny+2SK9G/r+4BVlptgP6vhIIX
AxvbrtWCljxCWZbjmsvNGn6AsTg/PnF02ZeLY0O4MXLBJR7yLkNPLS8O6LFQEFkn
P6VFzZ6KXmmSnE4yBkLbO6wV8/1BmOg1ibv9/bur4PTCrBnWCoprJ17bq7/PfBIe
EKsolXb4R6KfNSYN6ZIrDkH/+r9ksoZL5UCvXsYMDEGeoY6t2PGAHgV+AC7sxiyN
/zuo+9LRozpEiqGS3s+X1wjK3Fj93tSk73ZNSn0dGdgUvH7tAul7xPocZV1KstpC
WYYn0wj0iGKW9UEOUZMcxjArrsKXTp+2xe1tt4oMl/m45MErcwSfi9I5RgRXeyNs
ma5tzwpE+19A7ZtKEwMJuOC37tMu4F7leW+qRel949+AmlKionQYgDbPz5DjNNOU
K+oHXETGNuOjZ7cTeAYrYFimD8WJdACTtyvEzqrOo8CQgffLiOG/twNQVKoIiaEW
VBxYo8aHs/YD6OVCCNrNWhKjwNmQf1fMRwA1P51IrifacqyHdlk9Ql21EEVft/Hv
AhKy723Ugg9Snl4My0nB2Lkjpabk0hOQdjRHjyXIq1oDFaynZJFRGSyNLf8xFRRC
G+qHFLFWqszh8Cl4FtlxDDf3xMQGdEsGgkNm4X3vod1QZp/QzOjl7vorUBIN5Axd
57msge5srPq0qvWdp8CI+aceltX6d9vP/k7nYQ4qqOGzU5v7xt50F+iErZ73B9vJ
jn5rYYXt+fnmnGgh0+FAXEbsRcCObIE4QLhYJAnE8sF7ZusYe1u/050GikJu1beB
AZ23cv/p2bo03QqpGtk/TWDkRMkvcEcdPxED9BfhfPLzHXIyO6gYdgHP5uc0LxdT
StcN+oVH1VBBKlgL4oRrjPPA19J5kWGPyLf2YIxuKkWfGZYQgoDMWPAS1vqs+FSf
/ohpf881IsqxA3c1HSCiTaS6KwnII2tJnNH+u/4CsSYEJAkrD75JtmrF7Ly2uufe
T2yyy9wnp8kDITWdQEd7RyuBxBdxyDv1bh/GMw0M/fGr9Sfj1FKkdVLTHQd/1jYy
HdhQgslxOnkN9Yfn6P9U1esTV1VuYmnV7U7FFwNzniiclS9uqOoGiseQ4+o8nqoY
vzl1Lsc4/Xxq/0cGBRIT3vvRbXhWzyL0sUYPcOoG27Q92EERTJpyej9RptpGmWW0
iL2E9iUiJFYp5zOdZuatXrdmjM/mfnlJbYYPXaARXhV06V5xUEE0q3rqYez8NS2m
t6sG1icDS8i/MaiFMubU18ZtnYxaKWbwq07Qt5albVxWTQFaUxhFiMtd0ADlrKxG
Rk1GvGzIMVCPv4v1wymhMi5uTfwjL/Qb2rx1wpoODZmgaPyjjxkTY6pRVc7TZEl7
x8vDkMSVcqFN9tSxvXFybL2Eq4ZvG13W3+s+xI2WqPx5Ttz8dGCTovJFfrPCSpWG
HY7bu0UxiHkISKGVIn081mAHFBZ9cYfn8Q3NwxKN9myYkk0aDd3+A3d1wSgoNKQs
7Absc0+BfNt2R5WdwTC4/FBf8Le0OxxUVaDSr8cruxLNiU4sQXuiyM8jhvpGOzNE
4uc8GsE9o6KH/kdSI3aJDN0049z9eHKlK/vHGYEIjSHuODDIv0nWSnJjLxlq06YK
Ow/s7pwXu21uSr8aGYd32vBnC6XDwP8QXVZP23ONYyrFLZtdvkXqa3pvva6NWU7u
vwXUk9rBvMVgOOnJj6IROOsJi/IeKIjRtGtyBAY1uwbGeHcMYRw0Z9mewzltj+UA
j8x628VS/KHsMh2UJmvNyNxw7qAuoZ6IoIX2MlnjAGvQ7lveSSKdSCTzkwQV9/tB
j3bmsF1fhCOyFG2mY8Sn9lUhnF8rVJJAbJCdHcItdAJ+IlgRTIny8wY+FtuABjzW
8y4BTxO8lCVHmo5BSiHXV/Z1xqzRXKvNZFJn+gQYSmyLqfzmu1qTooZAvMv9LfRd
YKL1iVKs9MTuqmUG8nQMA3g/KvIM7js9UTV9roaFNBlV7BZPVV/5NIJkfwot57sb
pN2DZkMlMAgEVyJrQldmMGmrjy+Yg/FLi0NjbvI/kSJ3zDpGQwO+/YvyD7W1QrBh
NmlZWof+yTYfZ3KDvtH4AT7ZSlrMtQIQ7aOffbHYnefgE7xp/2CdkhJC4J3clLuM
wHiHB/9sxqlIbfgwvbQMj3yTKQgqhEmno7YV7ceR0tc0RNZLabJrgLPUrbAYq0CE
IMo+PHlQXrCCnYUnIsFfWbumalHPWSE7pvislpO+WqzsWbQqa1KFm7KCyhIWWaEd
sjw3QbTIIenRi1e9WySk2oANwBLHnGozWNsC7/Uv2c7MDDSbwnVah4FV+3ABlFFe
X0WtTHaPpZZHPHQhQoWofD4Kvkz/021u5s9r+b/6bbwKnIb8Z/3uF3M4IGptswlM
sfREqHOsEUV/XnSXnGJWIH95XF6HqwialO2h2o9NYJSIAz36gyf8arnJV+CEXV2G
c+nNe8UQVqv5GuwTW2U/f68xryzdhoOPAQqlfmW3+6B1SXBG8yGpWMxiNJVKpW1B
X1FG62lpYaqoFhK7P9tbMYHl3i0enM5o1qrYJwHPd5KiPO72IRZZSRkK8vp8aopV
mz1LGWniGX1/CcQmZajjLyE2+g2iyAZGg5tD1rCLh9Mkgigqexzu8qPmeILO7BHJ
Xb5EIvhXqlLaexZi3YcrspEJD+PJRz6pEQVruRrdoIfjqo2a5iUwfQx5Xyxnshcz
UuCM29fvteSWi2ZAkeQQOK9HQHDLtdvNrcFkw+E7I4slsWMcfN3XxSLcZ2jnLw8t
TheM+lqlsPBqEsA6oDwWxQWoHqyQe6BW2c55SEzwAoV88F6RFW1HCUxO4nIAi7AW
uAr/+MdP8WwosqnfbtovCt194flMpEuvjwGfacy2fYJJip74NofmZjY6Z05De6Nk
UFSpfTcVZrszTkEX4sHR7vZ+U5h0OzTJfzvwljrUBjpq/iZ6SZYaVEnmjWMMF5CW
c3hht9sjFpXiDUxhHSoL3tpH7jIZHjsL7+/xV+BE0qQsDLPOff2xrtPExqd2f7Vp
mxOe4xYlqYB1AxGmissm8K9S20ObZ1hqEXNbeA8TOWtJvsO83jkovzP8VRQXTvnT
d/ySneECT85R049kWKs7MpWzN929M3PZVYvAJzZIO/XC2b0Jv5bK14IQiXmcK29g
j0bcb/ZedsF5FV2HegDuH7R0mpW8/dYEMFCbAaRkBWR8hxEe2T39d5tiOKJ3b+mJ
vQzyc/Y6R68jm7I4bqqLwElV4R6GzZ5oWSDAb3A0JSKzEKV1CIrHuLQJEFvjPVSO
jW/TbXcYxZYX91XudCbphqXJ7dXZxMydM0eqgG3c0guT6/lMitjOHKEldyWZzfUd
QPldQKiyaM9b0zmy9MjKyIe6NvewqIDt/x0qmpS2lIp7JlJNfwPn3/Uwc3AuaoLW
O777FjlS0iJkoBCUAnHUzQgM5dkpF7Mh25d2elV24NJc5xJWIpWTOOTzvrwFKj9c
9sxloCfiJXAJfWPTztSn0pjNeAp1t5eOlrsYeuE/L220+CIkHpnxdyZORSApM3xp
shXOpKUH3YjtdUt7nuyaSbV7/KeaCS9EfVAGQFpLEDzceqMyR13d7+F0b90zKjpk
fTIlgJEJDUDVESOkrVlyvV/988ltaXrnzMEgd6LWgiAvQCX3Iy1TkFm/YMqhtVBs
JTImuElVLTgcVUWop8n/wU+GXJotdewQbJPxx9qUt2v0LbYKw/nlPwHz4VITpcCs
K5eEzavZHHTNDApX3W2SwlvI36ME0OVUVT72w43FjIPSow0W5k3gfld+4cxXHM7N
0HsR+fMSkIhpjGexU0JgUK4MpyKqHhZuDsHPojgJxr404FYQ71FEgwFNZS2YuhsL
FWdI+TOUn++kS8HTAvUMakYV1i22xw18gZG3kwtqymfQ98QJl+4MEzCCoOXqtKmk
bfv97LF5hMamjRg/2VEq2BHR+LqBxYiM9+WRo5RYJblVrLdyXgXRf4h07kqMWX3O
6nw/Dwcdtx8Z9reyRzN9jc+53kWVkGteLFNmD6y3fUXEsuYY2zbDlysNO3NJaNtT
JctRDGm3rbhIXhModQi2B+2fnTOSM6UOLZ1X7XDqtqnXplCeEytsB/XTA2DazTQ8
NchYV0NQnKpOvT3ts1bxJpBH5um2+yGypKWLbZM3KJFAmwht1GhwlYK2LH+64WEs
6+QfnWUL94ClS8xK2w3uvhQRAGIDka/COImUzCQfey1PXqmGhQWf79QT3VSWoAys
A5vWku+DdzsXYpjgr1XRurY/Bq+C6jGUhI/80j2LrvmGvmWPc8xKqzdi8BVtvtAE
Y3n5iemjyWYSmturF1h85QBurUvs6kWLPt2gllVuHqfMaV0ALpWkClB5JWpVnBEA
AoDax2j6zLFEZEUQ4JBx1ZCIl86DWTWbJPZc5yw5AiBh1h6p2bbb20KCWifc27Ox
dTilJAeOyJn76haXObuH623A3zN1Lzd44OL2SZg6FIb9AtQq8/kSXmFPLpuD0MvM
MNfTaoAZp6wZK4+Iq4kh6KAZMcGqsU4fntP8bG79/OZJDyg6L/iZoIIb1DCn+vdc
M4ElXy3iUtZbWox3/FNL+q/wERgbemHfFy86cX1LVXjtPRxzolzG55WpTToyA7FT
UluSc7TldhdrfiGcm05MaWQXYT2UUmoalp/nhOZ5opwcyagTR2sSlf/ZEqBaliPs
/YDXD8ot0k3vZDm6fPSLy7xuTHuVWb32yoAj0l5YqOW0RTpG4YjO7gIOMgSTi96p
AbN4HGZp0hxKXpDg2Bd4iDYbACFI3Vwyz7MK+u9a0ZnXAZIOS139dD/YnMu3aC3X
aodtdtHcjhQNMyJ8pP0fkQV6uAkAzD1xJlNVEJdVOe49WGcfT56vslyulsW0fUL9
Qg0EQPfTqIWBhBWThkmX6fkBlDMkt59LTWGBSP7+qnqkeG6dUVxfZ4s8nFlzHLJV
qtUYv0hlXcqwfjEJaoKzhQ6oItKhPTZy+mX8Bx69LLUPPkD9a+PZGG3jXSg7d3cv
BgfgwRcIThz/4cs3ietsj4oJ4d/nhXstqEt9u7DGXTHf+OqZGKMshV6ZW4FIW0sI
fGEn5JQF08xw3hunSoNW0YFhv3F6NtfycxSG+CU1+S7hUpqgD7L06K4/2V0ux2E9
MiuE89esNbnrFzaUPEB9pOk/6T9JE+QD3OVOBrzVIZ2UerHIPJgRql6thM2FhYWr
C7dbjHvLAgsT6n2BZHLMHMvlycAm7v5WLJk5BuvazbthtrVxagKozT/9T7uZ4Kpf
1u3JQUCYetPm3CEFZUhTuYfVRQ6HuR1ANhV8+Ocuctft+jZl7Lu131HNJJ/maT61
dWQG6YeawvcoDk6f6Y0vzNmA5RkXlVDZ7JKbfyyQ1XnJqimu64tsquotlEbZ9Kzq
+zTH4V3Z/jN8EEXkxHvB4VEuwQ1LUKeEJnShsEox44FOr3inif1z9I9LPh79KAcF
mxgT7uuY5srsuruCqm1tgY9Ti0pMoqMYJVO/WUfrYA/vaQY/S8B6aNMEEnynLVIC
QF5A+TRy1fHT+I+UDKDIWXNhAoSc9BHbk/1BkPmHoDxnLeJqZTkzb19EJdCS/ZvH
ZtmniJXDFlt/iz6UCZLr45p8FynAFM/N3N46jyXJ4Z4AU6McB8JQIX1EiILAIsHV
BBG+tYBHYKt8dgC2rspNuPQVcAEemGbbPm1C8AU9zndkMypkN0IP3KCzMrJoWEeJ
UZwPCxf9N4tA+cNGn7+45sDZW7SEamy6qUEbP6Jc8EjvLAJLgMWBSOPIxcs38n9v
wEteWOP/avldUvTYkg76MrbnPT61bxWXXTmjxutwtMRv3EMVZnybyLNzwLYtmCBb
UVLCGyvjIXrKaCP+yJSpMwV+ODbNEG5+6afWKq6ClzLnAApMo323Cw8y06P9qGVj
kz/BmoesyE7+a+r9/6tlnxzTv3PZj6UvpwDX/h9zFX+2gki8nJsrz6g26qRTcUnv
iDVjGPimb74w5YhQHwcbAtRYqHrENFnMbw5+SSqyOqCJ67D8RUNeAXXRHySun/Pd
DYjpQrtxXxbdOjpvmhFY4KbtG4KAUJeT3o0XBNgSRKrkqostGYe71yXhlh+5Drzf
DutQlry/AQCifn+8PoRWQx2IVOXVWgikQ5Y1IFYlaWf5Cx6tOMxWmaFzGMJHM+mn
C4wlaVu4sdnEFGnRTtk5eHrObYB9xDNNwPTv/vv3SggHT8Q5cEdFmDCvNY7m5ZLG
ewYlenPGo4sl9IyvXNZdDh/sjmC3ZKeBlHFQDtjh5bY+y46W4xBPJ0xYFV7L6SQC
4lUpZb1X+ZmneDbRkwk21u8xAdxqeHsNj4fp0bp+faYzaOS9nU1CcbtDNJF0BhXq
DtaDlVwAJ9ae/Y+i917eVgRPBkEAf4eXc0wcNDcn7HOZXDaQ5+gfXgI/w9T4cfsX
dwF9v5NCsPTAVNnwquM0TvcqI9yaEkb/lh5tXZI7+NP7WFVJQesH58RwT8ssHykF
CKMHYbpofpsc8/RdAoRgCfOX0XQ/IeCpjDfX/j2LX2qqO1cp8iHx3pb0Gdq07Wlq
hnWDapWfbUgHfPemfdu8ca8L+vD9+FhjZgxTWrnh2aS4pST38wLbNwKW4ya/elH1
H68bSSrYAFCZtUUBvtddK1ECZd3P3slfg/TTfTFjONTEAWzAVaf7zobq6mh7GE5+
QYQSG1FCnAveTNQMRta+upwD0Fovw06L8/tVBejgFL5NILKALEuh+0ES1dRTwD2n
lqaTonCo6iqt0XloTTQlvU9QOvFJqxbcSNVQG/XYhwVzBtq6H17LE7el8HzgXBt+
/lm8DUHr0f1U8GMtfFqBKho9A1gt2k/lg5qk/bjV06G+h5+mipi9/NIN/tENZFtD
LBhN/oeP4FbtMS8hP0Tcb93LKMwPnwfveOqLUgN3E7KSQ3EDvNgVPszgNxYBOGer
fMViNKIrh2O5jRLHjj6YK3tfNT99hoUpbTMl/Ra0+ljHGLREufL50m231MkYe5yM
5wnuDvdHS9/3QFVqugkF4E0zNz2v3DQpVYASAe+yDu/Gk2JJAPO7bhtV7b5t2gZg
+h6sBYulAAx107pICGMeVeqEp8dEJuXR3iwmj53FoYSbwLnBgK7cc0S193gzjT/I
Df+O5Tw8xsAH2DdoiH05MhZL649iyHSk1iax72P90aUKTUdG4r3VuASs3Pz1wtd2
z5pvxRP1Xnh9JtLoo2+IeS09g//7HmZI5RRRnOZO94/PGDnROq3hVBLg1xD0M8U/
G38Yblzl4Sz9ZH+lt29B1G35vj0lYjzEXT1gCWAAE+Gj4j5hlzRmWaqpBTXOLWdQ
V01XD2SeZv5G28EAPhS9tMVHD+A8FrJuAhopB/Bq3Vp6TLE98w5ZdyYTSBkeaJQN
0mXV2fZG8ee2dyd2KKzQw0C8wnPFn3sp2RXAi5tKe9WPYDAV12ENOGh7LpR4sLbG
LXJXMWA89JGz4lacbaqbbEAi14JIwR8oCHeqb/m2WslgyVk+exlWSGHNiD3EitME
QFy1dJcUdl/6lfX+F8SRBeFYFEY0wTUWX6SZb63HA7jx1Mh4pFZR/FLDNBcSl3wX
rd5ePDl5gz5H8fLfvy1OwDHqGtOwfuaffmNNKNGbl6cofh4mJtI2JFS1XzXERarz
kPwzgRbu3/53cHsc0roMe1GMTHqB0o5RlQgnTxeqxZf2aLoR8X+kFDKUYwlKLkY5
BYAU1zT704CH39FQzBxJG1ln7bET4giCYLhprsSKvsDSp3Z/SjmZm2i56N1MPlLi
cKRHA5BkNC4FpBrElK4dgpm4KMXIscEEvztRtKyKpEh65P9Vmu78QAmsV3KoNMqG
jHamv6/EVjKFUsEYaCtFklAI0sEYnNfNdLXkj/qsrZzrPY4gUuLt2tZ1JAsF99yH
7PkCucyV0WVBZHZDtLKGhtIVlV58h7RCCHOrklBsEyhDPDb6qI5cKXbVKaK3HjP0
mb+yJ1w25YgdcPwDQqjWArQo7WHy918LOeNy6XaSE9giDVd6EFItY60v/5FHhVGh
eNid1CFHyJZce6Y6DaCKUitAG+QNIruXjt2qFjeJhCILQm9Uegb7xo613/qaacES
6aD8MyettAHNTy9Tq1uG+u9tiKWVeBH/z+wVx1aypmD9Ks1jHjoBxE0QpeArxSbi
xnxftgsxXTcVePlEzpgTPcyEBP+19xShIinPmO3XRtt3zis1PYtDH2MzAmg868eS
1PbUzsWM83zfztE2n+CiroDqugIX2TyYa1bPC3E1qEcEPxzZcR+GM1KmGJzwQ8AD
85b5j/+njlEuRpA93tR3x5Ac997RMLcpRb2FOUpmEQjXdsFz2owfPGUTdokCi++4
8jU3F1szgSj+mcJvUyWE3QcGALTeBypI7s+CiSIGXYT1GzMyoUTBCqvnNuilHhYB
rjxRbivL0r4a5k7GxWHjyG9AteNgpWE9ClYMXT+VWGYHQBKZQnXnOZ0i44uZ8OMj
NEkAf8nryh6e4L9plCR4whXKstyLe/h55mQBwlpd3dXzFiCnt30SY49wK65YdLwO
Yy838PLbkl6sdoPtdOUmLzsAycD5/f2wVDwyKHM+tzvXeoUI0IsGQcmJkv/AxIiy
vZ/Y/rFc5bLvszS9CdiR7BaPKytSIcZJ/w1zQuQBXJrLRfbJLXouYBxpPCvZiOfp
v0n7MKDhT5RYHYoPGBDuYKMxWbZah0XhFEDFQuzalgmVitpgz7aUWS/bRhBvX9ca
6s9tt4v/97Sw6TNMolvSolFAYbkUeMJ0QuK9qQNlPz/yu87QkEVtsTInRGkilxWg
WviXYvazJEGe2dZINx97fgv98BF14AAi+klKhfzIhP/InJdA7vVbfAqHeCqJd84v
zvX3XkStUYTSFWlFjPx1tuxjqeRMk+tKtznxHOU0g8jBQ1ykUGxGAGn8GgQefwtd
v7JRDPnD2Q/y0y7E62Adfiw+66G8+FIJZeDUI91soWij/b5dgqLR7674D/mMKFUt
gY6c6YKdni3O8lEhe/kZNky+2wFjCGMZpK4GU5tBxg6Rz/2CXzpWAvFwAXDAaALJ
RIdcHd+hCUxn+MwGuc6ToPYgraJdV2XH3F8aS+BzH5UlMzkTQynBW1NRVUhvLwtp
5nJj2f7qyZLrh84dWIeITTgaDm1PIDNNiw6QgPLwbJqO09Bo9/vg3ROw8WjfCjTh
TkGsU1d56t+DtXv1idA3WN31sf28Sm57sCqHMdoKLFgYEiSqtU2Df2ho3Lom4cRd
R8Z7nEC2Xx5ildg0/DZZK7fBR6lY9tprU5C0ko4kWcccy0zrDai2ki6Fx/DZo2pK
fCHKngRGVaS/YwvtCqxJ8GB9v5MQ/Hp23gkULqIbBUmckcJTM6arEEgdt8beD1uu
WqiriS5oGDqkd3vUft9YYWOv67r/w7eh8uOQO5rU76WM5MDg6KEaXQv54qJ35PKy
2GpN+lzRppEcrT/MaN0Y+QdbS5/SPz9MX7ZRseD7csSfn44Uf1WuSERRXTRKblKL
J2T6MFTcMVwWXL5O+e8MsyExmE3qVlaiyx9LJDkG9DmgRbObJrJwjkxckh/VWf79
5iTYPhukwqFz8XXAhp25PRzvH1diJG0nlPWA9ne1WXnvtYbAMrauO5vjPgGK1PcQ
UhFvA8GPxPyVTfHkdUahjk1Nhdw1416XQUKXXrEVBgje0PNqe7E7siyhr3D796MK
WXuq7jnXutYAiYAbMkltv+8RuHkugFeHTO7r4Kx8DN6xDbu5XMaPWvmIS/9dlmyO
W3DrrOY7UETZvyBoPg8l6qnbO8OPAl+eSTc9YCXoO9gv9Ir3/Wh3Tz9VYNo8ZrKI
PBnrLSddanLDBdpcv3C3HsNgy8I5ecVhvq58lHkD3CYxgIt68k0l51IPYi23C6CV
+RRnwx7+a01ZaGfHfmrlhL7/cDzYYzwTnJh+QhoYp1EL2QP3PkVr7kft5aBbPwtb
qkkVma8ldp3SOjsPVlB/0UKSC6wxfT4KqCcCvu9CWYKkxirpvBZQT7hlv9xSOyql
E4W2GyRo4OOGnVrxedchPluX0cVvi04QVmLwn2y88lXZtS2ZfxFV7xHlgnxzvu/Z
TtDdTG6iF/YlZQ6C9iODVKly2M2c7iLSzyitViubM0BBHddwIVEkdKo3z4xhH2n+
LXYmJvUNgSmP+/ItodJ+0t9Fdrt27efr25mF5f/Wwq1j9VEtoi2r4K1xilK6Ku6X
FDCviZh7sJbcYvdtbO6DnXRmUKBbpHiaW7ab2tj+/XvQGKIvTM90SXti2ZHbMsaq
5yr1NijN75R4eAIXkwszMdBobAeC9TbNbnMlNop8pl/XRNoJkNa4SbC8WN5kbQH6
nHidsgpql6XQtblgg3kuZc0HN160Df3/EBgR5FOUnn9KMksPqDTk+7+M408uKL0f
YqcvAMV0Q02GfcjW/ZgBbqTMoJdUIYTZla6b1kBNkBuW2o/wIcpWIjEpkMBFO3X5
Hi+NfYSH/RQcMn21qb4cSZMuMt1N0FOglWxjI4zKYss/kXhsR8tQ1bYdAOVUZ9mc
t241d4K8gkSLYCd8p+LLQlafT1njZqkmMApEMyJItZ4Z8tIChX8Hp6FKGqTwXHqG
LERCdGNBz3BMpnCVOVSYMtr9y2CSkv4+beuKMU0G+vJinbavknZNcx1m79eBlwrA
ukSnegIeWD37gNV8GRDYYGXrE+C5RpykMQp3cw1Yct+Aeu9pO3XqX/boQ1iq4Lct
Eepf9wrpJGdwudYa2j3qFq5n2q68sWakrwnFeyBkKylWNKKotB4HJO8yYAd064s5
VUBrudV9KmMqKBOCzAKifiikPVOXXZXcLr4c4fmAFMTfYqVkR0TMV+gJ0AfH0MBj
+KoTbn79OnMZhtXIdyq4qoSLgi2zDVkykAXlW/lHT3IguTOyIYbMlMnBDJYBxfxT
vE47W1/bAEmJK76VKXvDkUSUB+vrxlSpCCfWQOhGjTu7ka5BI9SD83Bgi1TSZjQl
dPl+iwIZQ+15qwhwrsxJAm2nMX5Q2Jbc24AAHxBlRk3xMhDrg/Rz8RrXlTXOP+Xi
sD6DWpo6Gfzj5pW2+vWszev2ftOW2VaToSWj7J2/szDMPyMP4ewn/JL4WhtwZFZA
1nX7otPe2UPcw40LoNYsqYCCPIKi4YV1G4hTd5sgFFM45NtSL94RZgXWpHnN8EdW
v39sX/lqfUsEbw+/yLMUXc46tIKtFYEirYL6Cubw7dRh+j/3Sd6gf4mA1KdVRYZy
tr/ivqXQN2oDz5r8S0P8Abub1Kph21+2pZiqEOTnqt/JdCLjPi5nl6BvnwZLYuam
uF2CHeVsfk7ELP4rdrQbpzH7772FW5X8pJ8Rb3UUB2sz5f1zU7NhIl1X67xDipTo
/Ocud+i7zB74gbe3xe57ltw9vqwi4XH6cXxmokMn2gLssAigYOPgG4IlD//DNyNO
Ha0UGQOBrsYkk4TDgQhcZPL5u8LQBoWKy+d/2PzapqsVu/vCOUM7LZC2x1W1HVPT
iP5zm023gXJDgbsI1Ho0HNSLTjT2CFEiai04gM/kapRHPKea61JVHJxuG1L7nCi0
XJxl/no6nXVOzIqLiLMeybeLO9J/EI7arJNscUgaia6woKtC5UDTqkfrACOMOuEz
U70hQM6ayYpAYmAzrzWO1FAHaSq7K8F/ALxevTaJxUrqZi6HeZdP6fFi1HdUZMlE
hpcguBmLZx+RBbQiSkGG0MS9YtAJV9/QtsWtpG+FJtcTwP0u0O9NCFedG2Zek5fY
ALhnTtcufKFCOBEx/C6OqRhJO2dP/yLDiqLbHrm1eF11JsrIUW8wxG554wcxZTmZ
g0Hd8w6jRoXeen50/t9Lix5rM7/pSIBqbrWLfNnWkDPFjJNkfrepuuq7QS5INYA0
pb0C91tvwijFsvpT6hSLwzKIUu0STVN4TpmDJK754rOp8qD7ljY6GHxcOg3IjGZ3
rjvidVT8LeqvM4yGBi3qYKlKFbcYn7LMs9OcJyIuULmoJ6Gsv54CTm9w4evPDAJN
KW0l8/jryRrBou9jDurYuSeRIaLT4j+q0HJlZK567pDa2MADnEq2Y7bPL/fGVHdO
B4VWC051mLiTDi1puusZZmH67QozBudX7u3WBos6BM8o6gfpRDEl/mM3tBM8TMQm
JtWefZWsRR6GM8NcRTKdmq7tGLv/JnZZWh2kOpDh+AMSNyjHCG+29DKzZdiANL50
N+esSw7dIR3EbX0admUq3Q+T0C0KBRqG2pIf75pYBMhXUTsMJB9rHn4cqpC9wvG3
sPg5zN0mAFhotxsb2j2G3gwIBbDaOU4bLr/UYvl7qQnc1NPlpA1zMZKyjCECIP5f
KMg5662BJlMDff/JI5xagbfotm96dzd2BDFJE9pgFJcdY8ePmaFzXaGuwscSDoZi
J0agnG58YrDyUHeLbyWq7jlBvYJPJ61VFWP8rdx9sbpWWaRPjxS7wuDCBaMU5Gau
Rn52/g1Ut6x5vK7AXAG9WedUfcizNAsbBDtWbOM9cDGLD0Eg2bJsS941c1E5f3fy
kcJfNXIr3vbfyg1DMRvQwoAv1CxSH2n04nX/K7IR6nTEqaVgWy6d4eF2+x9GCpIq
EMOQQatSasq2LGbPi2l3WA4vNIDCq14iNTmdreANWJDAa9hHbQi5uAlw6k+RWUjT
5RPy7qLEvPTQmFhn066iF+jYKjDzPB5IvNM9ZBaZFfB2eAJyt/GkYNP9HxSwEhv9
xQ+51bj0WscSS7JZB2aTlYDzmlrEM5WXCnJSyTV3KJrq/qZ37G54tpFpW9vID3I7
qniNvpJVIl86JWwp0u3dEimrSGm9QbAvMQkinvHgnurypHNNtncEm2MJDjGglihK
fRqNBljFx/VoZkjLtIcZB+B+J+6V8sIKGyFyVRHEE7/xoGA5+3y0ZpSHOxmQHNhs
2V+nANsAz4PGvlle40ibc3n60COO/YztQEEjF6m6uBJ+1qGkSChLP7lqWr4THG+x
RhYkWVnWDR5EeIHb4vKyBl5vz+elvl2zDfrXhpuLfuDITX4I1LW+0vEQ4ux7FF11
MHNEgKSknfzw/ng/e+Tbts6X4zVnZMrhjr8e37NAQNQnDQfZtpw/sgY+/wX8XFM8
GslA0sgKi33XHtizmUaQv1+sR4U01q77rRAOSCw9yIFlw3Ae54K9OuaVy3m2vr4A
X1GBTdmJOC+PnNgSFgWf21GqUBwaTDVUuPsGC/8L4SDgz3tJfobT/QVc+ErrHHiz
PYNJL3qgtncAaMOGBjKqJO3IfFAh0NJlnu27dlTpN1ooOqL2fE2iUbcgA7QNIda9
jHi4E8sPeoBge9ZAxetNBDOLdhxu5W2+heBYWKtrXf2Z4xMpRMv4K98sZn4wb9dk
nI1aqkBZEdT3AJ5Kds1U39SBcbCp+dazTu+8zHxDFd0rxgXmh767IF9iAqclDbPq
fxTxF1UqJUpeT7rIEqkvU1uOzq9GvEvF7ty1XETX4wOwU/Pg+8hbTX3EiSHV9lV/
4bjEbA5N7hAVFIWnAybyPoYKOhIw2uPClO4FFQFGZzWxh9b9uCQZ9/9q9bnMNgt4
l5zk438SDuoB11pLDxheD0muYp566FsMOXX/jEKa0jg4kmJKrib3TaTEmUh/sAOx
ZhoDBAz2spF3bdGGyEdQ882V/KVVVR7ujkdo7NzlrQF8Mp/BEJNs7L04un73judt
zuFbQKD1+6hP+9FL8qLhsBMpOYc8ULSvmPWmBNd9IZhEyajq+mcCRoeeirUcDvOw
Wl1Ok05HE2d4z3eTZYM3kHbwVJpEm0/XcxHGl/QyAmSPjsHJ0E+JkI/rSC8BCT3Q
DYFLKK9wnVxK+NsizLAXncWYnFwR3kSZFTxjj9LCvGi7RvhzKYwcksgF4qngZayK
FeLI7kI+cJbDI5sY22cueDuvPe7QoeWaYRy71cJvVci3iGyN403EzvElCRvlqYuz
sqJ68NUjF0VTO23tqr6Gbjj2mDCd8fpS3riFDfw2BXgb1ydPSkXsa3C+J0jl5VBt
rDWM/S1ts6nRqNuXoQmwfntoaK/ySdIr4JS14anecO+NnoADXys1x5UGFNC3vVg2
flqi1RjTQ+jQ+s7UtIooWYUUt2bj62JB6ddAx/tmfRBkm6eNDwhwtknJqppvPI7u
TcmYv871qGKR0RaUvhcO9n3x5OqiJjUDkEldRG3CA0ouDncBAhhA+nkoDkFzmrFG
XadjaHk94zr1STfGGbxq97BqfkIigHfRol5a763TxZ0AuUk7fPYnHbFZWPsHlPtb
o5ryCQqadzjX3UcGxfHYXojic2if/8UoFC1QZm4wE9Fx8Pd7uryJClNmKcJ/lztx
qRmM3sdrbk1tXTC1lufpmrMo5y+Sa5HLnbBhSpex+RNIWm38KcvjR+wQdO1tTCgU
ALeIqaDg2s6ApkYh8ahx/7lzM8zooDzaYQEO4+lN1OvCTugDMgnKEBKGjPZfsbF6
13cs394S83hhZPCA67GrOf8rVNFyMviAPqJB6A2rkzJGlcmN8VYrvsyqjeG/Q0y/
N1BAsYllVPF8yCvom4kEOtqPZBxOjLzWpMiFT9IQoSny9lyj7paH5W779b0lR+u9
JzhUKRhIgEzD7z7PS9dleIx/caA4PbqvsXbbI9bD6cOormQGOS/qa/aZ+2/hIvp1
AdEFHNjMlXwYksEhXt37U+Sp3LiZfqOIghIgns/qE5KXbvlnk/3NyFdZeb32GPga
EMcyHfKKkELpDAPSJRnyA5+ofJ8BF6l0lXV4N1RJJsqnzHheE45y+t4zlh0pH9dl
oyLVlIGTigXMikTWweO12aqpyUIfxTPu4dQseKEahdu9GygqsnPX0Yvorsjo25oj
OpzT2Fk8CPDC93RI+OYfMs2/yv/SGqx/lptn5rUrtI3/6d7/YGAFgiu9wpsDXSmE
K6jpB77xFviDHItLeIQFWyDGO5OvCrgc+i2/CS4Yye85kNF+OtjzVBC3hReYnixJ
o5X+02to5F2aTlq2zUoXxLT4KmCaLcHCIMqDaReQt89kbkmc6Vl6kHXL+72DPgvq
XuilCz3aKc+VxVMB8drt/yCzE1lvG6ym0Fs2J3HhU+Rd8kGGVwhlKYouypUWCxz7
GTNbPdzA+csLfZY/kZtNPQYUsVeaQdoD5uTPaZpQhXr1HwZ+lF2vptVtAJEKVfZa
Dg6mG0peNEJRREq6dQ/Tdi8ETYf6BuHOthOo3Fx9SkES1XXlY/kE+CjkGo82N365
fDtc2Tm8Tmw+0ErMireuDrGye8jOfrwzrCYQ2gJq6yp+ZOEvpvEoZ7SS/4rg/bid
d2CMUgrX62TlgtHT6qrFA6NWAr3NVNRqK+/Qd1r7FQoWyz/hoSFyFveXGNzk9xYW
so0pIjWkMGLklDzRqzZ3ShhwWMr9xpCwCKaY8n/ghBH/tHczzhOVO7QJUmB4KNzC
Nvp54Vyijb/2P0qmBwShC5TTBrEQBEGQtMd4mpFFOnuM4y2gQRx7UsZJ4AWb9JTL
ASmd/5KkLYGNuxZ46lsyZhLb+UbVXdU+NW2j17XvmQ9Jli+RwemZ7JjwSflXI17+
ApXa3jsxs8C82L5DwUZYQaBu34MWj82CY7yDv8jFvZO6h3AYHj24sJ5Vv1dhVWYP
FNfSoslhMtLVAa2WAXkQd1lpGIvIo98spPqN1YKN2xaOER0ST5RiGGAdBfLdAPWq
UHz3pX8NoRSDOSMEwiSz9V9IkhCGopTgx5g/74eRYGAfByYpsleIQ2tOkdZ6EEwa
sBYqutsuaHr4gSHiIVfN7AuxRK1AUqf6G0AC60H9ySXVrTtE5/3JDIwgjwWXUUKo
rRq6gKhwV3XYS+XxdnrYFbGyidak2gbim03ZNHeQ6c/J2gbwOTULYybamZaQsh7I
Oi3PB6llvdFFl41EViA7LTU9Ver4og83Oz2WOeeQ+5g2wuPEpYSAULyxCb5/RurE
XKSvSpd30Ni5NQmnS0KvKg4NmIQ9fSRf9d1f0lhl19dGf7JAVYke58gYT17AfZPj
iB+5UBCSqll1MKWdm4bSLyruCWNVVL9wHAaKGplNnoGhjx56SPvr9Nx3M8rHkMZM
wRauWvAloY5OSC8XlT06xPvsFSjdGJSXaVo4M5hD+DarKPb+/6QRLDIoVsbzB1RH
nX0PjqkV6GdHAF1+K5PBOjx41CNsTpvTjm0I0mv6iHI1Jq1p7RGWPtQIP7Q61P3D
ySi/rt7wN48gtlIixVRoNtxT6+iAPKZ4elrTzJ/u9a/A27KQ0mdorc92wf9rpWaf
A53/PiUR8PNTBOMZCgC40d5F/77cOtmeOvvX546eYhExJa9MsD/Ii/3ajjA93lZX
Xpo5gtqP6MvhYeYPHh4eKG3U1rYz2In1yrp6Spq9hWZqhf/88LybSCexPmN0z5e6
XrsdQ4oS4/mDIlYOYi7WHKzYIHZ59HMqUroI61UGaYKFgf6K+mCo2qC1JIr4UBlV
LgjI5ICxmZ7eTTUFMLGfC5EYy17Y3YAZ6qCAyr72A67bzF54TQ1lwaZtV52Zdu+k
ln29Rk/dG+/7NhG1VFNIKUOheZdaKWIZDOHo+8pnqnKFjFG1om3xw+HSUIGG72Mb
SpntMwF+NSxfiX8kVbkXKgnbqnq0Dmp/QVSdMl0d0VYTMpA2qUOXIwvQsc9sqFA2
N0h47PicH/99PSqxaoXpAubEv5SXt6LRaZ8r+i+lF+Pm0BiJoLc5Y+Jkc8DrTD1a
oKG1y+g1r4NjTruWYclwBE6y4varx2jHDZogFpmhlNg=
`protect END_PROTECTED
