`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mUjgGcpoVByOibPHWGGzzu0lED7MaEYbrnrzkpiWCvfYQEYfoh6ikm7ZaoiucxOI
2YyI2P0E2+6r5Ef1RT0YdGv6893RgXo5bZSTx6iyxlGKtUh2ZaTjY85cF36oC8C1
jxmqsZ9SUsTApbmHnaV9kDlovB+vBrWgIot+sWnjmcVcFsrxwxvj7XKa80rkf+wk
54kTguFHeTW/C08sRTqcQg15xpf4Jvfi+siPTM21Fwx25h5M5O0KNvO2SOTFrzyj
ucioFT8aGmsCHlexTHQak3ZocrH7z02BY9WhOad/Ijj2PVc8Hcsb0VCnV91TJbG4
37BmyKuDP1XdjSYYk0S6M0SCQCxMFhkxKrNhzZyWfrMP9C8CYYoNXO6qrZHOHJJm
q7Q11TmRT9zumH/zyMXykx0swPD5QQyWIRxWmRt2SnAEwqo6+FqOiuN5Pe8r+iRa
pW1sjUqIxKUdFgFS9jp5k3TUsVLeytR/3RAb7xQe40TI/1j1YajzBEkOdrGdDrcy
aK7STgS2505GcrxMRd3PSsftQwKLT45OsQRSepBjxVCEwMiI+NUaOH1CiZevV4JD
FidgSb6HYQ4jJYMbCaM6dbYW+Z2xrLflKMl9jsFWWPxDirTLG0CrIVxHbTpAwR8+
+cnKlAaQywzhL7Jy6JUUT6OwBSQSKrbW8eBipxa5+oJk/gu0XYzDebPBgITTuWRx
6sA+nDjohZC2q2UrSKcEIE84pU0kTKqHwbWG06TKYQ+LA0jLUxHbQ0LvZKMGqrTd
AUfi9A98oc0zJX/Zzti8qFRb59LCEy4gybgOCUmcrO5RALcLtZZS6tamyPn7FnG/
rslF9yCpuM6uOgdaiW17qaTNd0CIe84RBJmy9vevozfO+5qXkcxDi2qfqsgWI+Nl
t0vlVg4CqYDE7NIO3h5Ip4RMJaoOwGOVPkcwmDqNE43kU6ys7wq5BXIbeky3uqwH
SwtLirW/Or6G6Yqon56OITgT/8a0G5EvF6ny/voaT7RQqi3HHOcTp/HtLk3tXdhV
D/ihGzs/bkXwMTcqjtCNgc3GLn34L0jw4o537aKqtdxETE47dvu79o9SU/Xc54tC
Drfci4t9R5KqNMFVuchvps6Bu5K64ocpGwCOZUZPbsWRiy2NXZ6McrjeTrG1my91
Gcz15AXEK3+kc/K8Nr+9s6lQBVn02SlyrA272HR4eHsshgnGgIdEOOjnpommXfEU
nj1ScUKnjLy6UWwnMn+qi9Ixi3oyni4hTUUJrUF5XpPtwUen8lLTN8Ax9nIo3WJ+
iRPQpRbAylkdXMtGeRD2/8nUSL5hD1mnmxzravQnSuacibg/0s+X3OMn0LYZMqhS
J3HmyRv41AMsXKxdqqo9QRs9SRDoFlbo4ri6ed4SK3yuiUFuxo1vzT4m8dSK2tas
6OfidBLeKqgltrC5G6askb7u1FsaEP8wmjeniPuFKpfZUUIGR3O9Egz6Vmk50c/w
h+ZTJmLUp/SAC9EHLGlg09mXpvd93bdqsB1A2IdA1kKKLDba8ZMfoNfFGjghGjLv
7ARafHXTvmlBIdrkWOwJU/y2dWeZ5H79UlwgtYKqryya1U1kV611BMDwhJk/bk2U
xsVeoItJ4p8YLpSDLJL+ilYcszv4OY7CRuGgpF5+E609kRtPKurYY6TlGkvKQhbe
wDrbFxps9XBDKGl84bbKFAw0x4nt5fjpbhJDIA1orpdoEVqx/owqUyCoKrpJukVz
uvAiNh5ozzu3KT/wKKNWKdpnJ1xf/zddMPSjtGOLXAGJ01wnDoRQh3Xr/PQTmYYd
3oZDsqkjRuvBmEo9ZDi3RT3oFQgrjQCKSRakbbpg5+OvnfjiuOyBe+Id9fjz2ycW
cx+Hr63njAnfyYymvq3VLtLSOBSONSpMPeWwhFuNjE+dlpzoVAYMM21+M/fGURY2
PSvLa7aLhn63oXCie/5ybvJfCxC/osbtUi/Rajtt5a26cE0Kc4lMJ3OO0TgppAOM
aotIG1QLA8aHx54KLWuAa4UpFd63D55F4XXagnCw6Nvvc/dnNV+g+XpuhrTl0rRK
X/29XN1wErXZzzo7GI6F4aed3I1kTP21WodeW0pcRaxLdeTOHFg+xFXugoRVHX5e
DTv8oypHAmEGNJaMT31vQw==
`protect END_PROTECTED
