`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OethkXdxrwW5P4eyg33upk5CbXzVyO4CO4sULx/Ec8ANRGpPg8PO1XcLEaDxUUBZ
7Fe7HfhuqrSNGlH9kbGGQwoow2OY0WxNc+VBaScKhxAVbOEtamnz+4c9C31jIT/y
TEfBcZICG0l5+QIjbxKgRg1a9y7JXc8S+7gJON+pBiWGcunClY/O8tMCjzpGoOmP
5BclsgjdaPV/dnAiGnoV19wyPTdVAh6LCWDzUqAmgZeMZ5t/BQL4H0K/YOjfA+Wk
LAcyrzMVTeIZ4yDUZtgtRI4pxaXi7qw/RvfRWGaCkijJc7s+7qshsD3496N1Nmhc
G6imx1nBh6p9U8rwFKL8uxLIvxbr3p/o0FDN8g+Dsb8GeQjVOW/LFDSY8p1dNPgp
nqe9iKex/De/rnd2SfD2uaxSFfbMg/pkcH7Ke2y9FkupJvTZ4RUrFG8IlRlURYp9
tXj1mffNkaykwdWvMEEtQGd6gX+5h46ByR5jZHQpWw+2Qog3s1Vg3NUOlpdCTHV8
`protect END_PROTECTED
