`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nACfCr7QdmrJh/3s/VCw4WQ2xHLDjzqITIXEv3YEpvQl9eV/r+FvCEjyqB6TSyuO
oRttvvtR1TAoqE/u/eXu2cAQjtcNlwASO1sDBjZR39A/HvR6q1pW/Nc2/1ymBAQb
EJkDPYd74JrFi77yFySsbwMWbT8oP4d86KbytaxRqjXsEbdIxLzsv0fcDSF4oIdQ
3xR2IgC98JNBvNdzELK+2ViLvObhbn0Mh4cdecdGy5tMgonoin019Fs/UODn7VpS
Q5CX8fV6i05t0kSp/4NSz2zbN2doxu6hV7Rq9XeIdZA=
`protect END_PROTECTED
