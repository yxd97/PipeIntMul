`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aTJCRw9OIg39lHFWfuUwqRCe7hldjomL5u4F75V9O+sU55qHPN44VCN9FlFhSeLj
hNFIM9NwVW+rlzO8eOW/N1Go4v52z1kdkDQeGmuVGtCVhM7tAqFq9oXFu2Is+bc6
CGPQJeMxpROpAdEicZWD798/5Y49eOCPX+Mkoom0lPJoGEMC83t0o96tNZ5zckr6
G/GEIxdFd9FEwc4B2oudRRaoSh1HkLiu0s3euKfcsCCAGA0E+5StZF5ay+o8q25X
nbvAJxE21bloKO7J1SsMWwR3d16pqiJxX1D9/rQj+gquv0kPzconn/QXsfVLNx1i
LQr6CkqRQfxrtEfUBxrXNZCSGLDMpBN3mKSKRqnX7dW4kzjwR763ZRzKtICL9vJQ
OL3mX9RWpS6PgjSQ/x+G9WqvFSBSZSNOXPswdasv04UrXz8+ecvBQfZX3dst6/mI
KbHhzpUSH+6rb4J05C9WtPwEUgrHjSIBGSB6Se3vbSHHHvlEHM0b5UwL5Tw2If+A
r/+vc7+vg3VS1w7pccwxcezJKvO8XugfBH4vxcpcMd46CxAjLRl13Vt4doIozaKL
oT5C6GU4dZ2a5weepSLYwfZDVY4cWZvqeazvl2GuK04jmYdlocJ8k5z5kjG+i/wJ
jrItmQ6q7B0Yx6KNMZDDx03b2qRnWkzWUbD7YFeDNfin026nfJPwNq883d/w5Z6y
aW6/K+S/WYH/V9BHuv2uMwQiZiq2x9BAjnDTW6+u42BHbbk2jzmgENzYIdl+YWUr
3WHvuB3GYCAJJhd5TQBitimly3o3h3CI6agy4xUt8NdGxbSzMQkMDAc3af5+WRCT
LxEH5MYLuiPhC/GWxemXs9NKJRX2PkDv9SOPP49nzect4wK2F48BWGP/AQXJ8dRn
QC7O5kQiOOWauWl06lkBVQwIhA4ZmrWcHa2xBPZuJ9FJmFXL3wHvRV37MGItmfDV
zpF8/7CWd2edD4s596vOSEL1gi9j66QO9xkhhux3a7+J5fgcbTBIzIjyY+NyrLuB
oGHLCJAnzZG9mCN7LCBugx6B3Ohcah373O6lmuj+jtgkxZ9GGfrylDJzAY5xp2QL
KqN3iLg2INY25XhMx93lLOfNETrGIsxdwmZjLJ2tb3u2AEd4lez1UKuRK0nEgR8C
q6qtrqWfvO/9asm4zI+ySZVsUUYte1y8MfDIMGdOrj4ceBgIGM8pAkToiJteMsgI
rg7TJhezpBW8YuUmIWNZ8GQxzVjD3KGQwBC2fTUUBuNEYDT/wfWYjfzIRW9nE1WU
78AbORWto/Tk5cioQ3Xsp/Y3mAQasL8NjEFGYlEcgL0k5Ax3c/ShLvD1/07vpyup
HD4hJDx/L1mSZHBWN5mpgdfvXUStnrzJA2A17rlGpH7PoNNOGDkWmiXhG4rh8wvL
LctHW15nFbCmq61C9fMOl9I97V7Rs7skUFCq9mFU7UO7IupkG6gAhRceB+BSCag1
Sl5PbY4GvjmyZVveqRnvFEAsvwVk0P/4XMWcDHyeYu9q+fjxcZ6gtne+TShgoOcL
3AH1BuLPDcU4LubmMXJy05cHHoGTY9X8CAg6IhvN9k9GkEX6RZ/1tL1Ixe/bpKP8
gGT/VrcaS86TD3ZjCVukcjY2hRJOo9YeR38rS14EPBfOtm4TfLcJILGdm/kV0Iq1
USPWyVSnQ3Av31U2DMHO1lku7/H+2l6Bd2eDMdqZBo1WeMvmFlex14RBAxyO/X7P
aq+B4qusk9p8gctbIKqSIuqKKB0rrVfEnvEFAKMgEWPtKaEyu8VC1n2FxOuNFogN
trA6W0UKQ2oFsdRtGKxS/Q==
`protect END_PROTECTED
