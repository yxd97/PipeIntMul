`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wZHh8Rod0IZTlgJ3wZQNWPkW4xN1RMlVGSegG7qDWW66dJMh6rdgTq1d67wcL6Nd
XyzAiz1kFiDxtBz3bK42n4fC6YNICeodBxmHJC/kmHsAsEWEw55R6csaQt5uhzE9
TCTFiDm9cv9OAUwyHog9ja6aDQsN28LJN4ufvhnuilvf3rHuQnioMY0KicpH66IK
Q2Nw9XpkmK9AL23/lvBxXOrnW/NQKnY4Wid3BojoJot+0ZmUP0DCozxjY427h8p1
CiPJaDTVNRzLWcx3+/FP0P/cTWLDZNKh9SQsxhYNXwg=
`protect END_PROTECTED
