`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aExTQ0oucbmGw6NtvAD3zm+uxMQ/ONniZKg+hOTc2tkYazvYUMRtPEezmclU3V/i
/z9SFc6hrT2+0KOPcaZq1/9zg5CfXiN9jAUsj00EiTHaT3HOEFSyWI+6WOf/O62g
zWOohimqgva18l8wPyvGtTUvZqm4Ni6a57vYewFr9BxfX7pDOMEiQG/5cHg+jpVP
rNVwHfd8k3YViXYpwWA+7NRX6l5YEoBMD92co9s3u1GdRSIqWMDzoEDTLdYe/4uq
cDkE1lLdg6r1+8R/aR1lI9U6N1LRKPqVW55frStExVz9IEk5w1csqEasYv3pwJLt
WIU67gZuluPfDHJJVVS4/qMJ0jAL1CCW23q+JLKIdbZRQ1PsU1XyZa7sBUchRw12
2GyCzt/ikTjYTbkzA8QpkWQsnH/fmDG+J0OyLd8CaupyjbHYSjoX1Z5m6z1nrkyR
ss2IvQ0BiMqrr3RQyIlow5Z6fPlfffzA2UlkFAaoymy+HFLBkXGHIDjda4isuMvw
d59R89LHaCdiISH1M3/bXGOIh2veK5hBZHJYHQCBA0WQI8uhoWnUzpU0lMCONMGA
HG2v/gypMubwWdcH/7CbNxPLLk5rpRXTobfumHyV4nDGlwJQLSTHkMn3Oe/XvnZe
vKDZ6NdcAws91T4VKRL0Bnk5HZwUSahJksYzJzYEYGOTGzVpPhn+AfvPAMHcCnTU
F0p77iYXBJOcvIptfHOAV9cu5YKGgRTmiYagolkLb6aQzlOLl210GZHWJmKZqAVm
QnjLp8M5ZsuBYMS5I3cA/MCUw2pKSY4crwBDmIjxNMviM1peMm/VOzYtump7Ze3g
SCOSySY8T9RZaZ61gPIhZ/v3wTLaBH08htog8uQ6MQql2N2fN2AWHuyJOSIpkvJV
bvqxkq4NURwUHiBiZoMq8R/z4bIeh3jmkgOGpTq/vCHl+MSAw/Fykv+iOctFAUnt
YuF/tScBBSCX5dZIf3GGAW7BB0xQY3UwWztjWD8azONS4xDvhj2e3LV1hp/WczEp
D/kGZnwWtr+21VoxDGlV53MsbOfdjk7KDjsEe8PEgagawB+STHyaPeQ3NBPukR7g
y/89mmxsGwdSANsBsNz+wdPAVRKlB1BP8OMR3skALM9cyG5J2EGGJZDPtFitLElm
khbugqji9/5qDujH8A1DUQ8xEs/JFc18ndcshFzAMa+UeY1Gj8LJ7Q0ecR6+XHz2
VZJNRsmrjAVGlC78yAIH4nsaVj1VyXnANMKMgkGL9dCzARqwv3Bxbn4L/RfmMbxO
rUXfj+pg2W2y9t+DNwA71BjVAhw55w6WzbyvtN4zDeWEtXrGeff8z2PV2FKYrFZz
YQ40oznicKssFiqTUxwKD2SuQIsbrztFUUjKXD5QOEBDdKyW7rkYENYNxlaYcjQ9
58L3auzDeQB0WQV6Y1RuFr707QeobKJkEoPpx9jLbnUTdZrq2f7nX+dZbcnq+j9a
5JdyE/5LlUcHiiXRUJRmTicTgGMzq36ifLY1LJ4eYigC07FrLfHhGaobwi7YEevz
jVFAPD0TSQ+frMaNXK3aICvym/EYKBDLjzGX2I2vOYZGi/OzKw7CxUBhleLyEyBn
Zq1Fg8drGX77PgUU1dMlegVBiXDJJPaJEqXwSomdzDKv894RpoVMpyGHJ682Ypl2
BEkR0ay0T2BcXLg95Wz5iTWEnv3H+347QREopi7gf9R7YbddQDdBJmUFrTCSV7Cu
qUBr8SOp4p93Ze3fPQLnGFrW0VrCJ1jYU2b3nqtr+1UaKdxrL8PXySuUhu77UBXW
wd8vrk0o+Ld+HfrvP6yiUtQcueZ4ib2jFoTwH5t5wsEctvifQwa4DSV5Dqe26WJM
cdY5WJgqvzeGzZx/FTCAzPj9T5qTDJC2Qu/KMyicjNzF2DpJF955tEk5NceBQ09H
BWA2IehH5LgPbK0yGiCkpF82qzbtr1rq0GnXd2ond5D1eTJOIJyNofLpYKIPqrfL
BQc7Y3j8s+STft8v0j0mULmoSImQCwoWvup2DTL1HryqQaeay9ChVAQLvwzOwyHx
E8VvAOKgOVsr+mxTjekHROCa03wf8IOao0thjWDLKyIOqvlahojtpESno06Gf665
2JK7pdBGOO+QZWVJibWuplo4gyKnehB14BZAAI804EA+8KGtkp+WMKINro8LG2zN
A3J/CBUrgZ+5I+4LVF33WPinM1YoiHzFSxYxo04bp5eK6j8U29NxxbJPTMzPfBWY
PRTfwpLyUJ9q3gAVtAjwW8PFukp4O1+EapN9aiGS+tsbIpZIgj7UGy15R/cVv8E2
62gDeQEzRqZ3vzf+P8CvKw==
`protect END_PROTECTED
