`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsgsdFIu9R4XdpDjTi8F0lknZHT0dBL/DyS9FbT7idl9Wi/8xQGkYk4k5EcKxoW2
apKab0jekCvr59Eet1wbUT3YGhErh+dcUhtqh5Lz8+kB8EJboNLW0zMU+0E1ZsWm
2OVOjrJMvo4O7F5k0LHB8XaixtCiUmWbwdq06YuVsY2LnmsdtwDUqozHucgxa4vO
dUh6BWx+iSGxkx3hsApCpY96TVuRMfmiQ1yDRqusKw4PpwR3+Yhpbe24EtTUDq+7
5eNK3WaoP5am9l/JY84+bVndxuvZoJkeD9K2iaYhLItNlMKKc6cgNfNY0EAu6E9q
t44TPStwYpRW/nDrI2srMgxnkBS4VXJKVPAWOLkbHtnUjp60Rlovu2cbBglxjEF5
Vr4UymgHrUyH/Vh4nnbJsnEdRkKUBcJ31LMNA0j2IdqOsTC3y52Gaij3J8QXJDe6
32BVrDZWFFH1EBgdRBdJxzyPyH6PnB+BuKRQqVfh9zA=
`protect END_PROTECTED
