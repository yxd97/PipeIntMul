`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mo+PXD/qQ3bf17PT1DvGVW8ZTDPGdCHCjKHWY3rrAcZv5FHAMT8d57lglvHt20AY
jtrxy+5FAQq1I9dJKFg7SOk6Uj6L/AUFQRnbGJMORq+w9sOOIn+aSUQCR5CVEPQK
P4rUEUI1iQOeOlomLHJ64mJ5dERqObeXAC+I3QficGfVbUvsjbjWDD7BnlE2CMOj
IQG8NWyupGMnsqnYrg9cADHHXqoi6rPmgU/uksRokKxo8XT2WNEOSJlZg1nFO/9T
`protect END_PROTECTED
