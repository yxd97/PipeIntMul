`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C53tcftXA3+IjHpbrYdCxZTigfgKlS2m9XETLNWLTirZ/It8yNAvw1OlK19ZjXhX
LzA7l2P9GPifK9E1+kSSoIo6419FPIlK/amxu5arpUrY5CBbamAyLKmh5b5QY1ez
5UNpvZFQG8cvALlL/g8T7oqxLgtWC5zVWtBfBvH2a9RFRaK2srEG0U56yTKl4pB2
O/R9RbxvCHTgiR6x/JYv2PIC5WtoB1/P/v7WslgmoXDOksE0DHmuEENV/nD/+1XA
QpIYQF808QYF+VMmgYeZ7epifBQCnGWt20px9CZdcDGn6a5VAWhLmzT81uyIlnkK
vqZyh4eimjQe2UmtgZVP+rBw9pAYzPWOzQJVvAua0dPXgiBcs5uxTSZMBVLE8XHy
nZHG8HJ08PdE+b/7wEFdaUAUS752W4+rGbfBan0BvCCFrmcpxcVRD5nR0L0jddvB
n2nk1F0OuSJ/VqeULgx8g+EuS4gf1cxhZ6t1Yi93/5aUA1fDPEEoPZBZQqOUwSIS
2kqZrC7aI8YRrdAI3hp9uc8hkgk8nxJWxskFv69Kd7waXuTYrSJnCgT7gayoczsG
4KGWCTETR09GfprrJoq1HQckjW2oKJMYvySpJykhRVHh63tQZnXOiuIaXAl8uGZb
gm8Cbf8iuDAqSgC2oWnnM0DGduDX40evBVyUZPNLNBuH9vYL4vonYMWpe4cugbr7
Vy5HPmiu3mlvIXk5gri2/iYFxk2AXRCkucKv9LuAmm8XP+kwIZj/3sBDcvZlLKMl
q3WuhPKsVvXcotDwftWm/hMvzxCfdkecS0lkRhwTfA2tyQXeKLheFxe6fNxTWZ8l
AsLjQVD/RKIUxwN/usIKQYduO5sP1f3rK4bh8Xyhi5xxixsden9YcGtbA5Pwcvl+
fH57A/O4X1qI84gskhtNYPyF14+ReWUNItkoNfCpLNOqMCrbGhSdOtKOFQOm8Msv
lSA8HcTKg1hp3MiBH1+TbCNMBSa/uL+FIJxFOUrIWBbx27gW1/V/uQ6QydUpIyu3
4Nf5Dx7D/J7lFqf8GCANCaNjl23ywi+NsImsvk6jD+u9NKkrFtYAmbW8UrzP2UwL
2yRgxV07dTlqO+6JOmxAtpJHBIKKpI7YgjK042ovpcX0Tpb+bap6ytYi0N1KhetJ
cUwUoAgeEAx3m4S7SI3W4/Hv+YTQ61Sos1/66FfR9cqIvYxI4sAIh1AN9fy7tSgl
Zi6jF/mHmLS0JMNQPRTgOibE8d3eayc/SazP8zQ/V+wWQE5aZj9ecz+aCsHd4y3c
MKkqk976mF3yWkjQlR3tIo97GsSNR85MwgdGLjVJINkRtc/wb90fm0NcIZpXPX5I
L09tN8sZ/g32hXrisgKk41aS7esvqBzHKtBceNjUA3PNWEWisH0o7mokacGYMFex
2TFUXNBWefPNMgIyfTfMUICJcGrhjzqbp7Q353zAgoRxQ+ikuzaYtcKgEhi1xBvR
5REFBOYBsuSNwfOMvWY8ANKX6AfwWF0WSG4IA8ycAcwMWvosV26HQnPydCqV/Mh9
dxIxeYY6H1Zrwme5hsYywWDRpvuv6JNpSq4V3krzD+JkSh/bRjtWLOJyMs1FOy1u
ZrLYqVZXTz4HmOr66OCu7vMBNaMyOt+kGDpv1mMqwUGIVgA8Jzoi43xQAicmoiLK
3mvYEX8rhuPnxVzfM/llfFzGy9v7ETFvvoGqHXFjwfNKR9cuEguIGUn4d7lfzAdd
jlPqPFhlJvU6GPw28T9vfLb+KD032oqKKyPJUEE33JeeToTY9vOHvbFnvybl42Cy
HSbniQZdSOH+nuRwho0vZcqlsTzN/1xRYWGGOKuoBMSeUO8jN/gHMtAqmtqa/kdG
dvi7BHr4yXfDtAgMS5l4n/2E7G5tFjKbdzlgi9GxxBY=
`protect END_PROTECTED
