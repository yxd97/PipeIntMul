`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wCtpaiC5IpzWZ0ctRRiTljRLKR4RnNjLfNiLu1jUErTkz6ehtmWSDgvT0wnCgl2J
1wtVCJ9N6HNTnNEqhUgkRGj54dE3gAaxNUErDRpBikjXtiA+Xb445gPrRsGaupd1
QwKLezbdl18qMF1mY26qYn4qC3zOauz5n05Hiv5dtK8LLjibnvqYtp7ftp9hMu+e
UhtKhxiQ9x/Uc2K093FAgnr3iupZ3mzDv2enUxIc9cdDeBgKtuOlFR2dYWQFmWFB
Tz1S7UM1sXrZnko96SXtPsYn5gVWnCVI3w2n158jzHITAvYW5KPevKcFSdFGBvll
XmJMExq5Xsmwejgqh3EM2ooI1+agKmCKUs5dtNTuqhtWwMPq9oOhlvq7DdDj/ga8
Fy/EQLYwDbai1yg2tH6pgNzSFAWtHmODTwyaZiFaTWWFqcJPPqNWWaSRQkI4Afb9
0wQyjIHoCqPGiDsgw0aO6ahO/0xfiOUJ0G2MI7WBnVPIA3h8o5sUKRB4BgdBhk/r
1fca+742o4P+1bBZYqHCFloSRFyXJbhI1ZqLNVpdVPi8h4Tvpo2OMUgE0/16PZTW
1Hub3/vTHVrAehuvhneS87oEiLCG9eXREHRVYVIZDHO+1wSaNZbrPNZV+Lui/YUb
5Md7fivQAIR8r1L75mYQZE1V6q2Iv3PCzTHQhg9h0YpZpQTKg2a0W6m0kNar1UQT
toBL/JUq/gJ68nkYf2DTG6TCnNDe1GrHIgnucKGYZAWdT2bMATTkdI81XdpkL6DS
zaFfwnA2CDbhCv+Tjcop7WSoDDdk9kzEIzzQcUAbTf+h0HBZdVTjjkDrdR4LY670
GBLXG6V9Y+alXtJOxJOat0zkYyl9H7gOLWNOk2eVvOIPYIIzQyemt/6GliVR9Pj6
XBRbi0AFvEvFlz27A0DhKzqjPZNLRgOLZx2n36FhXiZDsqtPCOZUy1V1WGNVS9tv
teMfTrvBlUm1+KAP9MT3Ht3PT293/OLTj6hx8/9mhmNXcaXCCMzluSm7uEhD/4NO
1R/sRUkgrpnNSg/qO9qYeKlZd2zJOe58yrK1gwWeNSVmwCTVKKEHmbl+x2yizuyx
xXUeoq6Qb56h8p34k5IldeTHx1vz3I93RzOAjK4xb9+Qc4fkz/JInjdArkmTir3q
ILG9VHUrEt6fq1E83W0fsR0FksGal/XzL4jUqtMMh8VUSnAIJ/jgC+35CmBw5vaH
pYcWTy+XQzeeRlgEiIN/dO1jZxZVpV97J31GLsThCFVVFfG+h64DD7ZS9IdiWXbw
dTvPMmMrNUm8BMy+99hdJRgOLjSh/ho/kkp4pjsZFAHwDJ2fC9MYd6YMFBBBQDco
KgE1NhgZsbA+6aGw8Qb3icECSNpKf0n8JdKeSejh/0z8IFW1xChFiRgxDbYUL6rl
FUc6/y4aJUaPiCdXoZz7XnXicLWV6CHQ8ZEdrKOB35lhjLhOu4bgtx0jdKTqTW/X
q3hxsiffx+HNoieBZyC79A0tDi/0AneiZbxeKYumXymcUOD7E6zIbaakPt/vkQCD
51QyUjPXIabZztHFzghXcoXT4L+66Q/5H6uis70b6jc=
`protect END_PROTECTED
