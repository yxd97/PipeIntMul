`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i0+GxsJWEjjLSfdKEepIdZrgN9iJXE7+7aztNeQvbSi9qzNz8ZlMvVE/tynect30
6/EooJNIxWY8EEfOojr8ghcCszQB9slCb/koFWfxoah4aehbfCqTzzVHYbphN0TO
OLj0/GW1CJWDb+Ti9m4hgwPS9zVmQ1xcwT6rZrOGD4Vv36wgJ5JDLGTixmhNmBwk
1UUkLL1dFOn6/g/WSyXdLM0kAmnmkFlL2Llml09dtfcXcFpOkw9OvuE2wReJhMlK
STfjmDd/kLJwdZ7arT622fGjQxVz7SbGByXYrpF8e4g/+g/8P8e3h34u4pl/9/Hg
2a9MFLa5aa62OsuT7XsT4JrVVU23VSH3uUGs8Nl/1lP2ltWvD9h+nV+bc9zlFojg
bcEGnXW95WZe0zo7C8wu1RxPe4ASgvGrKqkW+U6b8d3dusTWGl5STLh63VHZ9AZx
3P4pEY+Kynu2FQJXTWd/F6IvzVzjXiz3uuSxHchXqhB6rgmrKAgJ8sVEKFkwpBIc
2xshpa5rF7bv8kvF/zzurvrrzOcK/aJw91zBIhiE8cJdEJNKPin4SYOOaeRYD40S
rhMYUQ9/9cI3gPZITbX8I6A5eV1UNIhjMFJQCSQO8L/FNv+oDdtLBCdxLLaMNr/q
aCzMOTIo9uJjCLvzkEgCYrnL0IGYGuDkfaWadV6wlJwo89Bhiver588xBh33Hzq7
b037+fLrZB/IXr/g6Rz4yTmBY6nvKqH+uwq/UUlOT1y0ASZ8TeVyPUzD7Jyiaafy
Vn8ODpY3UxZkq+I2vH/TlzyWzLlbGU2mYUzH08DrHsthphqqwm3jRdriCs9pzAE8
HptlzHSqkfX7lnxdmq8YjQ==
`protect END_PROTECTED
