`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9mwM1kCb+0QVIky+URl8XQvw5hUkCM9kDA1tXU9Dsrap82DnLFG159ucIOHjC78q
02isEU+a/Ob+qAwBUX3asSIoKsnisrN+pCcI8lQwWdsB6tzctb2CGPMHx3XIP5pM
+xBYfkz7/cM5Y4fdBTV4RhXj+bgQegRy9JgsJcLc7/0Vt2Nv8FSujK/40K5NiL2m
c6vDW7LI1iFUxqkmWvq8eWk5W0mh0fGUKQn1hyPkjZVRW6is22mWeNW4QzIQtpoI
leg2rlXRLLvv6nXDS+I8TaOW5h6YVEcERu0DbDc8KvTWem3unMSNbgPidEdWMog/
DHkunGxtMmrSUaRQ+phSdEo03EQPsHkaQuJANV8GkwZlC20acfq7b2wql52iqQD3
cyb+iYXhIN3sCHJaAfaRZ6J+And0sGD21QtXEMS2Uh+hjfsCuvmHiyP1Og5RfLeC
l+62eEcsYNZ6qxEmPRIXtBVvGwyAQ62knZnnoq2UdZgeN7bPrAa8wvu7hzYjDOcW
jYBBA1mTgpNnDUxLm3q3Ns9c0IrSSnM6C+xmQmj2ZVsyxX/Dn7RKLFPu3suYuU7n
ny1an2BIYwwKjuUHGxM+RkXlB+650tl9H8fZZuSYLWUCPH90im3uociFcGKZXuqD
0I4IIIuxHCOAywHwjjOEQ8CoAYaoRIJ4Gl6gilBwpPqY1jABs3Tmom/r5xDdpVvo
mwIlgsqfQuR/7HUnyII6Q7+XhCK4VrboMhUq+qdIU5KMlPdbX8x/EKmMja7gNOzo
2HQnoV9fkg229LmQxbPcnAS1WhOG75IUuqbS9qh2Ql6NMCq5DgX2NsVAYOgnjT97
Kk5vh5Rz/zD5yI3HQzF0NKT/Z2x7PUm95Z5IWr7eYxxzZQ07IbT3Et6ytjNOYvX3
FCwct4n6MoJNgFRlq67J+oK2DN9aQtmKY2ps2WnYm/7UD6XYU4d/UnootjhYdQ0N
IEPZK6ZVSzhpd+cDMZ9JVBlFoAXUPufDJcRFHpgYH8HQamvHNzh+289AZJuOmjPb
oyLMPdWEcV/NDTgoLWyYIib5Fxd3Ygg4j66VARGEfI6480xf6bV2BN1/mWQxRQ43
33yTwDfB5yZnxwR2PlHDFiNcATwpdX90tuhocGD7K1Q=
`protect END_PROTECTED
