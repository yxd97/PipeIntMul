`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WXLCMoEwtvnkLu+C7Fi+eq/iByQN8laifEBuuHawJDiytZF32NM4QOpnw2ZTCuBb
Cn5SWRSVTsQiPeQmq2rgOB331ZzGkR6hr7s6Eao2WhRYAUc4jL7OuW8IfRInAbqa
Y1Wjs0yjyS9nZNB2mdl0H+3Zj3oAHPsNx/moQkRC1Cz2pDjZstqe5/6ayDX1fEOh
Ruv4FFfA3rp9WMk1KRBKx7xY8BanGaXNLM86a1eApryd/HvaNnIyNoq1m217ri80
ABwmQgBjyJbxzfdOL1Nr+hcmsaRKks8SBTmtVO0jppyWHNfewKpt3ibNh6j2AY9A
tA9icDN4o6qEtJOd0SL+k9u2B+HY/MBH6pmpr1VHnw3yQPLrXBvz39yZ9JuzbwvS
X6GFTVbwAEg/pYK3Ac4Kci3bGdJdQ2FB4YyF3b/FQJy4fGDBdElUK047f8JIp4QI
TEVvSzVHptqNpImJtHMKedNvqHDTkBwFBx4wGCHyfojHgAuWFFV10km1hqplie84
oHI2hgiYcOjEPWGL+jfF5pf5NFUQe5iZ30Oqo/PaBS41sqq4UazwiLoCZCLM0yot
qUo0LBAI2cgD6pdB3ZOYarT8YT7FZLy1c8X8+cFqzRv6pfaB42602a8OAaBIyi7l
FjecXPy2TlydWtVfw0qQMicPxux7WJLgbr9+fiElZINEKYXuGPpScEgyX1bwH6RJ
rstYb5/Gt5mQeBRoX/0oxkdY+OJ5atYSDv+juHAkIVMxYGh4NwiDdV+ngEiznakJ
hpUEkyjMwn76UVYBegSD5aAzB7lVfW/fMeop89VXRx1Wib/4Rp4zH7raYq8DGCNG
AGKRwnyNJ/n3Rt262xq37Y+dd0jVE7NyMG1giinAVjXC69Z1JFbmjkGUwA6iAXI/
hgia+NDsc15vre0B1TeBRRFLOV9jrAmuFIDYuD3b+nzh/U7bTE5FVT1GVsG/TECS
t/d2YR+65fq/pjbGjuh05NcwA+N0wUtmMWS8k0KrlzcmJOx7nzTgje4JSqBRev9k
ZLasI4XSJgYyLOZfbJZPo3Sdep/HlOpsy4XEWddSg2LyyLBUKKUttmhH+atphsit
Vqk1iKS7HHhGf62u6K2hR/2hGIZX+hOYQ1Nko61CJixz4LPXdKS6qpisMzMvgY9E
wBtm9abIDFb3fBjZJwad6ZDDlWPEsBBdLFzZDwjYOLa2mcCsMkwBKR8dtQajpfOr
seS7iDiyNSu3wQsrRAPK4W5qwE0NHuDk24f78oPuuwIKATDDyavKce0pkJ3tCkNp
XSHOI/0UmVzdvscU3cal9+Y0Rab5ZSRcWErOXYyiGle2ZNXhNJSmkBYf8ke/BhfZ
0DVKQiU1NduSojSIa1ZfDQ==
`protect END_PROTECTED
