`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YqzXyqefLsvtkt5SF7TqB4YMurj0VMBQomH0nqZq9d97t4V5ytoDSHlNBBPYHdHZ
JJpsttPCbAeVrdaQb1dA8S53SOrkfQUkxi8Ssa2u3MiDDpS1bvh4tiqwzoHABsA3
N2lY5FdUsr4wBFd+dqDonzzayO0KpmqUHg6D2qXrJcgKcfLak+iRMIvpBRR4dauR
punZctAvG5AR3k/PqWFc6hDe3uuyjqKDKWgH49SoR33KayRlFR6x06q9vWFwPW3S
57EZrBWAyG4idPQ9CTPc81kCi88p94TkoL4uJGbRxqM6SncdgMsqhLSHZKefsM4x
pnyMuMX5dPLMOm7m/59nUJvDsD+w04VhZw7clggwyzYjQRY2UKAKaRd4WS9Z1APu
1X152cIhuHlvBKWUSCZTmrNo/icoQ7r/AsMNEyMtjwKxegov9YPmPx7Z5A1irKVi
zTASZjZrwJEKf7tTF+ZWG037i4KPmYbLg9yzH980itLxjvmliHxhGkg7+jnmCZXs
7wmZVRlVANgG2JkpvlJolkfQkzNP6d47JOCn8M/tvUxX/9awWIQ86Dj4k1O95jN7
6L4pPaSOIy+bdZlplL+jTKLhf8tV4GpNqexF2uLy0e2cu+1CwjIXlogILesG96tk
QUC+2waZG/IGYik4JvH6Kq/U7q9mD7/q+egaHrFbV8c=
`protect END_PROTECTED
