`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
poacIkdvjx8QNz/mdWfIJ7Dvlv63jiQOBO59F0QdT+p1qoZu5nSCt1vEMk+7KO5U
PcYhZdiwqO9J+xfts+PYwh2bk5Uc2xr467aNMn7rttFpMYpo9wIBG6ECaCpckSvx
MxUCd/lpHyKcw+UTFKtMQjGyHT/RMre/9U069ErPQkkxEAXcBXUGmgUDBm8SyasG
2y4kgTm+SNPZqXdrH0fEpWNp9SXnVl+7E8K5PYHFLr3nLkAjfxApugmu1H4Yt9G7
ILApAWldNdZcyd4DtaNxj0kyADFGICLDXJoXY0aw8n0Z1FJ/mWz7jjt7vrkAc6tw
vRZKmlpz7avuOebQ9G4HH7d85ZWStw5/Z8rj/0MsMLBCRtKey5uaeSGUjySwPIg+
eb3KQzuM1eU3kLY5q5Nm2vy3JCWo3efjLZAScPTePgekDka7ouHllIUZDdeyQ9He
Ef/FcY2EterpX37mzTnTLvdxY0It8O+/kRmxcdKJGBP9hnkBhVZeqkzeGz0VoZlo
OWOf8Solv3NzMCbrB944hY+pRzYN8ssidx+zjEdGhefe0c3Uo/97stFkXNS5huaG
OBCGdvxZ/i5Ay4qR5pj33rq8+jdlFGCL2ZNq7XOZdfJ/LDzmcu6DZi96XwZMIRcj
3LFZayPyD+B6MmnxEjnXpifn4NZsc/bXeYGiv9yzwl3++d6PTqHOwU0qCeA+nsWp
05sPaUtnqpyQVTnoIV6QR0+8IcknHGFX4tAUzrD3SRV0EbNDdfOBhZREMDAS2jKh
MQ2/v0/5+P9WhmCdtqAUbRhNav8+UvjsUo/jr+GU/aZU0uhTWXMDxOjNQJX9nARS
aqbAB9i6J6M6dTd7vQ5S4Yz7Ii0NXgAeAgdMufT3D/rjL9ZGbVWHlyI2A8k48cEQ
qZbfjqegRbcvsj4LygxctBgH6DMl5pH21jnpJnJteA3TI5GeHcrBsCxhyPBXeySQ
CtRNJUBQlJh3wTD/q5Y00rD/Vqwilbl5o3uVtQmUrkIqB+4saFZhmfCMMP+bPV7e
q3pTYUjgsNPFQ/G3dPWuPwEmOOmtGbSip+fy1KDeEBK9JP8oRBOXTMFO5asHiNs2
lxMFb0g6g6SS74kW1dF0gRhWXg9oBJjhOMwSusYrVV81EM878BnnXdJ/+okXXAHo
7Cv31U60LgAtLVGVCMv5hq4nii7o9SenSQ58n3oOVYAWSazzg2UouRr1UKu0gY5r
3z+i08J38SKA9qcWQVfNKPrQlDD36rdQQCz1a1f4J9euIcLRkpkdh+LrSYfHQy8h
/3vXorkm6GDbnAyNEDJeIr8QLgCSLVrM+PpEOa6IQ+WFNai+W60D3cvcOpnQt70+
rTLfoLtfpSqhG8klr/PaB9rJNUzsdiDd24sGMGouwbsL5oLSRj4eCtUzRJZKOZSX
iUsHY6bqyZM73V6JCyD+0pEe1ezhjwxSArdz6oJbYVo0HRhBWN1XE63f4CKyMsQm
uorxh8xAWro/CZoB/wrU/b76yKUb+AIsUYmFJF8YWDvUIz7KjGxKC0ial2dxhg4e
zjL98asIdln6Vxf1coJJH9oUO74NrXjieEENrulZQQBaRSCeKsd+Wvi/q/4H45RC
S1VMkmWvYW2Ld6Dp2xLj+su3YhcwvHvbH3TP0ks0z2mN/sj0eVehIKojzsRvqLI3
Q6ACVWh6b1Pqv4GJQerogP0PKASIurwPtncrzs4OWfEfEhNec9f6zvUN/FSV+pJP
6yHvX72Z85YJ+3kATDFtLyO3EKzIihEjPqDSz1BRCfopG+NzM0Cii7wK/DUiOUZ2
7uIjWNCn6k2DuFFNwld1ataIelYPWLRTK8LpVnkTXHSeyZqDPaHaj1PK/LOoloqU
2TgvSDYcP46BUgVauKhPK4p9vgtf6FGyqaF8GzqUdlXsIVAFskkPTnCCn5DhV6VA
+Gg7RDrIbcgMqOm3VBjzSPYuNwOWM3qEc6YD46GXDl26bqz9ar6gJPd3/YuTo8Z8
CVrT9XqA/5DgebMZJS0snanefloxItS5+NGwCcO0ydalkK4nFYqbfNPdwQpsoZ1l
9Dih9mNAWuksrhsPoDiNhbJxOlDoy1lVSzEKfo10BL3Uht/urknCMqo4Pw9UlN9C
3U0bw+ODlV2jeJ09Gsva3VFb12OLa8GI39vb2rB7NKXfobhHcm4VUPndCdW3Fkox
e7rdVoMMNio4giumU11AEK72eePgF/m5JpIsP7pzSD+aGZ0qsxGrLnbRGZYpFZWq
d0I9FLKqjATBIapGdw+s6k5gtSEJjU4Cj1HfdNyi6oN51KAj+LmmY9PNmGnGkL1l
pLH4zURbSQ5UtOTExzGDOIosG75g1ibT6Z9kcceLwiXBmptNgXlWD+138QyxwciC
`protect END_PROTECTED
