`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MudMoKJ0aLY7QYpD91Y++ssbGFqVHdiuk0HG9MhxqUitASVDI0F+VZ2sh2/M0YTN
oTOPK+R1SPN67LvV7X70744BnDj5mgakqvrMICoyzadbgEiXixr2CjDPWZYjEux6
+KSEREdflTO9eBEa7OCbRp/H0hrL6+xqsMVEH4aCgFZj3YH9FMfWbQFMWryEjfL9
fIkMjbK6D9HwOD1tvxgxEnA1nFAcWocOvTIzdi8TNegtv72MPIebagV3RAKu8lkC
bDeq0u7d8G2Ay+yuKxjJHg==
`protect END_PROTECTED
