`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+GaBtvFUlU5Ky+iX6zwgJ5H/PuztVUt82HXw6xLGAxmoq+1YKA6GQzd2i9lejyc
OfbJ5XKb/eqztAhoD8MONCgZJV+l249bU2WySX6c8lnMD+RmWLZxU/HQ6DVuqdey
w55lkoyb86V5KYxcxT5Rzl5JNRXmbRwnZawcsRHGd63Mv3Mpf8mNUnYAtnId1KQe
G91lCdvPpLd9i1qt4SmBvBeSey8gnyBHbtCr88J/XEpb/wtKkqI70ROfYZ8fZao/
l4nmuRVvGkJPly8KIvJDSMsge6hP9BWRaiKmeAkuTOPUUARVv6iWjLVr9QSc11JW
4FPXVEp+sAXKSIEknQHMc3ASyz7Nyji4dQ7UY/fRDV8SLliicXddFOIZXPEm8yiE
QVLgMXahmMjAucJhWSgBT6NK6/lzf23pbuRo2sRtvOFyD4TACyBqF3QpfzmbPcO/
`protect END_PROTECTED
