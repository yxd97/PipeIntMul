`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1CNwLneiFlU9fx+B4NAmhn2CRMDbDVOtmSZnS+67Jh4//6sXlSSDpyVTYAl1owa
f2r8bPqzJsMb7XXTHtM0gD1JfVfEgLCAx0HWUs9MV3GiYXnfoadUgS04bTMZtoth
OFNe/TFqBwXTiiF2EaSrTU6i0PKz4svgaMa9nS2uZPRM04cmy+e8f9wkidXEQ2I+
ggh6vZmFDuo86KDjtRpybJBqGyPhN9cZe0bCQkjCdUmuACRnZ7gya6CV8EDPLGp8
rE13hc6DYJICf2DacUnJEcKWXkhYSFGZn/oXTXC80WSWkO62D0xUSgc548x4IW/+
87T6WFebZMC0PwV6cO7V52PIP0oLO4P2EOy4GE3D321HumIIidigZhtlMEh9LXtt
ntvxnxLrk4HbEGcVp7Oe8g==
`protect END_PROTECTED
