`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPwO5rXSma3AwU7seiGZ+lDv85hOrNMJuRShdVWv4nkihZ9u2nWvrzEOWrm0UZE5
F/JCQhIhrB5+y9hLFbQDnTY/pqxaNFDmlU/4lvuXteZJZMcUjX30hvsgbosWYFeY
FNxU7N448e47LgjUFk/vmioFTe3hJnjeaYpINMg6ZUG9/OvCUrlttQOqv92zOYsG
nQoUo7ZotWyD7ULzTBqYepvY+0+kx1AdGlopovLjQ0ybNVNmipzPI9CKgvEidYUx
KlOgR6Az+6TFc2xHhgKYDQ==
`protect END_PROTECTED
