`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIRt2PjcK7cacqfRSWx6CzpcZP0X9DNhBtag58nEO+4yWaJoC5nBEYcpGGPg56SX
AhCaiL21n8riXK8ERVAIP9D0EJCpuy9r+WxA8QzgEA5nVfrhsEtk11WzhVJWcg/p
rNzWAVLMqyTocOvGbrAcMoly9NSyh4oEvuxXpBWNmFZLoKscRm5XNGoKPLAIFe3B
mtRb1CcYzMpTS8DqRgNGmYnj1mLHUxbdWdZBCcW9gCAIm/973VOoRJxrnQbk/RDF
Uhl5PCpaGSnXCmmaQp2EgjDwZ13/iI2FqZvqf+nfIgSHOShZ0o/HNY6pBHAYwHhd
H0U1U/ROyO52vSNJKcrx52YjWWINpF/Mn835e8W4pZTv74qXw6PSL3+ttYfUK7sA
ep/RBezmncD7TFVCKQLoc6U8WgaccjqmEnQie08DnnS4Y5Y+gfmAlX7e5SyLhQ3S
RCvEozHhF4XKjTsZeW0SpV7Ad15pM5dJOQmFeDZYMrae/qw/MDwZQib3KllPoL6F
fm+SUolKFL5H4wdVpZ+y5gKOrGlxMqcWb/0JOzfj0402q7LeQc2ObLFKaEBkeHzV
ff5ggL1y4pIlZ2+SJQTGUzSBtBwcHWGgNRZBS/VkQRMG4Vk49HfiNNgEizjv8m7S
/4YS7QxejR1kpzNEnbP3+5oxEBC2DTwR06lEaSBjKJSVLZf+f7ef6ROa4vDgL+Y1
kSzXReg0wjXW7R7f8N3ZTv8qePlUBnvfnLqs6kxaEJp6Da+KlYyAzZS6dyV3ywfM
fZUFlVaig5s/XGIZwxCpdMiEDpMkFf5WidzqFeFQP5odXJAJ1PGvF2Wz0yTN/goo
WRPQU1+4ZYM5uyX0aqRIp6zAqYZQeqURBW7EUAyIbsH3kizdTmI+ol0pdUerfixy
ER2t8NR3O9Lfryafnf6z3Jd1vrUPAD9I3HvKGAS9OPXcaEOppg/KTTj8mixWfjDZ
S+hZHOMlW4IAjpKv+QEvuUCrqEhPMpJDV5YISTRQtonF0660GAYDL4y0/rRpeFb8
FI43puctecq3Q0MUs6TO07l//UgMSyZDS245S7kR/uA=
`protect END_PROTECTED
