`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DC4pCVcZ+ooG/pp7G3D/CXBhMjGTWJ6ws7umDediLBy/DC7r+IENZ/72Z/In2HGH
Eb8UUcvPomLOO9XasYX7prLsTm14RV+wwE+4AXCoT8S8QfGnKy5G+d3rc9Hl1hZf
W6TWQhfLJEpO8qJF0cdeeqMzO9vJ3TqjEk77gFcSkK8QDaVS+j7pB1wbB0Bh0IIE
VSYQZS5IDQKz9knGwBJQR6I3CZ9tLSu2wL3MsFzHWM0ZAz3G0F7eiHjHhKLfIbMB
aC7qRjKCpYJwKn8G9pQoiluucRBiedEaZbP7u5Q/6khmm6mE5GtFZArFRJ+tqSyX
4dvf86/t0/gRX8vLgUTERr7P2lLZ3j79e8VaLqn14/RTFXkoeLQTqQ42KhhnxLjQ
eypVhX6kBHgGQUXZLJAqIA==
`protect END_PROTECTED
