`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2YUIBmYBXtvHnHyXqlnkweMAcC4kxDV7+Ar75yN9VtZiNYh7iYIuwXd3W0NGiisC
dHOIibEj+vBM0oXbRxnbwN4TSvOtrvP9HjiAx3kIsSbBEjn9elTX0zWomQjayWBu
XABe2xdWyKPJYuaqMA8kzPWVyi/6T9A6WBPyNsGcZlG9UG4LR8zINyoIY7J2Ejz0
AzTIW0g2eKvVaTMIL3QAXlikyLbs71uQRNXLqx9EuqjT3bJUc7D6nX3TuFBcuctJ
MqBsJx8rGFFzGL5snty/2K/L3YfHFfTpp0DxawSIiiVyrmrKm76eQBB20wH9lFpe
NZIq6vS2s59YWrsvR9QqIBGWTpCdBHU49xJ+K5oaq/sNU4VixIHGhj0X2uRYdnew
`protect END_PROTECTED
