`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oEZxOxhUR8CISuBXX918IVcOU0tp//tgALf/6bsAAKBwRv7L9l//Ag1pQrkGRNDR
2L7RUo7yc+wUWa68yIzH70MFn+vE+6gbX0gc/AGM1gmgVD9182ZAueeN407ekkLT
pm3BAHba4nBz6TK3O+hv0TIno214Pt9MNoLcJUsCOmfVC0FVHUeiowAEnlxksSb1
w9XTVpmQBLnp/OnXR4sgFnvaOhG7CwSufSVFGAvlRrzlGDQkYVt5tZ2LloYGL4aU
naGeR0VEP6F4U1nzas/sSXQNq87xOzhzY3RbHpf2M3B6WzzmipnPYgkewb/Bwu3c
ruQ+/tbtAvxUhtQln3M+RA==
`protect END_PROTECTED
