`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iD5SXL1YTRPuVa7xRirOgktdBfzJMNbQE1XamcAwzODPV1McJpYxObwqgPtjCN87
siB8su7Jb+uAUhJJmq3o7Z6Yz7Tx2NT5XCvFXGLdQKK5K7YYXuGsIhSQIMViowpn
yogde0uZDFh86XqYYnljJjlRi+c2UTQLCTKay9yUG20RJgNJqZyYJR8N7yC1t1NS
tUs8GTd5tfR1Rc8SD5rAy4O3ShyHTo2HKvpdJqf2KFuhXoBqph63W18tdgXyLZKX
3R7zeJ9Oj2BrYQ8+5qTrxOdTQ0n/TooXd9xoPr5oiVyVdqW3KAiRjyaC0PX+77p7
XA8XE4hQGKj92noMM+u47uInyYuDuAwYImTddxfwOcTsPMiUgt/rM3v7j08KSfvQ
eXLBS3b+DfuThPXR7XIh0iawXhTFu4fuzY2KF/6D37KBSYAln10/TbUyKn4S9WzS
8tEaKZra+lK0akQhm7hV/g3efnUEnFBJSwonPvFCMdccT+/ZDSbIS5uLGEUzsyZi
+BLFaHvGV1uDUeI2eGmSqEZjT8nhVHhmyYGrifmhYL7c8MA40P+dia6wKLN5j4xr
aCSdMRIce3veCye0QiilJFMJqdpLDk7auTw8y5lsUmGqrjGfuYVG/1Hyw6SjBwbH
KwFoVoD9NCpRx9IYozq6T2nqGgRa4py9p7GMjtZZ37KLSsh59UHV+ehVnqU/c5Sg
htWS/1AHuXz4LUCO99jX1/XR0tReZAHEsE1FCngzOoSO1830AUm9lerS7KRNMqxn
fK32P9xRW3Txn4Na7PO59dLyKu1+NZ1agUGyvdkPf4XCpJuiG4t4daniaqVF1U+5
q6DrC8xuDgbtI7q0nmob4PfFksWDMKEV7nXdU9NLOWh3WCze4VdDTW9kvOLtaeD7
fKw6FmVg2K7bD6zGgOqMzhSnCUcfdR3IS6C3uck86kqNs0J+8a6uBjWEtYFq7jOR
OwVkW5gDxt5Bypm7sF5trL8brP9kDVMQMC/feUWhTZCuS2B7R61ZYI8QgcnyX20A
sY+3P3hVwfnoCxiJS6u2rtdozqkjrjbWz9VJD54FpAcu7oRaRkpxTQ107Y+Zz1oE
uNplR6AnnsdfBVa0AmUcPR/jtq3UNMem+gtg+OEpP78wxfYzQJO4ceguVVVCh6yR
5ODa29umcqxqx8tFP8WHhHnziuyioziajC9ffGEcm5lkidko+LesrvZf4FltEZVm
b2K2CQwRgndZQXAeCJYk/EBexko1OiLU/Ry+NQB2etxEfci6eRWezkiGF+VxgD8g
ht7YuOhx0ryXZLam4pJ6JOk/CcJaCIITFGnNbKrMy8M1O/Ww+wsQZvmsQC1Oyv4t
/K1rl5uqTLTIpODy9tHY5fZtJCX0S947REnPPnLT2WuvwplhpuW6a7gIrZHf4oyH
aDMCkyb7zcfd9G0nIQ5zebCQyaIliQH8KV3ZbZoEIclDsPNQOrpauEqD9JVITFGW
kpnpu6CJAomS3LBgRF/+cBPvgLvkmaCqgRn0QKiBjvwruNkETz1fcS+8GJ3vet8a
C/p8QXLyJS4dhDsxyv4OeZKc1oC/a9pHnWHRXRSgrYz4K7zdxmwx6fT1J4T7IGmX
rP16MiXQ8oofidRU3CKyuMa0sBaMZag2JmaIqPEah34Ce7jB+OKS/vw+39iIbYi3
OdWMpwd91UmPlV+BYUrD6qxxkYythhQYQkxxZ0h5UkUSDl/Su6f4vmDgZ2k83JJL
VM8YpZXRcUgtoBd42DjE8N91O9klP7Ilzsaom5fB1ba0qxkDJuYsz5+3y5mfe3dZ
5sa5gQVa8vxj+I8Ef2SHKJYU32L10ksN7EJ8ZgaflO2jmCEnEmucwfk4wLr46R5u
FNV8mMYfEFxiQKOGwY3ZdMkbBmydkmZeKBQBLe6uYt39ULRG0RH/ek7/WNpPR2/j
RJowSePCEFbbrBK/kVt+mGdN832obP0ArjrmivSoepYkfATkY0ACkaeflr5N5zNU
Xd9c8h8Cy2/+5I47+dzXxsooGgCG+dVZ/KQfSZOFb7kXMTgB1mQ/Llq5r6AbWco4
i+qDcTFS9cA0glmK99/pFuWCAo3/9XZFVkOfs348AxtqgNQwxr6Y7h7nrGUxtSZi
1wudaJy3Se6pxivg3EBmp+lW1f64CGjwdQebkKrEpniBAaXHeUYtXiw5U2WDgaaV
5uTZssPmj+QK4EjyGYVRMPL0YAcmIGhk+rWhAYiG8t9NU0k6N0qNevpbVq+eKaq7
iqzY7h8ng1yuMx2BPV+WOYKEyg9jDEjE8s3rrMJLXAqWcLnIsZCuAbY6SyP4+YQz
1b2eWPGvutm08UzAXHfzc7WKTs/uA7WSxaTBCDpQA4avItf4M6iyEOb3nxIcecF/
Hkoe6J7rqnGLsGGQ2fepowkVUjMvcSw0usZqn0eDBb4jhG+96doA0C5/h5T01PNH
xyDMqr19BzYhgDhsZTlWt+f2Xi9Xxl+XgmvSM9On0ZZVPuoJ9OYqXMhyGPNM0OO4
QaVi7bUk4OxXXItdDCpB1cA8t6ys0l6bkr4kxe2OM2e5XoZkU7MKa/D6ljcSdKfS
tAmI4FjzZRmDt3XHFwrLpfVqH9Ws3YLQTcLZxUDdXyMIQkrt5gakM21pgM4Wv0ch
7mFOiCgQolfesvNoFBB7ayC/3fJhUxrzsKAqGgfOxcZ1fKsaUzZblTOYwihsDrpu
Xs5K9XlhfL7a88J2FubTb4xQ7rB0bB3RSTc5eKA49z5M3yk15mNi4Bwmbt0y6sgK
N3iaPZvzFaIhmYoR2Ic+OwXy5DTAZjwVv66SBl8jGSDkmUttdTJRD6kVmrdbCztL
tZLjckJdH/4TDyQ48hBPLQXu4HkYYr836V8qu02TYBCNUmJvprXrD/YlELtrdlBh
KFbaUXAjqh5e9WsuEAoxYZPNKGHVznEGQRcFSsgqzsTlpu21hmHjNP0K/8zHwfeU
fcvrsrwBgHE0P8O/VQkh+ghOKu/gc8OHah4gAe8fvNNko0qlnUxboGslKZC6gyci
5WzEhannOIE34eaeM3BiGiHZ0MnsaW7BuxoC5DlzrnDVkxFIoJPIsJLLJg0XkaJk
Ra8D2XjlrplKO9R7xXAkbOFwLCSvW2tHam23rLaPeqfTZLMMgmDT9xmraqripAqh
ZpY18YkO0pX2MooXhjgTbMqqPBbOIDZcD79xeI9nCJA6m48dWo+JbyVP2Wl0CymT
QIHLVuDXINkyZZp8tmy9iO8Nc11/NkPBJI0DQZWLmp6DR6uwGd3HsaHJQFffuLtU
cx8htT8bqNDcF129usMe8g==
`protect END_PROTECTED
