`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRLzTKc2OjcxnKLbOqDNlMNs8PH13gUq0QlkqxHuRZAmnWosLXClNUGEPq1D7Slw
qccHZ7VuhISxhs9dBlCdNJiuZ9U7+r/cfFYufHjWUw6x5IFybXv78T5ShY+zcOxH
R8gn5BOTyl6lR4H7BdDIzvy9rmfmhj+QdLvmRkwRTiSmiyHhz3sysHkxzGyE+e/f
IZtrNF0IUgZBRaVO6ZQVF6L5TMWIP/U2rC8eEexL7bhVR7gemnBGg/16FL/tfFt6
V/QuZcjJIRH+NoB8XnrV/GF8YyPOQ0qNHd8RSxBJ43VYxI9c9SMzRLn5J5LJuz3D
VzlN2scUZjMAat2amkQfZVWc3/qAyHgopCjHSqCaONgRlZhu/CUXpYJFcuOP1jCq
CUrvbiULsl7mDiiH5l4ljZ9soD6Lq5ZAoxhpm4l+/mBwIrQHixNyQnUu06AU/srY
t7IjY8QDCU+GGJ/lBNoP4/QY3CUlp8bCKbRl2I6xnodeFj5FnApKA6yRBrH5gKmM
Jk8NumML5ZZFgCiq36R0sWjCt4+O3oAgMOkM/qVepqMXbmQsWmxcwOBpmEXPTyQf
mbnVXLtBCfdnPkUeHaXwFvhAePZBUMRHT7b53ij1PE5IfICOJr1M11CMkKY3wNsV
OvO3hTT30rDc7ebbCNBnO6WPRsnISgoew8gF0ZrS3GMSW0HrjNo6doGwSuAT0Ab2
nb4nMkfX0iEAcZZItq9eLpDixdjqctpMvIj4K/YUCTxXWk7kj7nrcQvvPG2ezoS8
5PY+Jmy8qpnjh0fuD9BXdhTJxapS2Y31z6cyHs6bEpjqXTGPc5+OokO0ltM2FdPh
ERNDJoMyeb7EohcyGKo4YR3nid63TEM6nPGjIDUEhTk4NNS13h3Vb25yLSHKTCQ8
sqHFEfy7uvD7QnY56PUKQk/F+FUozm5Xh1B9MX2MCO8WE9+GC1lHREdLnFIDIVGe
U3E3hItCZfhiPQw6A3TTM0xm7xA9EOybHtizmsDEzd2whOa4DblvZbEhcS0mw7ZE
8zUEBMrodtxsydGm3r8jp0Ffx5lVQPbwZWuloBd9kWDmWLGVy8QYcYq0y3EVxz7B
Z6YqumZuykQMRIkTSIVmg6EFAaRWRqigHtiR2xYAERqIOuD2LToVTx4HKoHIGfAD
kpZkafw+PuOKVhohs0vI84KZqGuYMdTe/TdJFlaQxq/3S+xaX8rrrUy8mE0NTdCE
E6jXLff2SykWLo+yf6QuDb7XVYYQJUIJnrx8ZdjNASlmW05YUsEI2HjvnBhzQhjL
I5tV2muYvyW2NhWP1PrTFciesfvhzep9olPoAUUss40Y6oZFBFcxL1aEliurOQhi
0M9bnIWjZMuOQXfmb16/IfcdxWjDr45mbisUXzdyFlB3N93B/wxLJ0c8rIjJNkvx
a0B6K7JH4Vys3Z4AtsylfyVsnEBZTrrDeydWbalSt4PjoUmfKOaSYidSA7voLs/6
32KJe7v2fuqJMP+CjzQPzCMf5QNPWCI3Y8JpxFZ92JPgqVNxI5uOC+dwYL/XiTsC
a54qTMSLQfw5q+UCawJcEiK7vl5WtA/OsDj45VXCPE55l7Vry7SFEgaEIqj2v3Db
hSJjdOa9oB9YRZRS8BvNm5ELNqXgIwumRK4klo34nDMsGA1Pzi72mlb5Yyf5D1SW
csVTZQy44qcRKQ0YTm6EO9Sq+xNCX+gVExqJxp+LsIX4rRmx35ijArbQv6tcwCvH
kG0zmInfR1m3lLL3D2TJJOGMyX3vykzukSWOnCJ6dAsStI8TA+iuWiSNWsh8tyui
DNYhK7cDk7tEtNUn5uspEvMgUZSQ940XqEbs4WCNvhVnbieKQTNZaaR9xTQeIEvS
GGQqyArf1Mv/+WpUThzvvnROnp4lFizxHZiXJg02Z+dc47iqQpe/ydOWFu0AO+Ad
QdLt4/pRyCCxRbHhqfs6DOtnEihEOnf9/JPblptC9nPrU5swatWViQCq8gT0gqsG
76Nm5yQ/ORndEoinczp5cfSZmjaZdmPeVSXYCJr2uTQmeh4NDCPEYwToGxc6PuTn
FBKbxGS3tjmj1pwO9EhNqj1bjT2ynlzaqUSLKCi9HOG3i16Kp99xfno1o7FS2aLF
bn4nEzFDCiYVOUPQZa0wMRi8RQRgiLtv+OhC8XJi0AR6r7312I+wyuVBlngaIVJs
CMzmc23OjWr3czKg0t4vfn8WLaHozZL0vXnnfRf4T95Q3BgXCRBJBiS0+5WdsRO0
M5+nNTHVTGSSOuamYeKSLIHdT5FR1DmgMgVkzDZ15hsVliWSwwQhzJRNcunZj7XE
+cmjOLK4q2tf2/uOtr6aOjdpYdj5cjFDpoZAbWb5+VdxHoEVz6pdi7yLSHNLIDjw
0vdSxLivO2vuNu5/EF20y9itEghcffBtQQQw7yRmlKAbHmNDV3ZdB2ZI3WdptFgr
DByAaEHiaipJRCMuuz4ecCUe5NNZ/eXkGXj1hhnn8hzgzVHPsimwdSRH1WijFp16
hClfQlPtwOk/9nEUmFocYf/oCu2geYQ7P61aFdWxcyv6h+xq51cfe2+fx4Fjr/s7
V9098IyPKCT6UZrvyAYu3cpsEDa3RR0TcDcoUALoHDgQ/YFoyAAYJOpkv6Sd7sS5
amkGPo3pe1SeQZ88eB0OMQ==
`protect END_PROTECTED
