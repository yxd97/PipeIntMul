`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mjslFprWmO5raRde7OkYg8QgEBHepbltWM8NmlEB2bQwnP0sZbCtKSCpzPIk/FUj
KXrpwWZniSdCoMRZeY/J1UrAQVwGMTFq6CogTgbnFoWxP1EjK4rM00yv9SPIqOgd
38VKKH9VjoQGPe40+zPvK74CKNFFMh/Eay7GWCrhgStndTZnr8L5etlKHnF0Z0CR
uuM1Cz2xDhfOKCshJs7K7YnO0EqH5cEuJnhFQFIFrzrYooF8Japp+G6BSHkS7/xf
JDEhMZVbuzWRBINA/c2khBd3tmFOIs6QOM0AO8mBIwNvUAeLEZ5X8/KT/2eRwrv7
sH9ri79G/mRTYmpJa6cTNfN19nW9jlx9Zc5NTntNmNlcM/JwS1m27GwsOisETJKA
hFFqqaWw1P42LRAk57dEOcduhRe/Zzh4+bIdwKxOdo29jNOFR7p1Qa3BuxiPC2YJ
++pYf1+QHZeFRK20P2Rl3OaxPhcrxy54Q+tF+JDB9/0yOFj8bLepQLXt7tFq4Hph
2MARlj6bkSGUGN+7r5+fNHAdaWvryuDvdLOKp0Sbp4zSyOPg178zgEwNnuw9bd0N
8qXv876vk5Q53/QT3pvlSqiPno6hehEeth2pVzjut1PMkFXH7rTzB92IEC+oNDDf
qzHuwL0jC1+35K/KVDC2Lap3rIonfEl6vSbSHx5uPAytvFG2tYJV542dWcSibxG/
mUC904CWuEhGQZ2Jctzk+NUXMgXtpGYFB2rDPWjxdcqA3AP99HqyjY06/qU9F9YY
q+fQ+UdbbLOLYpNPFq3Zp5el7G/NiFQubmnsTIALmaUMftSSatjtt34c7e8iW2KM
6Bemx9N8q1CfgE8zNi+ck2M82aOj+ZXp1m1gbIKzPYNiZ2mg5as/mDLGTDV6nw2V
+nfkI7/c4mdlrvg87aOvT/VrnDRadFY45Oaeijzyt+iYNRGSyj3Sp7ByaKm0MCs3
DmOaiDGB1xzfIMQ/w7Y5X21Czi6jekTY9zxEm5bpJFvMdjTQCxKVOtPCYEtMulGG
G8ui4vFtiQolr1AUo5aM+/uzTGW2ikIncoimR/wSAldnVehDYNfM1nqwnCBb0WZ9
8mepLBkRKDkQjRI8E17xXLF9hCaBccojh0poPDm5RiRqJlUhpu9LBNLGuWEB1Y5p
vPTrZhxdzjzegQRbUFwtG4tvG3G57HBpm/VJlKgdGGxg+j+7hqmtj7i4qDM3jXGd
QNTvZbN9iefsTM0L+vq/zefOidGy/xoW3xYlicXOCShw4mer9Vl3V58b7+flsqat
lgGOhhGyexNonGOl1SR33rgfVrcV88JKKcx2VpPtDvHt06/iUaclAg7UjCKxL83U
Ff6Xf9jQ6Ko/MPkdH8jweiNTz4hUHh5lkE2Zqz+ATK9sfQ6aYYQXx3FSa5dG3FkV
L1NIPEKbbAnzdntfX36/a2He7EP+3Y5V+piCY6M2bqML0J4p4fC9AhNslelKw9KY
u+i0Tho3YnIyIk/kPt1qgS3F87KOIqPExXWWTS4YO2EUMKd7IGDpzu4s3f1I3Soo
LfZa/oXofhUG25PzyPL6q7z8645NcAo8kwnOZY+l0lML2TdGzblawGzJGsFufHKX
2P0xWM09/Grc8pqm4KkKpqGeCrVlrvUbcPOTtKg4T5DD795yu6mu7RdYFKihiysk
N3ilxLgtRfgZ7+4UOgjvTnHkOM25hjbAOLXpp4GjJ9+LwBSdAKnMKJIRU4xvKoFj
yyu05GdTXVp8/JDTPuw+i6tC6eY1z105h0GIKEQMyk9orL20Xcg1iUOksWMgvRn6
FFR6Eu+FJXA6te9F7I7sNL0wuf/RjyH0kbLVQCSCH0FoG4fHgHqr7a5RTwSGvxFO
EFWB339twL39Egn5UYsdH71Xlo4pZCRaKR/FTJlElOLeeU8nOHUbyLuPUAqtJEXb
mx0vZ9BgRZVk9vjRaTqOkBkwYjjohifhC4bK8+BIGNbcvzTihfbqlxgrbMRJyGIx
aPzdsC3JmbIfunG4jXLfbFXb47qHqd9zu0uF+g11b4TF2A83k4wDaxTXah+p224A
Ssq7nj31aw1tLUCaR9hWST6KvZewlR/SEboCEFlQzqKhxjzplQZQUFmsOBvFBDOB
gefc74NqTCgumAzvsyQjJGrrhgDtoXZhbaabTiu+iBcxXU6ynmsBJyoXZC3U8Phv
MfGLACUsPN06Nse0Lamm8B2L3/3ZP+fhiAPEUXt9ayj4MyoNuMPzrkRnHasMGWA6
4t3Hn5hFAhnn2jTMICBA7JySBcJjDX4s9iahtUdcYvxxDT1UzfLqlf6e7hbkensp
B8PisfjZ136xq+tvJDIEG/JrtP3+btWf5P5CtFV20FxVey0XdH+jNYIPNu2WixWM
hhf/PGudKvcBuombjIoEPlRjZubZsjBJUL+4XXAcvw2I8WKWmMkhER9R5WIahpRV
ZMy4ilg4UzZMaJBsogu8tGhwd3apfnh7VOrAT0cxlqTQWewLkU4CP/g6VkY0sLKR
xhYUOPXtedgipru3Y5J0cxEE/yN3YPc0SCPwrslzo/YJ+N0EEGKN8V75Y31BNwEb
gsi22v1QH+iEN1Xl6rlGTyhLnvMTC9VrqXFHukgKqqRwuVU9TDnw1BVv7pu8ef/m
AMatFTai70gcTAV6yp7uu70lZHh5ZIzjKUdxDyI/XpxWjdz5dSoq8z40Y3Ny9yig
kSsjJ2vLz5G+ZpWN6bn0165ftiHVL88aXGdq5+i8L3lOcwMBxYzTcOjOgf5ZYXfN
cXI7uH65mVF/yddDilVJtz2LQNtf5hv6d+KenxaCG4OvJ5P40KcK79AUhaY9XqP3
S0iGydz91XluREZl2MscdyZVqwvulB/zuPJMviayRB6GXYdhf2bFr3SHWclCsgfz
+m2UWyigjB2YZpHtAmBsEVXI0UKnBA3lzkjqZzrgpJgrvQoFajcgxr5cPUgOr+Ze
VbtPeBjkBddMO5taKz7YRGezNIJGb3n6TSequh0wY/xyAAKHVQpiMVRL60Nfywjm
NLkJIaL5/0Fa0TqlUXQSAO6v3GCsBhr6OXDGgLflnjTC/sttJqy18TU32gVS51m+
fRwa0pBHt4p3BoEsVPjvu7WZS4sr4I8bXsT5kAxWGtYxR/1Wikx5wF2YWsz5BABp
ssNJ8TWSIYXfclmqL3UgO4jVh/X1pmgwxY6mbefvAeQLhRAMyuxSGFOc9A6LYZix
TK5m60rW9uuOM/63Wr1GnOlQrzzACrXJ3pKCy0ik3PfPJ05uYiU4ZHsPm2AZS99k
haLSiV9TzHfG2VgHz7gmudT7wi/3gCAc4e3zR0HITmnwnEuIOKG1wxrosaEMxWGx
fOrFUZxLWIkvYwAIzx+5tEMDXZmQ5wotN+sv5PyJAyhl6qWlbrnhUSpYOv0uplnu
eVhfFI2bHvOq6MQiANmWWBF//cmstejPikwq+xDj6U8lnJG+q/PLctUozesl4ZBl
wEhz6R8s7ibJysmMWuELSuICtm7v/ADEHsEiOQuz2kK74OrdCrVvQE89k2bVCQ+3
xPeOKvNuT0URVudUUZ0Cs5TIwNQs8sTQftmNyU3Ad7DE1O+p/O29Nis+VOwt3adO
tP2aNhgItLMJXRkFF8cjZrBz3vm9T4mP318rZ0qTyptnALTYV7hgDrHcJUzNsxgr
hITNMJTFacc5tAK7+LoQcOw+LSdVCLeZkN0I1qcMvfh6n2FzUs3Z+/E4cPPB5wpa
yt5A4RQJFcjBXn9HXzFWJqYxk5gRntgkHO9/R9b1hOXirkjkhrwVpGDJ2jlYrLZx
UHonDKNAHq46dkLbsuA5rijPhTZTJdbDtvsUCA/Yg7HwOfPZ6xzJ5+bvd4XK9fjm
0EG46CkIp6JER4AuL0m4yt7nApznuXfKcmywbUKOpAj3b+KVzXW5GQg9n4vt+8k1
1MOozcQPKN+LTRxlF7uMynMfCqQX9dw50/Uk9Z+5jtQcJKulv1PYRGeQ7xFxUenk
YCMoY++2qqVPO2SnZH6SWYBV3OVg3YiBZ8EBOk/O6TTK/B+IcD51BqxlJCbriY7x
mRfwJ555y+g7XnWdrhvGRnG6DVvct5P7kUgX95KE27LBggqgBOooic3L4RQRxE1r
69wEOkMeTzFQ21PeNxWN163ViQMppM57zcHfR+crugoYNPeriQyhIlLwtKEGKv3C
wFaRk/zhXGXAZIo+DYL4c8U/xUEdhBrf6o9wlhQG7NTHMfAy1i//mQJzUmIyWolm
ZnKQmGg7zV5C60LiiekRVcrvP6VUxXRfJesM7rtD8q9lt5+ph+83fnbVqldkLtHv
Ci1uQLznodtuMVK+zwagS56V74b9noqDXUDY04YtVEmoHhbKf+B4yN5Dhqh7QGf1
i419dcygA8bUcJt0M1wXNIy1cRC1w1Yl1K/MI7+1E8hhcCvAxCd4uwOsZT0LfIen
bQhB3NnDJbvw0Yw3PN9yF6cjsNpWT5JDQ2wqNfXR+ZIx69+rtjaNazFmt0Tye9mS
yW0qxNl/tfsdhPI/oQK6a8jJiPFv+0xlbppQ7tvbG09U6FSurnRbs9Mkt1Oj5/Dd
bDWaqQFkOXDDxiaZv8vVyIveQDnChgCYL308SwE9QGqoVueF83g0sHQYvHcgpvqv
0hKwi4EhIZh8swYdiJJXqDGPaxInOV5MWYnVuNOYqnZXeY/dhYJLSpM/WD+cXF8b
Ubd52W5Ol6pU9bwVeRAoem11QxaqvxZZhtELZWDOeR6oCrbF1wjipQmNnKgM8iHV
0DIu1wNATwBCQTsnYTC27u+WVO5PEGr4leKOOvSh0r3gEBf1NvqcZkdf5q6qibc4
1e8A7IWepIUv39QEd0hSzggPrP25qSCtfDFWSibyiTNazE0Sj8kuijVbzdlDz0V5
oU3sSPMj5nSvHX7BYIfzI1po34+pmvSTlAU7PkLct7fDffKRd49NGTmKWTBY7FQc
8a0qaJIERFXh9TbYweZMf7NgrZNvjZBWAOPjLCeq6e+EFeVWJVFWPnj4VbqnAtC5
9RCyZIotrAi1iqvdhU/k5Ndl0exGRBvlo5HpNBFAvSaZusmDBkCVj6uyAbLzYZpt
CxinLrlgo6BhI6mMcBxLBHpdy9byUvy07kU18EGInOWlIzp7u2V4hKFsBwdRC6MT
BUuzZL67DP2GIuf0Ke+n/yaR9p9ltrCl8clWahVjsFgQSCibonRdWTZpaqsZp/hg
bS8nxyjMEEwRVMYEYcoC1odtRPr7iJbyE3JQTvtBmNShJ8oZfQWZgu09Cu2KrJU+
NbFDYLWm6y46J8Z/DMFzYYBhoIzCqs55pIDl3G4OfMiu6qGU5hcg+1jlmZ5EmhPU
equYDEfE7TX7YSyWI6eZXLIbw9KL/uMNAA9+SLiYE31S8gUlhS8F1gafXUvhtSK1
Cj7Ys/5b9c9LmNhl8obTG+E93DYjk70cxCXYA6RhrVDZMrow/yJ9nKMCqTO7MLIw
jbID+Xmn6zCmB7x41+vGL5yRj+yIIHDqhef5tO/PpNVHcPKguSkfrPejnn1FOmr1
zTPyyKRjyUVMZzqxrdaqtR0UGGSSMkkrRtxgZ1f65mrS8epkgU1T5zyYRtSjwxb9
fi5T/xhD1VF+doVtdtlg6hykKDka0Lq/+hEedGOYMYGOoWkD6pE7m73l2vucVB5v
H+mHez3h/zS9ZruykyhOAHd/ssTlz5pp175lgcNItALWEd8i0o1mlIrc5icxeJU5
usdmTSptZeu9QbmYKKGzLdJNnUHpbGs7bxkHgxOL9JGNmOg2Q7gm8WRPcdkDCjZp
6L1M9uW3MNz1FxJBfqr822vV165xDzenrrFuXkCzDwWKktJSSZxRJz/F7cPLw5ua
wgJbSDgxDKNEltGEOBDg1WpkgiQQHZhPPJLFvlWY0CXMjluVmGqnJy9NctCnIdmH
WUOHWgyYj2DrlT6YH8esgnR+n3ay7uzR4yvY6+1sq7TF9h1g+H9aIbElMzwvyJdh
3gkglG/0y/IYR/Bjqm3JOK6h8gK/gzby7ftaqVmIZNglLTfU6FsA4RxyXj9jeBhF
IeFlCv/efKD4FjBYo3MeyaB/CHj8cjkE9MorrvbEHkYwEL3Xx66t8fM7YezorFB6
n/JFdKOAmyrBWHXzH6vt3He+VKouTjhQpoZdM2pH5/P+BDhgY5iizaVyhif4IrzZ
GsE+0opKDuOBSMebyyhelDBx+g0EJ+K56j03DQDb0IzeK8So1iu2w40ZAMmRXSGz
0bTKhSWZu0AC1lvwUEjCThfhnEa0DF8m5oI6y1gQ8+dfvSm+xJL8L81b1KAQlxVc
mECvmizctoBCwgVW0ZEnuEPtt0nao3dcWsOfySJsYZX+A2KomDkkjv+gMDwq+q3t
k88DFTpHW3ZCed5I7VRz72k7nwgGodOB85EG9I6Oc+8Yi5Xeu98Jvalov2uDZH5w
EhWDtwyQ/pvwzVgX6nvEwxR6zy950Of9MoZXAhqzPzluwuXxTNUACiiy+JdsDmPB
TASY+xmSMz2r/J9xYnVdHxAglh1n00UNOftVbk31k/aqF1vBhrxg/rfWhZ3wJSOs
DOGu++udnNWFG6EeAxGAADz34AUpLOZeJA5KMjdko0ackyaPIIL4rJqs+wlAYHHU
Z2rMu9kMaNzIPvj9i9iiV715Hqvp40W2VU2bt99TkmeEF1egY6Z3ei8YH2hD3a6X
xKMh8QzdcbXaidDIiHozLsQ9/jjJfl+9aPcp/wc4v+bA+ZJMqStjwIb/MtI392i1
OjzAkMGAhQ9Z6PUcTIo6TuenH81WQvtKaPL8QuGUzBKdwAMPIYOvW0lx4w+8mg3p
kccYk8xAcbVvxusygAEagE/k2dj4SheK6VfvzHjc3GBeBP8wMOb2/q/ZFFRZIMFN
aeU0dUokodBbH+qq5lxh/fgp3BxuYT7rGv2HPkjD2wbnngfuRx4jhO8beKXZFS69
lGMzeblixis5QU/+YwlB/wIc1bpVgtQ+D+sq9Et6CUUYxiwtj/+6ohhOz38NMuaL
ldMB3SNkfDOVjajbr9ut9xKzTsxlQ9D6tBi/XCdJiYE8wkiAFLtt/1jWSdc56q1P
SgMF1iKVGeA1fa8zddBmI/U2aUwevSdLvqykVTQM5VGzd42yB1gLrgz3BLz2OyPK
stWN1aHc9QQpYmMfnEVCUTXzap/HfdTz6RGh2ybWQgrkh05pDGheQ6sRCozRfIsy
HOK7kLi4IWXX7xhm66b9pbiUsvzkCOYX9Hie5wkIsN/jRaXmY22X04lISZK/bwFu
PGyn+UqYytWKuYyJ8Vg/hb3pf9Jq08+bY2YRpOz+plzA2afzR8H0AV2lSw2mgcxo
7csQlqPjgtSMjqjIy2OyePl/h+mN05cewdyNzvJERZZ4Q71S7SmwsKgL9LbGTyGB
rVAn+rHEPOuONMDQoRrQPm+tGvl3EYGGmpFgZBCQZV6IaYHnDAtNi0WDz6aOF/q3
78a8W+61PkGuUPVbqdwhbYPkclyCI5tIPTWKAXzRz5GWC3szew0046H9xWg5WiK9
+404+ZCY2czC7cLwogBHAf3pYRcgieebXmBO7M1nkz7DMvmIC7AOaw9HLvETvUZV
qvv2NNQwKgFNIT9XSUSgc2hXi3MO/GWpMZXYwDIq7O7BhuhLL6HFv81mz92ayREH
14bjQ0oyeJNThawGUVvd3dVATQKsQ+h3oI5MueYtnly0ERDfEg/9yrUvWhQeHnPl
CSx9SfoCKFGOmX5AiarSSU3Fva8zGYLpY7OAneHjFo35sJzEYD2EmaxSkFymFf+i
uXixVo2UmbwaJW7l98m0WwHGONkWebDfC6rGQbjBRjZJT86+kK5tPj8k/e+HwWPe
sLQNm03q8uRPkRXmlwjmlqKUU54OaPXdZR/ZHfy5lo0Y4JfatVMEQPSaTy54FscL
gxYjlNNXry/vdwNu5Y+4EXkZwAZQ/TcSLWMCDSbCxFX6SzC4AZqXaUfuuwnWvT6J
3xLpDygazIvqTIzCy+UQK0TH/ALLk5fLQWeuXv5TpfqSPKjqwvQyu/1ABm83+eSb
+RgOviX83vkiuRNwV179DnIrl05UEZzYBC+eT1Do/PqS/mUHjGOPPvQ1zRGClNR+
jtmTgQPx5GXGR6hpC9/t8VM5AMNe6gFriH69hjqIFeqvI6tjJ/Q/LVAumE5HvEno
kOVL7Qt95klCU16Bzp/CU87TW3eZnmLUV4mec4PwJV+cXJXgQydFptAve8WDshIZ
nMdvP+k07QTploK3rgIv6j9+HL4V5xUpgdDOLHAIeiMlqwCJJpxb671IadbGwFIc
tyD1k/kZZ01ToZaJ/rjX8UBDKQRM5aGA7HWTLqayLs+tnhOa6JGZa5P+UqUd9UPH
nqitiBUj9gP5ibD5TSJkKt2QIDW/pK9VpTR8Ne3n6x6SCxaFFKqgfIzbS7h1097y
Lkli5FKyXAziZ9QoEvyk6VMSoSPEdnDTrvWfZ7JW/iXfP3o/ZJI5qmtSkAPFFLFr
qi2PVkgbtluKhZFDpIiR6T2BPRS1xzv549LdO860D3oUKgNI7ae885yS1bZH4HY8
bdyF22Ps1YvssKbH6ZEF90vRfsZPZjMOvamla098U5TqfgdvlrNeEhpSKjB95sKh
JnAHRvusknMojy+CZ8ZsJ1iaZYkrZaVP+Sqv+KiAoHPv9AlHwfIrrufbRm/bq6yr
wSUbZRrWCwUV0vZtfT4Sr8pvlHp5iFsnAYGnoKV0Z6dBzdBown1LRn4Ge8oQcB6i
AaUb91J3MFvLrG518I0lGHsmEY0zpias/YTjcZbjovppOLlqKa2ShYrC7i8h/ONS
M7FiudJBbhVVw/up3WIrsDNqMtbXUTBg8A3fPbUirsVnlquKcpmrV0gyvuKQ9SAP
aUEjfR12rt6l0W5pkufnoZetEMzxgG/vc/nDOW+9V6azYLgONIsmXCzoHGQCQNrB
SOx4nKvr/X/iGihH/ZALVYdQGG50opxox/9llr8lhXTa0y7i6sVd/lzL3dhAYy4v
nWN4fZs+Q3kDedaJ6petYj2i6cff96IfMIOKghKLtdtGtjLoGbji0k8bmNO2juYe
DmP/7C6iC0Lh5BZNFra+TLqVau7Z5cOHRBNTvu0Ct5IIK2ZkSmhvfIvfIOUC+JbD
KFKq5DOJ7ENCDol7ek37/E/usXXJkYJ5mRKgaRHQJePWr1x0JsFHAUhGjZ/mIxx1
wCaa0w9EiOKVnMbMHdQEVCjwYF/cruNtjNC2giLb68Yp2JY9WUQXXxLO1YuOuoQA
JEYl4lQ/QWQnHotiGTRKBWnMF4z2ZUdBMtsqjJFNjRht/cgznLk5AKIFdjioVaaO
UyVB9tM1aNrgBhGTIDNMHLc7uwCWO4rSrCflz/lN9nLI5wfPRFrhnRVz6FxfcTqw
UbNG0YJifXQWy4F+PxAMn7vL0+FT+ZFnxCIws+JrujJzjQG3o4/oiC1Ncu4EylOL
hGzFKO3RpCtZUUYg2JehvtDcNYoR8W3uiTfOwpF7PHQQaBJuw+DMtZGEEJqKWuDs
w9+LbTPGrC57WMoTU1t/1PUYTOb6u6zvnKRj5aOBd8BCm7F+SwblbwcCH2rv9lQ6
ZUul/37Ue++OrlOcj2n1Cz/TnPf880PO5pod4G+EkprYpKCjSu8lManRDtNbPHt9
4dLRplK58OetgI95oWbIfVpyY4+qlK9baTN4ys+B4YDIjo60r6qJt35W6VdjunR5
b6DJzksE3QqPMJlpNdB0NzPRmtWfFVf890KTotCu0Bgjw39Deh/Xrgt57p8WdoZJ
XQJQwAPNkkuYhZjag3YQkLFlnTEQbIRWTwn4yyMmAiVuO/WjMh25nTSdOtDnP8aR
1nwAI4MzQ/dhhRoThS3u6rnDUhPF4shMyVVNq0avI2Hg4Xniv/o6Ezx5/B8xTHBi
QVcZqAKhW4rVVtqYw41tJyvdzCz7oA056mnINVpKzOZvyDk/PSNGL0B09avCCXX+
ErUEgWp5M6c2ZHYoVzY8MoBCHfvQHOD2MSfb8oYsHX0QEbzplpweDCukk807f1l4
qbY9PUhlujVcwFY1Z0uT8S+45Uc56BsANmZKUPReKsD1MPwOybK2DrLvFOiF950d
35WUl4MAz0CLOXacNBu43TwTEEjx5FTeUMlqRZwfQpwfKxXti5RFw9OjL0+mhvpn
QCVTaVUskaD6Aao/weeJ1LCMeCQBrmWG9y5CQmmcCvlOq2bnSIymE8Slh9g1wv+M
htK+2QS6e7doEFxoT3xcafJd09e8gNnAqCnYe4T7bdrcEUOb0NU/1Bny/ByRyTvE
ScjVM6z8dbTuZhEIw2Sc73Qk5UnNKjkddWyW5BxYK+kC3zJAMunNysbXJWJDXk/w
wbnOQBd7zCevjQfLWaiesVt4EuIVTDB9/jTC8Rl9U9YGc8bF/eAatBwvloLhueNn
kgzfOGUIVQ+nTOZu3FLfH0YvTkMrrfey7idM8nDyRxPYLOjKj7GmJ39G5i0H4LA0
aQE7QrjOszy22095PdfcfoIYy7FIX12hvOvXBRx/Bz++8hvHUMs1G+fxz0hIBs29
xpqJDGhEac3du9HSDre2kak02Whve2Vy9NBvIzfMdYOQiphgV5SXOLsljC7WkBL/
65yYx0Thqmtc1wmyLCZOrw2r6ZCCZydWMfE9V8TjG+D6W7BwDhtEXNeiyctITB1t
1um+utNzsNdquBmkZwnddkw+5LKpPSUEyc0gBBQXY8G+tWN2z6CWzpsTZKJMY9qx
b0TY4eh3iqXmjguLRgj731MkIDKvkZuYrvxPImOOPAOOawO997wFZ1f47ZFFiIGB
CtMETkYc7t0gUqoJcUrDNCIrv+XuRNiY5udbtpMUtwnAHoatBZxwnfGWJy3rh4hn
6EPgWe1vJMmc3IxHMtbdRdBi0SbKEU5tA6m/MFWyIOyxmaLh962tQLETAMv78gNH
VzsiNMs0edf49EPu/eG9HHNzdrK0DJRVIqRj57w+VYfPXlGewoHP77QbiQ45rk9p
zQXg7qX1lCsyNkTxw5Ou2cNCzOVdBlhnzCJCwgLSjWzsQYaeaNaI21yUGLNAzeMd
W42mLnlGabibe89f+7GzYG1/44E5QmbcqcndnFwNRrwZrR8PBI8+APlvCy0ggWJO
+x2kv+tq4MRZWX8R8LRYHQh88nPOrs6OQnF+OgrMlPEexLOL+NxloelGqFao1JyR
vgU4MBvnuildm6qGc2qBPzHsTvIHGpHXIaj5KvDoW7cWvDwHR6wMD1Ca0OuMLnfi
O+cAaGYTF/VLQaWdhwv6tgRw/kz8ozd8WIoZNJxCdI/YE02aYvL1CLMdgTEFxgpu
eoUN/iWseLxA18xgQw27jdUNa0xKoThk1tQJvi6jFBdpTwYKM2CViIZJrxTyirOr
gdcoSuLa0cur50v/yKYULEc0PIJU8iVQogAx95ldS712yP6Oypgna/ahro/Nz/RI
uOsSs9CNvmrf65BoWIX6EUkU0WiNrqK0+0xwl21yM19i+AghmNtFJBoKW1s4NwG4
fBcDZYYG8sfFDRhRisaCD8tgyCeLXaEf9LjVni2gPl3QEd6c0CVZnIBEQy7b42ym
WE4KlIT53HDEGeM13+E29BHNjgcVtMK7sRCc/uqsMy4ue6Xzmz7XJzgDR92cRtXF
zW1sQw8Fd0BEpEiv1+J1BY6GH7KBOqrXTcoFcan4TRuhUlQ8FZSCO5vSlgCbQ620
1gkqU5TyOYXjhrAJuNSMZNkcd9ZRjIcbAuEZOJ3lf1f9Kq09808g60mNr7LYww4T
m92JlSj5XL0Z2yUXO1T7lUZsXAOHh+5uyjHfTHiM4l5Xy6+eGDj/DChieDQ6wR7u
G90llXgqAh+UcEyP04VB4z7WKM6nby+nyHviBupi0ZO+ZumS4fN/QukjRkmT/YZv
rfD4euLkyc7hLQMWAHuSv0PzS1kSqHw4ldRtm1ckQIzVAB1tZxchlL7+NPbg6ges
ncheOCZeZLSa0CzZv0ibJqsaHIlnMgYO/JrFdmpkMxPjHVTryn35sRkxQ0TFqhSl
objJwbJz7IFp8c5BIvGN7vb0VyGJ/bAdpCOThSl+QBCeK1ji+RU9TPNq+IlbVBpY
nwZ5k8rPR7g0jvR0KHljzbeUaB+jgb9e2bcxVeO5r29yMuB/CaxTaSHyM1Wj1smX
Didstnndi8ce1LTCvMmDvwu6nXEBcnlkL+kpaect7y1ryIbncXHHR230NhI2+0Sx
g/jJtMYEAzV7n4x+nl1oKBDuynXKmgoKPVj/eH/p6XzcXfhfGI2UC2ZcQ+FBTSxq
fJMA9jJkQsLTCMmUYKeGUmFrG0BWSsZ3x9f1BNwT2I9xiEQeYlwB8XlFT01eu4WE
z+euw//6tfLcFBAdNUXIGffxtNSEPnvv4VTIcS57SmSwDPAgBfVyGXsFhyxFdOh9
UDjErDCNgQVKVAfAzWZZU7JczlkSJvAcXI2CwBd0EsSQ6zS4jNooLWJ1YoGNMbTD
dUkjNmBMXCQqPw4aMlOuGxvlnwnY8uWGkNjvHnCgktxI+A4ZHP72Y01VwbP9yWE1
e5s00wX33AUMJejoC7d4nyZPSL69veVeSNIkL929tyWOSr26tgLnJv0Zxd9qyEzQ
mlXWw4E7Q3+W3xslowCMpuFAgqykwvmq8/ivpyNjj9BDLg2MVQm6OHG0eySzVScf
ie4EgFRMVg0XqDRHRdf5Iu8lHOKML6gKpyd7GmIAeHy/J2mc/gYa2S2JsAWuSyPr
fmstpbN0DDLVEmiLpxOg5C+epJq2vBTSM2vppsS1PPpyxCuk8xaM7WUup0aZ0nNb
hLKSZw0QKNn9o9HyB4onHV3XNUjoH1jj9EFjphJ4Zl//hB6ACZ6VqKb70+tmiAF/
LOLbjdF28yd7vdvbI5LNSdysY9jtCaXUzeNMO7efnvUz93/X32dwWPjE4swfKX6V
x0RLrd1rzUoHcT6Y7XUj+qConflJC0KRwbpAC49WE8q4xetaTOvXoRdueEUpft1h
Hq5tIBvzVcD8I/tMDylSpQB5u8Eaib6U5k2EFWqyOcAb2NIrm1XJ2b8bnVnQslrk
EgVdtmmA+1B32SeGIo6z3uUi8RONNfyunXx5fEbo+pkoY/00TwCC6876pXIM/mfd
Z8wHha9OubBADvGEbJUbXXXhaA0zBRkJ9tQJvVAJ0D05DTts8HNnNtdfDbICcyyO
e9dfg2XpPXf6sUphEKdFLqMSTnvTzuOkLqtaTJ5oByc16vN/6QDRw0lAqAg21ZfU
qyaJhIqcMAApGvzhMjmVL76reAWh/vihT1KF0PK/WMc/Bh32VUmf+gDHNoA2Ib8B
otZI8A35Nb0/K9m7ra5RUtl4Gy2YmmqcVVJUEpyk/ZgPU1PgpkkOsRpVj+EjZNiy
6aqVJN+QDD0BkxaHKX2vfir+UM6zvgXIX8d7/b+gkc72/wzmgYSLTsXFhk0I87D0
b2mNWQN+OGayieerhNp72IbDLZC9Nvp1R+qJLuP6KG95NnNW90qIfG05mU3CdA1M
rK4wJ/YG9rs19GtSyghG8nSbD2o5NwOinJxZ2wPgreitQ+IlIPBosTtMsUTmvQt5
+/zGEfqjkj3OqNHS16XCX1oxUq5GWgP5ylXQH81ytJJ6Qw78I1wTtfO2DhuiDGkU
TM0z1aNs2UBJVLSyY+X0YCBi2e7PlInO2OCkQVks+aJSZTMApdyXf+vzHu80j8lt
7LjmVKji6Aquy7RNEXPObFIAYNez/dI9Z1VFlr8iBC/vnw5uvK/EUv+hj03ElKPN
c2+wXyuDQifD0n3VPrwVXsD6Fch0j7SpI27aKip6U0ls0NC2C4rcbYrksLNooQ0Y
F+ZliE8+563pxKQ3Yz6Igv+H/3vIN5SeDsHQa2TvzAELfifxuKROt7DCVCAnt3MQ
LWQ0OdWg6jCUXXq6Y8C/NJkueUS1NiurnsWVXUVs7+k0wDkYbjZXyxcvb/QIzKpF
QONpZx3MRsYePp4oXd2uoLp81vbSyIYWOWTOCBSSqISh0hAyXMZa8kFNsePEk5Cz
X0R3hj+VIoSgQ0LpivOe4d0KVX6ig0wTH8iMHendrKgYtLUwhHIJxZ8wU+wJGtgN
uvaPS4W3OqQWUgZtVvKeTCI6m/1apap7xPnXtvLg4GSzYD5Abq9Fnyrm3m0/rnR5
wlSPognjOmb5Wlhg+yW5wLlIdeWYOgTayrWsHdu9kIhozX55dY7ErajJ9XLx7QZ3
unzPIWHoAtafmkFIZObsxfX1OQk1EPqyW98AjBJKEsrE+UxDotTljF14Mu0ADxX/
dz69v50SknarCYAM5o6KRCECitLhp/glwaCzXbrcI2GrohyI4ZrlDJKCNjPUkUYL
zQJjjds/+TReJmUGZtxp8HQv+S87HklzJQ7V6L16Cpv4KP7tzt5zUuYbNb6+VHOd
Mts8+xUxSf1ESkV2H6jkgDXk5AfIM1T5NcI0tWPdtgV1b22WmP0arj9GQsbAbrF2
m5pP6GiIJXYoTnh3f8m1KoddEerlAnxhWqaUOJMu1lnjVW2G2+cCa4rkNKKmH0FF
htc/3WZASiMbFBmoKHPIXuTo3Qdp9abiNq/SVqgatPOjJFpit34BnYJKXedlZTgB
uM2OdN0b4wQebLDitd1RKFHdWbfyv+MYQIqWsEpKXQRwXXUZ9vMk0+aX/UCle6qU
OoDLzlMjsqCXTC8MBZ1e9AekPU41g3K8KasWWXV3bnwjuxwaVOLJfe3mlYb8e4J/
ITXzqQAuwF3c6qCF0C3T1DiAkgf7uwYQ6P2AbkuC/jkmzJDWCa8+/EXIzjTZ6sKt
bAWmWtuivBjwd17gyyRP67tHAkMYKny6sUBq0M/9Sgoek+I0oY+oRm0Ks42ur/5S
zY016L73IyuFMi7sLtvaJWs8f5LR4hFia/N2QbG6iZoSBG6rh04HS+GELnuEJiTN
lCLPhF14jSDzrLwHTK8VvfOCZWt/iZ2kGaZzp5sK0ZlLL6uTTX8UfeUKQ33INQek
KAkL6LDUXCgwhyJWYxYk1Y7bS0u2KBNpOdzIDcHjeuOhDx8u/UOL7kF3CE4aMXPd
L+PXyum3RqutzMIMGRzgtxIBxanf3Wks63JhN8kSC9zTlvyUTlVYzwiWHPcnycQn
7kphw6/q7TTi1NHJfMBR/Ywv3CEtAbxdWYpOnLFfQY4ha9xxB4VIm21cHi7mv5jK
pmkfOw7L6igLXNpic5ViYqJZwFVR3SeYVRnTk4ENmn2ztjyKx7/M25Vj+3iR9B63
t+71ym4YrQA6bpEbrMNbti8V2CoK7QfahqhrPkRBR+Ci87COhx2aofGxAEgziEAm
CRX/sXOAU3mdnNZb67Qh8d3bqPkl2GA7gctWFhaRPg57n9/73No9zhNH+UdwXket
s7MNJMScxFbeQUGX2K9TxbcNf/5gzzsA49rmngpczJeD1/b0KU4DXoxNJ4RNg9De
g7qfsje+zIZXt/TDgzctDE5NGvvno8Oib32pSQ16+VHv4wCH7XlHcyNSKPGOc7yg
B6kHT5p+Hj/kkiJVWVtq+g2zLSX2yWx082UapZsPk3g6zwLr17HBmJfwcQmffwx/
4PS8MJfc5SkV1UOrBBd7WqxvMkb3mFUMdceL1j7NRgE9iwKp4rc+sjLyP4JvRELn
mXu9+jrvlV62Refi3dgWVcxpQJTwfR3tuducxt0cHweCq7Qa99efQ3NSMXxmYgB9
8Ja30GN2QIEQN8VQpYxuFFgEJIlJTKP6AP/smSivx7SAzg0yt9o2+phRKZ0/NIzj
Bp9C/jigQ4F5XM3jGgnOHpxmcZRl1SvdmnzqAQsTYQ7zqj389ZGe4YrlqCeAUlwQ
v6SbUBH3wkNCiwpzK+B3QL1o8FcPnvQdQ8z/mbyfPScvfyqfIRYfydr9g3QTK06T
jXbcE7XWS7a6BTNqpQ2++sUPhdjX+4xPiIucV8dmj6xpZ3/SHsBBi9p90/z3SaoQ
LMF2SXJzsnojk3/5+q3Ta8PBKNuBHVNfWdbldO9JMjx2+JwyDRZoGJ76q0r3FKBy
6eDjxZybDxj3hS/dDZl5iiglGruHHUP4s7aUUN6N71TqfQV8cFypnQz6cvs+S3z1
vWtqic1GLzWs4i63F7hn61ce48D9cX/FN3K5LhPNN25LcRJFnJXymfEdY7qMVEZQ
Toa/jTZOO0nUXFwqOngMUIPo9T5hhX1JU5ssipA6JJkz0Zq+KrD0W3hcRaPb47Yd
MINnh4EOiZ7wtIRnKivJPMSNy1I2ukVx+x55REcbQhGt6QWnm+cS59mXCzRTbt/R
v8nZ06S07Num8XKSa1g0yvMqnFESIvdQ7AQN/kyla/8jzfqeT1PgyNGGNwNkp1yl
kpOl/m9q8DBPUd6JYG9rkbbP/L7GOkiDIJXraxOxO9AtGiFins9jk7dojGC4CzaI
t9jruhzI6efHpTgKyjRvKpQJj06dzFjzwPYujzjorVqmpQAaXoXssL03n0EQyQsK
dvSfr/DYl+uRRds+KCK2MyR2XmxxQd0AY//T/4fOwprO7APDghW0ew/DX+5EBuUe
5V3s3Ju8r8QPzKmXO9kn51+yHfepQcTadb2xrrhQxYgbswCI9jXOhSebuRyZFoP9
ZddMsogG67FAO/e1yuheQzvPkYwBEgp6J4WpjJudowdYdYU03Nokmkl8TSu8NOXa
puUng1XEkGYdGWGjrVXARVieT/XTzcreSHt3S2E7RDl3Jlvsu8EEeStIaRwsqzgY
IpqGRxldWpfJqbJ9ulH43xtvnR9y5Zjm/QTsyHTF+LMEFRMj/eDqwN6SJ5qtu0MQ
ci9AqKekz7BAJXFv7LFNjKr0DpTnqeCuhBLV18ihRnKOtIo7yp+zmNdvk6yd2Lfq
UiGPhVtMhzzTAVVOOGff0i2077LXgu6wENDPCb9Uhgc3c7o+dtOFhXAMWBJwdId7
1VKMuyDd/C7evwm2NtWMV7qMY8zKIY7hQu0KhUbMYJ8lTonvAhG9q246JRC6N4ge
lEeh6Wtbnc4uECDd0LvCxxXuRH1MJc78DHYm3sKl3A/xjQ2AJLtb8VGYfZjqVwiX
psRQuwBLEs+dZ6GqcJ2YoHG3BD/zVaquUHD8++Vi3V7ftq7QI1Om5fDReE+eGgvv
p45hYiAaskYcWXPWMJX90zL2qn5UCodVzY97FkspxG+PbPA3W/DE2bs0A5Rjity/
ImN2nX9c3LnGpMdmyLkFIPvf4ycS6bA0rym/J25unEiuqnWShqvQpyIkNFWmU3ea
6pSeP4iSFCXTN6xTK5UTPWCOkUT+4YmNYI/7VPMXeps1B0lhG+/vJMaDk64tZeww
idME34ZUJIiVBxHiL/KNB4GZgFq+0rhxU0+3brNNwiwyLy6dOYoUwGLUi2ztxjAF
BRZUQ+osDmhhT4Abf+3y1CL64ELgFnK0KBVlK3OY2x/s2DQxQMPAXN0imN+0Y8lB
fGMs1bubPZpQp1XuxA3SPFB+vr+tj3XB5dflzISlBcTDMyljAU93p38MrHWxRbRr
QmOkwsvnegnaTufeqUozTftwF6dGacW18nkHp/hyph9FAnucyS/ofI2nhU5XyhZU
649LyvhM7cgm3nkmYdsuPxG13Q0eGl9iJHFRQ6vefcqRgc88RNCcslWZh4WkIvWq
Ta4MYUhp8YT8krWxGXP8IGBkMYVDPsDfh9As7S5dj+RIQkOUWWQJH73ktm57atyq
B+YusPfd6Hrg4YeJ9tvqHT7TirfEjdlz3J/9fFiEKH6//IKEc/qkeEvjwAe01VPE
4RRlWjk87iHutGmqOw9jAEdr2CffIja0OZgSzuW737gWCQf0uEP46UVZZsfoGUSb
PYdNwf3VQgNf7Ea6SqCG5sy0t6283iIE54Vuhzw931Swt9HSV6YwnyuDhXdc3++5
xAouf4FDKI1gaMLzOdQS0UrVKSONvpZ30YJ3LLfYXGpf/J1bZEYvtNlxwe6wA4Q3
+sY31u+OBoGsQGUx9K+X8s5VlUNcl1sf1+ak1riXWnmT8rbmd0a7gaVDo6WIUkr7
55KqVJMGubRTQBJAnuRRNzADpLJferRzUhnKUx03MEWtoBgxcoiuPcGnuizW253K
WmTuJm3Dh/+J+Ld+MnIE4e5sxMqJ0Rl+oCfE06YLz7lQG8HWCfi9ZrJERbZthmt7
stVITa7Iz5HZf7u/4wnjkZF8mPoelkFHmyD5/OaVt/jC8j68+YgIrkXgEwrtXrUb
Hdz/5EUcOldJrZOaTOP66X0fgUWKZFBRUdUjRoxAffTWH55+46Ei+dwSiIVTR/eA
Fv1Ulp04/HUDGio30K72Rc8cmfSEVb1T53Uwh/BLqUxC6ItAPFLOfkDC4h6B9hIR
MX3uaON9gCDx4qq/QP/fe4Q3Z/NUBrfLHK5MF/CUqEHsww+690WtEzq2ZauO93Sd
xEj2oHDbpgoglY33SSykMxnkKkKTWZSht8wtz6HypoFbG6AfJ41/O1AQGHKSMu/s
qe1SpuvtKaf6vSReLdQh5iKhBhAThC17R3I8dIYRZFF8Auz60ZQMHVxiqKsKE58D
J0e3pfIFH9M+6GJg6VtoJqd1IxCeIp5L2tjcrUgq/bRwMa+dUFesscPo+py8TyN/
wizbIkIsa02PJzTWg6kUfdM2komQoEsC/S+9dSXLRWSj/X7tgk5qydQKmvlJ5dsH
nH2lKmTEJrDwSzeLDWOgmG0HxoNb1ExTB3JxwedhbvD71NeqVMz4ZrS+u54MY/sj
OltqlRozPcRI/DL7Gut/5J81WcJ8uc3cMhdiEF+QHA7rm04j+ZO8pNL344VjCABO
HINuMQKWEeKOn+h8Jmk0k6bMUXDbAlHKn/cbdPdmHImaM/1I0JpLMMNSdXMFJnOH
OCNby+evmE6zAKEmE27NnmNNzLs4Ow+gESOfQqUMBgbY4jhf+8NrYzsIPkCHm1Jy
0HhNIOq4Y4Lx3OeO3hI4NdQp8lMwKlKRXiObzANcAtZxSfnifhqJ2CDPk7cmmBAG
2MJN6NMYVw1xbhDCUQvRVfSaBAz3MH6KzQalyWX7TQ6lpCUfWKZvIxMvDhmMwd/A
TweNESz2q7VXs/GmaqwyJNBtt5kp3TVYnKlKObDTu3ZcEdij+0G3/3LBYRYACNCG
6IxQseVLHKpDbDz/zQaQLFHt6f3KNlXL+Nt+RLJaqCjOUQLjtefTaD9jkaz1wRbv
8340P6jdJYo7exAYrMFe8JsNvQxKtX33Cvc98pvDXJsbtxKculaGUMPpOUzs4Odg
vwyMqbzg+0y/AAzj+Wm5Ujz4LyW06cDhsnqtjZcs9Ufl/akLJzfdfCDAfyz8U2Q/
RwPX/tuavUn2xh3iAqcBg1YmfRZq+DkUdErbCIdZQJT+9zQDPen1sVlaSRaCSJRr
yM6dxU9o3c+D4b51ncm8zazXTH8OC2OeF1Few4tqmaTJv3m5VQb6TEJHnYlqZVzn
dppYNpwlREVu1xC/S+A98hmxRUzMfGKZtdQT/rfI8PNxnoCRgnu+L4tPRTDRy/lX
Rlulx9pLsdq4/iLM+O6WD1dq4nkirbQMVFTMennA1FcObtt85DnXTImFHx8LE1ST
7kcGpGrU29lS+jNFQRtIJBzYUt+/Rq0oSmHIvrfrxa0FcoGM/yMGvlOlo8lDJZlk
dD5bsxvgo1Xlf7R3BPvGumYHbv6SENUInrYgSN6Ql4S00tEN2ebI43fIqPgtEaKf
YDleH+LjybDwm+H9iIPaTynBr20ahvWikHeYG9NWsXekYKdJ7pSFHn9VGvxkcqEO
Qo5k3zQNID/QBVuo+v+uVt7EfZhQZy0ySAiUskSg/pSzLsVsF5W6G+ooo0PWX62m
iFE3DbTlUEGnkmXnxoSlCDAJ6cQ6zQCkc4lCfwhpk9NS7tVpCwZFMT6FgwV52+DH
7SOpLckr4fHRF/voywumAgFmPsHmaP/mNK4v8KqkM4LU5ltyHrWGTSYPkViIHvJX
pyPlbIshsZaJRH2hVzpcLkZfF1gDXeho/HIa95VO2Mm+MLueubqb4cTfiD3rCYXI
dhvxL6Bf/IjyskNQ9zpdkrlylSWvXg9WPF6MutK44YvGZmIFpmSmB9CcmhPZ8YoY
EEYyV0xYitWv/673Lz2veJUqQuB8ivMmr3uKYw9OgeVK/mfUvhfwaFOYmK5RRRIi
lEg+LYwS2wfBVPQRyF5iakwXAGEokUW7wyeL3DiGSfIvunoVMb0rZI4ZZc843lYY
0qjUbrvEh7723ZqXWR1prAjKk50WbstVe87drKg5+XfmFuRfPgppjJ7e3ZKJ9ymE
KDh/RO8NNBBizR/Wpq+jdRlHwRrkixtE3rSlthQmxfOg8ZM8wMll3GekgwM/waOk
FqcUCIWFBM9Pvnhe+CY6hwianoWmpTX6HO3v7XDngyB3HrfYuCKW7rhPNPCRsfzB
T7hc950EKGLknflutXepOX6ob9HtJV8PdlLyReuYyeW8NayXIRiXts0KIfoA2hqQ
OQTBAOcaSwtwgO760rPLVQ3+ex3ulV6c3yGgyOGKRJQ+QJb9BxLdMcDH3lLp0ec6
dOxNJD2+7gewgy8XDnL33oDgeo1XhfjSO6Y0ErRvWYayEGHD/tQpFqn7tIL3f1gx
UTV+VKry9isMtDFkLV/NAcrQZXbhyyAxmZcLUYFIGZJLxczWCGwRXH1IIY1jkTya
ff3mDi+UlY/oa5VB9+cW0sdqBgYC2jVsqz6Js37+i6iR7msxCFQJVujLqxEElqtn
iUIhrDqNX5KfSY+HwIYNNTQenbMbcyhL7rS+kkCC9K1ZDZ8gbhEucZNUifIChAVd
LT3TF6o6waocJEr1OqiSHnKR0YEbdnqIbIcsP5G6H9JYJr9ztFk80OoQLpbAXOzG
swa8mRkYhYjYUUGURhT4R7yv2A6PmgrNG+bViOJircPV831hHgZt6tQw40i8SGwz
hKywbyPywc0mLGY4TOB9AZHJbToWc6hDQkIO+/MreKAGpYVeSKb+4zYbMbkYVsun
Wbk6KbvVw0ICUASR4X0EqAKqBDolALyZFAhtqJtil62owtjE0Wz4lFcq3f5+nu0H
tVEJU+LrBMEjwTLML7qfAnEsSawNEBs7kR+D5mb1yG/7MGZeM4O7Ga2V0yueFDCA
cMZzXBKtEs2s6nrA5++ob2Upg0KqD/vDHGC/Ucw2bvWyeZva/GAGT2wcNpr/ig5p
bh7DIbEOfAZ5J1/uBIxzzugf9OhjttwNCoiP+GrdvvsO3fKnIEu5boa9GtxjfrfY
o+rG3gJAJm8Y0SaQXEqVjwvf+anpcCims4zWZ3kyza5gL5QH8KjLAlC2hix3nw7G
zQdGws4Q6HYWttCNn+Gj4XRa7wU4phi/H7dO5etv4i7o6s8XkRzoZGqWBrR8gtto
3vrJcNHy4us1j2nJiTE03rWrAlZY1zoIRZISATK16ayazEjSmZutyIRdSoETkraC
6g/cFuT7woxN/F7HTSQbziuLzcw/Yu1otrG6laBqonqMQKyc/nsdtqbeZt8M6w07
1ZUEIDjqgk05o5Yg7it60O8Pl3eK0/MHSMKQm8DWIy7kw1NzjlmoPhNKhspbIYel
AF6k6qFwYKJwrFw8WmXpuT2kkq3z91HvX5VUkODNEomfbVwN3/i8JQmiZZAPmhf2
HIMcR2gW0PX8w//UwPGWaF7sAwkGmooz3TVkw/CoBO0/GYFYYU+/gjhnpRKix4ls
FbgfANYAukX1KyPfU/TzUZoU2cRErTwql7RVvsU35g6FeFNLQW2eNwlcA0x2P+5M
wvlpDMSEouqLlzcbJLrS3jznabf0Z1fNiGS966dxQ9VQMNG80YqRvYTMhjiNi0FP
FFzpaQ8H/i8nu9QZBarxMtioWiBRV26Ww/zIcVzJ71kIxXALHjR2YfUWtOHKKUQV
/6RuCgWm04laabUid/+xWQ/PhRgczstqXIEYm/uUHLSRPEXiBg2udH2fpnsLgnVd
9MNda2VFNsaFwJWFKJN8l8P+ifvjIeAG00djBz6ekozuHRadGUV//v4cqeVDVnaY
S+LpmI+YJmve5ji4/NkNMNZOINAkhocP+nay9lKTL7lyt1EULGENQoK0cAvBkPEs
na4EMQdocKZTTpyP4u+QNrzDxgSq1lneFvw+GcTz0Lm13TBdTFmSUfyhjkkYP5rR
MHajsOpB5aY4YApnWOkL20EI2hg8aX2KfyadsnJxfzQrn1VZhbNRpb+gisGvS6uR
JCGFa9qxsOXOFHgxlei/Vt9hUZTj/+ABOth92DHNDB9PZSNGPzVmyZHVxNtfXgjE
BIDdsKV8KaFZOJCgUMJmgedT1JUKFtnuV0TwP4Wp4AmkY1trnqeUaxsAYncU3Szz
wF2e/GU7jyD4dKI6yAYDnC1ZGY5AKmVGpYs3ktAm60sPQHa1s4g5Ki+MrMMcPbIu
DLerHia8JUAHfw9VutjvBT1zdRNZ5rd1gfEVKp/lva1E7hOjV1j/DgoBLVI7LBMr
ObUxzojovWTEVcSouKo+rXA7fd+buc5V5G8EJek7+xx0KA7fqY/+jWMPCeeWFvLQ
YAqcBIqTtSjhPnNn1wCJWZ0aWmNYNs9CfxLhSyqlR8qQoQeGwgM6R687b/j5xBUZ
pHnW2hAyICGgO1E6TNXNkbzV0oqTma/AtXyfLCn9rwgESu4h3YqN36LDNsdkNEvq
1ZBXL7EWXgs7eUkuqpW4y6ujSjnXNVV+spFftJYe8SdJLn0U96pNef/8IrtvvuWY
6Ei9pBzBSnaFjyJYwKBXMTqjbU70y1rhTJE1IwrNbCHVke2XveEEQY7PzvjtAyWs
YHysdQsjFPQLKdVNehXzfa5IIzZHrdZUqKFB8qwhY648YBX0M6/rtSswCS3WYzQG
tWNMOlx/pNPA8KcPQCKdWK6ShrPGuK9ghAhUq89zUdTg5VuLnIKhcDOC+11kMQ0m
2XZO32AD3mYbptDXyjc1UBfOid7dtuGCtDjYnPy5j871UmlsSNJm2hL0TvdaLc/h
wEckoT8kpxlx0PHyfa9QeiCcnThlcBRg8fWFLpwUmafNuLYH1e7EmoNVMrNYPAFD
AviGUISJgoI4UmQ07j/VhcMRWE1b81naJjcEm8lXs0GEW2/uDYs9GVJjXGecIVp8
p4y/nCxIB/x8VVvzKPDg01uWusSofCMXFi2UWIc7oGuCgr3vA9DfiIA6geRUeNs3
s+ArSBE+MXPXKZAT4vPHKgdGn8ChUX4Y2ELaGiv5hmty6pYz7IzNKSF9Qrv+OAyu
3vN+24ChK+fQ04rCdTj4e/mNhckBAK7MvUYnC3WyVXGk1y2wQ+v11PP/INxQZRob
PxrJFPgrqvwp8kGu/OlOUZSqPIHBoblP7va5B+i91EnFT9ivs38B10ObNulKyUbG
ZPUkkNdp59qSJFK+wzSQj2a/9fo3vzapgap8vrhMrF5wL+mvJJ9DToU3hJUY94Vw
thnclfYc2itfT5wXXGogFrHZRbh2DnSusXsROQOF9MrylG5mECzRQQC58QkG9TtY
CRD13wqUAfVPu17QbXKICCyXVNx9QS3ibt51K0LRNZmrJVme4QjvDcX3H7utzOG9
3pV7NXK/Yv/gErUtKOBsE2QFoLuHxJe6vmvj8trAmQhQOd5NQkZotwIrQ+0PTfrS
+rvGRMTShjZ8EoBVl2crsQ5WBalzVpVXezrX62EDBRx8AvwhXz+N9YQa8PGJMnGd
nU7SLxyiXEw1WiDTJnV0+ih+bh9soq39U6RFkjlc8zxsoXsI0pDS46TobT7qIvG5
oVIMAEWxNl75Zxxpe6BK/JDQRXhlw4VQl9FFQSLD5ZH3xKB5AC7UkBcip0GDAXOg
w79TNBF+ddgLpRVnbmlWyXVUNdoA91wwRYHamM0VLL/EYiI82kbNAD1Sc1kQDGQM
8EhxP6w11+BAaoJMatnDJlzJWi87ZVIAyQxaJrUrrPJdWDkptisDigdeE/XlAgIA
eVJ2QbeT5/0uxy2whtMk+YbdYpaQLQfcsFRvoIjo5I+LwjLa6pUBABaEoob2U/Ub
PBYlLKxMlJtx0DGoZ2gMmG5R+R55Zjj10nJHgZdbuzJZPBEZ0Bi7tNdN8GdYvi6K
cQMjFvOcPDFfvt5hqVBn+oEF/Yz+8rjlvmp/OLauMokP8qdPwv4SHnCDUYo+hff/
6q+v5l3gZ9wsuJV1Myjz0i2bCjDsltMi+PY9oXMPJxE9jSmpLZFBlDWVekZIywLE
6JJDDUnKw8oVuL5I+8ncHc09Jjq5YS6Ux2wMuJkP699T3sdHc4byOcwqZryZxChO
VaSvzITZqFlWKaipHmiSVOOMMZdNE/rRNKbkfLhDutgokG7jk9/rMsSG9b7b4s39
ZpAXo4+owAfnk4c+ozQInFFOZ2XM9A7P9eC1ZissL6rpsDupyXwrwJg//zVpVFH/
6lradyXg/0T6wF/y4ad+p/srH2M/S56P4RgvYhlpZtssxkJzp49Rglev2MMa+aFG
fh/hQcGC8u47pZm2O7XspwGxp4VBvwP577qflWk5mp8tssj8LTkLExtVHkHZoALt
J5e/1YSPzHTS28Z/4uAs3EyX5mi5Bhy3Jh0ntXyZuZkmk5lTT31hfAeVxlLo3RWg
q9fGkLk3PVx3Z8FdrB5I5yMQPJws3rHZ0RD+4Ti8xuoPlmDp4XPJxAR5uFokLXb1
3KTLoZAJBBQE0DGzCgUfE6jRNnMxFLshJvaOIDOfs0CW4nk4dcDrWQE/aW0cQsEq
hSQlwEVFWqShfcm8wpN23wKG80VbXIxDQtjYzXUsTbWMbdfVq02b388mkhAmEQy0
F1rfgJbfpDwCicOnHa9pelnyDnH8fqjcv46ljnSTRmgOD3Svbi5r5LNbhPPbxrNz
tZ9RZsdvarnCS41ouoGTqVxy0i5GLOSErWLmzF0Ml9OH2hiyuAat/J0ZSQk3UC//
nQUq3Ir8gHSY+Hq4xPZE/WlR3wRZ6z5wDxL5DXUdQwzw/yJIhoS4UP3x8T6fTIUH
xbYMrc7OUO+2swXjw9fPEbcpn87EJ3GHMZzyA6gYofZhkXyQks2fzQg7j3hIZ40S
vrxhr4C69sN87l1dDakr46R9PQvmhsfDtf32Vj7rkgIsaTKslvCB4NqGnj6MYZ6a
AellPZS+ueMmH0PwmbMx+uQngVx2cpaq2HCoFKr0E0JZr6Xy6T4cOr6X68ewBmG6
8gNehzGzyrJgTv2J2eaTesMFsYFfhFNE8pMCNIpYx5Sc1gOBusSPIsBgeTnI4+jw
nO7YuaIzX/0D2CE5JmQsYmmqZy5wb3UkSBWS357sbtebDQDaHcWGruxQPV24FHdw
klcJzokJrgN+3C5I88n8SBj8iVv7O5MnwK/PJQp7SuxdVabHSRFtIYRwR/5HcgXM
9aK6vQmX2Sqds1snHu8kGutoXnLvwKs+S4tnQ1gEzZIFPFK/o36xsyICs0JpSbrl
yqzN733IRaai0mTN7N5H0JRxRb3yckOLaC2S2QdDL/6vARp0KtRBflCnS7MZFOWT
6gsqjXfsPhTolqX44VMz28N+E4SrR883v/8bjmIslV5XumX9SU/RpCFivLOali2D
e1kUvntNxz5St72NN05m+7IgSeUxwbIt26z3FXe1tLlTmOzBBSx0ts4tAeV9RU4F
PqxtljGBZ6DyhMRLcoRcsPEDrabGoogyuVY2qQciMRkm/5p9Hg/O9rnaLvhVkahv
AT6FiKo+ts+IvIiZ1eU8tCb8sVacLALcJw9sRci3PVyNeUDBKBWT51H7jUsnHrLm
LTAS3Q6Mlr0lTxiRyhh76AbHVcN/IC8LR/yxSpjCHnIzJycHAjFi8PPf45tjuHII
S3BLYcexgh6xSUDzKEWgn5fgaApR9G0MOGZ23SSmA4BoMv+2wMKyRJ87yodBqrUg
aTUhn5YxZEicNFIBgop0Cx2jACF6jG4KkE5a7P5nBEghBgdoXubvMSyt6Ep/5Dms
gwVejIUJ+PEtE7kDnAH257s5bUF1KE+cVScdkvRzO5r16YW4A5KJZHSvrGB4fRbK
yyQQg7y9K1qSVETYitGkPWZWHOBdxXTssWs+8fMZBq0hUsqxEr8J0CIw/vRo/NOX
0WfkpV93sJ1e2mgjqtdfvANSeLtH1x3eLUZNTO6wpg1xEo6MwXhEPXHwpiXG0WJx
yQdXlYR1YymqaKtX3qX4hh4U+K6zUdO4FhTxI/umipXn6pPK3FdObMr4bOeS0CfV
HGXvXvbTkTHAdeEECOqFkyzAPW1bB1tF9pBoGluLXp+bwlcUflYsddJisrxKj0MY
v9U2shUUito87sITjD/NkiApSkJ04ajw6DPdzdoVxvz6DT9zK2DuFKIribwxY5P/
ShhIIPyE9F1gjpWY+BRlaQlvM31ezjytnm/fK2JphuUkVzsjFssY7VQXKs5I/lYP
Pko6YSW2Aji+FqbnroTk2PZ3TSi9XfA51Z/tZfBhMKrnIau9VS/O2q6vqOtFHW3w
tGk3XFlzKAVlYL7ggLrnJCg5kwMXCbLZMK1f6bBSI/QoZB/0bJ1hLVS021knDbVu
u28nPHD2y6of+br4rwJB94sYmKbfMm5xMlDkMTQN5a7VPeQrPzEPlslLe3tMtSFF
IYw/8KOD8cpe1cz4VRa3NiVdAVYFyGW5MVvO0tVkl3W0tK7piTaEma/9wPhGPnaZ
qlpMWwRZ7eTyDn+Kg6EpolqC0Ri+Zglr358JQQ4iTIcmuJ3fwjt6MZLehfnAV4kj
N3P7krLMcOIi4qiPEK400edDO2NDsHdq65uZYC6N0E8bbCE1BRhNq1QrV1NDvart
TVRyEEIbW6NlCVZawRNpTaXJyMslNzU9K1w6G/k8W9C4P6YWVVN8IhdBueym1LJ0
gxywX1aiUcopYwDIkiMBBG8wCOlbeeHpPXLDVKhMF4XdgFEcANoyVDDx0BafdyJ1
4NPz0QIcqZZqAWHpmLTkl8E09LKMsn4Ew6EbyNlp2dsZPfamoiKz4Pk5dHl6Cnky
SKr0pWXMBFf3bWmbfF3q4oOCkOGMQjRux0JqRl+fmV2WESuIEts2zOT0E2kx1xB6
HrqiqoaSFYLchoD0pCWsaXl0r9fEgdgJwc+kOlHnp687UbSbtpYaCV1Hdn3XJTaN
o49Zu/TvSqpZL0Xi2PY/CUnU/ZVadABpqc5EwNGq4xH9+T6mEqh5ZP/oWrpaQZ2B
bkZROmutfaRc2/zAyztkXCrwVrcSU2ncTZ8aE/Vd1Kgbm47qH/SprXO/7YYamwt2
YzBkym7j56+1F+fwjwshem0mUYvrLW6rJAdZROeIRlLTN4DKe8sPM870CYO0+ZNj
IKuHrX2wAj4HpTAqAn9JvhNaooB924gEpPEOS15yJHbdaMzy6DejDSg+EMAN0yUd
xQty8JoQMFdOIhISYlpRTDfcA00UyWJKPGN6UvMlLscP+gPYUoS2791LCIW7hvWp
GFtpI44T9TWA18OeZHTa1XW6rrA/1Nq0Bz4spU7jr+4BhbxqjDOVArhW/ryB9XR9
j4+fDCZrwzdMycKmaSedCLf6b8quR0inGHiWZpzPXoylEEeytyu0XsqGgUr1RKkJ
KVjz4WUWe4lDfCPn8z+o1fdAQk/ZNXxmXhK2cBOfY9jolyrFGt1aflLmfQ6BiPxx
xbaWXwzAj20P/uJMaCBhMPAkyaXgDQlbze9nyVf4J/v6gWRbhNh58Iwgv9l4QQFB
5698ATJlKhhXGMYdglfWDHcgTbcJsEx6/7AeKYAiNDpjxIN8b7IJLQLrngmLFTfC
ekJofVJ4PjZH0tSDMCJuhYxHCQjIrOFWKRU9iSP6o6hDKCE2zZMmkvKCwNKZ4zo3
EgDMvfTYA+ZacxPhU2wvBT40mhqRIL17Qah258Jrl2cTaXaD7sNtbtt+xPlrwuka
20jnlbpSOI3XifzagFa5j5G5fB2Uv4IEnViUSlkW+r2M1+HFtXq2v4fPYEvOfMMY
3wJKl1BQ/iffsM6tDztIfF6o6XHpA0z1aw9N65yRj8oFGaebU7ktdw83A8pumeeq
jC+PYxe6Kc4PqQDgSA2rjheChhNGfypMIqSfBWkwgV2ZiUJwR1KZGSw7c9zG405y
+5cjXmuSimOEwmpS9r6ggK1MwX+6FoYbzaaYOVfRH7/PICGUbTMD3pOx2D9QwNL8
JkRyVGGEthKjg+nahkCGHw==
`protect END_PROTECTED
