`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2nFneuzX4B1JjZyX+pTLiv5lq/MR2vXHsGlVtJV3599A5i1NPU+6+5hE1ubPFkX
HoGbo07ASaBDJihE/aKsOQOPhAObmLmV7zEye9RxYNcJ+gQF4TahipQMbqtan079
W0i4aOk63KjulfjTPlxa6nPyPt1wUEg1PGzviV0of8F5J3+56bt8d5ddL4Y5YAgO
qirqWFhon1g2i+7WaRcpuN8mZokGDXyEjmet27jSqJu310vj0L3zAksal3G4Emgu
LFzQUmQ8Eq/1dy2k4euOwF7V19x/QZMzk3gx4PDL0GKtvY4ICvVqJCXYEcJjfmYq
GL5/8+NEfNsDabtRNd6V6LCN2XlfyR29MnVdUJgpesKLXMAu4Ucser5cwAij+D7W
CZ8MT/G8q59RnZ7wPF1kdMMkJYUM+SxvDwrXu8bbotir6hERlVB7dUdtpklu2JRd
e0qRgxOiEukUd1a3SnF2+CAY9Z/dvCLSDtuKPwaVItIGKChBrStRSv2tHgi1uc3n
jbT4Kv1K5x2dwkqPm8Lt2L/8qfTdlZ9GcXTF9v0/C4Zu4pARsOg3uDlkBS6ZOK+K
sCN4oSf7H3AM6gLEJ23Qmc/ni7tzWoP7diJ7j3VHws4Zt4676CY3dGm1oLiYbTBY
LuN98Wl6h5ycWef73NouK2AYDDc0XHloqi2yJ8/gRxWOO/VGt/GTMWsLq+s/Wf3Q
11nmY7J9m6FyFqTl9Fha99r+PqW9rZycrIg8aU3gvjva9XTA0XpNia8lMsfchDv0
f2o7TxKed/E+qISesKyaL/bUGB0Z+lnDCu5ycPEem/SmFL0TPU36Aj3f/p9o35T0
tiDnRTa6atTsUeVpW1YfQ5jWzmSxZEX5ie8EMF7QNc9lBEFB/15G6rZX5EqUgec8
qK2ZGEYjzpw/k7m7FOOE81AQK3q7bPxD1jAxaws5MgCpuXyC7stlU1rkDbP2hap1
4uGGqUy0q/90lJw0fOsTDbrwo4lCeofT6B1X7itR9DWniivqLfTiqzD3+6pejhI2
kJ4aHne9kcIzidQx53FgKcvKQ48ohI6Kiog6rMkvzb3ZD9C5Hqw1S9aLd3Ij2+PA
DB0nHq5we5WQgV/dd4p9dPl85uAIJ8pFMBeoI0GELddHyfBveN3GM175SXpk04Cv
K9/+P0bDJQOLaPMt9WbuZwsOoZEp/ztDzYgQEujpG77pCots1xYpoUrbbCfOzi9E
FLaX7+yEUmDYChOu/iPRE8BvgQN7VRLcGKjhZMSnv1279b87tR9DW0ul7kkGEXZs
ut0emowFv7BsXhy0fk73GaCvJlnruT1Z7BClquuz5zzQMDu1koCLpNfkfYdrIcT0
aN9Jl1JgRrpr2lt3gEsjvfiqSZnYtW9Nhx1lblDm7RAaTyQii5QtO0SMdjyKwRs0
STRtSZe0/egfl/snwaOdd2IU5B9IuPbEFFQ4cLOrPIuJquy0ZmeRQWBuZEY8KzA3
C/gBl56ulIZKdYWYimF8EZ5f0KRS6H6d9w40PPfFZt6X/k5x+sH5R6Pihx3qMPWP
GZNN2Z05we7MB5zH2Uwhqno3Cd7TTL5924wJfbMfXpEFK8KJApANi+/6UG+XcNwc
oyY5psXp/qgA7z++FCpm16W+k7WJDfNpIbDs+6o9XPW15zSdlGO530C/FLgnqZIR
DvQbmvmpdEyGr4DS1+DVXlul2GOxquKyu/PZWcRP3zn036rbRFuz2ZR1tEzenPE0
Q8Ziy3WiqElfS6nb8bxTbXDg9hifBDJsoY6s7MEw3mjOB8XVaP4WaPZnMFndsIqA
isZzA9suZlgM6E40xi79xjHqNZLJwwTrLrk78SLXj0CsLSwQlnrLOa8Bsp3bUos4
pcNoEc3y1f8cI5JM4w/EpLPHveMy32m+oEly37dSs+6/N8DFIXaI1dCXNxI1iVVi
jPaaI/NCr9KdHoB/42FMtAdA1aWFy34SY5Yfuj870AT2nGWnGWxdvVvwMa1aTH/T
mxshWk2Fk8Pkl85syEU7P3B+gVietFLF0MdegHveiGyuR+b7LEZYKy5eQ0nghGbe
LD/jf+Fos3oM8GVQddFPTyrwBTw41xdEuWX64SqzqO++Ur+xrIgGQNhuwqcqbeM3
THj9o6EOBB3bbRqdYtAE3s5d/tq7uEZuZbZ92sBJb+RrYkPayXGCqotORWWkyuWq
RqYe3av6senlbqAgCuUk/lCbC8QtPVptvrDdDECqYF810tGqvIG8W4kgXxI1dBlr
v0ao3iEvYqlja61rJHl9o+xIEWi8KugbWGGRKUMwqTAyxgRABQu7aJi8cER1B/EN
nqOIfiswxg3ltfKkzH/Ofycf4r28nmJpLxBmzgybVpQpm53ipCemj4Ek4YZOuLVR
1I3LEMoc52TuXtYcthdeQYvN6QY5MDkShZ6hobxnBRkpK65vizkHqGXzf66KDFEH
1wgHa86N9xUvxQBMzMU/N3VdzNgapl5Z3AfZXDl+ENnqlPPgo//BacFuOn5AG0QZ
XiNpMBKVSdP2PyCEYGyXB4jmtTwEvS9jxmKpko5VmXd6Aqn4lDtq7J2zAz8Kii0D
TqMi2jmuQgimdisyb/Ix6rCfM7eERwKUWsS3H/7zkLMjd4dUSMNDFNeVVxNR/3Jh
5tjRBlbZ9quwyVef8IJgZjOiTZ8ADEwRJOftd8dHOI/ZWYZUZ85W5t6ZranCIqHp
AFdcMYLvEgZY1syR/Dm79Bpaiy8Um+EEHUE0xBihjqckNtuf58wxJfrhLvzP90Vi
MPQlFI8HbRZ8cZ46Zku0mGmDEv/GxvNpF2tPv9h8N6zaJ8N0SgUVCY+E9l74YY3N
WqhgfcqOaAMBcY5St/uGPi49vM4DC7egCbL7uoZKYNvXErV10Vk0AvnPOq9SJj8b
7ilNjAiU10XfDavG6UdZ4OTV7J+pF8GKHSVrytajuEI0pel5yW8hGMxcCVNCmqIQ
Gqtanm3vIC9uKPbLYiKKby7re4GffeUlhTgYzW3uL9LyPPVHae8gkvr36g/4jrfu
ce1N1LEzWwajmkVbta2dFzMZHMNBauqE7ilk9ftxfGqM/S70VBKB8sSNKHIEr2EQ
5odks74KKGzNGVBcRZSwW6ZlqWUPDirmu+IT1h4yotqN4cjgXTT/txzlFnFvS++P
CReHsiM74fPKU0rLO0q2KHErHGn3LKXn0wh54JN+qHcwFOx519uffxNNabd3NOvT
ZzXHOTOnjzmxiLCven8W2/qR1Qf9uqf9wItPwiWREZxzfJc/X9OAgZODFpIxBlEE
E3f4DjWPbG2Pi/C2PrvPSWqYxSFr/BIQj8NJcgTZBG3JCUHDK80tVFbm2Th00b5D
4hIPENPkyxYSsxfokaz8EmneOaAQoOfgTnnd0Cy/1WnESTJzJP6ZZVKTD2yakrsE
A30255w9vaUYKgH4rSw+5cKIYW7VQG1NMDRAtnGQyyDlS6BfhznOeJAdFEAc+vHd
TQA99Rzs+EblpXOPdoCvX/un5AQk7U6s+lZRTa0xzsY8MwOOiYcHRoSp4J9EKxKz
JAxA71AKAJktHp4gi8rWlFI4i2V0ZmobxdjLiNzFeqB2oNuaMe42+Jq8jUnpJh5w
hdWRX9qu9YbSd0YRbvYg0sUeKgUnQ2khscje66gHB6SxxEFEjsfiU0WMkicc7QGO
sJa6MpI0S67XyKXvXq6KOeZPFnx+CHWwFNxYxwcc1MfvSpphGbzcvqNSOzU7S97y
sYpDm0eWh/NpdVLSFzMbckrKyFXBE/ETflu6ojuLX0XFwRXIgENrDgpj1z5ze6+Q
2fDH+x0AfoIl3ErWdk/yuWDcNXzPxYHDWgoCHhbXbEgn9e8yCWM9pxlX6jYDlv5V
4m9puiflKPzBhTA81FXr+7qnK8ZH0hxLQy0g8wVg6c8lMcu7+T7X9MmH1xrNYy7J
18answCDZ3J04YWxtY0vD+lyhpUlQ/TdcDj6G3URoybVjZmTccavh02tt6vGT40Z
hY9GFjJD1TJjiPo7oZ6zYi+Z0TjqxMh//zs7OH7KsrxTmfZyC8mKqtCq4qjfb3BY
LKagPJduITQCPeiJGCb5UlEMgSsyCO5f0P/q3cUSDgDjkJlvqeU0BLWFBXExzrE9
KkHrnJkx7G/YmV9u+5siFjWzF9a0pisSJDFB1EmcKNaJRNQzJgGUfx3d90nLkZDE
wGvClUCI3HqzKeD7Z5u8w3R1DD7SyctZEdufbbuwosGI2JTrSaFEFqUXE1hyghk9
fIRLTQd4Xi9jviOyChwm+oyk9IzmTXNtzetYsKWifYSFXvRjFPgIgQoA4oe7L6f1
THr/9U90LBJBQqcT5D6TTH4G7+eve/Zhm746T6RuHEVzo97bpmoR28WZ4kjMmA99
6I3KyFTEAYTpXqdA0wowu1DjwpBdkpFoWl9xvDowAd4Jdti0KxxDyMuft6oMKWCb
eHdn5sQosDCihR0O6ucrouuuI3o/vFvugJuZ7dsN6L9p+g2ZuY3V2WFFs249kgTE
Jo3bHCS8ka0M7IvK8mXvSt8OZV6WMXBeP8Fa/xqrdD/z9ycnuuEBVjESVcq3Gm50
fCidQMc9Kxznuf6ncKtxEUNW57zn5pkmFT/WCslbxbfz0d1mvs509jz+N2j55N0b
amc2E1Fa4hViO4IE2y2xbv2ky2DBUMLlHdmk5il21eCsFV5R9rGlVyR9Hsrplfbx
P6Wg9CkNJ6yIC/SXi0zAztqpIGknOdgWHzT7wVRJZZlxOgPBCqnK7riZhoxpgPqD
aDeM3Gf7762x9urYnEh5DIe/V+d29p9M9+AfGflihkaXSqggZV+1JYd08eCbUo2v
S8u+0m8mzXU8l0vSU4NLtP2G2+ZHj2HOyaZO0gmGeNFbSwDzCsusEUcNN5rve9yF
bflZ2r+7+WIG0PZq5xJG698LSBgbPIVUseQoM9tQmeq+5wDk9VPUQAcHl3tAJCpj
6vAj2L0O5eVdFpF8BN2sPdYBmNz6VKb0hw4Xw+2UbJvxiD6wK9YqGOEVEKCd1wGj
KDyg82odUAcSpD2myEAMYALvwZqbXR9Xoe7lJlFXzB//7Ao/oreHtF/J/o7WbH4J
wPOQMAyn1Imrb0n2AjWjz1iGpSeazToMguweI8roQHE=
`protect END_PROTECTED
