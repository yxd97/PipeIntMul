`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cJ/vNMlYmvJLJ7x/slNpJgau5fvW/vcztBnKuZUTSyg2qG3M6EEQmEduQzXpm+9
I6G0r1vFBW5hkn+J938WTxMPQEvuppHVvyvmFv7AzVwPKHOHjuj0mzZ902Jp49l1
QN4MKQiAa4e02REXZJrkPgQcau2NeGnziCqdplFnW/oPwH7kQRvaXqBSyOUPXLMe
6GLNUXfFuHhDukpf+m7I/jibJTMR8nKJwEaG59pR0pkS3QrDiQowMCKsJgzfVbQY
PhV0EwhKDA33lDFxS6JkXnVeejsgeXGiF7vUH4AGb+CnLWox/EqvSBEFfm2z62Pg
MvYujlBnISDij3FlnA1M84+B2fHmqffU5mfSWRs195P8kgjoMljV4yauw/F/4TEl
irr/9qUSfd/3A4NB/vkwiUr9PQeSMGcZSu2AVrYu7n63id25tew1R2pGzADmK8vf
E5Xx5oElJC4iW5xCKQHoIejKnC9MozMUgXCZ0mTXChHSog+4V0uJ5VDHtUrLm3DU
`protect END_PROTECTED
