`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RiNhsHwyTz3KIf3cGWBVsT8Kn0QxU4pxGuH73zFv+9CDrMSzo0HGAePi5M0QAcWs
Q1DDDlFmG80JOoXx+Sxu+dRXFX9HG5kLh+/SHoXenYuKPQLRnORw+CQUTVcg/U9S
ogd0WVF3JnfiEdI7mCT0Y9E/BbFhI+uhyJEXNhnqEXKd1dChWs60DAWMvDP+mg3R
CZMSwxyFJIy/abuisuLpArQZAYL1p2kTvzlfZkIkBA+XqVYJkPaH5iinBrxQmn8d
Iez66tCFMSBu1yP+1Af/n+8KTUAv0w0wGEOetUb4V/Jd2awXIkLdVZ00Z2LXm+B5
YB4LBpqT2xUkYyvJ07pdURZsXRdrU46k8PigtJceV9qFcv2dLjzKL7i+WjL8Hvaz
ClZw1grITUvAaBQ7TAf4Ir+KEuiFEbfSeYrRW9/0jGamB5okAfr3UaUCUzia0L61
tMMEhtCyNgH4D6w0SM0Behl9VotNyTkEsTYCCcEQSRGohmb4LRER2L/aqR8fd78V
`protect END_PROTECTED
