`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RA+apSS3TxHmy/vwtG4LOArBMurVhAseB3VfHsVB8ev5QvnkLPNAgOZOUvKS9FEJ
niZFxGP8ijHksY0/ghcTImse5ZhbsaHyED7eXze0Ft8bU01bpt5vBKRzG6AHeFN2
6SsD1cRcirkXpcsOo6U1blBEfXDUddIvdiVZo8JmxMNlXHEZqqRCK0FfSqQsATrY
8hzDbql9/e18iCyIt/N1dNeIc+rcy058aTWjkghWhQRNU1rs2EPXLth/b+02Pv76
xYDHyCqj8DF5L5m4dvbbidK54iVJO9tiE8KeId08ZrA7VJpKl6ZvvXKIznmkhhGV
V8w6U64miTm4Al1pHEiDpNOVmeA0vV1vV23JNiOSxleED42Rv8yh41SGvKpBUcUj
hepPYDrZQqazhWcz/VfdF4TikXQ6kpDcPV4yAQ/xieUEnu3ZhVXtdJo2I8OrvlVG
VA8h26x/52TRHneV1srkCys9g6wHc7HM9eQypgvT+nVg+ixZ3vUr6UC93hMgxziO
rMIxp1yNi7WMSCAF4DkFQi1TAMbIWVasVRmeF0xv/v52wFdt5wQNSPYNUy9LCSba
PQTF2SYAF2bPpAm4CGEH9ybCX3IczFownlYPCPiIMEXah7h+8Yi4y72+3x1bkwtr
iseEnYp2xkRe1ZyZvBjVhCFAqrLvVzPmdI4AVqn1V0vgl00b91HF8D1QWaHZ2wpJ
KkJhTpZPe31z/TQaWQQJK8c9sw1IS0GgWCGcMfUOiYnGlHfXuB5/1ZT7956eY0Hb
1Po6jcW8ZiS46IFGa5BohZ63zvRUTCWu8Qdhz9EkUlKJff2DmjYAz1ZNjdv9QOtB
D4pDyuYy921afnITqv+kkVQZkuXBjV3cRbMnpI9CoAaKlAhC4dxxaVQ2JsA8xyJQ
kcvACh+AvRYPkHuibIz4HmV6ZxFGWoJEV4T38R0+svfywHo9JyckotuJ9SfDGVoy
2W/NSYpiIo0zKInA0IgmfLohSZnWbmwpjCJdiOe8OruvaQBRCe2KyVW4m872BGmo
gVzuRMk/EBdiA7bkJ+1d8+tWKSsja3jdhq+LLOcj0P0g6BROlHDqC9sxH9jT6S5r
qMmxuZV+1lQdwA4qCG1xzs+nDYSoMwVT4/fLotIZmZvbH6V4i6unZ4kupegeGqhk
PmLklKT7AtHLO9SUPRxYo7mkgamUej+VBb4F8pixcLhLfSwIxMiu8deBBrdWyRpm
u3ihmPYdYULk+Ue7pSS7oGROp0ZiWM/+YRh8scsU9IZsKKzMmp5UhYTjs/vvUkic
zI5VYk1FWnUknB8/zSDfSiImSmJqv/B7IaHpUllaG9j51YXouuT8rK1rOSXw4wB/
NR9RDV/AkA1xxr/8Aj+tR6lO+g3IlFho9u33oaboDUy4goqVvLcf4j5wh03S4vHd
pFZGmER+z/09PzrDSs03yffOmzaI2fNF6HiNc9qZFCc9VCvCXd71ISuxySvpQcne
wEYJejVk2m3UwqxpeWYbPZPYTLkDL4SBASGGP+bqQEEzK8kkT8mKN1+JaJbviJUV
Hn3DH75OOnZKZYyMlkR02Cptau/qP+/++YAv44qbqGoSooiE0hXrgmL5bKDvYkVo
LfqzKbXZxEwmFdHZAbMlVzXn/IvPJPy4L8dqqFw80tjIThD+qLsEH5lKNkx6NNfT
F4sSlY3SsVeb+HEEx8YggPhaK12e7Tcj4LSmEUcTkEYyBN4huLpvcrNsAq1+rOr6
+lwTv/vtBbr4nhG4SNr43kUyJ6kQyrDanjIy9aDafSFIcPU8NTPLqDiTumjLi3HJ
XY0yIa7skBKnHHs5VECuOW7wyPJJPhi9mgrXSu0yhK7BKeEi1Y5WcMgQ/Jc1Z1lH
zi2fm9KGF5HnzLgw+aIIu30Gx/JTQl85PrXvCaL7o4epSEeauqKt14KPcuewZkvi
BFH/Bdhw7MJMME3p/NL6JAijVafQrKG+xI53ikGDeYuUdbo79wiHjrGNGe1bpir/
JmLvu6JX4nL+E16zfRouXH/al+Bkj9gbqYeVsqiBfr1ykdJXjETT3Lz7f+FcLWpN
4LE5OFIiLjpJGVFa7vMe6vfCRxC9Lt3ZCM+dfOsUIGf2J/KsDaAPWdHiKo0ZEfYK
nxCgyX1UpN1igd8ah6feZWbiDDmElSABUKdNCEDIMlyDZNbIOcp1PFqQDLaOwMwd
ZJBjMKdgN/papjU/ysq19XS2bmQl8W1Zkz+E+U23FlTn7INvBOgwW4IJTPajw1A3
/qRAQfky7sA4W6JeDynDEXjcpmPxpAHDVX2vhj617MOJyAqVoorX58ajIJ/yO5/x
vIHULA++xVzFu8Ch6PirM0XakhhZzLsMD6V7OwQU5IiH32KIyCNnAlN76oNbEd+/
fhSm5hewqyXaoB/JRrRqFCKm45VHuUhzNbJxbQAt9laVCgcOIjWu1HyyLbj+j/Xm
MCB7jxTf2zc81VlCggHn5iakeO69KM9nm4VcGbSL74tq2ULLqQFD5NJpg71H0TIf
Jf516coYD3UMSHmbdEe0HhJSA4rPRlBFQzYTxlG95rrDfI+w9Nr3xPVF6dwc+Hxu
y93PTQ9b2ODh6MXmXyjbc7o/K5BXpFLtiDnf/626wZ77lLtWald5OEOu8+0pDhyc
qIlBtzpFxv92D8MRkrYNOtuxN+1MpMui3rnVaPVgfBmLtRLmzWkcpni8UKL7bf5R
/T6JVwjCsltln+4eVuy+1ydOqE+uZJfM2txuUND6WHio9fujE3dHtsQ/s3Ach+pe
QSMEqEn/kC/gnB0Q30qYhU/QCi5IelxQwBeZICrWhomCpYHQaT37+q88PBIsRuC/
k5PwvFpkIHBUXkjnC8WrjgAKlaQfJfqq8+TQVEwrnCGZaSIjGESuAppiKWqgtLqT
1l4Iywg6wtOo2+Lv98i2yZclVh56mzSuvnymaOV9jhUdVE2gD8h+klFWPmOGEVq7
ZKTnSDNgAFRzT0HuukUCe6NakeMmhxYMBDRMewbHMU+Cx6lS6gL3WRaBVUAP/Ttg
AXDwF344sVM+X9X/CqgSYDRE8LrB9CIzN+1a3ZUjdqqtwGAfrSrUq7wYu9LC2/of
9kaDBPjL31P2sNP/9dlFj3SZOkMw47VSZpQO2wnXXMHKUPSCW+kkhgmUW5IAIpm7
/NZd4tLWtJ7//ccr9h5T4VS3MIbyWZ24412R3UqGiF0lWm8LareX1/coUasVxZRS
bUjSuXZzlNH7kIxaY92pbsA22/Y1FT3nzSqQKgCSWKJxej83mgq5tqmbfO50PAHB
fyFKbU2EHCkBSoPDUcjtKeAQ7+ANOiBYZGzLTTP3bniiGC2lO/krle+1AyyEX3kq
waNNyCoBrlzbmpeS7pdyrf67qWVFpBKGBVIlUwoicKVyV1PgVSFNomcmW180vNaj
v1HuHocOCqdtLyivZoiHBcPsoVMRV8jFyaebMsnF3x9wCxM63pdFIN22/m2qHaPn
gmzLIvsX0hy0GowqEreEj63l0kuUYhdPkf387mapvpeB8tl4EDmvUha5CORIWcwZ
PAvNSVpgM40w/ctQQeLluX1GIkR+Z6+L32jXxJuh+YNVSTNv8V0UsogVqxTAgi6g
OCRHQ+WUDZ9uwcvwqE26/htkuaWN11lqMLcnCb64fyRvXzhf4E984eYYdbr0KiAa
hbFKA+kvMZmXTe8JLs1FVGiCI5SH/q+RMs3AqaWQ+c/0TW6/Vw1xE5B433I0AtFw
rmlfdtof6TnKofkiL4h/uJ5cGwCsHLUYOakbVkrX4cgdefmvNufnn8a1pVdIuI3A
fB5b/k/ueZgS/9OD/CAM9GKS/AdK4wHbuvATOJx3tE8xLJDPe6gV+PXbBh5xByUA
aLUGWJ///sYxHkLJ9ItyciK/74Dzl1P4+XMozAFsRhzDCm9EJTc2EFfpSijXCqb1
HRzdoh3L713qGhsquEWQKXoR0J1imwXMXRAG3p3TXvFwzbMLhbhNEvkElLZ+EJy3
lcOwgSYg2rWaxM0qVK7A/CoX2z6Po6RJL79kkEbVmk3xJm0VxypKe549e0m5l4le
mtkZIj/iP08dSrqeWxyKzkACvot+KvkH7FJlff9Ces4TcfLjIirw2qZMXrFQc3Ph
cB5c5VGvbqXFqgiAr5M2p8PoH2DzEChs9nOkdA5ixDD8VGKoWbVQ71kZMe5pK20s
cpBMQYJuvkRWxAxxxkeN/ZEJVvphVfeTXfJpSgrqDMKVUhYwOvXI0qXvv862v05/
SPovOrkegcrtEg1Oj+RFjMNP3ZOlRlbCMtEeeIGKoKVw4Y1DHB8ptkeDmPnRLItx
yR10matkahp6SLht5NdUbXaFtGukGYuu0o2C8mu8vwjPKh9/HbK6h/ZnZTeOmSBA
tmU6NLRWnEEAA8PLLh4oHD5ff5R5KjJFiR2XGV4DyYb/mrSPM5vXB+geezz8eEtU
Q3pO1stCDxiUYYyCZQOqEqNBs/EcFa+LWgNEmaDz5bXH63Tm5+jxigFZgRnIRLO3
loK6avWDRBRQgRkgYRYBoyyUr/3I2VQFAhMRud2e/xcEYe4nG9YenVJj0wX3kt7w
MJUHSrpBS/YwUQObxKYq15x/qhptZJKkbDG/BrhWO+LMg7h0/7eywjtRYsC0uvbt
hSjzJkmbird0508f6qXRQdQVUlqWqOzIl8OdQOEa/HeJ1mJ2gnCwHf84wzWwnlmu
ZAcp5TD4nRmVvgX/H/WB1Nw9nlxPovY+W8XLvMGyYFeZAUuyAG4CaoMrUAnMZd4V
MLKO121PTVXyuY7jySUK9KpmM9bDoM+dDqdF9qtAbtX+KLoRPFlP2CzPikeY7WVq
W44r/cvN92SuU6kRrYFvMLXA6fnY/dc4Hct1fLPEJPC9iUYWibWMMEJ1EPfqdNIo
09IMGc4+p1hFdm3mzvzuFfNjbK0TjBU5NMUdPKeoRioqHnty9EM2FuGTmX2UX6jR
Vk7aaXX9jM/dMnLqH02VEqBToIPuRq86s/INxlasYt1l3b18Y3vEXz6y/JkzazHq
bI1fyNxnvTnDVj4NzYwKnkGAvVko8Ho2tTAfwOpkvWd/mby0wKCEEDcV+REk/i6Z
EV4fC2Kbrwbv14NIPz27XM+tNFTGOeW5o53tL0Zqp53CgRslQXSQJJikTaV9wXrI
BCMfToHszZEsS2q0k5LJaQqqsAwo+wzETeKAEjIL76It9pufLJs6Vv+NCqr6D5Qn
iPbvQWcgkQkreYBMcnrTqxaUxLNdR9xoxtNSbc/FY+q0LuS6Fu04cMPC3fPbubSc
O9dj1kPwNPRgNaIcasbwovku9FnEVlRwR0TVVZoWyTtbUt0FhS5f/wxWOtE3BlNK
vuMxfiLND/ShHMZvjXr3kwRpXVmwcqbfUnXErgfe7Bqk9OE46VpbyimZ4/pXlR2K
x/0KjmdpniJqeX6NluN3VH9twy3zNTqNZTI4bh5gzG81UJQPsBwp8mzqyUAmK67Z
GoSWgA6RCHspJJUSzuA/aqAKAzpBwuC2s3XwJf9PXWoNag0Kq7fgBKDjetEClfCv
3JpYVuyBOJpYQdXvU8MflCCNgtZ3wAtqnt48z1wabJU0MuFumfGBG57Ug4OCgUHA
llOwfgc5D5YZ5nNxHHGo2MX4ERs/FR538lplU66N66J6fGoPFNFqevcnGBfjs7FO
3YWs+HhJV66epgNFMF6nSUaco/Ytl18z6Uc2Nwm+YUQxWpleXQ5/tklwoEz977aw
uUpKnxUvkXKxIgStcdTxRMDFmYbUs4aG8wOYJmZ5tdLkI+k1LWkicrvv6kZ42iy9
DArO+MLV8lZo/RbuHGO/g9S1lebuqe7ux38zbdJ7dOfzrDLYhUoaWK1x+Iwv76Hf
md7I6SVTOR6b3CUONvhhN9ntJGfA1uQsqPp8SVOLYds/dLKKzE79hmW/8g0QUvWY
37PrP9DUaMoKSasEnbaMqWjBs1AjWMfjALRwXzNtWSaZvZVV2kC/6MIrjedM1WsL
xx8UxUP7UZ1+ScjP0Xfft5RCuVe/XmCswU0VwSoWef08rUx5c5uxiNVfIlOzhnzI
q/KE9QBDbtBdV63CByqCv4pj7hDSfAigX/CGiEsWjjtGSbJ5jt9r79fSZnI50Y5n
wDkZm/6R39+THcbp0cGaPps3x+G6UqjYRS0EWzK856pHeoYxsSM+aQU7xT3h7UIR
UQQfX6i68Ndt+24Z2kIuOn1VuMW72+sdUb3qZQuv3ATx6K7patKG4JXV20Wj1Non
7KeUyPI8s2xJhh/PaXmYzqknf9V5N/e1vNzrI7qXn0EIXUOdmjJ1yvXppjTSE9i2
ML3H160ZlU70mcmBJhPoDT4cLVfy7ncCg1vw9ukPSvfSoJbtO0QtSAcKzSKYGGOw
/jK6SpVESA3BYeTC90S72Z/a07XXoaZTUk71+6iaNKzUOpVXwUtnRvRVsnMTGq93
roCZDd9dApo/0xD9IH5PvLP+y2W21nDj0lNtJn5kjH2nPY03aLstZHTGKTfAbcZ8
s89TsaYEgVQLyl4f25v1FMXo9H4D9WQ8VZ8M9uGzIc5p2/xJeJf9+EjuqKIZXItV
AItA58dPbyNz6crvX+fbHmv8itJvNbk6FeqjK8THZYzDpsh0njbpxz0rxWVItcdL
es4eVwVyygnEsQoXo3p5KRZXeGwWovJ90ItiGrKWpmH1IdE0v89BOCCio2xHJ40m
HsA0sISyHWFMV24/z/ECeqSvGChSFNCojUtXs4y4OoSDkQO8GB8Aj2m/JK/fgQ8i
MrEMzXJmSQU4pgszi6NGU/pQ+m7QWKrWcsjWj3NcUAB2D6jOu8+mv38L15EU7DuK
Ib90ppeu3147Q+x3wImya8tSjDA/Vd7MneIQbDkD58378h8XeJafRQ1wca+nnTs0
WIKLEaRtaEaKWOFcBNOkwrpypihydedWyKKQbqkUlWrbZti3TAjffvRsaDaVhL0D
I0Vi73kIVw5yNa3EMYPDeQMUPGx2oJ4OlK9PRtzVCjUrAJq+4gDOp8QFx6TR330d
evWAgJO/gIK8jlbqMSERUmcgQzK9K2DcYfRgWhP/JPznCfvApyJ38xadw8uWr57B
WYfJykkUTiRn0vO8a5+UzQqbf/gIIdyKEinX89eytxCSuzLEU8dl6LB1q9MAVCSr
OEBth0QM7ciJmbOEw9khLuGWfBXCUhUjO3jxaMQE1chfrmJu31wSymsL096YWk9r
FyLyHEJmGsHOeJ7eyaQqotwBxslvhPPYZI7g4H5CnGs9dAqpr4gKAQUj3UQUAUa4
/teoelRp/wNKyrnm2whcCVw+9hZ2kI240fIxhQSnjVvw+4B3YK5n5PrHCvSzfxoC
EzcWW/sLOpk7b2MnZYMOtMAFDtpHum6UHeKOXObx9hx23Um7H7T7R7A1RuPVIylI
ElyLDXVGV7J9IENR1hSXLMCM5mtADjIoaDLvd4fsIUEjCrrN+IF3MEJoEphGoJIk
JaQ2tS9XeKPsAWupCWW3wrYJlNkUk1psi/dwIiTHV9Vm/WevTHNQIKy+TJPAQ6S4
7KjrMFxULD7Hgduj6rSgt43P08PL/xy5XsOQOy11zjC+Paetb8xrybIFiOHx32aF
TXFG1tjt4tqSsKo3+HJthy5UlbWj9FoVasUxT/5+uz9zboGP+xN8mxSyX8WsSfxT
kRJAMgcUlRda4RwdbWzbzMQ32SKxjG92pb4zoWGZ7Cr65eM9KbKOaWfs57mItGPu
d4PEUjMWNVwr32Uw7LX0R0x71HMjtI+Jz981pd2t1UC3ZB95WveETkwuM9waj1hF
Oe5lf8LLxREAFEOS/EiHLn6txsbaiF3D+ZCr0GApne+8eMCaBhpBOXOjhKQeKpng
yckhgpjXqCYIhKoqKs/Lc4rvQiUVO8ccGzTlFa/QZuKw4pSD5T+PGLgV3p3sf66b
HHhwMjryXwo8nhWL0bAMtLd02Eq86QqMTuLJU1/xhfwhf28rXInij9so5EV0+PBg
5tDQysw0xLHQk+fG82mSS+NHSgbM0g4DfFTnxHkUTC6QVfbf8KE+xJxW5JHO1oM4
JkSyxgu5srT8x//hC16yfd6L6SSkvHZw2Yj5A9DpQD9V1Dziea91FvNpQ/J7ldlm
3u77r9Y1qKdAG1zoUjZa26hqqPyEauHrEKF3tOj+VOVBlOURUC/Zw9PPiul6dpgX
TQJKOuB/jMLYz/XaQflnSlnl5SV81icSF6Do1EYfBnVWsEp/Gh2IdStwAr8SLHs5
x377DjKzxKdEhewEkvxp8UmBpGTXqwBgQ6JvDm5yAFWOlKvrD2cTWMkJs7z4Zk2P
HnjkEtdlgSo2CZwXb4C1xUbOcHI2Ga5hQrC+S4ouuV4uzZpHRtztjty0RlrDDOy4
mZErplg+XW5NCYItpapiW47j4CWD6gIVQvg8lLBHsFP5UsZPKW3kdc4yyEysDzw6
6VTRF+8hx7LtjkP1Jt5kC1F5aVUcm88mz8gomlsS3PEJz6zJE1GFHZ5HseLHLSSX
GdO1l9Hlz7cDGYUGDKjBq9d7+ocB7AgT+ky63hRNGVQ6jiL3LegPGYNjNWeT0wet
GdA+oLcm1DmEQbN9Hd/fbowNJyrm/UWZ+DGJdELv/lMCruNSfsqhqxU3GXIQcbFX
LefHnP+g6PtJsMizAfmVLWuS6b7rAjIRAyeOtDtHQOd6WtjEMKSovILZJ4GtgHWu
UO5Ja1vWayyvAVWzsLQinr28lmz70LjvKzM0qS3Jn+ThUnTbtcwOyDRuxlyWDk0R
ESTqYtjH41pKBGzye+Ee0toKq3gbdfinPpMUk9TyyWXyV4x1YxNT9fuSv2lDOYsU
BlvgT8jYeieRDdYXRmzUIxD9Eap24ncNngxjrdxN5yNiclvynCOV1VOLrF3KT2+/
oUEQ50VXhCLmDTBxAfXpwE09kEO4wWpcd/LWSXgnA83jZ+gA/49YPuE34EdaJN0k
rMYGsxWGRnXvI1HlCkY6GAebGTrXLEH+tvD1F/cZUibw4AIxAPWhTxVl7dqMI887
stlhTejsu9OFHSiQhA/SzpfK9hHiwNVYPuAk8bKLuiNpjYKAKgcLTCMu4ird+Op7
VNl7YpZ/cx6SGE21rXyx/743mlXdnazvFCLMMEcv2KG60R4NqKTouKC6Q2fH4IrX
fLyvjaXuM7oZg8010LcQHp98R3ccT+VmTeXmujoTFYg8RZFM3Be3J6UQ3eUXe3gS
ClL9qBvBdCldg6I+4rjE3InZFqnVcI3hxjsp6p8jFiMFNfVNI018VFxoV5mK7+IN
A3VPkEC2uhOim7wWNWLdSQaXBsRNL9EaDQqZN82BOkZlCfd/fj9fpz9G9/ZQTsfK
JSvqTd7sXykzmbn7DjYgfNWyo5takxax5J3Q6LvBR8cf7SKOvSRX8MbMxOghgwjn
5wQCUAgOQj7xsBwhcmSMYlgH5/uTuIYUsg2sHju67bPPfwHy47L1yaJveJRf5/BE
43XZOeg1oZaQqyNL18lvanF9S0mNDFQ7tyhjrHbhLGWp2YW0q/VALlndpO7tI1pR
3/Cu0TbhEb36tVrtxDiePl7KZR+xhFVVGn6OlS7wMiBnRa+Q7FNURwa0g/HRLw3z
cl7ETzJWIC9bKzIaOTdEpIt8eTwDU+UJQtoZuCGTulEZMr9cXSwBpzWVgnSRR7z1
TFiNNqFDzqKd8A5IyZPC1MGZ66LYjjFHba0B3CVYBSSFhz6Ct9PX7gMhMigN9mor
2hRaL0D7vdGRkIi7nsx3/En3Xoqw6pp5Rh6LNcHRTQEeWmLU5AajzEfSZzKi323H
OQGQH793ZtY/e7fbzXyC8dKaUV2thXqEkWl5ncyyKfi5eE2fFx8bG8W26W4nvmGp
yrwtGve5b1i7zjZwPbC7vB4goOxnBg44tKFii1A65Sm+GwTuL2Q7oRrOXgV6lsYp
pKn/A6E6YDqqqAboQosfmmrGRJrw3JE8VRtOdMjLhPG86AoI87hMiiSiG5ri+vh2
PjoUdVXMAJrTuueOnqBKSHKLXVVRpW38s2ubRj7cJeLgQu6bP32meCB6IUs9F8vh
6/AZmBcMqdJRd6LocvPF/d/94NWxubReLGz5PUi4bAyAuBVyZ+endjKITOBl9fHI
3SyUeJhQ6KlENSIPnlIfMfeXOlGq1ThQYC5SUQdin5UVGu/oHDSoNj1RaSj1Vy2a
pnSYb980MxtLMnbjEBNL70qkMi22TAA8EAZqe1HGILJEYYaAeGfCN6RtdbaBnTlz
wxMbrWCImMvq755jA8dMIouLiYTbzruJY2zC0DNjZN96tOjOlYUF+H4BZCDQMHCF
QnJXAKjlAMD3m+Jtby85UOOdedsYSHH4CpQXStYiGDN53rU0Qv6TAwrp6j7k+yl9
cp8kl1Dgo0OqtYrY7BwQSa6bKMkIuKU7JIHN8IeeeNOQ4UTUeEJ6qtBSae4lA1el
nqIWc0MAaOVXlFdeow89isbYuS+qfaSrPI4i6AbWcdy/Qt1HC0i7jN8sqCDaH4zS
B51TNooseXlJNeHrrfRJ5MR88UQxactH207V5hvME6gQ9LnhqK+cY3aB/cnUJmqu
qKGTpRgf60Ii/f00jgMEH/zPDxGjLzMQ3Ugoz4OcoUB4oluINrWY6EbxGpecdz09
uIqMO4pBipP42kFR22eoeppfZ4ribts0l6LB0QDgNfMc3U3b61aEDuvaHziPitOn
mej/e7aTNabSRMgC5/+QFmj98k8crVqY/7VqiCSPMOgAfCgDuBBWjXsahWhNyBr4
ugq4Lh18zOzBBS6RWG3skAztix+gx0slXQnWCVVOiWYr4u91bNAwnbEVAfGd5i3r
F6w0xafkH5lG8EekfAI0MFb/gwCs6ZTdhXK9HAujYDvaWGtFzDfoUBnU44kNEYyl
7sULofc6IlO6YqF4YynooGncykvcUIwtzgSOwEnBlPXOliDNC6G904XypBQFmhq0
F1LLi0rszhs4Lu192ErT+YkJSZaMcBa91qSU/Z5R6P60IduOZF5gPZjaDZ7ykGG+
yHMkiMTIWrCJigsZXU8Q78NSSSOS1c0Y8iqnyFJVp12e8wnzYLUwXgDgR7NGhbc9
xgMlJcrPyAxBxQ3pWz7P6yNaeWpgFjrXnxZCPOcCwZ7Od5548wvYS9Q5IokUwKCf
KxWG1aBRdNvcu28280BSi262jp9/IBHVCbCGoyxiO31+whKssTeAic0x2UFs4VsQ
Cegf/dDjz+bFV+wSGhd5KCKZ+gS8Spr23mngixCp8a9WTQi+c/I37qifgC/CFmUH
UmhpP7ASa8jTbV908ufjjwXLXzLWqmL8lxCBVX1qwtIh1vfhkhF3OPAa0hVHttww
rx6dEDGk3RSKyIMFZc594r/goXE/8WrUx8hJld3DlmOsBopLCzQJAWvQGd/Rk9vN
PNE4XBz6cpBNynyoiW+kh+CHd07N2IG4wcg6QE2kTeaReU1iCyPL6lM+51nWfecE
EuaxUU7RnlzmuvM8NvOKUe488eihUadpFg7IoXHr1YahmV3WzbhlLbNqJogxZ+lg
k87ujBq72mSRCdQqtmbJKF+CpGSBvt14dz7UUlkNaPnb47xPDy2fxsL7X1CmXW24
xSf6AKw6rGkkZdNnC/1Ppjw5e6jdqCZGAND2B2AmsT0vY7OKf51YQdFiwkB6YAWT
R82CYAf+ZPuCjIeQmsST+JYQ+kMdXQ5YtEQGbQNTnzPNDpajklczJSeyWVWwr2jk
VOqxdxcEZ81ea2X/++8ExCHJFwf0WFucEj+tyEbuDhN/mg9cSUKKEDUAu19d/nVH
pd8GYVOpTjIlnziXoSh3Q4vZTzvsoe5mQkj1W5BoDmg0G8OJRoCRUWrPBj/yQ2mF
uX+JsNhbHPJfGdbCc24d2Kcyqfwy63RMudOioZKOrLTlscWmvVItk/ZeOPHcN0qo
mGrA76Y1WJC7VO3nWG39ec/aePguNSdEKo1K2POg3w7QURj5Ih/ri3mFRj8qlafG
77TJ0uMfcBL9GaxkC3oLPW/CciW3/6CLIKxYWui3z6OtD5zM0c1WY/ZP5Yn1FEhb
mxQ9qfpSoxNKhmsaUazDzOSJX1kXHLC+zCjwpJTTtzkYIa+dpFBawTwaSE8GAsv+
Mvj7htVqv3ZDwk/4sdo8j01z9SxChykLBQhWinTpt271Zwu/dQkq3r0NchIssda2
OROoK4/F9ObzNNTTUMnVYCydsjC1HTsnQogpqeNr7ReVDycGWtOw5lzZSxpXYZsO
OEl7vijvcpi+KyCNhkUF+tAoF1nJNnwC59sM0on2koO720/3ueUsseUAHL7VNVKS
9KUI4OHAZO5q1i4HKQ1pMtZgE/MVsQVNahWPkx+7h/RE9TdY3cErkgFcl4y5mzTh
Yn66GWRWkEh+lowW9qvWQK0tYZxKxrfeURY+8R1855RJfKKiGsYCPBLcr973yGeA
7sFK14ChRbSk3PP2V6XCYg3QAfyqofLg2yTQDtrfE75HH0CMjdMD8oFkIUkja84c
8WdLdiXZKdpAg0PkN+9PWequeH18C7/HA3YmH084v0qgdzm+rl3maX+KL3bVYen9
qk4Al7+CUNPOHVkAa1nsaHlzbprpHs6vWBlWp7HQNEsLH6U6NBTG1i5osLQWRLLb
+5PPdQ2arDVSiF9g1T9KqyR898Q5zLxi8Tf9+tQ/D6zjCQPgtcCImDcV0u6VjC5s
It6KlwBnj0JMkI3afATT91EXUflw95kuzLhuSvJw2CQ5k3U10SfaYk0QVZNFbyDq
M7MLLr2cmzgzmTB+iFcEM61lNFS3m2ZYOl2FwuGDN900MTuHxaM72vexxcGWPAxJ
CKygn4jqzTv+S78H2R+IEbWXT6uTCdoE5H6+8ivepBd0Y61I/uqMYIPT35lW29H5
b73T03ZarIhAu+9NJn5jV5ZIZjAkyqfnCiFQY+FepqPVRoxvg6Ue9Gmw4cHWoDWB
yLpM4JwCeLxQimQv6WWMWyBozygojwfVN3r8PCH4ej4MkwY7Zsl87leHDqNHxBE4
WL96m906sYCy4EJFQzwUqwZhc39uPktHmkCfHt6xlp0XTABLwriCIS9hQAylmUln
RIvgk8AnAYO+FD+tJDcRabAqh0e1tHKLdZ/74BXciFAzbvC6qrco8jX0vBbTlRj+
1kboGNQa/dxQUYyjJwHEMbapujZxX8NbADIA2wMzfKOvPY0wiBG/qA8WykgQwPnE
Ra9TWwgMVmJADa4Jqe1QQ1hqYCS9kIDYzoeIJ+uoG0QWw0CO4tYftVua5SgXWii7
lNvbYj793uohbKA+0PD0lCE9BX7xkPrbNwEDk7VhyL5kTE4ZqaLwpM8BmQVNwdJ9
UHkA7ZPbcG5ewp8BWPbPq2bQ+KVltpNqYrVTbWaeYWLAJ/okGW3wYbVBCUWjT7go
s2q0k9aMhq9Z6r23Utja1JyUH2GHEYV3fVB3blESFsYZ1Ykp7HPwfTjhwIY8yWEq
xMltpgVtVz/f3nS7OxNcGxVdvc4lBDdo/rkiRLiTcNalZ+jlD2vKi3hhjvsBTnBw
Hk3+SdKThv06VECmdVW8pJpQoTg9dZ4Rf8jLS+iKKqFTOGXN7kMRK2C48IpnUg2q
ycdMbcdy2HR7uGTnswnCjdW5PzaE7wvnLwRQXf6JaB/EPOkSkWpHG2tvBj6LSf7u
7RSBZzHrsyjd84viQijDCBVO5r97lFhZJSSPUmy0wWSU1I7PAIu6wHfw8I2yHGTF
/EEhJASM+n8lHMalQWKoiRxgc6CEWB4i/fxkTD9DPDAoiCTUW9bv2kC8Lv3XQzCh
kBR3YnPSXip6M4NjXB5w+vCLRhXRJ41qf/z1upPKU7MgAXOu88horDQ54P3OlN9l
FWas4ZKCz0U99rV7ss1UsNfWrp8gs32BmDwBxu02r9766xELNdlGsHAB4Y5DuVOM
p1ovmtXUAeofHJTHVKFc1q3VWOQKSM7PQCztbsj2GU81xOO6gtN6n3XuWNcNuXaW
f/CRIOK6VBlsaxUVZkTsf31lzBQAxDXaxUvM9Xtd8yoyiuDJzBO9bUPxE/euocmK
9rvJ9vwLsXDuk5mURy6WUAXufQ7bO6EjT4WhRqliwVzWnCI05S/WtJ9Hvgut/4Uf
M7MT8p91nV5lIJu8EkGQ9/abNEnEzkdrhstGzf+NSCoTtYkRCGSCNJBypeV762A1
H1Fto+Plm7dcCW5quMCP0GYYHjtOSNujuackMaUwau7ENa+qNq2CWSDYVdvXr2/g
1W4xiysDYds8y/iTmwGd27zh3Jg0JaHRDZtXojELmP/e3ItP6E0TRgER/rXku1np
KiwQrUmpGfD9ahJp5JAjQQf6bUqH4kMIKZ09YfaElrtKxj5nyzP819kLFco8VMm1
caVl2gHhLjpADwdZ6Zu1QBexnJZCa4NNHqF9TucUFC03KBlexiiI1LvLUgD00aWe
vjBHyUiQu/lsiV/ajVqbpcPbKiG5rM1FQB3q8iNbR+sc0HPJTIF+Q4RRcu2XDN0w
9kdpcoh5AEjlmPZ8Ttjx+MRwsEYpJGxUzqNGScWsEqQrJDfoDpHfXQHE6i/hVt+Y
zgVukPmjiVyUfSBB0qk78DpRHK4AMzXy2dvkbn7Af+WjhMTPPAVP4J4QO9y9VEzG
BARe4/jvftFVUvq9CLAM0WMqqXdDCIyGvtAylbmtefRcyngn/dKFnCXIsC+9A19E
5619GRPyd+CTd5xgmf+XgE7A9MRCSpXwG0TnVxRmbOqyyzfPZi15a7sgqFj/h5GZ
g36FYlO0andGWVjENL0g0jvGrB4ypoBcai/O/TbXuaRz12zGQK+kzAVHn8AapqHu
faYIcQwFh7dQCRd5y2WOyIQtHqSsszlyJvhOyfuKpZ85b7N2zCGLLnUWDXTtnoCe
13VCw6RsoQEoUBuRf48bhVAOH+C/kH6KQ+34BJErKQVX5Cujcnkl9/WajS9VvK0A
qubOVn4yJ+IzwHYmEfP78kc4XBOZMnBM7qsOdR81+CHNgLG5444Kuadv/JOm0Kiz
t9tcV8wiHk684kBDvU4Xn6w3r1/jzPrFWe0eub9xH/PSGkWwsY58HbpThThZZb12
0NwcWmEPw5Snri6dXdK828FbQC7Zv1cvEI1lxVhVDY08QMxm4d4D/WgjgcbXenKF
RJW9yBVNnlPP4mrJIq+1Kp6HMqDZc7zgI3JSTJM0LpTYAFZPlLW+grVpncDB019T
d9Z0YahTz0eWrHzQTjFqAOWXc0N8hh3c69LxJUtIAmui01A7dgDg2D0Jo2zrXnNj
spv10KgaE6ZDlPrgzbCeomwexUEm4rsHLGRy7Gj0UegAxlifv1BkptbsJIr7zRTN
IGub9Y1jYgyFb2Cr28F++Fry4O+I4/2PmlVt+F/cOuGXVzG1b5WjZzA8ZLQLJt9M
Pwiqsv6hEfKqYL5+3d2nZmAPRO16qDBcdnk2c9NxfP+nGp61tpohKoX/sdXicg0x
EPHhhbRtW2yTzQCANW4QjBcBYbs4O1mZhRLY2PNNtWe/ibMje99PwZNaGAbzUit9
Twtt+zkel9uG7ywlUvXRKlgjS7kAObrsckTwh8r1DTEORRUZJPS2hv+OGiTrEHP2
y9SAEzDt2uQVDfT1amIyvsrZrSlRbWhayKcBrQKaJ3EUN1mvFFMfChsFlnrQOSNC
LCnud2n2aDc8/rTox5ZGNUoD9dRf6U7qGaSE09cwE4xkYy/4/SH/KDZg95LzUgFE
yTzAHsc4IvHXSnFoPYKMN861nlQ1NoVBCt144IH9dRBCl/G2nPsM5ZhHppax14W6
b6pDMGHFwsifeds/QF7mtgQ+bU5USnRl4Jab5f8Z5IlarjhyLw4hDyTy9fE3D8qV
435VIqR5a2EaHSXWtc9iqPP7F0LqWH9nIgo1E7XBLhfuOrNZ/wcakiqJiXiaQdy6
3cFZKluQ3/OdHKMbqXuJkFR2iXz/yM/LDuQvd97CgiHcwUX0sIz0tHGbN3/xJNFT
IBrUEExukBs2jJ2j5eKGwgEFyYGR+APlGVNIFpt8td0AMU0U8j5Tb5tCAqTf/0Me
qs5IsW6LLNGm5MRAP9WCOjIZkgoxYny+DsvesEM/yd8Nn0sjvAuuWi2+SgCRR4O3
0WKqg+VEaDTE+ldOpU12a5UbBKG3gQUWeQYjWiqzEwkiK3dgJQQu0/4P1T+zjdyx
cxvn5AHmsG45CKoIg+Ls7V2s5QnYf7BdAkSb6kBaW4fuM4nFUE1AIIxR3Y4O7HPU
jUdmmWIEuOjFL22jF3fmNWD6Eq1WAUdgU3HvWyXhhJiRNe7G+WwsAs0bwHmt5oqS
t1hOjDkDECAX1wk+Bmd+48ItlNbMVbf3eU9pz10ALAIdlxRJ9tUtiPZHEc/r2w67
4DOXQH6AXCVYiLEm5oGjtTdEBkUAkzH45GOG2j1+7yYXVrEtsTDA6LGEvq1n4KmT
vGJgiglMpnw/98vNjUHJGI/hIFiDFOA39ojpoIHSEPpLG9xnTru+cgk6QvJx9OUw
VGvTHdqjxg1Ga1qcSddXZg7UOuu8zk2fblKi081F0Y/MUQWxENEqoYrR/tM6LED9
xw/RFpKdMzhDpCE2g/C5eYNh9zQOdxb/rc7CZBnVjTztBsuyNIYKSL/UlGyAm/jW
ydn6kfMyCI5UCf4sEF4dFdI1pvyhQoPRxSbJSovS5o9PIY0Q8WhRGf3PEaGFaObz
GZsrq8hOwqbRTsgaWvL7u7joVPdwthm1Uctl3RTiCaQcmWkchPlPlqNmlaFuWZ0p
tdFZz7ndIuJeHOzI5H/Rgt0zR0hPLyxf1taYWJfwFd5/AXl5FxAS1c1fukD4anfn
Ho4mSiTtX0i7fzmJeh25D4qRpkB7AVBj/ywe8W9MADdc1lx/CL7KhYatPiT9lc5R
BVdPYg3A8XyGMowDmNrHXLTSZIIzSACH3JlM0PGubQYFe9Uba0rYNwRPb6QTfi32
woJtPhO1qP0JrMPMI1geYitIpkaj1ixoXR09eCO7xd18kYwXVcYdxS7sLFv2wwGB
gsGzZwgjUcgtxVJiBszJnDPUpPe9fDNsjLbYQdtXTO787KwMJpdTbyvIUuYwY4z6
BPyq3rMy2a/Wk7yhlLhKvywh111Faxi8LdWRPmvAFX3DE5FY5499UrhYwR3FExGQ
KwOO2a2Pg/d0d8+1zD4S0giaAPxlMVKyplVPgu9MyPbbIBOmlXe4jVd70lqfR2wV
ekRvaFA3rCO5WdsudCD4C2dXDKkzLb58XFTFTuIHHYuoHICTahZzbsAuyDsP9QeX
o2Mzu6yxt8LHKxh2h1jwy61pDPPPYm/7pE+ssOAzJZWO2HyTkpPtrcjCxQsVCupN
BJ7Upblz3o42Vk4XdsexK74i1tadsHm8sYMuBA83DPahRN+iNT3zoceB9CIXTolP
pEH4uBKrCCiLfLIExha1qxzOxnAuCNjFT6kyk0kDMmP1cIVUhZw/VQVtoowdehBP
hd53wDeLTqqO5hZLyAkG5iQC3VN35pvXzrHKpALc+ac5VQoWvDZ/GVctCnXjFZ9Y
7xatk8d8AejIx+//izZDp5PVMpazHJ1fc3jT0CvmiJTnpWxBnrD6h2JTWczw6pOn
wjsvcb8Sv20yxYzGLQSxCNpaA902wYIFmswQH/w2V7XdcPnpoJaPHPcRBfyktrAF
vGncvqIsD76VFAvkonoR102uVXu4goK1r5nwmauJhdmzkc7itnDTtTrkPJ+JZxi0
tN5vqRTiAl8iQXCidO6UCFKko5uphk/4kCmBAN9Oh/cN62wK6oDlzOI2a+kwO1Nj
eC00bYgrWVdH8WKoiZZcoe3mZCgBT1lWGe87YybsqxKBD4o32kPh4kPRywrAQNbN
nt1pYQ3qeuLnGiHfkF8uzN02Vicp60zNnM50in6rdN4KjBSqE3kD5lDr3RROTuBw
opePq4bCNVNiw9nqOY5YyiLBqb07DNIv/DrlH5ZNqMGOlHA1UKfZPqfOnAtyB8Qn
B21exIXBwMBqdMEWwJMQtzXvAa+1uKsCZi1tgWbt02H+8sNlRwdiNfdCmOQBRUNT
aQ4wF+9AKUSeeIcsoT/uv+90RI5FljetTnZf4DZ/HRSIC0GZzqlaNdzLCuBfJjdw
NBCFWcWml4D5q9xiXamebHR2weuYhGnb7xkhk8xKr7ccWdoe26DDcgU8jis4d85d
8MfI1tPyzzhozypVAnQFgeFqII2f5apVFGZSZfvW1SMraa97UPBxM65+kcLTTzOc
jh3BQRumJDQ4w1+yUsg292WtjW9rqVP3FavQc2y7bWWE6GrhQQsh/G3BuUjenKuC
FaIYRUq7dkZWGu7KbZL+cRBxLLwEjkdu1vAvSH/FAY1Ea1h9zDjR7ZQwhFxNsTZ1
4SrkCsDkQ0sQRlFwlscS9TVrR0Sjo2VL/Mfb62wPUCZ4yCthRgUAaSMWNm+yGL9n
o3TwDXohN3oNiOFqqWTN6caGjyErfMDRj9vOMbh5gxHgLOo3GwFSNa3FQ9lsYvBm
5EhSiTc60hDMvaJsUuzZtduMkDQqzsCq1ux3yNhGX71rJUBgy4JvyfJB+5yU5bIT
uSN85JzyA8lAwBno0BQq9emJZ13IdItDJam2rip0aD99t0TSwRycDvg122T+dQAv
AlxXkU0xaMKt5ISG2bE5b5jmbLZBNqIqqyuhBk1LS5zSgf5qYxJqAwEwhjzzSkB8
KgSKDqY16b4Mv8LDsmQoWVzMVSmadUxMrEqh/zNSm7XYlpH7F8Is9TXZEiorCHTc
uCoR5RdH6r64GP+j1BSWWcuUn6u543RfTQ2HEvJwztawMGY7crtXEcc3kzKM9rl9
MgMygN6DxxEkgB16xp60LSzpcMDSS5vWoaOmE6ofHuGW3y+G7STYqIfyQAHcarRQ
AHCA6FUx79yol9XxoHzRrPNSz22R3Elgcit2cklCxi9csx53CNfD0p6qnVFtYPo6
9UcWJjqb9Ji/xZmfokdGkszOBTvNq8zveEHRbHYCLsyIr6HXv6RgPpqmXkKOAuIO
QQZudxElUHAYZ8ugMNdbMgvISAL7SSbkMLOUURgeQAIxkBh+6hG76zkFe1viNu3D
DJwM27oBKSBxMaEoTrpCim4vYkihAf0b6FITZ9fdAphXZc63GGQbj/UmVentzA0v
pp6AICe+1lBtXFT7r2OHPtaOCWuyIMMtiFhkmtD155jBW+YajFG2sKY1MCRaIhBB
jW8zIMpjItmVfoKIzoZU4b46wcJK8MfYqqJU4slItBOTpWy+Km8thBB4zEoV4Oms
UFNfONEOBioJab4LQ3a8B/UqL2Rrk/y2ow71JLJqg0R/stZBDoxAgwtcMs33mMxD
ka0Jnphjyi4ULjyKz+/wTwJfFbo8cQDmrrjWcYAUWLLhM08jOSZDmlXx4ftFdmw6
ky2Coy0/7rHDbw2ojjJEvgAGExpqCU/vl/fUNlqjyNG7rol42Faw/L1V85qOtJIw
8VhqBZ68cXyIdiNknoNQfHCuy/i9B0qjdiSJ2tgOZX/ye2jqslAvj1ydcpOOibR3
DqJjDuWyfSFUS+MsMd2Gt2hpLoI06yk3+uaOwyuOsCWC5q/XEFXqm3hLpHDhQ5E4
sYOurh7XiaNs0FgVtq/xcC2/2QGCXmDOiDruzHJQINxqYgDEgj+t1m0WHnr5bCJe
etP+9tZvtphKkoaX6PmrjyVFwgpma8UydJpqKn26cQQgqyppDvUZLtDnqQHz0Fba
w0daXVXQ528D8oW0rHRvosGcmPepnVnXtO4F4a/PJ4cOq9ueIqQkKA2//GoNTKPj
s2eW4LfSHaAjWzuSAb5glQMqHTgwZ7rqyEcC28Pu5dup6WNp3LISHDP7Xrazfs5H
pZUTjdcfyZT1pl0PG/Zi+RZz6HPex+XqabvsC3KLk64qOkajsbUB09T143YL7y8w
JSa80N9YNs8wTreVqcn9hU2hN/4f69C2f5UkUjzefkX6pFipDlL8kzKRtxGBOhqT
OsotPEAG+N17/hTwPDbffuikAmyrLc+W3sFGYcwKVxursacVf806/6gNc38/RdIT
1AYwC08e/RBQoGWyh75rfS6squT01GpqlMHjsmA0V0jf2CNP0rfAToxlbUSMSQDE
FzC+gKpZClV5J179Gz9+f1Hsmf8vmVzQd4dr1MMyVMS7zz/MT/l5smY/pbPlJbNc
gjJD5VtkDYkgWgzEJWKK6Q1gR3eELlbUfRPnk/MJaSRo2vh1HKsbcz5l44dpJruP
YDNLYoReUSXgEw66IMQCPZFsILWxOWhUBjze5rxk1MmmRBezdldd9EF3F+MPMK38
VlGtaXvkNoLLc60ED95p1PxYVOclwCtxXMgH5PcjK34TlVoRkZt5wFPbgX9D3Mxu
IT5qpfrLMZ1MPu7lXneG7v2w6ta4ABhNeTzQTnFHO+5boSqnyjNxNEn4TvAwMXim
SZ1C5xfx3p7Fe3VqnyyWMTOWUMc2XalVM4wljXSwLKloYp32BO7r2w4tafkI5T+E
ykZnMXguvgMANXj6aJSw3F4cceMGesylKO9trIcOFsCWRzXoaM0BcdRxjgVP5sqj
B9Y2+3C2OOXekPqXct6bCdqGoZWjmExHZMx2n6oeBPrMeWGRBcyFzN7YR2OgfXue
wBjOg9To1cmLSedbM0IXwpWAWy3zEoUDvKps3VaxBIM7m0CuH6B/LW8ovbQ7Mh0v
dmTKpScGLDt+zuApwTkJYHYVPIPxRTEtcAEOKoUI2Bz4h8onKkTQ1GG6T+Vx6wGk
5ootJPBgoPsyoNATyyRZHbDztPaDs74baIdJU1UhxnlFezS0Zmxow5mr+rWkOF7T
Tm7fCbrfups57z4+sId4+wHLu2AlVI11IoeSrrKPPY46L8t/pf3pzE7528wiZ+C5
LEmPjd6BET45rK8hwDQTaOuw44SXspeY4OBeirXz+YJsmIEsazZCqVA7yyBnCZY7
BVhdwSuSpVj+tT0Ok2rqwiMG8N7HP17jQOi2r1IXXX6nRkNRLMbsrsECOPSyHgSG
mvL9Hz8RCwLRYst9IvDlhpCLngM6wdxt7nnqyivcuBxO475IkvwuifB82nGLrJzB
LpsYRMT5aD63ZqlktCWmweDD8WVaHEa8N2SyrN3mHyZL+HwHB0VsZjQj5ZuFzb5I
QRq5LwyuILD4DjjjIENYtU9O/EkDBhMz+ekmTNys4+Frbln19qtIsiCAgNi5rD4B
wrtxOD6LlqhjNgItK+s7Sd9sLo5hQUC7c2/vJzi3/2RntYdE6zdYANtoqo5dCRd8
7Z5EkATQgskKoeXm3hd5KGqr/8SM7GMw6ofIoYicShUZi9dl8C7bymw9soDSgpU0
rtdT12/p9F22pj2sse+Vw0EgS6JFzAGohEFMOLe2vhhkav2wr0wtLO/2Wmi9EgEz
EtGJfytWVwqqxLhCBBT0cVdJjpLArDsGmNLhWveeWvyP6Lce2CaMFJNMdm4qVbE+
v9iG9DowdH6/uOxp+rMeKkQ2dOGbiP4OZoNFaDaUByJfsGhD4Qe7L6MR8M3vVWPP
Nm5yZeKcCVdj4hIALanbV1yzckrB89S7J6sXdM3kDnma8i+AY4q3zBgO8RwgR/N/
P+elkUed0MslgaaUSlnErMWr3n0X21W3CGIGQPDVUikviXAq8rVwD+Da22MM/tZJ
QT4opXKBA4RdrOMNYdSLcqNjJkvcwp3wwXyU1z6VUfVEyX98jDY1O5l0nBV7DJaq
+WLDYA4oCpRk7ZmYV6RNQRYEWOFXiqSZiRcL+hmFCyBHG/f0rZYfMUxWCFpSoT6M
lgMatltozfgZKIN2ViKmvJihQFTFMFXicfoTlgEtdr4MsBO/Ty8Dk6HJpcgUrkgU
cUGPTEXqG5rs3jGWmEeH+ypqIM0ypjpA8fVrxotGTNakl3WzawjL50pGwf5zIQlo
UfkR5ZnVMUkWBm1/DmwqYjctmwrfaEEbzH4yWuAElfcughdosLfnPb25dTeXOCZh
klLj2bMDPZnW97KHgkMilV2vpZ9uzfHzJFousIxtUYjRRZwJQz5wDlNgQA2+z5Sx
ni4GTz7HklEdlwyxy73TSRgJDkdxHrZOIZiFSvJSnQDmH5lwqPkaoIpWnoI4//uL
iaIelQiwGBek5KCwF43sbp8p6eqnY5fi4/f0pBBAP8Yw/8a/RbEqeXt99hpxAWlC
ZZ0cKm43+w4vb9LQ1UlFihNKf7eilAwmwJPTH6cYOhdpMAUoE9okCABrpnclcFOh
4qKD8ssPel64P6QV03hr66CE8MDc3T+3f6z3UHj3HhpJQaAhXgM7mvy5zXnjDfN8
Z14e7lQCmxMxrlSDXZWVelL5JYDOqtrYsJowQoUfXSNp/WDBVtVKzGISMyzCTjqI
uzPXLTr7bznL1vWQrQuhlVBcXT1qaAR9rSpsz4ABiJuKc1taJsGxFdPMsoUUeOBL
6gO7K2dM0HcpMpDsNFD9woUcunPgVMCVpcjjGkVmucBtEbBRkH70spFieYpCjDEP
ReDDvlMsPuFkU8hGvCPpsYjJIiS5JKodhnZ1vw3TpXKSeaVz8zC4mi2nO14lhRjP
yvthDZIjxrfN+7XTg8CDviiW5q2cqUuDJ7hzRHoseuQ5AO3YCKSD0BR25P/aFTkG
DRocgLAlOJO1xB//E4Xz5igCwMrxE+wu0bCNxU8jDxd+55KpyNi7Qzgbe57uGHxJ
1TbyEHtCpkiOfdXwjCid8DBFm9b5y6Qzi8Nd9d/nLV1/pje4kLR9iwdQPumGGTij
yYq0e9CMO9emJTQ89iJ/lGlOsksXiAa9nUX2xn0V2EZUxONeBRjpnEHpJpoCOTFu
iKuRcqQxCm0jX7L1GKGn7wS7s922pS6EB9QK0bonF9PxQp6BYHe5qYdj3Ld4YVm3
YxNAz1l/bKRRYvRMowNZMnWKq2IKvKFU0jFm0gLtt6Q/unaP1IPl3didog7vlV4h
yyxQcs6vPA3yUeGLuvmsilRWNcQMiWBvfqatNHBXoINiROt8a7djO1Ncgpuip613
HSSIgsjdIGI2yyFWfaQpHTeEwOaW3UH74+1pCmgetIveNFjDQH3euSCPGXX/ggmo
pH+6IepxvsjJL+hBRVDxzq1WMYy93Wrbq/26nza7YyCSze4cOmgoc4SVq+G3JFkJ
nhHZg7mA2LmHgmv0WJDMW9nVyCvd/Okd/hWwCnwjF6ThcYj/S/r9ryt/jA1RwmiA
MtPH7NLC0oATsDDEiz4lja3JcO0vrt6h4G7EoVGGBMXtR6bnEQhseri/jyzek8cf
vMiuKDp24594TXSNyHoEZOwmoF1+Vz7l5e3MoPjZRSrZYl3q4z6rJldnscDK6ujJ
tCQvaRIFSISmgyyxabtlO9qoqDinj9Tqp7C2mI9fDbVNpGu5TIOmz5UcBXVmNDy7
CWCyLRVjM3xw0b5MN7+JZraVIaj8e0CP2swyjkkPUguAh4zrAxiPFVvq2xuEKyb7
Vrt78rYVDiZFN7W1Abx3Bf0auheaMoY5sQjZh4k967FVOszn6UMt2IK4444za6wB
8OUS2lEroXKZvv6lZSCtOmV6GR5hnWyXAtaoinAtrPfuib7ym28K7EFda+y8qOKb
dueH+ldGL16lkYZ6ji/l3bxQQm1MWKWrGLhU62Ll5VLeP+ExzPtDDM5oMvDnHSPZ
octCl9w2IXjvZEMbAjxiV/h4RUmYcejViOzsyERbo9rdQRu1ambSFAaZeEziiGdU
3WgCUtbcVJ4KUmpEvHqsneLzlY9ZC3HhEXRBZfAAgxPm4pLQ0YZA0EDbDUKL3G0H
GNTOORATHvoTkMRYdt8WmCZYK19DLmRKtXHVN4KuTpYFdhQbQpb2FuPcad8dIPmi
k6C59absBTeu3mMlHr9pQYUJN6Xt95NlHL7wkO/cipCMb1ah+XMLRCyI5aJdnGuI
Tvq2zkvgDvSy4sDmv7SrKUotO9TEYjHmZdXMdQ6KxIp1kZo+/Wd1JRTqSG6mXzkF
zWjD/IEP0hzsj8LeuaddK7QChQr+tDTFgVMr271CBGYt0Xy8xNoOlwTD6wVUrcdH
8C1uUzjRzJuLi6raRVnU4xD4tsptZYWlviIWeFUQ7+xe7bzlkGZ0gPlpKAtq67aw
6tLsYsW7LsAtRGJYcnNG7Qj+dNiNb0YxvDoJ0+srzFxY3ZYqvg3JKFeKI1gotHZl
fyW799tSYj5c/id7T8GNHj90YbkSXHi8wZkPewgd6BW5darSAAEWRy79ELLzkyX0
s8pgR+gIrA4830Ubx8iRJMUz9XM6dbjpIr8/kv6qDl4h5qeZ8XIfT86g5JhFgQSr
kfCzkFRPlEcWDpGgE6V9InGrKyPaAUXLReRcs0KoNfiJEf/Hts+erBcu3+QFTDp8
X8wSnG9vt2QOVbG2itwD1fYB7TWEs/UHOupWsfRI3hjzSnh+Ph0qECYty4jH1Awv
z932uZTclesEot9BwER7ZhQkH1dhRjzi/0Cp3QNfyQEWGKhH7qfawZI+9aDz0Piz
emY2yHmtDC9xTACWEORvrAVL53ghkWAgRL0Rm9njU8q8IxrIn9EgUZc3oNNHdLJ/
V4ArrekONIvEn4j1HPKaXF2OAKykvbC8HNvmawzueR+jxZgStqAFYN1BUw92DVlx
V6MOhQstqGoUSh8SiLUYh1vq4RE+mfPcRrXQViY+DQg3jKgZKMYyJQfvGOou/r6D
bojSl0ydpgHN/6+YEwSE4kEBeg5LImmxeOZb/ZNYu06SXqlgES2afCvtR5U+ct07
b2XEHusuc0ySriDkHiyc9djktW6l1QGy0FJ0jEC8UtNOsqlGSjmWfHxrM9p8chPp
q+V9vBqRd7Z3wd1NvHxWooxHElfkI+vXv5XS2kMjEU7WShWBodvJ7lS0C/LxiO1g
JPfXXyXVhOzoxxBEGonOXoi2yMOW6Fqs/WmcjlIpwV2x5ceuMlhhNfhaoutkEAj5
l3i/ejXGA3ek3tBeMBTiFXgSVihWCoohHQjqjfN5JWmeYuoqBErApu9rJHHRr6Hs
nmb1S5LzDTsvOxXcwXYvjOiovi5AWRoYwybIZhsqUg6IqjXVf9rCSQR/oYxN5Mzd
03wvisgpLxtj2m10BXodriFpdA0mx5PZaLF90a/16OC4gJZx2QZgv7m+1r7kJ1wC
vgCakF2N9QJCebahH0uEkdQognNFD2Lye6EemtcctuSJrda8z/PtgVN4610v9seP
dzTKuZbmKeunRLAzdrdHZ7Gphz+tdbITLHBwbblx+jLA2/FtccyVTTtvS19wuDUv
wDSZLMsVYPWP4LTU02CrGTLbUlLx5QxdbDsyyHYiGUh7GI1LKPSWRaid9O51IAvA
QFn0CZCuHmjr1j0oCBZ0azIvdB+7MeNyMdtPq1yc/p5nAzJyqOi1WVItn2rsMinl
XJ973S14+UyoJ3FA0zPI6qtIMmAOgZX0tuNRDXDpWRvYN67y57gL43slfv26r3sx
KjAnYXJM7cwZsyGS40IjqBpk/7ONiCctfiCFOhjnGGAYNbYcuDW5h/QzmbK0muLY
tpoc1n9wZwskFJ7Ymnduh1eWXycA98CLoJJzM2V9kpD6elcwiHAYNnqFdAO4M9qp
1CAIwQNyJfwvVlBk0bm/8bAa/Ys7PDT97mj1Eg+j04HYX3kqzKxslKjy60Uf7Mno
X6JsPJKcGhhyh2USCorbxbOC1hsyH1/F3xX2+9O8OePLtMbAclEEuAm+JsjCzAbT
o6baNjdIlBP/UDtDS1RJEZnm3Ft7MhY7Ph0ynLCwAT0KSY93XG3rj62SQnxsz/+e
IxEo5BJpnPzC2Voh6S/GJbvhxGiWS/jd5E5cNVl6MOMs9x+666UmpV0+SVL5W/76
Q/jKOX69WqU5K7JFKlj+AIg+WZsMNRNKsAyhRfWpYRL1xM0HOgKSQmotH4QM11Az
V3jR6LcPGbKq+paAveE/FW14txlol93esBS2UxRrUrYXGjztvDjvI8vy0gllDeBL
eHFKKhYPLNp+PQDVyR+4JP2CvxVEjo6UDbpTcJ0yEl7F/ZmDHl00g5F4hnnmRD9U
IdObvpASjvkvg0qdgYwxV75MkbrPey/CbXAL3ROo7/e1mVW/ZBiZPLOtPog48Jud
kHeWwB5ZdU5s2KJrn04tuH+oTQIdvTN43MM8BweuBSmSUmBjxYIBPr/+ZK/RCvYz
C8mBiPyMLj2P1dd39RZSHxpFlFVhL9mtjLgeSio5PSd1t8RCpP4iGm1cEq9g+XI0
+PDI/YwHPZw7jGs5DMNn7DtG4T9g3XT7CpxgEJ/1Ohwnv1C0ufOBkUQcJTl2ku//
AE5xiSoniFo2wNbaTMq2qYBFhYSlRPb6WPbOHyXWr6mWZfrrmSjL58BbG5E7bwJD
xGszvnBdumHUR/X7SYdHZGeGtVO/vtsyr+vaFh+GwiOtKpmYq/R1JoNqpii+84m/
ZkouwRb0BJpPGHDgCanVUM8u0jZysC9Qj8v+a19F6s799r6oqGd08FgDFI4bJp8i
LDPnkR5xv4MRkUI/5sFgkruWP3r2sbiARtSvQe1IFii0oO1+zjn99KKV+mCt4MKu
J0bIBO1/F9WlhMxYZRGzOp0bCek74jLh4po/3K5r+JbKM24AmClR9GyhC4Uz8lDe
lFkpzfxZKYNogNhFE+wXrZMev+z49sQIMEFndM1Adtf0NpGAcuFXNgVUP9hiexu+
eJmregl00w+874J4HjW7JgruacRRrQHoN9Pv5PN+EHDRvH9jP0SmQxqTkLZRaFCX
Zgax8ZLwuiFGKP2s1qPP01IMNJrpzjt3Rr6AN48wn8pDg5klqwX3zVu++w8HCv5F
mOmNkUSVuO0ZMDoa89blp9wUwAOYSiBj8/yN6USwqfMT69XELoT/9xHbIrNLQDgO
rG6nJ9MRlc3tbanv2nUzJ245nST4PdKxIcRfrh1KVSFM7CRGn18yPLTPuL1wxRW8
jHJ5EzB1dXFTkhmhHWWn50lfcxncqrwUSPqJD7SO4E2vVA9BYDRyk10jQgbXtOft
7GketFAoZraiCTxsGFKp3D5Cb6/XFngXm/EpTxRknONavmEfQ8GKmwPNa2zqCJFV
Ztw2QBLMAp8SWSyQ+LBz23ffVX9wf9uJGD/BQZZQcUF1+W15xpnP5qGGxdir/n3N
7jBrtcv4lDiebz7QloX9GIxiTkRl/DnTJ9tgHNlIiJowHaiZCNbM/ju/JEigTb/9
jZIFwErYckk9QHFlsN4hy8TTfb1wp7x+wie4f52+H9d3cqYHKtIYhYXQyDOf4CRs
XmXJ6pCUMQ3D9wNhhHctMmcMS8AKcxob5EHru1MLf1QXPriwSu272fuqF8gSub22
urDJJ7OH9cCEkEOCcYSNvBbrV+zcL/Hxw30OAOpZu8IK2gldJrjObcHx30qdwvrj
rdxP+DBQfChCKnTJpOdfN8tiP17NY3ekCgEd/LJgI1rZx1bgsbHOLDevuF2ObOWL
NoyYDhpcxCX3vl33TO9kvLuYANShB0nbVghTINDHtFr/wZpT1l1dasf/+zzy0G10
Xf3KY0WTnB4YgCAXrjoKDH4LlQD1KxBAzvEG+YzlPBpgAlavhdTE1BggTnwJJLF/
QWwu3zyWt4PvCiS/FP7hewdx3znK6dndwd23skha0rujnTx+qBZZyYOiCzFUs61J
ysUA74JBGeQsRnHwJeF/+uNdXfSMYYg7EE1hSqtYihHwmWopUy4jZ9O984T2RJtv
4mOPPkSxAb3rHzbuZl6q9uluggVqwdTcaf4XMX80prirmsbULZiVB0cy+kJuAAWr
+njrg0ZZ25nrIwJdh7GmvXFe7ocHMg4bI0UZJ7JecU/QMd8jJiUhNm4gFoI2cUr0
enW5E01JiUFRfVjTREmavA05ZbT81RvrJQ/UZVdSMNWiniIvLwn/3+vxIPfLZuXr
jL78ndchKhbq2qtwn8N2Uo0bLWg11zshJ82Y5cvEGqfmj6oY4jklAU7MPG0YDW4Z
1+IsCtus1juLtoahuqE3poew3bCZOOiiV0ZA/VVqfgUOpnSqMqCTk/oBaklZ6BvH
XjDKe1S6iriYDhl/xuWexdqOrxWfK6Z9KrMyQA0V30Kt4yxZ9P2GxR1Lz3m6jBve
CfpoVcdd4XF1L4XVxwWwHFnuM5uarwKoqE955DjAMq1J7FNeZEjOa6JAEd3wfp2G
Ln1/F0nlQvDMHJRv48eVJ/7AR7QHshKGUf5jUXAWIZDqp+M7VkXwEXBIbrvHkGKi
OzpeK8fLnchwj535PQ9FJ7lSmBwVJYEhqxHR9ZVFD1ozxIHOWVrjDs7YFchMd0JH
q5fi3fO0KwpDgcol1zCJ7Aky679/BPenTlgkSrAjlY7fdHwJGgeS3AE0YiTDIZZi
8KdB5OgJWyAVy5T7N3FYmrz2hnhByoDK0LkbgnjSC4a/9Z+wOwaiPQ4luf/2c44C
oyArNoHaxoE3wPqbzKaeU3IJVXCqLGDdcYykGgooGUYfQ4BI27wIH5LNEZXs1TiX
ezp1gennMLpqyPJwKUy+C3ZGRqoUYN2W73ga8R03lHiuT0iG2NF7TA7RfcY+Dmoz
+dMDCN2xXF+tX8UWgzG0uNHpcf4ylyCgosz+nIJYkQEuVpqhSWRF9c2rRXdpJVpw
S8arRMTXSjGo/D0bteUIq6OayUrmu0iQU0YclZNKb1vU9VmBiMkf/RuUJ6A60TTG
QYxOn6pKWLya02SkGcW+5RVtaAztxSHtZiDTkzpPgtglFa76vCzkF3VBP4p9CWDx
XjxjQ4U7KZwYl9D9v4RG4qynJ+lkBB5MAtycEq4hOz+fseUVUVUlZ9KGRYV1MHEb
3sHWN1mjxJ+Fd/iaNpZetf9jLNEh5Q4WIx5br+mY3uETUCkdQRwbORukboLX3whA
yb0LhLglTF0sqcjVgRfpRliVEGIfF9PJJyG71FhhdMVZOJym+lWercB61htG8Xe3
0XRlcYK2pOdtpREDpSobFhgDrI3eQmkjzK6Gi6xupM/5kIdffet7z4Yayyt/65pC
e4feaKitbeZajRixYKzfVBodjyZuzm/e//tCR0RGURL3RwscClGpwXE+Y+UoggJd
XH42XwhqIfyRLDYjvZX66HeAU138Totoc1347VEthGN/Pth0PQFxHZvNskmLPevn
Bhx2RnxZN+fZmueBcBzfdXHCCvW4zaJ/4ixhisq5rIZQrmsWWy4z5IhCwXjpT2Rj
6+RmwmtjLCwSW04p+0VC43WbA6p0L085xdxbatQelMYRRoA0dbZOyTag2kdKWMTI
QgFRdBxWWLLNVZZBcekPUwITA6qqon4EYPTOV7U66Yxjd7SKtcZze83b3wJimNtW
Qnj270bXryRRIMHcxX6l6rk3mXwChmC6UxSGmg1pbIlvIpVm1SikA1bfdseXxob4
81yJkabx7mX9x4eSEhNHOlVs+WEKz+FYwHgjMCUmCqFEMnCF4LkAeE+6LWzAzH89
twgb9L4HMBbtthUcZN+V49+u8DIUwxoMnr51jBW9p8V+uK70STChDUlq31UIUbja
mPQQxw8ftUQyddMAWTLii7WRjip5FzzqqzD3NmzLIAr2Q89PksR7dcCVuU7BwTX+
ZigYdjVlfLwhLyxCHA8ZFSWb++dV3ENLGoGRtu3TbKOWhR9yz/9q8XKUO7UUc9G+
FF6x7wTPdWEZngsQZUQw4P4kh3ABx+E4EHzZPCbT0zCzJLhoGQS04vQzPtjSNHEi
deAW4uU/ZID2ghGCxErmdLdy0KbTkLsIWO0+ilNREfpPlrRvt74T9Umcp7TgvJwc
/9cV5xz4R/uZHx2vDOsg6AR/yJN3cWUKFWEFx9kpiUzglseqoHcE+uvgDuys45pb
XopslxYzE5rGHl7+XnQmEd/mbZKBKksGP3IXD8+u+eORSwShl6hLj+rSCahPeH/y
60FnBbsO9bN1V80J3LrDbKgynWZvazJsfA5weHEdMSbX/cy/JcLxSbY0l2WnafNW
VjabW8zNioW+LwoHdbG/WU6qVe+zbLWBho+aYabnWa93GKTaw//XkUwB92rGqgHA
73R4M3Fkcl1pjoeCVuUKfRD/CGI1jRPJs23fD6n8JruLZNNFX5uxWgvH/THxuqfo
//pofbSRRjufGimiqBadp74BhxN+6w7dlMrBUgH573sBCLYBvG0/6lcYwzFAquOv
duyyAOHTH+lm0VfCFyl/5+klY84K9Ne84/GuIunvpV+H3lW2eQSrdwH0QvwGdnC0
XC/R5K3HOpAeXqWbMj8D/2jiQ9iJa7YUDhVnd1DlLmR/PIydov5q88/IHHjfttSy
ZY+VBRwjiXVrJdWinxfJ5h/ZCkibMTpSz5VedhdymUJoNzYpzbIKZIpQAopp/rfn
0nwae8PNDwUHnPlUAlVW3tzpJnJxNiX3p+FAOrYaNIhMf9iZMVlQTnsiH6B0h1sF
1znyP8YegL3ug5fegNx6xR/NUJOFCk/oQ8tTwe2452+uLF+7QAcL/wqT9gVF/Ugm
EEpz+SH24uGsA6la6WyVpYbvOJQkJEFidbztqqN9xuCcDY2PvEmz6LrErC1AjUxx
4ufE4v8ibLKnKV/QsIvp0QA3HtGqPiIIFwAi5mTOxW8U3i6PEFuPelGi/1f3TG/4
BIq/qy42d8kSSY9sUmBau4P5/IVSPGRMHhsgGcG/zmdxLRUnY8b+ASKnjNk6SLLh
qmc+SZQNuuOvz35nB6FgpP4AebbWbhWLjFH01SrqrVQvsvg+HVSUawpdBwveof55
cmUJTjjmmXwWbTvueENhlwJCwYOA63y3W2haf31N0yd1p4icQ1N0PdX+VoRDF01F
9zttSZLje2qm06vCV7IMkFrtwXHsBedenKxRNlVzrnXVfwdltMPMm6XBe4dgh/F8
3e0HXewZpGpJ5mgBU6rGu9xOnxTVdkbbWcTBaVjtcQcZXPTZov9RSMZ7G4aFH3dE
2RYBw31goO4egkKNO/Q+r9Xp89NfkLoEQsrF0duNalBzqYBHR2dqbtcwoubqEqI/
4y8L+tPE+X1Y6wUNjFLY6wd39fiOvbMvTTZ9ngoRBI5/aWWubT2t63kjrfC/8luI
kl8CEFRufH7TLoMxfUfLvxbkB6HvrcHpc26hFFcPWRM8Nt2x/7T5N1MNJ8a1n+iQ
aqGAn9jqeICyNKSppCh9k93uIvRQXcxi8roHWMMUz8Y+XS5Sfp6OGwGuNxpfBiVs
8xdegM8JgufPaO2zSr7wJQfRrE2abOC0fjMBJBAk8ttJze5KW1T9tTWC6uRoUShe
gEveVRKTesAzl2LgwRUNQTdHqlSXBwbXTfvLSqV5nzgA8gQupPNuCGNz6W2neRLX
FU4GlNrhBZN92XNKJXiZzr10nN8TMyjke5S0JFQAYTdcDLClu3MnuXN3RsEH49Yn
OEnGDWL76u+rx0sbHcjuFt3Sk1oWYOQNPOeTau95vt0n013VRv2+wk/7gHU8Sx/g
0grd2agUqid5Drz01Q+CiuCfgdEbKmdakfjZD7i8279uiP+EfsahpHvOTW4SYA3B
WRmCJixaT8/3XqgATZqsWRn0qPZQnEc/Cr1+2Xlq6+RQ5LZxhkOzKYBmBPl52Obv
Q09pQnWfYYbF9cJm9nCZNs4h1HNwkUe1EwEnqMoFEj/0lfhGOoFInssc76aM34ky
tahHj1aXB5fzZHdyFe3GIESAEblYUxyMRo+16uOX/FFlRhikbhTtyfCbxCkdC4Or
iAg+7h8vMe9fH1YHTwPd2YBN7s79bq9z0OJAGbDCmkOioYGhctQlC8ILs0Onggsr
Bt4C3m+82JcCCtuLml5J7wshW5hV5J67sog0B1xiYtanFmMI80w1vmnGTGCkmPvG
ij7WPdjWj9z0YscwNLz0nnEiE1dZkmRB9SR0ObgyOVZfkvyXefKaWrwlVNiHhHba
L762MKUTCM2sKD841mEIzuoFqpICmbPD6ZQMBUwUc3x3Ngwo2fHjiRBMi9fkyYo7
eATtjPXKvDtEjRhpSxTfmubZvwHAG8KcGHoBJygBtLoJe0juywAulhmI7rmxOE9q
W4JQdc9nGmbsieqTgeVwNBYuIlS7+JZBBRmlQJ2F0Wk6Ld7Kaa+qoTnxAsj3RZUO
Kit9lRA4Z4DGQtnLLUUW70s7EHdrwpVnENQYwW8I3A/HlAl/F6X9gWX1LkxroJ0l
ahYg5LRYWCEISawBeBRdD6c3JbrzpQn6ynNXykBkdfoRwBnoS4Zy8gGKD/uWb5Yl
UVnOGsI+3DW8Kgolg6+V+DNX0mQCRDmkws3B482Beio3N/3BXlxgs2sopVSNKXXB
hfNRHpLcgibAP3Lwbz/4S/kgloNo86/dUjcBR35zfcz5xwb7yu9hU0Y9o+Ml9QgY
9UzdAGaQX9Zub8UASlUn/Cfs/KsYZxPgVE3vLiGNFlDCFYMPxQ+k/SAl/JlcayjB
SzCAK412uYxO+AGvCLxdSNg9d/UcqjmU3d+6tT43dwF0SwCq8CrlnRDLNgoqeKPG
e9J0hO9thrOFLBX+33QxXy8Q2lb5/W9x/XXrF1MmCko5aH4dRWgqnjE6DJ9lvo5I
nYGp2ywg/ffsapEFg4zIdVesWhb8Oh5CoXMQ8haroYOQaOZhXw036jK18GP6EbsJ
Rr6oa6GGqb9Ass+GB28bimB0XzCbJzUbWoFrDOqvV3lrzYSIHglOZ5Chxcjaj7c4
rZiG/z9W9geRvLRrPqDR9ALlYdYwBHB8EF8SLN/7DxBsS9FRnd2EHxSden7VbSVR
RGwuFL7JmxF6onNi1LHUcI9S3/67ZKWo1d2/vBvpDyQufzqFvUzSkkO83f2WdfZk
zKjEV6du1vSOc4os+ih+10uduhCZNnEkv8sjsUNdNpJGqQEeLw09jTHqDwxK1qhg
ynrDQ4zcrjbKZ+GqDiSBd5jqFIuFMTZjKSA+ZIEuT7suxNRSLDCjGp/iYuKxN6et
m9QmlEfn3KhGtwvPnI91anS9Rbukx9xU3D1/wTIdZ4ZMr5SiX/bSd9T9cn+GdWAu
V65tbk116pOZOI6+Ggo5zManLy+GAmLUlPV0ljYya4X0DbMJOIKrZdDFE+Ef9Kri
gdya07VFrP8LflWnEyOnjg7xwLgN66qowsXyu1e9Z9WRcTum2+tpShMO70DdXiOI
0hagqnblAVsqIKXzfu3saYa0xaj/O9Mgr5+7rDWO75sEelN6SvqrjcK9um5nKXMD
9RvH4tAZle2eab68ZHn9SkZ4vixwHe5ga3QHstknPbCjb/o8kMiJML/2YsFHV7Lx
tQCOAssOdwkf0mnjXOZTOywehlduvPjk7oc6QfK+vFw9d9ZzftLhN6hzB6b4L+D9
c0BCV+4+MLFza5wky4eNRKARMtzzGFIAz+YZw+uP++o1Rv5Lzu18qHEmSnQ06pjJ
SnOhhnjjhe4//wRUIbrR893v2PjOKIT7CXiiDoVPnJEafALlu1zfAM9GWhltjMx3
UX3tuSviu3Xvt/Yahkpf/I6JHRcvIHtUkmFyFZXMsU7wEPSLmi7Jm/1FhEugEJsE
NRCMzYjjPTEIHdYN8kYp7dLm536pmYyFC2ZhMMs4Vbn9wvg7fGmzvMVfwXh55+ga
p+DAxpkCman8HDRhoLFKVMWXQXSoQmvC0pezJZ3k7zFzSj6L3YRzfBBfts2L/abd
uZlPDhjyv3JmY0+0bXdhzajV59F7sJ7CXiNKU/ZlFZrXiDa3sx46pOzq/7kWgOyx
RKzQTH6HTbssMuIc+VMd0at8aB+tQ7L8sVZ9GzAwYDb58TArQw9gipRG5hh3/bsu
0CDab5qKSDKqsBSheLq/Uj4OIP3S/Al7wLW1aTBpbmwLKsdKUS4e0CWcKh1MuBll
8tS7xf1Ip+mLpf+fTlLML1Oomuq/5k7imhwfCBwm8jsa4CvuWxdQTuy4N883CMJA
3/ywEBf6yH/D0+OyCD4B+Ta8j5mWbwMPTuAhecjcY+o1bJ3uLViViTULBO/G7rsz
XB5bIKIeFNlxnfg6AfmBH28Yzbjt3mfcpBEilaby/ZRIVDX1UPrDsID2aJkDVGfE
Sno9s4w/YJp5E1wsSl/j6NBAcpC/erpEAH8Nv4vw+El0+SfVeSW/io8oo1JW7XtG
iugeqEWFZ6Nw+wv+PtVOr+xeF0W7v8CmdJTNGaFaGOip1GsyT8hf7kBgAo3MMjG1
V79VVi1h8NWiLvBiH0hfEimEKvvnLeW59EQ8/8hoqWF720QTDkoRBAOxf/93QtIU
gxGimt4lSNfkpVyUHcZPFBR1+9/Hqd17Fz53ca0iukK63aDK9ctRACX2555oGwSe
C965cMAYlLQmcrySCybIl3ob3WgCmnVxvze1wh1armaW9TQRTGGROUKzuaWBe6As
wJCGPae0xOJu5O5za7lirl18n6Y8wzVfsMY4xJG5YcLdSODw5ROWPoYl69DDEOe7
kVBt0aN4K02SjBAeJts5Hkm4yTUoV1slhIyzKiLhckAcYysADM6g3k/knSg8fxN3
GWE317a6e01GKPUIy5eA/mukpkj0NT8WheuX8grkFupr+0XZMAq3VopwOVfEg4Rb
4XgZTyTbwFhUUfznHu16bDL0ziMehW+82/om38rx9i6aSEz9dUWTGCRq+cDrIea3
PlUAtdwfF//y5f2w6dz/HTDhSKQ5BnBGKISb4iuV5ggwcpli5V2KvgoRFswpnPmP
Rgp1WEVRUYUOu60xmYnZv15tP0n9TbDNr++AKtvLcBX7z4oJPJDnGXq1udubA5nx
0wBdSwD5YtPEADqtiBjwUoso30PMGJvJW8O2DGw60N+u13GWaWe7k5rRH9GTha5j
pilr5Ague3BMko/IkECKswrW4sLceAD17hdhVsDtPb9KeJdgEKpDgGSSDncy2CML
eZkK5wUM2czN0dzhDNJPlkEqiMDHp0jr4+yb5105nHNGwVe0bL+bxku4keOWLZCs
TZT3eUQO9/kwPlqPcVBznevLj7eoG9akbKUA8ttxQYCHcZZqzWfhpVPK4K3eaOPk
5M7C1C4vVAW6VPJQxABP3hvegWJOvDUi7j7BRoRuUpl1dObGrea1tBEQxWNnCZ+3
wOZ8YgBc6uPPLSvfG8FtVVaA8q6dvuKVN6LfPR5dKU2uwFMwwH5gBtEpaPzAxiil
kaczl1s1+xVklNP2vgKwlubCUYT8cIPX3b7rMYgtp+t+ogDQuahYVQ+pUv02kFhw
1rT4gpgigBxt1jQRACcuO+M7spdPLsfZfGxxOL9s1P10CgavVEwkpQlnM4kzr1Vy
KRsAtbWaJdPzFOJ1TiRHfBNlbZY8q4/ximp/5okU/h9UDdF5jy2k5x17akCBFJIj
wkXhKAN/RfeRVXxyv/kGoUOMzz6PqP6dQjUahteDUDfonWZ7jcZrTOPLD5YCv3qy
H6Jva+Lk9fxt7AD9WglrqwXVp6cZFkcRL709O3aZaYp3i3sdcZdmW3beN7fGyTN0
Kb+qeljmpTOdeOIR3KRnMN7WU9f8qpRkZ34xnWme/4p60uojZn065WS77icQXI5n
ofSVsQgIS2V3VPZUz2OsheBoGDDGx/em3jJGzHqyEVetyY0h+vJXMYM234zaCfDj
ezl7X6R964r2oC27ECZTVC3tl+QGtHDhl3kdJYwSZfEZ35/XI+aBooxB0r1PPjgA
dTSeuSCG3rUEai70HnY0LvPngv5Y4t6O+tLanIOrm/z0J4U5fNpQlXfx7TlsWZa+
zp9tGswUsBpIvg7iZaHJWRSmFxc9sLo08d7igPAt0QY0XTKS4JevhwE61s7tSbbH
smMGihM10FNgOMJhdJE4rERGKNh8nfmc2UFtxtHYdau3k89CzQXbk3QWwfM1fxJ9
AOlev/I4YPAn6Rd8Cx6KgtyYRrsQwO1f9a0b/gs3cl0VWk9W8yWUV3cte6noHCN0
AI6Fttuexwg75TWwjbNdfTgdkzJr4u40rD6igzG0M7riebis/aSy8ucHyx4s7Qt9
KbWXEjJDCZm5bs95cWrSc3GhlqqUHl0Gvn/raGvmWXhS2vBE0wZ0Wiq7XXtWj7+r
a3gk49lmS5ZpFhSHgn7B53gKvU9aXOkqsDq+Plhb0rEB8kIBfJeMiwd0mOg2cHmq
OkiqGuJN3HapjYVe4UVbgxsY+sLB6cDq58Fba9PkI3VvfqGDX4qJMEbtHu9U05Bl
bUEbvQBvpTrZQczz7ibp2W/ThPApLw/M2m8tx8Y/X6+e+Q2xP14iEVMqWSNqx/Ym
d8Tm7idqbmy5s+HTiNwSfnRCndQUuGExBXGZe727TmXwYf/6i0fExy6JjparXfx7
dKwrZaF5NDInDy/l4d0Da7wXV1/RK9+UT4NXE5HdDQrgx5qrtjx9b1PMFk+jGBbQ
RFoVIDh/bUW3iDgE4bz/ziBt48s2+Ie6n2VzVuwYIfkS+eub8LMzOiltgDizn02Q
EYcsmENFHOEuZH8iEZyAldMh0H35M/mJKzbrMEre2laJoQVaGuiKz/+V9SXtBaL1
ahquj1xq6AlXWUxyrq3gjOWJrwF4IdJijoYlfWZkSPZjnRW7xiGnxOXDpQQB/cVa
VQs0h2E31kn28UWrqBIUtSjFX6/jzH9frEqJVQCt8fPKMRX0Xi5VAaRyEhd1w1kj
RBRCbcByt/FSyVPgeiILSH5GyrKjdSd1X+EnEnHVbdEiY2Jxw7jlkAb5zkpuK0iD
whM2f2FfGivSWkJ+BznbkWB0CYZy4ZSFlYYrWgUoik3jUl39ZQbtWrpf0sz3gLAS
5F5jLFwgv44VjKXWcz9X1UrY5VFy8nX1v9l3cLcZE6dnElpnpOMncvH0jeOWRCzv
SuS0VMS/r3EcT/IO6iXfE08DBg4+scbMUuNAJ1xmNFEopUiSu75g1OYBHIFICtvE
HQmXFMGJW3q5/JLJsDiV47BNVAQKHqKIVpkDsLnstvIUaofRIMgMtnY6RYuo3VBC
iTBArb3BaDeU8YXLWJaHpqxAHgSKJZ0sgtTFaQdAs03cBAPfxqL4IAKUoeQuW9Lo
EwlOI6RsPZXjwctr9eg+SuXkQjj7Z9KtH1kJ1QIH5kmEH8V76e2q5jpD/4z8RG8g
JmQwUVrzSsV+dehTbrpGqWheu6ksSDywSHJE4nt8hjmik2rbPxiRIsB1FbukYR3n
7oMg2E+IspkZpsfllVMLscvpZBm/uo4o+kDmW13o3/4XXBrxSQFEB0g5yt3oefYd
LxcG9bSnjDnA1dPoPZ7Eyq4nxoO6uoctYVcdW1bQ3hvIdiTTtC5duONYqz0Y/j40
k8F2mXM8Z3gWFoouB5vF0iH/iKnwpPyEnKgpCLY/wmfMA8nfvRqdnaTKgBh/T0DN
pPB7bgpDYfkTgj0H3fBq1CjQqaYE/OZrSxFI0Rxn+Q1tT6NFnkKjrLZtXLuQpWsZ
tFQx+wq5K/4cu8zerCWfqHSgFw9SS78Kf2mGxH7/BVFM/D45qL5tL//x4/C3sabz
n+CWNvnQqseiYEbWrzq30oGngc17RSaPn9PHYmgzjfhRu1rO1AdvqnxHAaLuaVIw
tj5zvQCJgFtSZAhJAUMIbk9O1K2c7EULU/GfcFz7XC8+5vVq1QBtWDcVwSu13de5
P13M0GxN/H1wYQMLpjcLdL33cQjioxGf64jNkk6RvdpQLDLYkn8q6U9Izzqiv/oY
2YL+L3vLzbMrUBBHAM1xnM1ICiZVdMjflMNDmwbfR6Mb+eEo5lJSwUTou2UiqO+c
plu+s+4Hvp8tFS/SHo/neIMgC4spYs4SJmps6X/EmF1K6RqswXY1xgK8mRRPe6FJ
qG6eacU3gctYdTrJavUz8EA+X3vhEZt8ulvOcxd9qR/hwzWlKHQmvU/XPYTrrCNI
1zUfmIT22zn7YCvyK9QT5FF6yb1GdsU4Xz7EaO1DWJPAs09vqmLJw/XcRX1In03+
xVtYjwIo3An1VAk2q95QwQ/cMEFvJgLfXOSb87BK7cRQV4S/fJTuVSGad+9f29jP
rXigkqMGZKcwXK9zYppWx8biZVM2yenZ6aQBJFacmdeaLmg0BcbxljoO8zYO0eOx
DidKxt1Jc2kk8dYAn1neGL8+CspHur636wd0QRRw168BZj8X0XYKOCAOJpyShzN6
XdDr0AG3gDhlkHcFDzXsEjvFV5FTA369W/IKLM+tWDjNQOROQPdUC2f4lWGPF+32
WwITZKVKq+hs4X9bYYbyLwNww0/5AFsUnO1lA6FcYhEX/CYuxyP/IkGKbHXOxdVI
K6WMvKW6T9pPpcSbBmyqBk46UP/a1N3RQ9kTrjzNQvAhxNwtaqEqPXhGqac3f0Ex
KGYH/ynrfcgxebCOwg4fv9sUysSJQG23sy86EUO0ndrp1NlRJr3hDCw1w38u+wmE
j0i4TZ61PqL7HNXy2LkykVvOaLLljMU4YkDZ2SlWj4VcumrsWC+gRlFKq9t5Ejq+
GrI0YFUL0u3t/4xxrsmFtyDRn/TqyhK8rNetw83+KtB1s9scEuBhnwOtGJ+47DXV
5dqhRZ6w5bS+9mS6NvObqymdhF9vwSkdNSMLhLYs9frA9E7GFlKewaZHNdEuEgP+
nD90l2Ou2Hsf2b3V7Sdlp4oikOUCZSux2etMF+QzvGwOpm88P9PjwTBKgrHKlm57
8ykuSxTNqfZBgIi2QvntPj/hQgrLG/5dD6j9K8XzNa4qa1v7C8s0VEHwus+8jL+Z
a2+tvZ6nRsVxJdBPPScMh4FVUWDckCQyRu5CrziADvW2oKpa0lHynqsEh4AUyiLK
g8Rf11CCBYKpoD6GrWi/Mv/aLsiF53tXyXlkJYZHBdXRUrrtxKaH0C0epEl/G7Vz
LY5weBe1exElD9LUxEFolNXfpzOPvO39BaeRFaWTT2xPPDPOg38CeotEcyvBRnAW
LjulO+ypyxJ2nRIKXDLhZp3WoqRURAwnRfFvpNstsk2X5XCNm/2KgTtJZiH0AA9o
AfPAdLueD6/HwmKehMNtiZHOi1/MKZh1CJ596yAv90mFrcARNYdUxiLtb1HRv1K7
kDY4gHt7aTYMm8Gp9HEuwmg5TXHGsjY29rLBOQT+7z5miwweyiyFlOFWfwat/E/Z
ANS/O8IXtZWKxxiw9RogjCxTljorhrbXvZmYPYQTV+kIyCZFsdwiKtGBfyVCC326
NatH/iiIY++DkJLCs9yihNuq8sx3pW59E9yorvIEpOb86t8Ktesk9lVCWbwgaojm
Qrvr9p3r0YABp4SSXXQfrY1pQm1s/ME8bajyQ0jCb7DeOXCXKj9zWSQPvGcNrFEE
OFkbKsMBmW2chZ9x7HEpczXksw31BENL4ieH0M377ddct5Y1bj/nYUtOkjXw/7pK
bhGa7gT4+wdk/Fc6zUcj2/pVQ9g1r4lp2UoLyfHTfcb/iLxJnezGMsFFDR//tMu5
`protect END_PROTECTED
