`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VRqZGFNySQeBnbDaoDTQfhAbHrbw0gXm9HFpkDZdQbKlNtj8xEFXPxyKMKMy1a4
FEedz9zNsxz+lyZnq0G+enDFHF169Vc/RHvd2lszx1RBe5g90yKp/CX3ORJLJv1p
pYASbXj6YGtAmrDBoEmTBuVjAwJVrQDEVBbnxTDDeaoH1vte+bU1LZt3Qo8m8sRd
s8uw8g0R3fmKOmKDFsVZ6UFDn1zGgpyMY6iM/vhSOV29jIirHnaZfXCO27d6d2fo
K/DUwpTiRx7eW4TpeQnwBgciPxMKG+4CrVdE9dvS0kJGY1CaVohJmEYtboWHnLpF
WbOqORnL5F+9gTdabq6DtK1oe2UqoR3Y21VDOE/QtqctqTWS65URR2PAGBlkDGKs
M/WS0vw3Nhj40HDSeoWTg0xU3FV4oTeK1cmQfNEbN7KL6jtj1uk23y8T4B/dVUcP
PDG4qNVnuECwwRe4ntY3x/pwmfTjRGkDZid6TomplNoBZbenp1F1qoWiQqUTG4qq
emB82In0tQS8fFp1HtLmPjiGonvJyaCqtmRJt6CP9u8iXWdpzLwLjY79HXxlu3gJ
HE7ZefD96FGV7r3n3GOzQfVYwSVfru+kcSQe5XZ4ZaJVE3H+EAFprSOln8f5I/Xf
OWAe6WcGp/1UxQMCjExVrg==
`protect END_PROTECTED
