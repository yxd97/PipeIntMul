`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v+Kc8pJYF7QLSPPSxzPKWL6JfR52DXNH2bwAKqOxQABuYeywZXVfO27PnFd7nhJx
JOlvEiDFK90xNntLynhzmfK6pKkSm+jJkjMmbkuw8j0b97HOf/s9MHTtUEE62Y1K
/E/bNuHHNVLGMtpM0c/7Do11caWyouGn/5sN51gBE8Fdt6KcVa+yH9eJ65xS/4A0
TieG2zeaUnofJByAAgu4dAg5ebUoYT8q0aWXOnM784XLKfpl1Cf46d7KxMm6gSky
slJyyWgbMmXbLkVQPetp1Gb2B8OPmni8RfyEZusG5LA7jU4Mt36LIb38xiMMCXFJ
`protect END_PROTECTED
