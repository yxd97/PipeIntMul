`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9yuK/42mNSOdPD5pTRn2jM/ara0r1H1NippGigrwUZZd33UFF7OeSr4mn+5S4Y07
mb0eGp3Ov5vV//jabyCILJNesd5p9fBnYXVnLiYYM+LDmU2FP4LhoyKtm+vg0s7j
hIQ5KP8ySYj1L7GCSKT5Va4KIA3xpExfajZVFsR2fIJOrUgK7wgJP1/wWCcJz81H
WNUlhijPlGBVR8gBYV8wdcZpL/ThE6xDl01PKdE907oG/ra+m2efJrChhksF5RPu
FJCet5DXq+Hcm5HGN42ky4wrVbBkFCRuF0FP7ORAkw3w5m85nMFo0sqQbaZ0jRxu
HKEz79wIaBqNMRs1eqvaQN5Lc5zDtTtvUDBcmtxa1efzOT8MltM+VP4cPwa5JkZ1
BCZFz3BMGoAM09g1EGf5ibdceWc5l73AvBC5vvHytE4ik9Wr0ANm0ToWpEWW70pT
sllRgv39ogF0pHbewIME1Hgvw9OMNRl4nsqppHNwOegpTwDenHv7NPa+1MGfGPxM
BU7En3ae222KDfmtWj5yFuS/J3pW1hmZXHv8wEWQ8OFk4WcdQEMWO6RroS9eecoD
ibfVQ1IBuQPPoZgUcScSomHGWQBkmOFvWtRseNzrdtKh5k71tb4xVNyr5dhND3J2
+c4tUD32MBHrPfgoWPnHMA==
`protect END_PROTECTED
