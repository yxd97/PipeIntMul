`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGZpkuWKz3HW2EHnJeqoPGAztwHeRgQzn0KRmEJiG9JncfCR3UD6gyYaOHFbu8TS
0JkPzewjaFCCfWe75W+0jGkxcY2qgr+6tLtLqeqc40FrsnCpj+zB2LoS8WVlySvm
ACD5j9B9I2iRnS2ZiRvoxbx2zondlkjoIedzf49kegPKFlqlIxeOVjUI0Z1kH+5t
mhX3Bno0uGzbKsXgN9mXIf/eR+rPxinHwJu9E6qLEaZRIf7ORNX58VXbEUGEpT9+
Q/youyjTySZltyBvB2o/ew==
`protect END_PROTECTED
