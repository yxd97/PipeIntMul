`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YDhTdXEqRn1iBj6hKr54P3IN9U8fScATwpeg0SWP68W/0vyS17tQyn789EVyr0nd
UqNAV8D+QY7RSS+YcS828vR5MvYsnYKSaOoJAsGFSIPme3rS+nt4cvoX+vsiygUL
XG5Rfq3jxIeynWmrjoYQS7C3BUWaMa+xSDrT0GN46UAuvAHZ/nZuXS11BZVK1xsn
J9V/A98e0FgteJ2NqBBqQiwHBVbVCgyMzwqtZ1Lfxq5tUCRGF7jL3B86WWwwuQDk
9HW1j8EzgsTfbvdTvYc/v1HVcZKX1HEhUaIy22db+ueg4xBA6xAfFhrz40d+jIn7
iILzB/jF8psscuJSM/BVKg/8q04wmXXajHrJy3hR++Xi0/gQTlt4NLLGf17JyKlx
AEkiprifZSFT4DAaHFRVAYKyxW3c6FcD60uZE1JzoYcqjbGTIpAMRPf2QeJNnEvr
3g+WYr2B3fhNvYKFrZUfzoHiO93x2Pw0LPNEiUrFYYRUQlGNRX9Cxd2t/lN7TEom
ut91d6DJz14o0N3Qfv9VkrY7wYAiZ+FKflu1Daupvb5t7y4bqPK55L103FZhUrtM
k/M8JGzBGATK9JFGDaQQ0o83TdHj/tlCeD4MDMnl4XaKDVKfJAzEytJAUrjKcZTZ
bBRcw61LnZ0f72DRZI+MpFLDHSgsQSfoOyRif8qoy+Thy6y6LuAwGdr1GWFQ9LnN
rfgDHmY0x0rb3yUcGSiF5oQY0dy1xLFDeokW6CxT8oY66rZKrjUQ1EDszM1tKvTQ
hVDuuysoTwe6/HtlJtKShOJVambehD1rLogRoHNKT3ZvlYVxoERmQbFOi/rCkLO5
9DTlFar/iOwWH3MdpKt1UanLqiU/ZlnGH5nmqpZGw2QnJ2fpbo2syYyPSawq4PMn
UUAEngq+PZABKvGaZ9LsGmGz/jk1AKrBnx9gtuUDuUciOwPcuvt9Id8YuZmqzMWs
c37MN2Gc9cfg5daPxcdnVvN3V5RrkuIwLvLXBSX9sstPcAEIDBZdiBPmR8CmHRdb
CVe/DOT8jMzyZssSt39ICA==
`protect END_PROTECTED
