`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
880WYFBkDP7+QOUzPZeXkf/aZEnwbiUCw29VnjVI36vp9CacsQPtQh3KINRQ9o6y
zI+UXXZjWvO7cU5KXyzhSS/SAztqgc6ThYHVMD0jJwIcr/bZOUAO4nz/aa0RakSS
pNIuVGbmlhYHK8DVSQ/naRH6evAi0KSD2odfXqW/kt0EJ9/PeguNjX5sG+Lmp1LE
jAwcfbxYrrr29+81rv8oYgxQfOK66trWECqEPcdMJvNbYA4KC23TTiEqiXgrsT9X
rQUef3TZszj+k1rD1/Hk9rzmFZMrM0XOcGQa/A3Met8jrW7+L/eyaq3d+4/eQq00
E593G9S+gf83i6+o8iIppIkD6pISichbVePoQnl44Nm3fl9jrEYW6k2F9k5fn/1H
mWfNDy+JHQ/R6dDrXSNovo6r9zmknO0eKmjuZkmR4XnjEb9cKY6qFSLTQwD7IDzE
xvXAAgMAXANB3ZrHHOFBd0zXRGKuJ87jry0Ssb3fxmQugUW2lT1iv5pm2rtHIs7W
8BXbDGPXFlephx6seJ7Z1J+V4ZACZ3pUn4KlGJhpOuUNL9Pq3WXoAZ1BcU6HZIUv
nQC6LtNk1fY1tNJ+Nl0TjA==
`protect END_PROTECTED
