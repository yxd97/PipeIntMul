`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjK6LeJG0hRYxpCWSa7dEQeDZ2IU7eZKmcLm7F1uWmqFky+ptJ7D9XAnBMc3cRJV
akeuIPwsjcIuKDBpPlSz4PwvxjLajBqMP9EDSt2HvRSmWZBa09hoNgBn/BpkRqKX
X3C/vq8L7ot/A9hs6HiDOouLQbMffCrt5csnYSYOInatXYWxvP3ScysnfG6mwGjf
l99wdyk2gMijFWzT7lH1tTgh9P3tPUPnO+2+Na05ujzbJ7cH7m2vyfS87mQTHnsW
hEVOHhgcCVNU0HmHiYYODIRSzT6eOOx8ynBue/OMLE+PBJypSi9BKAuJfbIu0R0O
UzolmgI0ZyyuIH/1BEoXeV1s1MYZE+19h4D7m/lFnrJU5ysbpMBlzpOVjYKOyma0
dCTxluNDE7BJHq+aOz4gKAN3tQlH06QcnNbxkkEvN3TbGAUHRgdEvg5HDMPwyvEd
pNpZYBW0I+aH83a/aouunmLozNyvLL1W698ZmD8eKDBWXlxRcPSuZ3Bbi06LUwOV
`protect END_PROTECTED
