`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XKRwWdHn/Uosoul4g+mNoTHi1lzDfzPk3FnI+aY2ZWXNUrq8mc3OhVf4Oqb9kLlb
H7fBPH+gIYHKnCI0J+dmwf306FzRRq5pZ3qEERQl3RPUZK4idsGEM0WzLwBzyEqv
+4HzIgafFKeZJWebcJNEuy9dMBPdJoPVGcI+lgUVP8y9ybLWU7cLt+Wx5kmOI51Y
YdfAEShM29bA0gy1KZB5EWNsM6qyKgEpiMh16PxMj900wJ5OI6u567toETtHjGo6
A0cTmjh/4NgQJYOG/asX+NMRJpR3tt/OSSJ7J1zhTIyuNebLnewR8pWUDYe/KglD
zJZIWivDV12z+MKGoJFeUrAo2e3y7OR3KVaBmvUUFki6sySQSOBJiw/mPeKkaTyq
NIioDc9TDzYqbtXq6r+M5VSh6Ao7a42ZQqPj+c9+6kkIdYq/ePVttkcY9WGGbj82
PcvAC7u1qlAx52bPZ1UN30YG/z/EzPBBfqnxZ0nPAftF6tvqR2iyCxhumFQx8WZ+
m2ABfNN69I73kubeyIO/KvXfmnycrWOw7H/cb9pjH6YUtLfwDMcu92eIdh8kLCv+
y5oJ03G4PS/FAQRIBvr3LJk6Um1XJrHBJGVYvb7+FSjdhAtYFDpoKxKMrmi8MHYj
9Llrod9h/QhRCd9jjxbl0pn/tnzxn8c/V3Rfa5a4Ru0=
`protect END_PROTECTED
