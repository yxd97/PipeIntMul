`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMZr3qzlh+v+wLlguK1Zy/MyUf5OneI23yGxNEVfQ3QSenGLINwy50T9HOAXGYUX
rZS3+Q94P8eyS7QPVcJ5o88u4EXWQYkIUsjjHr+oS1BxhjRLSxyQnS0no8VVZR7K
+inb3f9IBQ5KYa4Ne2VP+DtzD49ZHJ03zXU1FnJ89937Cd21SzjsMqTxhb79XGVl
fLkavBwt+b6LBZ05VcMGzabAEW17J/YEtxwD53zzn8Oa0DdC11iQs1jZo32H2BPQ
Xr4odEvC0/voga5eO+hjlB1m45BVd0fn/7gKQc+HpBJLXJld4Q5fxJ2UY9QAkjOO
3YWKhJiO08wPd3BeFnNPX9DDbcrb7KkUAvTT7HZB/1GyEITEOC04iE5eQ7uwUSDF
Ve8E4HjuGpBLBUwEIAKT5UqsHkF0IT/aBWc5GprvGvRqt94BnjDNbtYdEjDbReQt
31PMAA8C7VB0SfcdjtJLSi2FP9h/IPDIiBIXzeM3uBnCWG8/bcGCp6URleAh7rN4
C+4FoV4Du+sBQyyE6VnIkMhFWfkkD8lu10Yb+I9sF47mfYxzZeaVQQtoVexz3bvT
0nYHDNlHSl8U6JQ7anvsS3yBdkv4R9ZVAOStt3jDCHwaeJBKheddeu0JjRGbqkV/
p4/v1A/aYtC2/aTV9bNe7jXrgE9yyU7ZyF6p1kd2Gcb2e1AEIW3h5FBMa/IT3wk4
MRiDnOVIsQr2EWdzl2a/i6eiPxnAfxTzA7aMxTsgpuuz9HJImrZY4u5cfxJizNJn
TC2wYaUGYE0xduiMIx5IUN9nJUujfCRJdNRIN4RTPZk9UCMhBKc86FYZgV3lxL9m
mqZ+zIB3O9q+XWHKYewZ2xyDZ91DY5Sb06Fg1gL70TA10bXY0W/mQSytDlfK1MUV
RwA2SMUJbVTDPtEE8zBKNH8gjLx7eT3YCEaQ2lqKehi8sOFPaCcKQZKq62fZQCOV
qKL8514kGs7+qS0qTjxbxlYy9jnwQxVZz0boTsoWKXHAkQbXUc7bDCjG8vM1957C
A8+ginxLrSqJ6NiE4CeFadkGcsj9d1U6p6Dp1eo4L+VJbpcEvGK/Ic7cYYWXpKVb
avSERSe+wGiVZ7bQ7ufEDEJrlLg2XjdsYSJduC6ppHymrK/BDrNcHEWJn3w1GLkT
dPlGu1nxDflyb7rM/6PXwPZKsdNPGBDNPv6rt+qmf2Fk1y514FNkHK8K+Fs+wbQo
a10+8rze/Y7HsRjTe9PyBSqIe72K17ecgKYpnZszSggkZMtFetQzretI2pIWTGZ2
SwF0rnKJC8kSLSuAZBmDlefhJcUiDW7imsn6wfB0IdREb5pqOgX068DUengSj9fP
CV7vwE9HLil4kAiZWorQSvPTaphQiLKZBV9efjZlKiROw/e71LfImUyVM3tbkQtx
ZmKjph3oUvS267PE0syqId4DxmkNisa/l8pnMcJDss3W2Iz6S7v+nre5By8Kn8AU
KIzciO/tsJYqijf2H4EdeVksjUgSYoUH7owAXpHtCbjyQArpV1JOr5P9Da31Plhf
yh2mvaDtSQafWE1mvMMb7pVU/scGumkQ4oI8Grkryo4ZqbJyQH9Zrr8FVVxd5fRh
1pcvUGsv3EN7+/lefjspAjrWAnSiFh/Bkvw3L2Pxfb5NCQIz1Zzhx4JbjL6Horru
MYFrWw/y0xKFXnu056UXfQS9KWMVJlmsxIKXVNaTtXB4jBg+NKjjDVwZwlN8e8j9
YpQn+UbexddgWhHuMt7Exk3B11tUWglQWeBXj8d8VjY=
`protect END_PROTECTED
