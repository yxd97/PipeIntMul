`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iZHtfJootVNpn5YBeRMtuuOT8cER2REXKsXctE2vtFlzUtOlD7sftjax8k1IjYW
U3ZNA6E7Bd4ovvITlTRsu02P0xRjT0UAHO89EvvMgSTWNp3GEQqQG83AlP05cg2U
7WCBL2raFyQ/tgwc6Hs0UTwiHLcpSgkRvx3eDtKq8gXE2uhJU6+Vxfs+VLiXuzIe
ZwfVsqlPcIH6zIiIg6KpJ9FTUhdD33TRRyU1ABduVOPz6HkltzgtgbjGy1lHXJ5g
BFyCNdlexVCtVjWDbaBkuX5RrRoqHVdl53jEA19iDWDjclq+ISmi+RdynLhKi/Ib
`protect END_PROTECTED
