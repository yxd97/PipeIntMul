`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bl5Enu/s8l2jtvzLgoeuO3C/Rh4Kiqkq4laUs+4cdJNAg/2wE/JWWIKpA2wxiLwm
awvRIaHF4fdc19c4d40l2J4MiYVzcjLnQLSSp4PRFR31azVTuI4Li4de/zAHH1G+
eixfWIWRprXnfpo9QTGuS0nd9a8IavzVuJ+a3ZiMQGEwfTmPFCKkY9YWYHGPW0Wo
AR9aycdLCibhwU2oRZVRRVdT0sPZ1jlK2mf7hJMhXKfnNUEcRtElxPoim5ejtT38
Tm3CaaV5z/mPN5qeEJop27eF8GUfvLfLMeiF7oLgYlw=
`protect END_PROTECTED
