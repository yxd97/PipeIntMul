`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J3vCnsRBH+bccT7wK6Znx7yWQpHdoOmwyv8ZaLtpYCxClwufdVQoH/9kIhKQzvMU
6yx0drNqGi1Sg4yURF8zXu5k2KhG6oFSbwHhtGPMYd0iZNX1yBT+FNV4tIbiLhO2
kwJPCFjjm1prp/ODLlKjNp1nPsaKBju9tcBWgMRiMZpzezusAGAWfYgA9WFrG6ns
ufbyfDbukm5AKdnccBLGWXnlkiBCv91LYwRbHDuoiP6PoPiWU1tGTx2ZEzh/eC2f
hVPYOjYzb0he1LC6cdk3QktJkjuKAzUMWv6VeP1KbFozLuSu+6AJKqK4PlIFDirQ
wuEINi/moKU5kyFkUYD58uJBjxyYV+5yw7sgtINj7O9f9kHn7zjmRn566gdVDDQ6
d+6shO2KP32WeEu5UKobeWt5sC2zBYSleU5NBfKmfxnISAZLzDTR50DXARs8JIek
`protect END_PROTECTED
