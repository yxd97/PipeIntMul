`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KlbyAuWIM3GF2FG4ksDNghFhwH7YbivE/z3uRkunKfTuWa9rhF1h1UkbqMwrkant
avXrXVIGvIfEErF1Cdn8FVCOcDyMp1bunRmhzlYP7SAPU3Sxx7WPimHXVFa/I6an
NsutRZVxFW7aKMQTzcgTGh5AOKPtBOccTRr4DAT6BOq3sTEPfvfmW/IKriiQ5clL
DsRvqmF3wyFJU3WmhMoq9KaMhMUbFg59K438Wn4F2IP7U86ERqhomEvo0TDakVCQ
RjZwyCIU9AUyRdPiimxdjcQIBVhb9p5Oo5WLV73+L7zBBpG8fqG4pz2K3GX9R4RZ
Zqcndc//8w3OfAnQZmltzTOvu6tuuTxX+Ar8JQjz8GGb215jvOmkchNGmCed0r2W
vqx+z88esb5IGTCcbquXuA==
`protect END_PROTECTED
