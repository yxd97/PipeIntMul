`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1trHDF9ZQC6zJQswV+eUkV+2UceQYmJ98zaI15SYfdxU9pdgGwiVyA6mFKCrLG9
/jh7OSk8NozjIzqY3mYeRhGwSdcA8+uUIDIrQoMrXpEdTrR2sp/EFuYqSA+CHarw
RDE5RjO5qV0KKfLT/jv7RB13feh6k9al3Kzjqc4W509YIu+acU/kcsoZH02bC8Hs
VzVHEKi+6Y5N+Ppk4pjzm2rzhm58jN2eEvF3gOax0UGVb1htHFdSOFGKvWryW9Vp
QVHHWOLiVeY132AIB0UGwI2938oI7lRG+F39CUa/DvJqnhpY2MgDHKtzg5wOaw6W
S081qiEYmEvi+miw6EyeFk8v4vDLGY+PR3PHmkFynrdPOhlCX/ACBAosbH1Us41f
Paw7CYvx+ediwOWnInvMSW/PCvdjLHHBJt8vNAsEvg26tEgEw2iHDjl+HVlxkvsZ
`protect END_PROTECTED
