`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vZ9GKIhFrVSJOpcSeCqHpwpWwLRu3Ic9l77TVTPSeb9nJgY3mLJZgkORPe5EZtuq
I2Tcml8DRYkQDLOipzfaVwWX45yF0bvZEG2rR9KFoWTkz6IyCUMKAVp0jsHxOtY7
iM18Z4oKt2YyquDWaJfd7euV2W+lARyhNA+YA3rOKXv2p7V30TpylLqcdXSjMGVi
gK2c2KSRT7GGt+TumPjF7n6g/FdEouQmkMfYKRuhDxAO2nR2avfmvoEiNldXYDum
6VH2BqbsCF3+1E7TpNO4HZxvpb4q82CQw8YZ0VGtg5iohV1D5AqlBiTi+A1EJ4gE
+5huoUQKTMpsTCCI/MgHWQ==
`protect END_PROTECTED
