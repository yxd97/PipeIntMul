`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTNqC4mPQalaqg45LOX6NDeMECRF76gVLISTfeEFIFkMOdnwovAN5dW6RHrAX/II
x8X0yo/88LMCzUParazJce+OGOcQU7xPxamLj36zU/SDCgzDcgrgJEjZTMKXHS87
sT5T/RtXLJRz3F4mcaGhdoqMZiEHGubIFjo+xJw6oTZMhHishVR78VAB0Y1BCEkK
Z0jkxI8zyYzADKlR1myoc4Myf8ThecWmfOvYLWBw7Cuv3UZQiexyUNyMQagt9yfV
+ye+scYVdtY5bhl5cal9qLge0ZojGvcD64/BoUFjzJMrfZe98VwpGjwBY+J1YOS9
WKhDB/HTQCvECOxCknG4F3oKblWH3GCYr29TTObcD7dhRf+vr8WpWCj+K5MrARrb
eCsYfrBHvyKLjjiCyx7q3JmcbSC4Bo55Bo1EmrdFcG+b3PBfNzClSwfV8Tr5b22P
JbpNYaxl4UQnAt0Aeb8Zspm0JTgpS1QrUHr2MrsmANUq4Ri88F3FKw7sPUUlFbXQ
ztfTCc/j67ZVK3E3Vs/CfOVwatFm1naOnJYdR5D52O97ipjL9BiOfPWdnKv/T0Qu
nb6OjDEjD7cwcojaP6DnJyID3HzZbfXHN4Fl3MYWZPZwLtUasG1VyeNPll4Tp3By
TvDItKOL9734FzYxfo9vmSIg3EA3EgXjOCjQzQ3RSiMDYr20+X/FkXmn6BMV0o15
dXI4IrAQe61FsyYWjff9VkYCgDyV/uk8hvmLR1mxBPnOzv8vhKSeUwRoevxHSAQO
cc8ey0w2WXHyaFiybWSWhMcgBSMR0KINKJWyN+aG7myAUG3mb+5kvWicnXgw2tdW
G4TYZeeN90+ilk/8eZpKWDE5WGBTFwXhB2N6RucozW/kYlLgOJUSwQ1gK35jfy3F
DiW2YO53p5/eMar1atl5PjaPH0zoAACgK7kQUR2aExTZ/pLQyljmt106kiyrJ0EQ
bqOOD4jXzXqvUmbC7zW0MYPB36IVatVTqGry0xF524Qkt4pCSvHqkQnXmFuYyfeH
gnSQNwLs/BhKdmoosk+gyLfm/PuBqQ6oz5/m74qPKTrSQm4Ncv+aMhWcIDED5mbi
okSjahc27P1RpDT9DF+BVQd7UX6C/wxr0FDHhXk3jcTNFcjM3TdxjPO3c28AK7dE
ROdD6BNuG37xE2qCF5dcXQkqn//3026zdRAaDCX8F5bMiEtenik0mB9Ee45B5D3v
s8BXJwSctW7bGz9g90VJ2HbTqzBY/HwBSG5IB4dHYzhstOBoB4e3dr55+a7kbWEN
aChwtxeMmSDPZJE14gXt3sldH6NgZA43HQA0n1v1FTbHKt/n1cvpXatK8f2iuIFd
WJqsGvFcFcysY6maEaOTSwf2CURllNLP0tFHwVCTfmIpJqfdKZ726jBBXR1umY/j
JLQ1bvgWQUwtGAJojpFFU+uVJeUcZekmoLZNbhyFv+4Y1Xggq1O2Tnvse+zM5jqz
u7vAwPxJIgf1CY0nvvR3jGceUKn6Z+JVXbQWkCdtyhOb2l5I0k6e397ex4buCwdA
qfh6LwQrbOTlRu/DO0JtwzmtFujS1x1nkIqE++34zAaGDhWMFCdrww7oMd5hP3o5
oT8NPNng11QFm1sU3goaFGv6ZDVTZplme+uwE8hEVAcd+vEkvYekPcHOCapbK/02
x3t/uh4WXkPfG9Ptztf6vvUkE28ErfQmY5S4LI07sUamaLRVsGvFZGKd5nHC4dv5
zNPUna1PPutN6KUC8KN9ew6TTosbX9SYRaWnfKymmCDZxIM+v50mBxt7GR4zCjDa
8vZkh2x58rt2R6UpLgRTHkoLJEK6kRBqdJ1523Jv3RBl0Ese0dsLXX+ARuvZhFGe
VMksIS38Fdj+qP7kBbxg1AxfgUGFXyaJ+3WSNv+Oo8UsQNC9+qZOAx0ndilF+wjb
8kP8f20uFFYzyX/4GMjb8dK4ZOpI1to4oocFrauHeGKQME2Mm1QylKxu9r8vCEf3
eO+BIC7VR7YUrGD8+uhcwWZdIF3VCqxttDuQndO2SXoQCGV8bbebf5RSMnMr6NaA
m125RewMkjj+vXYZEr4YDq+EN1liaGM17xYz5Wgevdqukbn/N7xZ/DOAysmZQmn9
pjBftnAPlAZalKpWqr1zTOrlaZFOso7ttEtIIgqOGcRJRlG43UpO/cJ5Nl+km/oR
1ycCuEulhFCLyhsFJLUgJnlmolqjI/548BZl++Yp5Ci9TQNjWZgL9gWhiAZ5wdnf
XcYJbSKQ5pGAr5ae0M5xs/HBAnp2FJtCMa6iYaSkiIzKwwlKqN/K1J98rMshhyvZ
t3R07yTMb9ZzWgqy1zZClaFPcA9yASdp9NSZ2kfIt3OUxrzkHdILY8Cbk2N6O/is
R/z+aL0WTvrRUSyPVr3H2M13AayDxYYRC/nFHO7atjDp6tBBzhy510q/uNi5lGFU
Iz3oEM5wwK7TtqWbA3Vay+m4WPYgysaDLTq1z13Efvm5Qn4AXfblBI56wUWWJE7k
Z0VSTX5H3VZnBab69djsNP8UYQMoBWvL3dncev+gc41RxQVxAng46KN96QB0o9ea
9AdRnlWeHDABjbj1BW4UmrkPb66tHCq57B2Tjioq6UJhWU/z5u03PBzJGOCb75LL
VyZySFT2ixNDHCT03OMmFnr/ywj/8Qw2alm4J82GxjA/5xE9e3dIoKSh40qbQK1Y
96xpgNHsX5I7WgPgcsB5APTQyrR4NCHpDvXuLcFKXLpVNR5BItnAsfdWBzn3/3Sh
HcTsEqOFauBSUD7T5zrs1U6q68dBfhmwYqyvy+zpzW0zlsl1CXZZWNNoUd0M8M7j
kpoCwYtfr9FHd63DRwlLvesIfv2ghlaSGWq8djlLl88K1dVKle69c1x2YubBAqV5
rfzZcMd8ekSictHCwM3xQLM6VyG5E/IWG5MQStkl2N4ImmKf5988JAgOy0BXchiJ
VvCIo7n+66y5zI5EIfv2iGjc/hQf0u49+HESovyKmABOffvTfsvpq2bZGRJALYUp
UIe1i/LA3kFWF+prEAU+wPSZ5TGu/jm6EIgXe7rktbxOpss5X+MmI1mkJLn5dxP1
7WlCcHQGDzYNXTUZ9OvWRDk/L0UmUMJmYW9DipolgzurqhJMPzVzcT5XFZQBhmSE
Lot7Ps0NzdHO6M6mNyGaEBkgNkCiei0c59tc8o6VBq0ov8TEPA+r0xAm1z6SbFNw
B0oCXjbt87aTQUxCHatn1yM8nVrhiwssGNq+PhpCA1LBYL/1TjsId7ueULqGdSrf
RHdqA48hWW1sAIPe89rtT2QGUlNotSQROWRDkm87VMrVXG0olzKFEvsS40O5+uAW
VSXaOfN7+qzttOMinPAu+XOjkA4adewef+JwFZEBMWKlnSk5d4HCNtjI5CU38P57
mgp/RimgWySm/tlTourbt9XiLITKUkc7vUusA3o2ciNiaq1hznUvYdQk9ay5Ok3n
u2tOTGr/BXbcLmMLJhFyOIjGwOcYAjg1xbJ29bsk52TU+1my5jI8oFBxLCfiICgu
Xe2uyRLQqtKnyPzlI2J3+N0x1x7scBXoypgJ2f2fqQd8dbrougL6Ioc9PgZomhKU
JSSsz4hFqymwschVlRF0leHvQ5lE1z6JTEFfmr0psPdIcYjs5OcnGbQF/6zSNjGH
A4ajZMxDRrCgeAzl2p7FXp6OeIp8cHSt4aelOjGJbZ61Rh7Pgt1+6WSPFKIpqq07
MKxtIsun3BdXBGoNn/HtGk8bKXGns8oEAWy6g6+PPnGZebuIkauWadx3fJvPEAbu
14vYcwIXv+c45r5hE6w3B8rNwqeexaaxli9OkCVlh1r0ENW5Ud1ZDxFW83c7cST7
RPiqTJ25BSaWLcYfhXlcZU4rg69oBeYNcDe1A9GZIjtZhl1SRSBD6pMqMfPdHP9n
jJjkVzHW8jfmPNa2hjEa3iYRuiMyNeL9GaIlXzjZMGI7RHl6g9bzLcyZc1glz+OM
zpxkNOx3E8CNMWUwF/Ew+diQZ/bu16Okv37lbBpsQyt5TLTPDzV1N2ZAMczgS12Q
7bQdKISb/DkS5AcHLCYzW2jxgt8Kcj+8dNWpPdTFW7hZfQP7plZE6nYjh3bwcDdT
k7Pb/crnQ+CjqGPoiSlHYcVfARKef4GvoZ6f4m1rqjkUM+4SMBPFx5AZRarGpU7A
C2okp4NpT1+mZVopO4rXoTFeN7Pbjaqmh0d3LOoFQ9HfBOzQdOvpPqAObk0sr5D0
XszpQlmQSiH9qYEa8eLQ2hQPsvxgUuG70iXo09Fxw6WBDjqNjSpSZrSN8AzXsKF2
Ep99Cvj+/vBCn/n/7Qb//CNUOExEiL0/wLjFMlsNfssTVbfilj+foMZ+tHNOF9uM
5DvWkgBpzCW0A+xYF/93npY5dfm1RZNfp+FjAbmjXtvKdhKxCkWza2+qde+S2wF6
SBaAL47c9UGMBTNFqyMzPm0ALsl4EYh3+dLKKFfuBILJuCo5YWUKOSsMGkzxGWWj
iAyVHIe6shIDlvGZn1ySja1ryQKkn+MJGI+eVU2LZ67h7ZB2FocZVOrHtnoypzcH
/XmVxbNCOWCBLTGgz9d0WkOB/tEmz8pAYIBHa42oCYGWeMKR5ZA51WmvSZeACW/3
z7wsB17lOR57JdFzfPwuft+Y5kshBHBFBwcZup3MKqSVNm3mSnLyOwJeSVymF/NT
IN/3TOffyPHV8asBoKUdBHaT40+1nnRGzmyhuQHEpjMneSlVtp+/RPQKMAE1IxGn
oHyaiP1yYePCcoTUCBQbE9XTu7mV7R6cYnx3xUUGJkQxXsQQXaWKXAmLJRR91LWE
dTCIWxRjIwIyU716nAeflKMW9XSkzmnFNiwJjddqRFH7VmLGwUHzNIQ06k6DeJTG
9ufCOrysOn4iTV3Ns3SkaB3t0smnaqNin0jD8OinTGqW47BRv4rMPlBtkPGfu/or
GqhA9SNBM0raLq1SyJBC3PqF/Lkmb3y0OEZYuDdpt94GfrUaot6uIv3mF0uiNATJ
ZuIO9g7DnZnV1A/Onb71NrPPN8ztutTqECcFedc6IQYrITU2bD3uk23u2x8axNGV
9Q5c3HMDynCL4+/yneBYY6SkC+Hrg7GFfn7iAZtG07J0YVP+S/c6EfIguVjyhZrW
9HmMfGc9+lPdtXcdc/jraR31muWyAQX0wUczW88EkEgaLGOD1Yl8cYtTISOM3VkB
IRggAIlovOKNH+qhYm0vZ9uprVChB0gBGGvfJmJYwa39+EV0sXRmriXzIoUjzaF0
2eBgz9d9o2UMCnm19nAvNHwf5x4jNDaUaCMk7m9ra80H9YmfORLIA5K4y7F/44gt
XA3MhGla3jrYDoqWi7KTG3IeJOe8OH0K3dNHksufVyfrt+EQNOn0qz5Nvpi/qwGi
+O6wJ/y1opj8UIsGT+vRdcr6BIDw+uzH9dQxPcC2sOrrAdeEf8cHK7xLZRdB19b+
m80fnSyM1+WPZYeyu6Zf2cP3ujLfOYgBJioxBSCzJOegT0oGPl7tnQPTjVcIxie+
ns/PoemYCE7hNZNiIolMqfLrIHMdYL4yOV9MTy1ZpcoD9DuCZNZvjOcd9nup6bFm
nL4YnLc+9JM9W1n0zbR90i6R7pA/8p7lxLZzYqerSizuMD+4tv0s5natyJvT/Mot
k28kE8R8o/HQWCJdmYeb/rL0Ij39oU/NfiBNS6SloxK0Uy1KWl8QrZhunMcNamX/
vY2hpbS7QlPWZiOWQZECBKwZOmgmrMxPxdqo5TnXV6n7bqwFQxnIuSGmf5LT9X1U
rjNUrdv32qWVy6NtSJkjHFtU/wFYcRsVle0psNUhMJh0Gl1GJbVUw3qIySM4Dilc
cjB1W+XXgmpVRGBRTD4y6xA0Kzk+PBrw4HVDcsb2pWI3EwDydI7/uO7Rzi+SwQBi
tyLPj+gUktpqNKOsqhzgt9q4IyPBazcB0hXoM217OoJANz6U3Lta/0fM7aYeq4oH
G4DbTXq1iMx7VBrxgAIwgt4IleDmYesAB3FzuHwfniIMee7pFYKhI6OKq3o0OuMN
`protect END_PROTECTED
