`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xNydqAsclQSMGuxgEvkEZI7oLsq+De8InWZ7MNOD7M1jGjVHkPtBdE/ZSV+A9MjP
hPTw4WCo1Z9ZS5F4AXpipTEyJkBgz4rz3L0XoEOmfzLxy7KKUC/jG0PF0IPSCDBQ
Qdg8+5JFQpXdS+GaYrKw5qmYnG+ubNYWhqXJGpj1MOt1A4wFIqjnJFxNVvY41CqJ
qnns1KxdiWfFYppPtz9sitRLuFaPEmnKgJNwO09eAJujgxTSVep2QF2zTWukxLc3
dUwA7dk4r6iNWibtLEX5oUd0Jr0FG2Xbuv+f9MBID9A=
`protect END_PROTECTED
