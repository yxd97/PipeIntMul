`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JdyTn1tfzKslNlOYvY5JRBF527YdkLc92RIo4AC7ifbDz4nF0qZcBafKO+dZV1Qb
R55OmOm6b2KBV2GoQ8+1NxbizPRxaHGisVQbQmh1cIcwAgG3dMJsJPEeHPaLDqaf
M9rYwN9J28o02dMl318u0LQAzshl8A+45+iyZrqSRn2K65Jw/woi8XoY4cgXGLUs
7vC6tKZtrL8cbOd+gNkOHgJhK1aR7tHmoxBloGMUjhctx5IgfLBGquj4Qi/j5/bh
DO4tODMS26ptzIQozFALXOFQFoCeZFm00rLC4O51sSspfz4ZVnJ9nNsGeJibgxrb
4XNRldGS3xlAFYhgnL2l9NXH4jkfFSwad7URFDfmprUjJy2ZOXFvXK6XvMBrGV8m
OQDyL4SYpYmZ1u89OUJZtA==
`protect END_PROTECTED
