`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBJ39+U5PpnI2TXe4Q61A2EN6DQl5t+xd6MoZOlA35V6VEECAQhsnTFUXErL4bqe
Nj+28XIhDlJv5qMuKQQUjg47VRHG59shVJgFTequ9ssnPO6bqIFkJ42AoXq68wdp
pJBCEaTJnofo03Pp2CMVatS2LIRZGJ1BaQnvzFgQbhUZSbI27ypPd3Lo2TX0Gp5u
ZoDnbkgzrbl1jAkh7HDIIDfe6pqYdan605EjSUhBx9u/e6+yExNAalt9yqCAsVMQ
`protect END_PROTECTED
