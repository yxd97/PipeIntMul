`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVdgR+fMjuK1Q3fIl2gZyRpmMja9PXzm3dOVhA5nMW89ul74WodZJWEnx7eNidSV
JcYOZ4EoGmEOw/Ttzqn/l3ZzmnGDlaRLMYrLJTP2WzNk/uwovl6DKKyzRc5NWE4B
X2glW3WOQXYaSDG5OdrAx8q90AGV04A+jnUjZAewZvfjjA/u6sSw6zqRCmz3bLrR
iHqiMkRRybU57sRim9y0XzqmfmfzkPAV7QbAqnBhWjtrpIy0OcXerI6/mbaackRR
lIinDa+7p4TMxTv/QoTKfTr1vuLfgNbKuqTRk4XhZ1cI4YEMSflihO2lVfaOiSQ4
GyvbKJb12E8aRauOokGhRJ0gYMd1vufQBxQu0FTXQH1mwiyhuqO9oQtj1oyT0p2n
yqeQfqyIdA3N1v4El29TL/seX8lc92ZhcsCmniE8Rtio0ivPjrGcDsmCZXVFba7L
eGu+hxucJm9LDiauprN99iksWtMydaF4CXux0soHa5dZfZFX6y4G0WSS88B0nQ6I
E1sT6QjUWncc0nkKCavTnOtHdpVCSTTXpYV/w9tFGW2hbpFS4f1rRrKRbD5C0KJi
4za+aHqeekxC+/QE4/mjyoYiihER7km4U/1oSap2QbcIVyNDP7+quoHUwO5h8BKA
HhHm2Qow3UqDXo6ZkctiFAFndr3uFIe04xqcyRfJIHqW3Hy61vjbTCtC5yet4eDx
njVaBYf2I1lXYV2qTb4Xbe9yjfKJRw5vD8Z46BcEQq5Z9v9/CzNoLISPyBrbGgoa
Fil4tUf4Z3OJXeeUevE5oMrrnZI94P7Tp29C0bom/RqOmfXi9yOvbsen14+wFNd4
rkiNtY9to63VecrZmAgpwpAWgU8DI9V/ASslL/vKlSoA0rUumg52829xGP/g0kDH
hVC5PT9zxxVx8c4d20gnwA==
`protect END_PROTECTED
