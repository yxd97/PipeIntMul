`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBPCWxIIJxMsBl6IInWxYjAVbOfZDin0g2ZrSDabDrzUFlEwK9FHLBh1eY2VJvpO
ygNUeQwRK/szElk2LipCZ9MflEm/v4JQBZ7BifHLfRHq0id6jCwFHcyXr44daoO2
l69NkNmxet1XfxMBBzxnw0De2KnL2wVfkUhpwnme8fzJj5sS+rtGIn96taM2wjuF
lSTL9mzpVyyF5wL+4x+NTr6AjpHdwuN794bPUgIkTPrKwWzh54/yIx9XV0/iohYZ
lusB0H3QDUmhmg0lS2BowYQiVDR3epP01Eano9+ns4XZ9QZ2T1Mszh4J6+1RTMX/
PlOj5v9Wag2s1eLGnxCqHwcxjnInb6rKR+WEoh2987AmhbFk0C8LO3/ET2/AHr/N
WkUMeUWJNT+mCRABrx+SvdAvT62W0h1h1Q6sGqEiZ4fZSuZ74ESEvcSS3/zOrioC
`protect END_PROTECTED
