`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T2lUnPthFbpyqYjh02brHzR4fKHb4DJV2SFdmiGcQFMo9WzqM2tZJQKst7o121Ok
cRcKXuM4CXGDEWGV/vX2zTSMSTQIAQvezN/lm8JSrHczBWLBz7BZ3vluJ+rSwffk
zAIQGL279WO2oLIQd4wQj2WbeBuwzwkNHjgb9UrXKaKx8vTY5CiiKI/b31b29dHG
4tnC2INfHv3icJDlIjtl/Yb7QwmVR/6nhRXlLaxtsnQunwS6b2s7W2zxO390ED80
dO3WzZGgiWB+ltymUy/lWfq/+OQDBbJqRdJtej9RGwW+fBDt88D6fbH2Zcu4BarV
Hv0uWGCQGJYwsUte/V9tr7yZY9NhKUlH/52ZjBQ8evJHWwJWmZrcoqUrKgGHdt4c
UWA2mjXNY8XnaA7l7tdbEsCAEY2gBcGwD/vvggeAnw2hEIuUFitjfXlH/J/imfD4
+xUBnxhUeIweS4e3L8xkl+qJlMOG8Z14C/cA7qhmTh4PNLzjdvghb0CSBr2aIGUE
oUQ/YZgtNvR+JM+/J2nxfHuWFYOjCu7/oMnCOU5AVdUB+YjlWSkifj6adkaJmuGy
vXlBaj5/P8PO6PF+19O2I2zexU/L7WOwPHkGOEwCSdJW6mQ2L3DexswtEpinVCcM
0K5bv5REfkdm/Oq4h+FgCyI/f6XQ24TMmy9a3nsUiBiUMFUm3kA6OdpPPF1gpyDr
nyl76LpUEh1Hz6pWoDL73vbYa9yTI31l21zK6h0hWWPq1BUNZTQwwHdPSW1LWPdd
VFUjLRfAknhn8FuWtmR+BVwfCx5JEhaxW3aR0tgmMJMDHclVICkv7FrDPh13Qbyi
0brs5Pdgo36l2RQ/d92eY4ORHfvly3xdfRikSCKM86tre62m7Cm9rciL2F48VRl0
J3/CzzB9v4jXxf9wqnlE4KRvoxFZ49m0229eV99GNtey+CXOW/xEAdTEBTrAnSX6
hzyC5hQ91Fr4C/zCkQc9WRcAj2a7wW3EVhbUrNY+S0ZnR8jEbyzkjXjYrqw6FQJx
ZYYe0C4OTaq+FVxGdCQG/VrJguL3uWUskF+jLpaZuvtOKwvOa7+OZATYiL6yomlS
DcfwOlTTeV0+FY93s1XpjQd4tA9SyY7rpp2W6W/Qtg42NxAD1Gamxe2WFSflfYRM
3huZ7x3OoghraKRE8zBMnKJo4lfK38fNVL9lKXS9tJJyO8w+25/dojNc4mrRsEly
boX7lCW2CLIedprwJLIQhv1G6v1YRfElXtx4wg6PNjfXQOp/ksd8SP+ZVxn0ERag
4cxG6HIsd8RIvgFLOlR/Bo4wDkDNQEyyyMH5SMpYxq2WP62GOEdTic3TTulL1dd9
mb8L+HUXvvXnXnmi51KLyCgooc2yOSYhyo67lE5Zs8kgVJI7W0ix9U6l3IiNEnY2
3TU9WceOxRJasbsxKdxn1jtR+Zs5YqZhZAIJl8p1ZLytyME3d7ATWFsrx/lo1z7q
ZBaa5K9Fq877Zt0viS+qUPOm5Tq2U40/2f4Z8WVU2oiG34ufd83seE3uK/3pn7JM
ACebp0Qu/rKUsNvC04cou3PdNveTxTeYbC+uXwDxZHt1TjCkfBQ8pPjme/mimyGH
DWOGMAfcuE/Wf0/IneWPg1hK/hTsLKWbioqtksx2JXTH2RZeOw/KgP7Gd4mRlbns
BPs1bDWXET2JIebYyTmlDTWQfYTNH3b/PnSWqE0G2AFORRuo1l/Vg03ppoy8ZZYl
RKr1FwUpWl2rYQBxk01qlIPEItM/8fXU7cweTL0S5svVgih7HL1FIN3zK8Q/Bpkv
a2OQyX80068GUq1WMZPhxzCYIotmCf7uVRFLlkyidjc60Zl/Snd0EUamuBt3tYpB
5Bp8r2pUq66ky0ALNlYKLb34I13eU/pt5R2YnRbSVnJMstrP8rJmSlwGjF4MFUy3
Rd5iGWQwkvtqGLEnMBswyV7FqOdsb/fPFPR4vgXT0F+RCXCREhWZYI3FZQywfhTD
jnfCOYyGp1QXjutKQ1bDGA==
`protect END_PROTECTED
