`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBPFL/0Jx71q8SbSuJx6OikZrZ0foHE539uPLEtI12Ug22cQ1vW8A+IVLUnf2HR+
iP2K0ghI1N8qrioTNA4zESyIEiVU1h3HdXG2Tq/it0xaKwaQ2x8ms40LeDlHXtbU
JcTvPvSx8UJmasUPO5XYKeOQbo5Y2y1IEFrhIM670ry4bKo18hE8PxveV8Pt3U+e
GyHqUdAzT5CSq49ERLclmr94WMY3M6IQpRlSIXjNn9KEkxA6oq8zNyer3K8uMxcq
jmEgObyCmfjhIe1zK5ehIYyIHgDOVD2Nvlll/1p2DXFTDhpPsN37RpWvmpewJ0di
IQLyWicqwsUyB1YHch+akGNLdyujGnHv6fBzr4UTqA7ZInyWFgfI8iIOPdS0Nsb7
ZFGy5yFZjE0MFWkxBtCuYZtQXlLQBSNmNZCKEqPK7QFTg8+yCGlEkLdgYfXBNHQa
hWaSBfOWOOniNS06N1ETjYThyr4Hx0OqYgk6sAp3KO/5vtJbHOsik9Jq9y7+b3pR
0RihP5qvFmQ6ZRbApz9Cw+vatmKRE0shsvKb1DZZmr/gTtz7yF82laAuBCL5OH61
vq8iaWdNHiL/DknoroLXLtskAKJFBzwzWh+TnjRSl1WQw+eWzf+GtKYygFU0FaFR
CZqomNj4t2c42V1sF3LkWTmWnSk50dq0eyUGVWLBsDv9zWKeztX4ck34hXgxha6l
QirZCgfTvl3FkvdZ4NORzoNxCOex8fOUj5/t034oVT5PqN0l8GR557XWJ2f7gaQL
3b7jEiShHwrhUcQ66La4QP2ghCLGsdy+FQ5m5QGpPvX8HOFNKPT3bwqGFfNuzfF3
gXi3bH5UC+9C0i92qBHRz5FPCLElB+IkF39zgkyT6tO63ICwRLdzLJgR4pryUuqR
ydIQn2FpORTUfdRp0Vbvx7Q9KReGq5e0zryhvbVlb8L6l9Lpb9ZeTQgrAB01y7lu
78jZ9X+ElwdNRTjJjgshsAgiyFhgbU4w5BsA36mpkQIzDOe8Bjr7K+Sv2zT4Xhuk
3uyF3V25UNp/C/jVC0RUbH/+CBTy3XnYlk86U7BBZU5WproL1i+8yeRmfPUNxgTr
F7bjeqQShiH41YEOQ24z8TPRaOEnt6V1BUPcG+uXIaGgAaScraes0e6MwcbArzC+
1+j4QfEANqqt8XADmjl0eo9yO+5oyjOv/DKIOjGtbGF8t+rYikbnZL5yTmJPg0aC
ShZOBT2HtCCxlRW5awe3+KGA1ctUrmjWdqcmzGm9zYYPfeI4Gyvp75NgjNXT0Ajl
jaNnOQa9pmlL+S8z1WIh1Q8UjhPbXOP0sKhXbd72pIaH85BgWP5O5w2ilMJnsPqO
YdApMqzA0RsUN5BMBg2DnxOhUcuwumm7zlHp0Xd8p/DGwczEKzfkWqjeykgahrUZ
d7G/P5Uy7XFv0iM9oDsu9joxmVqnx6C9f0kaaa3eiQcSMquLTuhwVfyLuTEye161
+y5SYpxqSsIsy1KLfbZ3qRMCnOyWqpoTJQTZJbFM2OqS7FwdUh9zTy57Ik7OZ+Ee
MwokWvfLp8Gb8tbXykVLFmhJ0CQOa4Or1W5+/iLYF+cxZ0BdLg/2nYch3bl02bnX
CwbSWQ0TxWhwsbtN+luKKqWWvqycvuwEm4WpjeMVQrJG0kMG6hGZ+vMU1BtoS5Dv
jbWPixof2d1XmeA0p5hLo0OBqMlloaj/AnQuHJjg44DehXZ2yBUXMMFEyhBx9A5E
PQUxFhOPo0FIxesH1tw9eq2Ao8y1L3oHPlajzfKQj+4ArN1lUNQ+fzTtiC//ZuzV
Cj+vLaT0Xbo4oBlLFi6yETN1a2Kiu9OAkoCQDOxKPfHiFTv1LUNqmWH8xsvpAbpU
uIQXe5qmFzWarfGcMjmkp4OtN6UPaNwTOW0ZgOJblv/UHiaPSVPxf/x2DU4Coorq
PNiNkMwu9GO3BcMTH++TT6oCJl3OJcZI1QKk3Ma4aQaDUSaIUhLsqw94ItovF5ht
gnc1RrLWNY8t9UKd+4MJ90aTcmthMmX0FejES+NzYfUpW1CYY2a1nNewl9DYRJPO
CVw1Q8vTsIehjnnZHOPnJTsoEEuqU+uwovhDLFqKFH667beUXyRHV76OVwNv4xSe
Y3ZDcuGlJOIA0/IVfZTN8b2kKeWMc9vLJ7WXYtA7w3geuJR4yvhHsdoSqltU9u8d
`protect END_PROTECTED
