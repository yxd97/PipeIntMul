`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+ukscg5r4vojggGXFSrTet0cKEO9j2UsmaZau94ItBVIbR4EoGIH8sWD8TYuZQw
a3Rbv2SgpIZpS7fU7LUdvd4mEuPL36M/pNCLKB4UaGQaKZximhybJ+HESA38F9xk
SazIVaMmmqnHA/owNhcCc8yJKcEd00OJdq89+L/TKcTrs77HiLHwz312ObDBYpW0
+duh//wCpvZ1VsR4sgxq8b84W2wIA4TXipN7+cHaa8J3/970DeunoVWfEiZOct65
/xxahiwkByv6mi+dsNC4FvMuz2S+POWf5BYjLvNt53B1JKe58qQfc9EidgkdHM4h
Uf+PpSb5u7Dz9N73whr7SKJgQsL343QiRNWGBCPH0HVCnxanq5weze4gRym++SkW
A7PMdkExB0gyp7ThcBbY+doV0dL1C4KZmjQ2rUaBka7f04o8FhhhiNW/vYdBhNK+
fXPW/mF3CakcrUrLNqsWhwMfnoUOQooSU4Tew5KZ4bjVrhqx/d16zp75tqQx4t71
pb6gREL11tIi8rERJ235IN1KTnSPuOW35odQPR1upuj1WuTTJJqbxlGxLpDnvUd3
EP18F6LxxBDYwYbeoOZ08Q==
`protect END_PROTECTED
