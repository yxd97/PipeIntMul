`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbxVCdEKHxe3GWcVRSuB6XASBigBPlqQ+nR4vE//55g6zc/5pMkC82tKeLXEVRNZ
NYWmLNdUe5Is6N8OAcsdnjA5JkVj7stjXUuNOCGXH+WuTnMXnn/XUmsQbMN8X3J/
G30ZI/XYnim9pgH86wB+IjXd1B226FOvzsd6aVJC+TtmqPMlbx9/1THlZ0sW/Tus
Vh+QHXbI7ZX7x5k4wIKrkZOWhdl9k4jUCnU6sKyD+znaJ3sPBxLbfrjCPj2QZjrJ
qs7GdpBXQYXZ314IxETRA6VvwFLlZiUxRLrdXwve4hmeigiZCC8B3BSwHeaP90HS
P51MckF0jrjCA9V1svQp0CR+i7NGookaeS+ZEkFWjG96cqPoRPYaR3MnBAtoUqVM
tx3fe2UuDD87ppsthf3ytVOaMrxAom9cgDj2EvtztoycT25JBZjfk8iw2MDNzA1W
575GX7VpuP0cHsKFGyqfSq/K6h7oXka2eYtacb2fLwoNiUX0HydG6xSCxIal9Zbk
AjveS+3JdH4syFtHAOEclzCn5D5f6vaHLA+uTIMWktnaSulDmKmbHBX1Q5OijuFF
Yvs6+vJxpH30RVZptSP168VYBjtMpK36WgLQimn18A9dIv3iJvPpgDyMVzlk99LX
DD4gkf/W0Ek7wVB/fG7WPiveLHX8BB6QVorzxHKrttn7WlKtzHQpTNpDwg98q0Ep
jaNGq7s1vdkj6t++HFbqVDcUtwpUgozizUgrfHv5ZlhGFvDLMAlMa/llks9IzYrr
idVQXgeIDMXs3wUE/eVr7A==
`protect END_PROTECTED
