`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AsZzYHSaikZWXFPBiGNU5priBE9sg4RQtc3ZAgTHX+dEKeN3kKqenb7pMo4rbfWr
kEFPds4vmsMThy9zHxcalAhksNrWHrTJqNa2DCpkC6SMegHRYtgj4Fjv00jVeewh
+iExLvyYtNqn+3H31PJVJTLNRk1V3V5/yRmrzfvonmsLPFfLhChxdr/nY7YmUXk9
K2wNDkvW+QSyeW/luQkiDd9vv3c4oMpO91X4grkyQi5JAXqbKlQQdRMyAjX+zApn
VjERL0dcuJgZRblX564XqnQ4ba0aK37SHOwqJ7qiMZukj7B8K+/J2wpFeobTC0/G
Q45nsUtS0YH+2Qj6qTmIwL4QJ8sqq1Gd7GhTAfIr7X4ZSBko6KxFrmhCC6cACBV2
EKUM+vpa8ywksFY16PztrzYV09sRRa8LC+HAkiLUPTG1m5K7Pc0kWCo1nQbUBR7L
PGfzEJ2ljhx92dfUNPUrwzMOOzuJB1nHztAUotijQu8=
`protect END_PROTECTED
