`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5J92oGCEY/k8D/eYEosf/FY2Iffi7ZdghCGhNeXKAE7yIeLwvqCobCUov8ZgoPGh
+TucZ+f0JLcZLd/Kg5nxA7CD6lxk52/zc8XXQKLTlJoP7K8wVL3pTlW+jz4PAvh3
Hx9KW/JAklDe8wrvd3gstsVeyuP6WgYF5wpoUU3+y0cERyVzEr9GugErRXI3BBxG
UZaafyGhaI9HxkJPv3oD8ATa4cKCeCThENgSKYvIUBU9HK5MGCM3JrtDJ2CZSVNV
GHoqw7t7RLOVnf8rv9O0OJ+VQn6b9vu6ywyjkuP8n8PdRuHcV6q6JT9W1bkUrqna
xBfg7KjaYGt6JxWcREQQPVOZF5PayuUJkj0lWibbE4IEVH3PAV1OJOQvFv6TB1HE
+h2DBLP3sjEuVotlLmzxtQ9aRLIBkChhZvjjSmFLM7eIqq/8uEYETDmSIsU9xzLr
8m7UKR0LkEDj6paaJRPFZqcIDJk//D7gnwJxQuH2NFJ6DKHRQhSHDjgO6jVd0rGU
rFdHZ3U6PVvqCwxnfoCqCZs8FfxMp9JGquKIW6MIgnG624CQ/mk4hxq4ytjC+EIy
jLEW/TZxL0wt34gq3xkdmzRN3UgeMu+URMguFfei99AoNL0rygGLfX2EYcuSIZ+f
sm44Wixh3yWf3008JJTGUYEVHvi+qIOiLYxFXmdOpBuOPzpDKRI0wi4gBtoPT+gZ
AXuezQI4uKPs393+h3GvYTlFvyQi8TpNCg44hD5//YEx/A/XKVRPdHE0G4JhNS/T
Cu7SFmMPMV4G2kD/5RlieIrEdre2T1XM1a98jrD5lFFav55BPr+qYVcgh7Awcv7E
m+ld7pn89kEeG7itUHJchE+mWstt8obs/v1jcJ2hyYJNqY2uEUldqTCFq6wvE7Dm
akarb6wsrBGQPwzcwdjCKDeK61lJeN6tYYOUETUEhCrsNQ9z4pJnljxr13tlEzIQ
+Dpy7Xlp/hlWKXv+uy2Xh57OZga5z+aO71b3PjRWB2I=
`protect END_PROTECTED
