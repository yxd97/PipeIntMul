`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fl9ciCNaalF+VRryf6ZS4CxKKNegVh9wDTNpLQB2BUmEsGTTy4Q1Jt7EGx91ethR
XGQi8cd4WbLSDe8z0ZGxFijN798vcwXXPskxkZ6XKb+AQk0PKORveRcFyR+wLhML
NH4YpjW6i/jd2Gy3PVawjlPsRhXc/0FmN9rpJkMDlr6uq/RuP4I2PqEpiaqjqI1W
2YThzTwUjQBDbtyjg/2hcxFf1v38b/NoTcyhCSyJTa0ORyLtBdE0hYQmAfREUUsk
+wGurAUeA6FQpKbPtnm9CsITFgHPDAxMCjOGIJhWqvhXk8OxoAvftTTB6O6wE+o3
sF2glYf+/oqfczolxBvajA==
`protect END_PROTECTED
