`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xULFqi2autPLnQkbruwo9vS4GEJYOCPotwgQwxLCspAyXZ9a3KLyVySbX/RZa1HK
+7NhSCVgHo5vmhqmaWoG6evI2GHgJxSyn6oF7fAPJ6vIdiGthQkfHol0Gf1UgJy/
EXa8oDjVIbqicHuOtQbgWDzRfnv87TFj6uc6YOWmMrdmgLXoC5VE5cHiGgItldUd
6H4Nn1EezelXtHyt9PjF0iwn6cBYJ5obrsrYk0Kk3ye1tJuw4g/88daBgrQOK25H
c0I+LqC035XEu+5zVBKcGz9jGq5ZUst1tmdr1P2AmyM=
`protect END_PROTECTED
