`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YRRCKVmtDusqrjw2CvKklmk3yb/K4DcRH8zOQxsoLl6n8yCi87ZrPhq2wn0CD52M
Q5GMABHVPjx2EdH+lC6X3LzchJEdygBGMjhYILHN9k7Paoc5knS1oBEqg9UWxYTg
Tb/BZmWSxUABuKSxfZI2SQ8raendaP3MFL0NTPljBAYsuaPkuFy3bECVsDLXTYb/
rJVOXY+/VM8JQIg75/PZQbhpzbOQmXfrphrA+A6jePxeIf1USyRYfckmAawEMI5e
pYPh/fTGmomegVi8uH+8S7z+7vzacWODoPVyOZL8GAfjpz5Cc+TCcEecYcGqFhR2
o3Hl2eV51LP1rLMG8/rIQ8/ZU0ZKmxdZ1RBElPq24wwhLKyOMvPP8TSv4VycXpRK
GKK4ZxYELk6nVpjMUW/3SjEWWJLOijLGPyQZDgAjI1+pBM2e+MHT0qrCf/ggoENR
cIHxVrPhu8hZn/R0491g5/h5HxkKFH21SgQnn9ieIdpm92MgXNvbKoai8TLrl/GF
emNpYGU/Jn2Kbd1tGHd1DUoHCqHr4M86Pp1sYrbpeG9wx0OLJK+LSebgBaF44RAy
ou1Xite/3Lbl+KOup7kntbeg2UmchJCmgu/qMfFPjb76iFuxFXhqp1NyJgvRlr/p
7krtwIB8rEcS5X0RHGLPwjqonvFDXNOLB04jXDvx+NFMFNyK+oa8z0FZEs7H9pqw
zV8cbmN6I3g6CccKHaAGvXna4dGzmWTlzRfbNSxzRtyiWtpZV8/U7F+YRvMvFxYj
YodGRkkrl8qfxjRvtT5iHwFL0lNg5oOFH5VUFVgRyRoH8eMbMylbijHJVmo+KuPC
F6g58ffbBA1WxGfiY2Y3rLDDsxv0YACGhrmRVGY5NfWPEmQ75IVCIOVwgAbmw0Av
c4zb366EnxglBWTAN6fA+BZW8bdrZH2qKfNiH8whpzebEsSY5EeaWMW++HFfUSxP
ZaDGZIHdO03MRKXgnQB0N+Abm0iWpM64ve/gzpqsngGyHATeCQTAuYydJYv2uVl2
5vyMEMrViu4RT7Eivlcia78uNmCAI3aeWkvSbo552cXjrAI8bpSuBsqFBbefTWZP
b5W7xxZ6gU5la6h7dHaCdXE4pmLAtf8w66JVSMxfcG4rCPSHS/yI9HVxrc8XJXDa
oJLXoTR7o6rP5HSOebk2G4pd9As6AjYqtPc5q1jV5XukcI9TxJOqIlJlwcLdBHtN
FLp+7ib8J69i8znGiFT8cRh9QE7gmkarcuCWCz0MGohDsb0JzNU8OZDHoSphwg28
Vfxx38JhWQB3ODpadpAa+vwFVdALdf/VkHrsiBMjlleukFxIty8/VW3yRCCIRvyI
/kzV61/IzKVizQDNJo24W9oc/tjbRrcjr4xmPDbrX1YIbPDiWegk3YFZVz3Dbr0A
tgikp2KvQ1soNvkXU+9Zwjqfpuj7mk7n+CFQXLbPwaZP/ZbIJyNrd6difU3+0dSx
82hrUPPAWlrw3whFjM48SEKGzCVDGs6uK7sfaiUUvqZBapsPJg3ax1WVJuCApuM/
g2QnaP8Cb6FiRPlgT8BOdlhdqsPeKYofXM27IZD2pcoWFUmHCoUNUGCo+t7hV3Aa
Ub7kiHqAR09OWwbyn/Lb5lWRMhGlw4BDs8L2aRQm0RN6FmLcohOmFU6f1dVXlNyH
yXvh+9C3tpDqQJkJ8i5W2xuK4G8Yc/D4jEc/YoYeapZhANsEiliJnjTlsd0UucI7
7QGNoAS9Xn6YLQlulHXylDGM61fMbv0SNI3PEjvkZYxHVSxAdsb52yRhwMj6sg/t
CubiqrMbjBUGUMgEJpkrOL8PZG7UMV+6Vij9R91lce+c9tngGQenOFOBZy6Ck10h
Rv5qtvTM2LvYMDT0BHhyijgVQuFzpcAA+caxGIX2PAgy5jjCqKH8WIBorf6WZp0m
0sggc0OHQ1YN25l6aB8gqvs+60FjnDvUKyQZg2eHEQZDvQSThMaj59XVSAR3Nf7j
HNF7Rx6wuayPlMRlAQj7QJW1umHqUtA7PBIEl0SYWVaguPPkkLLdbFw77xapGezW
J4D9WgRXHZ83Ko6xyMnAQlGe7g+KavgpdLH+Mm3EV6ERocEXP2f1A7UBWCSm0nOW
jhN2MoLuN6AZAtOh8nPKav45llewA0wiZZG5qtR/Ue6TDTgu86QBnAKJ3qDLwt0r
KPod35JdCQgeosZtC7opifFlTy4lRAKF06lQLaiv4R6HWmpCvypvKSGQs+QfQ8nD
PBuKWKPDxTm42B0LUUT4AxpzfOTLwTZ/9QWefIlSPFa2XDY00qsDMvwvCBSvooDs
mS4hWTCKiAkzlNp2cpOq2ArrlsyqrVr2OJPS0mx9Cz8kefbsLI403aH3C080GqZr
c1olJVoSetd09ywCmptbgq1b7XKcUABQ9iuwKPg25Y/sfkd8DO9czeZ78jlCyhXx
q9RkPkRVIOj+X0ZZ//DMTWYjMks9ydCWCWsqd/LL8k5n5FmSGMakpvGSw6Cvmdgs
hl0biI8grMto/aVxhHAbKwuM4oe8PuaEcj1prfxHwipPxpAcJkgoVXN7O+Jv5OrH
EMREeQmH58H/rmfc/mE+MAFxday7nQDngudG1faWtTlMjKZJrwT0fL1bOfCyVyMR
RJAajAs0tJSsOY63TkJmhP6jdQTmCOw/y/yti3gz8+jFW3V312Mutt/GWNy/RSU0
MiVn5bhEnC7QtmBxlEPeOGfzWVOp91PRQzG8J8FiSBmfvEFHEcKNHk54Td29Zn+R
gtUIhhwimf4b5YINOt1e+pyEYnp6p2fh9S0Rqu8Iv1iFWsoeTaBi/Jxk62BZkPe2
BP1A9bWKJSosVbUvsQHUr2yZKtPeTmlooyWL4AJeW1zT7bpHDgAFqWf26cFVJGAe
00VfbHsVR55tGbqx35iykp9bHVx8yc4dxwp9wYwuVHpN6IMFnBPb9AZUrISJXfYl
9c7ACpYeKMKJZkfwKoB9GKFCvAIawScvSB0be8pRx5ATREp7RlLOh7eF67KzQSA+
5ZtW1kXn7YQw96brEfukiDCY0tBHZS1I+a9XdRi8gd9anx47+kHdB9msjpPF1Vch
AayfqI4L2LeZyVmXNN1ZRgez1rqRXNqVw4fWpGKM7UJmwpaN5L8/dmebm6HD6B5H
mvo/g02WexEiHOhqo4p6vziVeu+DphE4HbuPQ2vA223waB5v4CnHwDlHInmPSogw
bUMLFlcqcNuiwwbnFHo5U1ehp8KgOReTu9yjVeRRb82P2sXPl1u4TSzkcTQ1PBVt
v5MzUPF/xJqv99zNUQfuudTvV6umLKZtDFkFqIPxlMHxuVM/nP9/cRpj6WzDjLYk
YEeiziCot3W7rVnohRdDmwnQn4/VRS/8fiKmpz1mJmRcsIu/KFK+ZUjU7xcR+TPm
mJBoL5QgJN6q7A7u3T9ZzgtzgjDVSBqmz/Af/kDSWbdmsQiqbpO6vpa6Y59sNcHz
bcxIxXjeoxfJyuTnDDHkdFu9IOO9bwQGzR5l2N3YUwIFcegtuXamCGf+m19vXAGo
srt3QWx15xTtgc2XCNivPg==
`protect END_PROTECTED
