`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4eoHHxTXXr7FpgNJS0JwyzY5S6eRtce+Pdn9I4GaY7fu9vW9+cuRhJFuxDHg0lw
9KW587MRs3Z3RJrM9Cp6SHKtlhab867DR7YE6Uv2GZXt0ScwegdWuG6aTVxtoJhc
Y6skOtSbR7Pvphn1D+pAF2uNCPSz2IiMycrSNnGsJOcklBJvQfGknMi5rJiyi7LO
fi6q42Yn8PqHPHe121+4maFVe3P8ECEpthWbptis1t8oxoBFy8zSmq71AcfdqIo4
ArMS4ZM4VEI43H0Jdp4T2ZAygLpAtoXVJ4cL2ZSmPZ4KQhTuvwB+/0pQYJFCl4md
cybIFN2V/sRTATGEWDYXwSyf24gjbAGNVxgTbhlaDbnHdO6h+85Ma86/zQIlOqHr
El/4wpbaXi4E1YvlTI4bb32Nfh8R2Ru9NDIV3KFAENaUYAj/4Lxn7pGq9ZENUchA
SPv/1hCs+ARS8E0/nmSWI9av4LmF9UVGGjiTuyTw7y0=
`protect END_PROTECTED
