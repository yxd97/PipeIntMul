`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4DyESy34bHdTr88ZvUGOQp5Tw4ks3+1sAMP95pIyPJpjkWj76SaXkiisltXfIB+
WdCf1BzlrSfSIlSRI5DM5ioI5JKEpHY1w3IPdW7Z2wAkBs5yVRUk89KN1bZS7fVH
Z/qZZlmHTYs5sJJQUbNFu1v/CZtryWAR4SZjvKs4BGcTgLpHJq5YM0Xe1p9+YY/S
t/TYgMyoJVa14J27Yz51lUUchBzU25uH9dtboH5bVDkAhSE+ndr8OnKeuOMd3Qjy
yl7bKa3YB6F8UTTFQD21Ew==
`protect END_PROTECTED
