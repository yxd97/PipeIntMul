`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i/pvrGRTZhaae3xWd1v8puhuxUSFE/DliZ7qGlLRtkntEMcFOfl3kNJsz/P5iMtn
fxKtFXJ1487syGHD0VRbiUyGrtz+SiNgxRFXoH1pGpC1arJYZS7WFMEzxYZV2m30
+QQemqJ5JSdJBD+mbdJi1EhaRy8pkANj/3Oo8ONlV98UhPE1a9AaCC7wSQqUNX5h
hazR39pTX/Lpc3zD0HLzVHgo/QjuOMX23hrxQGQuRPpyc5VmL2QDUEvAeJT8z3jq
pij/4huWc1ngIg9tVjj4udwqErl/V1rV2UzMnuHCpjOF4GdFQghr6A/FnLsGhRq2
xxf4FH50FY8V+j3wSpQEgw==
`protect END_PROTECTED
