`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Zz2KC7wA7AMaAVFQq0hI9YsxW9DcA2RXW+0ROVZm2w0ClabzbR0zTu/X5K3z4PO
QiUt4W1wPO5WTFizvNbVgFa5U6UdP0lKTCyqwfEdqszqKdX4iEWtCDn7KvtjKkHi
Pa7t49B91ecVKWLwujZicD1YAh2tLJceu1U9dJewsNSDSWcbwlkz2jGCZYUVVVG4
7/G8UkneiX6+kd84aBKNHeARQtd8kqHQJCW9fKYQTb8sFucxyrwaitjsgIw8Kpv5
6/uIeOU5SRAQBsiU3w8ZnJFZvdhF8ROvAZXruE7Y5qslAWwJ+JyJl9hpPEWvFBBy
kR7sxPNZ8d+FOB6FU0NoIU/qKpUNGhrgaIwO7ZLdiFV4uPD4+HuwdgSXSVwX7c2Y
LR2WRyhBwkAUq7Aq+zRv2EWwgS3IuRaJGDVrr+6KDHy3qWfTBjZYUY0gPFDRxhi2
IVMgodyLjCQ9CL0xQ+geBnmXWYHSeCPq08JKIU4MDOFHoKOma7CZyXOAL/bVq7ds
hi3M13ftNN79nhGa4KOH593KMr4NAVkJTZi72lpQlGB3G0yu0jBCvgJ9TSwAUOls
iCeE1NtgRETPNB0MOi4GRZft/S5l3g44yWsApe4ZEssZ2ClNL93swDSM7TvxWPNY
luKSBtPfPYfJsQ9ffAnRuZ4W/7d2gqfWA3lEk1JwtfR5dH9NcyPG7Gw6xEmeYCPd
IQ6bkspncShlTwzbzpWzk8YQZ9wCLvViOm9D2SsvqM3+16rOuroe7fTROXDADJxR
XmclPsPW//I//kx1gnvAtrSkwTH7oxRsVVGT1ThJmk81DylNGUUZBx0ky2c7pqnH
+O2TcIX8dUjNm/WDAhJ3W1EVy/IIGnGJbIlApTA3yBv+90TiISDDrUofiKzH5wOX
a2TD0moP0/9x2aKi5xPTjE113nEYM5zFqfGKwtqWJlBIZQAmH5bau7m1tEWwrQ2q
Z3HzUFnQYLWDYoraipdtzGfg6RZZS8h2XG638EOU2FQ4TWm8WqbAgLT2R1NVnegF
PhekYKO8s62hFYqZiJpKFzVE5QAEyC4r9pbHGJAcH/oRZzgzty0H93lxPD8sVKgf
`protect END_PROTECTED
