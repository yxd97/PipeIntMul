`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNwKVE1xVZavbjmk2FQG9Gq/kld7TlOSgp8zL5d+R3Z0qKO694x0bQDv829k4E+M
W6fpLwRJ/qiLkEX3gMHqA8VCvFC7/Yc4amehgdz7FM++hM+pnVoRtkVGrRaGkFQv
qPSw3OGbHGBayR/eA1H4sW/cLNda03x9PVPwLI3QPs3GzdFM0JWI6qK3WTKW9TkL
oUYC5WPmXQgdNW9tkFt28c3ONwNIAEEkPuPuOQ+xsCqxgJr4xoUAMEixi+KWmpd3
npLVWeW9wTwD2vWC3OJUu0S4hQAz6YGCNj2uJ7VvL8vW0S5tbiy6XQJLFfVDK7N9
nJSIIPrNAzBd9LhlMEsFbp5CG4KbBq/U7ZCf2L10V9VjddeZfEaMDpS2xv3UZyEA
nWvFlaAD4c8KzWjOLG+PDk6w4sdZEGi1PJe396s5xUI=
`protect END_PROTECTED
