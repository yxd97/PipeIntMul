`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9t/9uWrI6gYzHbbkbkKIxs5qsh95Xl7ORG1p32hQEOc5iks7Sus5/i861x5TBEHo
7alcYcNl9WoY97z6N6aCT2vs1E/in3OvZHm/MBSOPTZVyO8+SmkTKyZzWOMoPlTD
7kt2oCwuZcLoBaMuu+IhN8bV0V2SHV3y8l7zVyqPSmL4vRxvgNRaMlCG7ILE4Mt+
tV+2cf5v1qKpbFVPABxqivqnflsYhnPlt0vVz9SFAS0ul4+p1uTp9N6QORB6v1Rl
IAbUIAga6xJPhr29Nrl1DOGtpfwPmkEhquBCWF9VNBkWHkfQjKfm2C0W8Ip/30jQ
cBGN6qSjoiQfkRv0/pUx3iU4FrVr1ChFPy2Ewlpj03lu/eKopyJfXFyOq6TxaKqg
g9IE9wFgguaqu5vqBahnrSFTDbagbtnZebvZTuIhhrwyrNpAYcjp9ChBr4CbKi7X
OfvGM9pdSd46l0Hg+qG2zqcgEi6DaCreav9RQCDl4cVWaosaRqIFXmCHo/IKU1MM
`protect END_PROTECTED
