`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2SJm1dbdmwmpyUYwNlX79PcpEJi1+lLEbM3Kg0M47cVM8IZEFNuahM8/96f/XNsY
n4iSrSVpMl+qOJYd+/OMqJLIFvyNko0JMM8eklZqUjUWVKA8JSJ52fdA5M/I7wys
3rNLpud3DoSz+M3rkvQN7+yvWnOpMOrG1PeUijx5j9mpGhVfutDvcNOZpBbiFnae
0I+cpCPEpFCdcds9MtPjaBGL2rTDvKv8TK5S6ltQhpjjrW7eGdgY91Tt+kFVX8KP
`protect END_PROTECTED
