`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2TAK/UpvrZxKb10a04gfgnLdiV6vi6ROSkqOIAiwdQ9Iyw6qRxSoHN4pODI+Lpf
3+7ongiuiwYvYD1k8DNCl97WPNTjqNmXTVoFikHIAstMrMxJMU/jorjcbbwV11GD
mX76oGZIHdcYFg9+mb6PVWBFuyFTdJxYfp5vaWVwf1m6zXB/Pkw3IYhTARl6F3yH
Tm8s0LxdJnbJmWWxzlMGlnJP9qJPLycBzkX3Er8vPF7+PvEKokjv6UNLDqnIDuR8
eZQ4iFLLtjfbeJ5T3CQBxUMqmdlusDyyWQs0Hsxu5r/g6K3riC0bPsK2epMyqZ2f
Rz6KnMlGP9k7duYuEic6KIVLHHR+XiSc4uA4I6dPR6IOOX4ufIOXMg2PR+pN4yyk
KJPnrWMNdfcoBP9Mn3MRIWfbRLWk95B7Zf8PkuYFIxhC9A64isO/jg2dXGt/YAFj
1sgAMEO24HvPzYNa+NQqO8jp9er9AuwLtNtjiDe5kMcdqKZBuVq7PKW8ebfEdGW9
LHyHe66PVLXJGrlRlbwpd/nZK6Bazagf84je8TmbAtsTFm+dBhU/5ELQR3Ew2doq
GIOHutdndkMJ7Zbk+MUutE9qOWk7pP4hUpYDjOZ7Xain9CQLG1+z1ozVNHmkXmIu
SJvvx5vlZPSuV9MB5NcCswBW8u1HqcZRIrFDxzQrdXhbzYI/QoT+PpaoPSYDtJak
7xMIhTvB2zA9p0aoodVfHVmAnEpacC+NsvpPjck99M+RKVZS4Tbdh7U6lJ9hglQu
Rcz9JvYjrI8p9Rf2VwzuA9suz2IO6rkwfKm2zTi0FAJpM7wonR06JIY/Q0MAtHpq
CLuQ7a3TtzuWhsT1K8EdA5fH3258GYp/mkq8EtkrWci1kJsktp+Nk4REAQYKhtEG
OxjQu603O+ZgkVmJZjexrehpTV6QnzJ9Jj2gR5GMu4GzBaBsMbazZU3agyt1b6jd
u441BW5G1Jp/1tLqZt8/aOS0U+PohPoisAtXaOtbWv36yfRLzdqCXIAGqe+jiDOy
gcwz0xcF25iaXWrdxWeTJA==
`protect END_PROTECTED
