`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97GgRp41pQ2MHSKkPRKpweAb8uq5VeTwxrz/sG0Gsc74p2kyx+PtWWeXdYz43pX/
WHLYqpwd/nO/BIcVgzrKT4oslHFeQ21BRC2arYzAXrXGKrl/kICsXAXwT3qMVE9c
E4J07M7xUp3+xCnIygA3qUhGV85syB7qaYSidr5iWhLelTz9Tr8ZC8uMfaVZ+spZ
0GCz/lG3+Pgf/eFS6nHxiKWmZt+C/TH715xXTGHJ07Kl/hman76qPLNQeMga+IoR
YmnhHkgmByclhN5Ngo9xmRYtVeFESwNg7uRASH/bAgVFLX798fWxnkZMm1GN1T2r
9UNKirWrn/mT3JrswfqFpI/Jj+FOIBF/L5msTksMAsqRp7Ygg3Wrbm/qkuJ7b/zq
AlVI8d9AzQPa0GKWUsCTfEaxer8TTHV0jO6T7Qoct77ZzpTcdwl0qJLwtS+TzGrD
HuyGNj5WqQZNgIO1edJABKLYJdoLDbbYMTZ7u04hHviCrGsstd6HNlLiFb7MF/Z+
8SdERLrrb118W2MdT+ZhLP4vdtHah7nY2wdPxnWfksskCMfqxXasr5GlGa4MjOng
2RuOLvEFhZS62VA7dNgF9pRirWfAoW6bAQj97a89eUYxXoxw2P3s7GhuV1J5Gr8U
/PyPAAFp381kyUYH5qXt7XtviMocCUacybUs0GsIZQJKpAV/LMyq2ASAvKMnm34o
nc3GjBl8LhVf7zz+wdVdqDlYZgPbcXnZXBRLe2DeJYrf1dfCbF2qQ5bmIvAAxmLq
AD2wUl4xB7PsGkHZ5FuAPVzcvEOIxykmq/ueNJwlto7fxRoiBRKHvsKqTdN6Az+u
iKzVOlxNXlYxktJn1Lo7ThQgvfifjjFZTaWrVJys2SEVpZI3R98ZRHUaNm0kp+at
B0noaAUeDFoIU1N4ROq7GWBdlb++rFK9iwv7XrrbaeWcSrr6nGKPrNgk5YuW2jWT
pe537L5SRjJbS5gmYOkxmG3wXVh6Wu+oy1Wt3innYNQqudHBywot1aRFN/zugnZl
f09Rv1haIrEvMoXWiZeXnCt5/6w2q2S7yxKk5/cu/DReW2nizZq2pUaIIxGV8DYL
KCecgN6Jr+/xIba3ww4Zx8buMX1hCP0GV6D829D7ya/Ma38JCRKvXLX4lU+7wKcG
OdHBMNoUc8UpTlsybsL2ng28X++/ZCrBj4gpOwfsv2nDjrzT7qYPfdPImMoCykEZ
s/ySqQHNGMiu7YVw9YfkBW1OxqNC2BTQ1hANmVjhupogmhHj3CKymJbLCzaM2QPB
wNxhyBIQiC4uMoaQHV8GAuRsqv/ZXJv9PSqJPD4CJobah/QEeoKISD2ekqabpMFh
clRsdsMGn7CycIbyfQ5rbvzziYjS0SM8S3s9AKRmllRG20OCSrZMfHqHFpWeJYMB
NHPDJCCHcW0aKu7q3d+vYN46O6R9fWJenX92BxVZ99psSfOm1R9gCjgx6wLJRnHQ
cUi0j+4SZmlqtuV3CW++uDq6OKaUbKX5CY/h01CRaCKK8wqRrfV/hGHJf0oQ4fKb
VgznN3oO9wjLHfj3l7+nqmWn/9s4fi6ilvuJmkocNyy9bwgE8jc7lEp8pK8NHE4r
pnitCjYO0P6l6W57hgZDvQSOBXJnx9VJOJw3K+XsNYn103g7GLAOTGgYogVGerzX
KjDr61xskX7ZG311fvXPdQQhTa6Hamaoyxw6d57dX/EzHo58e8AlgDDSzJoMcn/n
rkT3lkxpBO4QfjQmGtMQro9YbJ5kiC75RtI1PGGug6Uzl6JBJM5Ld8JggyEmS3Oa
bUiaJ4GjKNzWwTMEKV78QSvD/TyEiYZ+59ThKI1sjQtN1ImlL3sEQU1DSZTX32Hj
DjK3CfRonu+l06cBFkCs8yEBSeCk6Awt4MJ78FUrJBRDUTgsrBRFct8yDYCyOk5M
XxofXis+bDAES8sysc+bqCq+KfDtYOFWcDP3I47b81zUA6m9EGccy9kORKV4aHJ4
n06PgKlrHI4IjPmxT/PYJNBexgTKB7NTeCnXfYIOgFTGEC9gK5HfyZSxDjPFV5sj
v6EvxjW70lgDzjyXubMKeBj9IXlJzCanQWziX1sFm1FbH7J0HksC8K3eNlySLa7K
k6djM0zJKS6Cv9vOE9uZNd5gIaZU0nmzmnOlZ8aWBG9BxoPiU4y6Juw+IOnZqI7s
t+6g+xrCIKvctN3669mx26vX4YKp5QlNXfaipRK39b+PsFrIXaTGRVnPYd0TBHWa
v2zMX1EXdTxJL/JNYnHV8LDmzzDpCZmsjyoScPUOY4hF1pz8kkYkL2DMh0qpjdJS
Fz8EHBx3RXTRxYTelHSlNRZMtPv6AaPF7nZINcMl0gCrkGc5jBFBjSmVswS4CK27
M7th0z2IOJOkpfMDJQJywGA0WKYDhntP+ETK3elxokBfCBt4xealGJUu0BFaFrzQ
E5Vg6tTTFRlMqpTOpCgtrJOaOrJzylFomXwtf6hxkeqaEIHEjd7wEgbaG3vJfwFz
OoBk8hjBheuDJXLY1pJoDahk8gOJ5S+SnIaQ9LuIIAQOsntbOEyXs2HPn9VDx7xf
fY6YvelkaeuAEphC0fgW7dkiK8pA1pNWH0S1Y9t5GUUfGsrheMgZ07/1YAcRy1pU
ZS/NJAQV4L3uW9nJ07SRRPUgbPXRVvOiQo62l9gkygaGNVEtGeCKqcCIj9b2tn15
iQpwT8HVUxD+RHDsrE8L60zUlIeS7fO9S3DcMedygJJDx2lI9dxTpOfZLlPHKZh9
i9PpEQUFPX7MSyq8rLRV5GrUjvaEWOKi86u1WC+cT2Pv7Td3Ni9nImqgIZM5j/KD
lidFZVCeaE+GsERUEgV7aHoMaJ0/6ZsQgxAF2CLGt2FIYdV2ZNP3Pzi9nPqXQ5Mm
qIZGoMWdPo2TkKMUPk9Q8Wy/GCiapFmTo8ezLH0snUxhgEVa6tspU0u22SAoB18f
ZlWDRoL+5yeXqbD5TZ/BiSi90n6XiQEQDaWmA6aMzvOc0PFTGAi9qhKzqqWV1U0X
Wn6a6yGTgvDhObfp6Wc0wDVAF49maer6BNCCmCnIFTmRdT70Wb0y8iL/SQ3RxSD3
Ab8GXQa2ogIShwVtAnck1olBVMEt2Es0EKJNPpVxwhtCh6pAU5Lcl3mOWBhyFpRW
A+jveNOLrpttJyfVrPSyy5kQnALgqaVvb1o1jNMLNSlzAYnh44yhlqyGwJwYA02h
CdYX287q7mG4G9l2SPfIYHaYR0uJacMrrwhSkmhuGTaVZL6/QC5YgAdGoRTvNd3U
+AC+M1/JumPB9NoeHN7cy4I9u37kqtvhBVlRxjlajEXUYLi6Lk0BqO6tXrd8Umv3
a+9Hk74ExT6JYei9+CfEfHml8P2uSYgJoM9JanhDyVwIwHZoXvyqXzx21AJnAHtP
ZfAQnPVWn1AV7WmeFZZ7ajqKYXfRyqm4OHREyG7yGSfoB1U21Eb3SkveyELnAZtU
Zz7fV85GvwLCY/Os6o9Q14lsIUnuCJjfjKRqQDiDg2DocMbCTBxEOd43cULXWkLc
N2YWSpbZrjcYq9uiLpqRde0T/5xdXSldZb7DdVNbCk1oFnjHUAwE2ePlm+ddOTLQ
Jgv/9OuxtPzNvU0MAqy6afLwKTYuWte+0FahcFtgEtgae7CBioNKyeiFNE0K25C6
qFzK0lB2ZHmxjRmpZcYrypT5vUS+iK9DwTlO4VURRFqfjz1bESVbVUOYXMeJUhjp
TArYb5MxRBTNMVKF2LgwHUK99VBPXdgdRvhAYFU1ox5OS7kYutJ7YJGR0JaaFrDs
5OITMW8SvFA61EUx4I1iyWsNtK1KNCD8OEje3+pYC7M7cE3A1BzUa7AS4aOuTV3O
xDwYSv+CX39QhLUcCe17aB7jfbm+FY2FL2ND5A312H9oy1j1XlWvt2VFhuQ59qSz
K8sX1ZvteRXaCjGudh7Po4rYakvRN0hLp5LG7Fmb00o4v7kOPmvCi4jltYsZnLdZ
dwh39GO9eUv0xSlq8pkhFSpE7PjBd/vOzn9nu8kI+0C0aQLOaQBC796HiC9uDr7A
4NV5p4YinPf24zfhnaPmdwADonn6e1B8344SahG5lFRJJGYsly2GNeJN5yfR78tO
iRO/e0aOXV9WRJ8+OwywonUmTacKzrQZN5vNYcfdsYu6ffCSXrSUuCRQKtcT75gG
Jf8HN3QU702dSJbOxdX+UKlKoswkPuSf/xtLgks3yoe5Sa5bd7nwMJZ32nZ5QOHV
/dj+KZMl+O+Zh9v1y4wbZ/H1z6bGL+rVAUlxyRjOI2ductKIbx3fzJOj/EpLrEgN
0Emi7KY9i/Z+SSWvRz/NEY3cwMyzyWuojOmDqH1tWEX1pPETWNEtB/HXxhSziell
u/PUhtudsFzrIfqFVdtbsc72pBRmF87LUT3JtiajWN2MypR6hgdgCYB4H/8cIHZZ
ThviOnLrRgmBfEpUWtTsuZac+CA5Hz0mbWOljBHNC9L80OlefET7FEZP/jgxMb9A
XjTQW0N8327fTHk02qFK0ziAzBnE9Jw3IUR8mvhFVX0NHIhJLBNIkinJ2KDI4adL
LYp7x8xex3J1MjiO1JgISiAP+zjopXPyA8MdCnEo9hc1KjhhN2MCPXmxjyzG/PGo
uDiUCkz83AFD6s1mrSX2DOS0IZg+qT9sfqwhj6DFoiSXWSU0DyWV7xE/eYzTjzVw
5exAYxQE7+83398ebJGl1YfbBrWQeCAgIcrVsaGEOkRDmkhju5AOfSBzVpZuIeIx
JSQkkeiO7P04LfMEbBWtH70EPVedEwjlPKbbjgNOQpcAR9HqaKoZsTaZ69UpdzC2
bAaRPikhjFkfAdl+k8lhKlmThgQrwblBJdqhkXUlMbREC7wwe208xOP2F1qL7A00
0oBrwyNFQglGQnHYhJWxIgtZ6i1HVco1Dzuerda4GOf0l6vPOFJ4+zcTPWCU6z2Q
iDVyuajUmI883uufhHky/yDbaKTK9uxfAi55kDNLaZGb22VQUOuB7YeuC7JCQIr8
7uXoAsm+T3ismBhpZt7Z1UMS6V8num/FltUnbQMIIWhsmNDvfaFGETrSgeQWMmNB
rBca7/xGLTAxL33DJ+i7Hnwrzkuu93J4mdRssVh5tlieK4VTIvwp9hus4mmseekv
cJ3pn2OA03bB3xkzrd6KVHGi9dpYIgdr7ULeL7TXBmallwS1ShiXREO1agdcrbSe
Eb/5aKYIlnry8FtEQ1hktbtjuWOWPmG1hocMkVEemBcrQrGBptPk1IYdrZLENQFj
gpmnk1n3XxdOepBn4UdFP7qtS5kFO6nNDg+YrG41MhqoGI2rk72MxtNsHYRG6nPK
Qqm1BUhbf8BKW/Lx6kUVM3I8W/fMyd+mGi8lxHuMDJ+uI7kb3yQUDbRQdFnKAycG
IfJEbV7czuXm+KMSG/4oEIqWFE+RxVinSAMWpsalPcjl8b+v10d7VB5G+HbDqW8k
n9yZOGbI7zORZqyFixFrEvtw1vPG7fsLVa3hD8K8EOBUoIODpbR5/nAz/DoGZ495
kW8ZjDbCfs1hE2qTDWbpjF2x6QMkyKAx1HEX2FsbUuAKARws6g9+AsW+YnYXXdPR
+Hbs0VRd3qrqvWZuD2PjIYWh+P1oZNUz4I62vwHDTWbmsx/fyqB1ipRcoY4kigfs
WgZK2VQsICuNMzcwHGVW24mXxW61vPLrNaEOvrdzH8vxil6C/KddBSe/8NxAOmdm
6chKOqG/2nqetkeQX5h+lVdASK/M318fAoXes2GhmhohqAQsoH3nwpmEQuDhb4ZV
cIsYIP5e1d/qYbNBZdZvQtzFlCTub2HrsaqaqPBAaEZPR7gmoaERgTsIRttyf5L2
0DnIsKHHCq6dIFiLKz5wH6ITF8uDAUmqbHE3H0H/yBeMunlQF9TKZ+5R0UiRtH94
OCKaIpNK8Ll++XCJpZYQJkqAp1UKITmzfhoMomcZloU2GGjD3JIY0TFXQSh1a3wb
xuJXBadkERilgLLlR1nbBQPmiz96wpG1Y5aBcZX8LA8jfMda6TGFteF35uJWaGf5
qI6qkt5sFpo0ayMaN03IVuJi+l+uQoJ965pGf8gBh8Ss6/2XBam5TffVJgCJw0qJ
G6N5Nn26Sq6x8+50qSNgP1KFEl7ZacBN8SOW/3A3H758Gqfo5JcUs8zomWj9DuK0
iMKmeF6Nbzgry4v76SQHLjk1cL6IrmO6BiG9H6ZyJ2N2JoOe29kW+m265CDcEAF6
hssA9deZbf0KfEGrxl9i0apUf4IuCkigUQBRYUHWWnYW6DukLXoOqv+r+P9ZhK5w
NdpyU8JYO+jb7YtZgAxzyzcFCDbQufpJ7KVUck9O02+yT/wJZ6nOEslgvu7XaVWA
XI0O/MgcQL7bRAp2mtqYkJMpVWkZ9O+wGxkBUxUd86OXfq56EpUmSbcDUtai+Fo4
sG3XhoAlFKi68zjESL8dwOHTGI+zM6elMkOuLDdoiADsPtMphmepxfIPOpNEKOQ7
W/h7lCqCxDiK8E/YEAVLS66VQt5/N0yJv2TATUkw1vMXmGz766r+jELZau+/Tn9E
I60TyY0QNZUXYxhkPiXz8xFxP85u7rOHzjsDrCFEdnno8VNVKhv2U33mU0J7plpx
1ehrs8RkN2LA9a7d1TZw6jR5+nlH8GylRi2mlOL8Gu+G7idxnJvb6j15/DSl77+4
gjJ7smDHR+6JzTHVgNocptMIPSlljCThP7S91AJ8BhgVsR86aj7YpBL0ZjbvRr1t
2DUNXZNctI6FcZiplUeWGsCpKy4LpCG03b5YkKAedLDget6fY8hvvTwPLg5lNS1Q
gCuIqMB1AsYD0eZ9UWYJAPTNrGIpC0y5WOE/TlO5L5zDXSZ4TjqakkKrSK+Pz2/I
iasErQJ8AiQLmBKhUBDWJqw+UZ/CiPvFLBu0urpV/os90RO/WLy0MjxrRpF62GdR
CH10Xkdu15jPaAw7QeHP3YoHpFaZQHi66rNbCtcBzb41oB3Sdgpl/EtS4ZZXkuZK
pW/tueQgjuwqEzfz1KmQrz+da5VqvpxsPfjaA0K2Nm4Gbu12p7CA9/9n8t/bn16Q
M0yk3Bxx0on9jEBQ8U6lVO3RBvZ/iNqR/LZFM+Aewyrfhb37zgekgOySiDs2thWY
yNICk1/DC4zSk5Zpo3BhCw==
`protect END_PROTECTED
