`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zJR1Ax7KIqipnEjnIErhbk2QQIxCnoT2gUQ1nCSdYmmb0i/DMWb4e4tRJLUTacGl
MOg/O+wPTH2iQ3Z47W01sElAl7BCbbNN3G5wlMLm1IrXx/XIBm/whGhx34gOm/6x
aGn8mTyBa/BHmp0Zr0eYWKhuEmilt9PGqJoO7v5ege13VyCOm7dCSZSt422uzexQ
jHnPn1NH/Nra8dEUxrpxKjuYWzQWQYpTRS4ebtqyqvcYgabX5UowtRgVdQ6muYqh
LYU7B3a/R0KKun49pVi3jLe+kC/CigRXHvD9qmdPUf2n07o5Z/ZlFrMg2YG+VWhW
+mP0Pg3od0MDNSeam9dAKSNEOvgSUgFZtY5bAdllYZx7uEI4BQuHkIUs6UFGHzXe
jCb457Rs1cRKPIBdKaFvKOHzKb+Yn5CGX4PMO2+MFn9WKKvNnX8Xh8A6unsSIR99
`protect END_PROTECTED
