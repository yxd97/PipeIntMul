`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L9iGFnSWD8U1HBN70AGHcRaeIPLXv1z6BpmA/2jDeHAa3OQmflBTGBkkpLB/1j4x
wVLZJxlsKbefO8wkEBdGfyhOVSg8uWb/i2fdE/SWxdQzMnvas2C0Js61gUHpjsfk
tiW6jZ00awkxhpA8d8mQ5MvIy/ccBE+b8KOMHfGXn2+uG4A1Z3f+BIT3Rae3wdfY
A8ODy2mHSM79YQxVZbeoUCCRhtw1wnh1hE65eGPSjs+LPzEOBwbaHzXqmzR3g3VD
thnhBRAm1glSPGTWztyGKMnDkgV6BXCpwYa0UVVeXJ3McD9lGyjvVRNS63KSbHw3
ZQlrGtl+LCHNLOE5sJmNxVfpkrAUvppTAeqj3clw/n8kdYp6hsWir3fAYLeA+dxF
xh49HfmOimxhoM/KJo2hBNmVS+YLvb3/g+D11NYQYuS0KhtjOZydHk25sIjmMmz0
vljud9//wbOhbCg8UHLMMw==
`protect END_PROTECTED
