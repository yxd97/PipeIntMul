`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZJSIJl5ZV8qzlfo3nI4Dg0sxz87tE9vVfSwizpIZ7YAJEJ9m0+0crJcL10c9yP7
F4lH9X0Ryl5pDDm9sJ17AJdxZ7wLfwCTLEG8J2/aukwMoBtgw2+aFtjHWsWDzlNB
wPVwspPJA+ILD0B4B3Y1VP/X6GCvbfv4zwcuKZk+M5MD6zyEaO6Z0UFd2XHmGs4G
pW8b4p/tS78ChRaNEt0LYcaihWfgj2VtB542UL1nZE4IqDRVEvqiPRPIvGirxMYR
BGQEBTt1LCcZXzLRmRlpNQU6RGkmszOJRcKnZ+RWdrMX6la7JVIwNB/RxRXPe5jr
8yb7IMvbe+mhaBiV20whjffUWo6ghAW2lvJBXVnhIyyebV450GMO15DWl1jvHRza
okG+xq9sZpQNcddAoDlSiul5Hu77Xjup0b9SAcn5bgZc8TO6hcqLL968d4bNTWZo
px2ENZ420/O4wU/QfQhX2BgDWn+0zT+ro0bxksaOCwMVg95SptgP72uuLv0M4Z1t
JSE4uVBAQtUuSsslK3qIByzH4NqF6l8q/xPzBopsERHzB39LSpN3qZSzHhWFS/l0
+gv/o1uiIng6C811rNWIk6Utt0HHsIUJJpcMVVcc+S4eVF5lyOZMmYU9gPZt0tfp
gILzvxxQrQtWuLvyAO0I8d+hGpYHc5ypI1rWNCc6uh3/PDxUZRt93pNZTSeqEFvn
uollIiIy2nzHib6ZawXZASPgTiU3pqZ54ahtIlLd4/3qTN0sUm3hmD/Rjj9gfG76
VSWh3oM/vm3pmLSLudh1kbaUErzszPzfEmhmt+bQVpBUKdw0HoCBUsvQdSlgoWzb
q9OVBU8LsQatZSM15udiNA==
`protect END_PROTECTED
