`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCAeAfuSv324KQhjLXe02n/1c/KWvKZ87F31z/9VX4kMfgGsfGhPoA1VYkQY3kyh
CgE/uvOXEIIyFbz7Rb2pdiHV5DORCrFn2xxgF1nRbPcD0vm8f/2WnJYfJdDikzE9
nwcnwl6r/T203rquWENxvAoEaRUkkTlkNLcAuj/Zwh5aPu0jjzTDXkbRQuK52Man
P5Br9jxFdq36h0QHxTJ2A6u6aenTEwmopIHcdAafPvmuj7HKmbGoo4RQaGlaiWin
VD/Dpba2t2FM3WoHo6Hr4FmfdnFiDRB2cOGi8gM9JcQFw0NUpERmCgq6m5bfFVKy
7WzWinrurUh1J7iG9HjPgwEoZ574VH+tJB7b8/urgZnh0G4JNoBTi/wlyaRhCWir
2ml1TqJDojOFNbit7Np2I+SajA5biIycmDQwGxZp9rC0tXwkMzJQCW3WzlIjJXi5
rcypWRsMBRVsD++9S9fmDthLw+oqidAEHmpx0hraGZQ=
`protect END_PROTECTED
