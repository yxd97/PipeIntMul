`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rr2F5HXn24cy6hp/e1NVvFjfw+wEUjg0258LoDvAoZdG2Wp5kgJ0A70wnE1L7dE7
E9YfGTWz525YmvFkmv+MBIi7zFHc5KcWi1sjuqWsYuC0RnotOc6Ivg5+3zeuR9Kl
opYe9r9/tVg6eWHOL7srdaUIMF8FGqbtFEZL3orY4Z//LPPk1A/DdJtYCzo+ccp/
AAO14dQx4crgyRHSUM4lMlFCYS/70fV1HWK2ko+X5arj7EJjl3WXCm6E8/g+oYio
`protect END_PROTECTED
