`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9ELU3LRxI+of35U9/hr1BKk/+K/DkEzJ4TE5BeWh5g60RsfdIgReUsxAGc1PNms
oUbIyZ6OLMZHeLUyj8jBdQiqOyTM4cqhaK8u8ruUWlfqGhSFtaddggEwHOhQhQGl
FRoDheF7NCRL0PiR+kjxDLpcFWgL0t+FQTlOTNGEvSfA7UHj52m0pLtr2D+o7R9x
ViWzQBaAl4apwgePtFtClxhi2Gzr+D5PL4IamGO8FigRz0pGFP5JE1iMwudIy1GF
2FaAp3TusCAHDoPGUVVGvLMKJcD0rfhLHYqTvEERbWj4o9fKWyQlzuszMmrPjEW4
97NjFzD+J6bYhrn/rcsm7PK1PFM29IeBmkL6/w4RroTJYpD5AQOta0IHXkzfdHPM
`protect END_PROTECTED
