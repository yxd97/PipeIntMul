`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ffLRYhb1TOYTVPC1mXTMXSew0JOHGDlfi7ZLp3Y/2YcYYPiPIZmq5OU02KZd172P
m6kM4+3+ZlVoJfT5dc1qAC09ym39L2a6FNkityoKdcyw9mEpYWUF/Od31oAo3N+S
9sgnHMJbuH2uPSxFCwJWXN/0u1fQPXl7sE42/3FR37xm5CDRECXUvYF5Dma8xtM6
5EFHocBqlkeWfnx4BKOprHnq0+xNT4Zs9XlKoZJFZvtisxOKSfiq1wZa6Vyf7Zp+
dDdTOBKeJ3ld4TxuV57LW8eJ901oFKZXGcXRe2+nnYAsTwlbrjEuF07Y3gXHUkNf
FBw4ufqBigQQFIN0kF8a7FTlgmI3LS5xmyKEIW5yLV24TAzTNPOXYbcBclBkPDCH
TJAW4G05Wtpz2GkQatXvk2zULAUVBdoyOejyQrBCf/Q=
`protect END_PROTECTED
