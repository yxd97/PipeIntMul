`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J/MLYG6t0z3kGTuZ2V/Onbi452SAbBiijj/psXCWd2TFsymZ242vic5OcDpBq+kx
m2lhLodkJoNE7p/BAzw9+zbaihwbApIC/HlaQdSwwN+gmd/j/HSVJ/VOeX6+V3Vo
B7/O1prPOX6TUcQ4NZ4+GDaPqlzC3iRar1nn9YiCnsvClRdZvD6Y4XLzZeVPKCyX
nEAdgIOHbaM7AtcLl8iZTiZP0vXAZcuRTJ9awNH6a/kO2aNVVPikowwqtmMAWNnm
7acL50HX5OFXBSBDkFy19t9qTK7PwUdNCFLGOG1GrcLL+Ul6NvEEltipl/Qg2IbO
h7DN6WqtdVati9g83p32tkXbfJ6QeD464axFFiGVVIiRW/dKqtRGnOWhwKRlCYL+
rWg4ej1tJGrITs7g0BLpejuKoosMnSwHUr/NAIXUgcb0w1AVpznqK4ear58pgw8Q
Wuqypw616hSSHhg78Q1cUuwYuvKJKISDkR5dTJOwoNEnJU1cpG1sWO5nTHVo6fdU
iyVwO5F9zl0+cMWgswWOtuoJvC+6byQw/V5HIREGELU13aPWPcL7AnyRbDgxrqMh
gEAFlZGd++bjx7cPYLaq5wTPRSumgEOs6afNmnrzzxcN4fFK9v6rEYmxibV23+dH
7KGrjaXIVjHJDu1NNJ6IHbZP1m9SMTirzTpXfSxnXZGXYv3jn3wzbhsCQ4g8SHpG
h90jmS56+2mXPn5k007fZ3MuO89VPwyI1MoXJjhSXvmpNkbufK32269zrFVLyWGL
oYmCGnKWWQ9oGiRjXZNP103KIOxSVlrSnserWuC5PJt6lz0GshCe98yPXyM1ecs7
gX35HALZsS3FVllgDCIHw3zW7u8sEtshhwXoYTMg3+a/HGgi5O3mFTxBz61z9pxB
J/HEHg04MNd13IyuYnWXrhNG+hgR4z7nAZTWWqOxltTdQk3di7ZBT8TIm0hUe2JT
ky+hg1zCvLJZFWACTi+hLCHsppfPfOmXwrjga6jBGtIJ50vlzix+EL5tpYTNQKi7
T0GZUDrdxPp0w4qcFFXoZozCcaFi+6nSe1N1n05wzPxgz7XOBWLGAOuFSDyZEHec
bt4edG6yeVmYZNaHEXTqpDcL5xrpyMroNuHFpsEeikOD39BDHku6kh9iKHtxnNAP
rz3ylZmO751y28MmAoyLOtZnOneMceuReBOayH0isR2AfrnYXk2tOswXWqWxjPQe
B3YLK+G6R7damLyfH/HlC4oY7WFr9upzsQOtGZPpQNXDQbWo1TB+g8QOOiZEW4K+
`protect END_PROTECTED
