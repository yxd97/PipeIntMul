`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tXxkN7AEnPKft8GLGLBVFCBfhM5EmPomVtvZp3RC+LLQ3Rv/QYUMnF0/LpE0ygI
B53c+qjDYBnJH9duR2G07lQPSyXQ2YqOU7RQ8LpR2VqHLphVYbd/bKIoLGoOy46S
9awZLF9YHTegEBSIBmcQNVVfD6sd6OwO3nx3RpcWQ1Lfgh+YDuhYQUaBCVlWJTi5
0thKy6IZ5W7gCT190RaGMbRPYQITzfAifbIdcsVkiERzvVdB9T8uoTJlGgNq0alq
`protect END_PROTECTED
