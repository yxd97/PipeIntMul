`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNkhBMa3PH4c7htPxojGR+eo88iXAoe05MtftZ1LH6PwFUB4jKfE+ynbM0bIFq61
MUdvLXsDCH14sEqw8PRLYnw8kAHSSHTJQ5+eQlEq9Hpr1c22vAifxHFJvDLt+ucp
T97wAXLuyONdbEMwyMwlama7evwSte8R8Aq52AvCbikB/2LWhHdWySwA68BhO80z
t4x2Yda2NIV0pW08DZ3OFGwbnVvA39CJbNLqKjUER7glgn/QiUUzke86/j2rp1s0
N1cOygKnwzUv6Q7v06piHD7hj2iSFC2HTxKcZBQps85RvMLCpU1Bl4ckTRqGwPlP
YgqsS92LylNtsLVqdu0n4w==
`protect END_PROTECTED
