`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4RWJYkGYf0XgmohfS1z4v+D2hpyw5YdHVoXWNFuW8tQe9zQ7dzKt74ZI9kl9rLGa
6PMtD+/ZNqBtShS+r/cSRfx5ZKW8S5oUp9OlUT4Kp95nM1yC0KbU5Qvz4E/kJZya
E64MByUN1FcDxSLOw9f2YeZBfVXHQ7iFP8XMw6D9GDyZvNfHk7rDxaz+5ZYqXS5Z
3knYdSp5KarP5A4O0+KBQ/0DdhV5l6PeaT25swJ3M2ezYjNjiM5COlFAJsJ0QQmP
60ML6skDNcJvCCC2Tg+umSMAdx2wdXtrZVTWPBtnZrKRqdCV7bMiFd2oDwoSHcw+
orFNzgwAvh8p/KTPx/HUHrOFv5N2mEr/qlxXzD6raTv/UfHCGO4tVOhNotYqkNhe
mAaTmFRH2wolOdmhm2NpOQFeCRYTqhVQmCPL7LS7VllACRAdiHYVwhAkmNXJCTiX
p5Rg/l6XPBCB4PooFDM1MEAZwx8GtMuNt2zKRBQK+48v/yf5ryg0yqTU6U2JbGQs
F2cjw6vRt76Op5NBfMDYBg==
`protect END_PROTECTED
