`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3PivG0m3Nthv6bTy5GhwkmjakIwn6J4qteJv8wHCvoaLG5+KXqr79bnS3X3KbFUI
r0E0MZNxj3JPPFBHHctCj5Uqg6dc+XmFWBNIyj9gm2HfGgNXyJqu9tOv3JyPhsOn
svrU1sk9DHLEKTF64QGuTCjFUKQ8WZXHDEmUdNF9IAeRIyrMziJviDRuZtTQNV92
8NOI4ZU0OgR9bnV8TK2GCuZZjQ6GQZc0QrNLrPGFK+zdtmF80YxQZEwjQSVQZM0o
El1C/kvDYe+diozw/E8l9vBpRc1IyJ9vjvPNwYVn4Q6pe+jZxAm19b0fpFn9bncV
UU7bE9ZYm6VmdhB6rB9RFfJzj5HrX3rtDh/2G/KDyPGHrEMOJKLjUsFM4aS+RU1/
2+DyQg5ndD7S4lzjHcesd1/jt36/hNyfLnYppOy6AoZZGEfIucmfINyy9Y8q2zZF
O4GvNGV9MV4pmPV7Ir27kk21G1RzW9CasbQdFha8ZFCozpUMWztuxBq7wXFTY2Cf
53h+w5dGMuBhGtPJxqIDY2LWWEC5bo0dst1OLeuwvFsaL3iTRVt4IPeZwwVG5Vqq
wCYES1eRc9g8NRMl1QJLT6Fi7BOv/vwBc1KdGewPYXjWOiraX7F/oHDFshdgeF8E
ZZ7XWuBEzXKwaju5rPq1c9cmbqMrnv8NJPvhs2b6I8nbN3cHMZsezjZDVdm5hb72
04ymljL0o+k7CBdh6BKVD1F85VQH+1V7L6y9FrOd1snrQtBcuVgWU83oIeSxdS6U
CZ0ehbTaHnKGKveLqP2upbjVVqAqfGdp/i09CopsI6yidd7ny6YNELn2K2iEeP4F
E7l/7GGsfDcDfR954aW/2rccEO2R97x6kYKIGJtCPoYgNuylQUnWyK3ldynbgG4j
MmD4vXfomc5nFhDatjGq/asCwManuZ/xScTzZpPoJ71iMs2JT2qBYt3MVyI8/Mt5
XDM0N/9k2hHUzb2zx4/gtGEJXlA7221lNktpv78Lf+J2C+Tmyq2MItdcnqfcq9vX
3x5v/Z+F3BbxrpFVibsusiAST9R7qiBMZIY0YkoZ1lPGNRN0A/aEgGOIM1h1YiAv
mlgVV0eccX/gY94CYplLMK8/lBdJfzWYNUpuwMSRDxYyzl1AwqgyZTJaRi4TNx2Z
9LfItgqadGpjRDYtaqaWbci255pVSQbCjWxqImHSzGCgWBx02nbrcZnOYqQ2Jlu7
vTEOyfn0IUaCP3cup8c32P/3TPk9rG2Gxf9goKtyooVBY8VJ0ySrK5Zx3HxkKTbQ
UJo5h7+eUqS0SnhYE49eqXExDCrZcvpio+5HyshQr6nGZ49hlxQwUY4ytZecWgAM
ZEbAleXa4iRQckAGAy+Rgs/13VGmiF7pdl0bld0TZyvNi3M33+PFZhAZpjcCpyaS
q+qtWOVma6SReoh2QVlo59IVLBr/0CRcmegoqMZ0/+FVisXRTPHhzgS6eChpzONq
y/czLrR2R3NkGMk9zYff4zuB+UyVAOTSbrjsYknj+eABypzSS7rJZPLSmNe5wGqP
i0lchgI6VRoI/TQBalATYH6jQozGGsV8u7fQo3pVI6Yq4wav51aN+j7VWzLmxwh+
fOlzyeNVyNHfuwxl9hxl12L/9XCSZuBszc2odNv9bhVYYopuYZfliXqdJQ7Nr9mZ
538dfxqy24vSVG/8x6DpWDCrmjfst49AE8IgJmhu+0TKECI4SUjJ1eGU5mbzj2ay
VI4qcEwFynSfzZLyshIMwpItuuPuRuQVedpgLYGXrEGJ+b0VyVxkSH+CzbbLhcho
yrJfaulzbhaa99JSQBcSnSTHea5+5WXFpt5YohorsVTfAFrVrZibUJ3oTF83bKUt
gjFpeDP4U2DQUOn5nXCcPyep9fPo2f2TXh8FOj5Z0l97LYim7zBfU/iSOi6uYSCT
F7aRCYWeRKjuWv+sNAF+QyuxYnlRUK5GVvyRksny4smy+Fqe4K4auyfUfqpZhDT1
RY57WhaJ6Y8zM5jRBxojOpEnBmYgA04UIZECVPVkXGQTJt9Mx7t7B3abIAJkj7OI
xXFu7siLv/6/B8TqS8+qv31Oeajg3e3YxbX/5gk2XMh1PkIjHBVGzR+48lOhjIgF
WmO1bpr04jlP3NuDBIFz12BvhgSoJNEvkaza0iPhlWBs67OOEXYuffyd8UwK80Nv
3KPdnGwNTiR3pHKCZ6LqvB2Fa8XIMTf18BsuIZHQtkiobYj78HsXYRNkIsbnkXK9
JB/zLpdhDhlg+rbSVDNsy/Ss/SmllTj1LehlvuzxVJH0Pan75c8wj3ZN62vV3pYc
sFuPKGnA+7EwdW0ZQs5XRWd2TXKIve8uLWirifEq8tLoNawVV/iCRhIOb+k06PKT
QKaCpV3kLX97g3fKvyyX2ap/5++b+qjqwbTwwmjd2ZFlvEJ74l/jsnRi04VNCeKP
IHjzKoVt4kTEutWWqq6bh4mceRGVAE4+ZFr4LPWRS5ouCnbUjI7NrdhArE2pDaJp
z5gI9MM8navqCHJ1ZRtissB3/JRL8xfPFjoKTGPBt79w5HTIZX82qW1Q10c17y+V
GKPkT2QfwkNs+zHl6hp2xGW5r77wQxvNcstGeiRM9OkfttzkQEhThtvVIk/lZMUe
SU4q/kZca9Ca2VwyUioZrLJ4sZZ/hscVg2y4QvfViKYvLQd9lVAIf5SGoyIGhKMi
cz9eqactnrdpJAesB2diEzwEbZXGwChDr3MWJhOVEnbAx/jCn1J7fnz/i+b0zs3B
gL+Dv2cwgjPwQCUFdVwwwl+fjCx3goBJ48MQeThtoEDUGycO9gKGZcSVdypI3a+J
sgguZ0Am1HjLgEaJlfQAD/r1rnWCB2hxWkHZMcFmHcIRAirxja+9sYieauPMVCkM
VxRJlPjL/s8Uru0xmQtmuZ8fId9MTwvF1PB3p3Z40RzNN+3Yjim4QqE33GFzxbG1
DgcOF5M9mvkK5vrBRvTR3dMimw3WzH34g6FVlJ1i8D48UZC3QTA3NxzL+sgdDA7I
JpN/IycWKPqgyIhRnB0kWifYWb2CRPskotaSyyWXUIiKkr0fjMUkPeT2nJh15mOn
yoOiaQeq4ajucmQzR/zhLB2Dg6Kax45ffmOl9GZDIaz1ofUozX7HA+PDKCzIo807
7rmQMoQ7fHJvG8h2RHNGPGLMquWwziZbKBjlEAe/vm9hgdwg8mJBSNdDBRRSRE39
B9+aDDFGlPB+PZs8mvxXV3oUzHXKbDTmbb2jeLCAA6OwPWr7IeqDZ3Vm0pAFOJ/7
+Ed5PZHVCi4uG0p8nn+UElAMaXT0yFWi9QixPL08wMSX6GVVftuz9fyrfAiv1k0P
C7RwqbMNAJL91pm0+l9xtmQRZG0iR6x1au++hgYqheHtCwYyTR/kUWIguUmJzyld
PoyJ/Iy+vzcWG+93So4wjGEa4rL8GKlwn6AVwtrP/AnB+ZalJwV7ZvVe408BANBX
ssFgwlZB/Vzh62nEGgYdjpGPIASQIpB7BffznOHm8mZzU05SApP/pKvc7sjfZyvR
G0dBQGJwyZ1b9KXMOeJWlxKg0uz3ZNwOnegoHgbYb6JKNZSdqI26QeyZRLnJbVO5
kepX/rS0jT4+h6SMZPtt/Hfja7qPZEv8Ig2PfPsv7xKXx3VGhOiVIYuEmEHbU04j
W5vD8gaimQOcVVdhoLdfPrvyoMf7ypGecjFckJNDMguu7cRVx+iqnvwDiUkppTZo
dyXZvt9r+sc+4RUPdPNVF69SL5XiDAUDJQDeAUDU8wrWNg3MwVQUhg32L/vey10t
A2oDEIlIayXHIkdnILYt+46rPT5+VI0/uXcNTlNrG/BI8spcOMU84NoL2IAI25tk
SKJmDR4k/wHPnZ+Lda/IlExBBU95NJFJKXd+cA3JVtjUyWnbasxTspUz1Vmwz4OD
vcXSNjQMjcSnDs6dhRzITEHNHMgSgF0yYIvqYpbRVR6/B13iNXqqvbAYjA+uGCTT
pdxZSXyYXsoqr1o6cvlGHCAIPD0vsfEdnFS69971yokfUv1couOeUzR/u4GO3puM
sIEsm8CjVlpDvWxoUETJkTF86MzGyrmusYy2MH2annDZkbihjV+Xg5Prxf9/fNII
i2/YSb0nThhcxiIsyqpUf51JiF/q8lHIAsbQstR2J6kYScRurmkJ6seRoiSH41Nq
H6OHlWIlaQldcO8D+NPbThaEv9+0ww4L2yYvSOCs2RifUY3QHv5Jd5VdDdkddSLc
S5ZpPCQMxD1qdzZyUiVafMblFJb6skdLYHRawHuFIUbeRmk5MrhoNXW/1VrW9Hxb
7LS4xZ9ythMaowxic6n68JIjxxBKzbNIKPIV4dqnKrt2fa+WRWvVPhMQROza8Ih+
aqU3Hv9/k2R/xsR7dPs3OGG7elP+wAv9EJ57n+ig/rkueT4J44VcPjYSh32Sjy0T
5ESpU8HvG5zkZ5L/iQDixI6NG1tiztOqndRauViUx3OF5AUJJoDc0pv1YQDafTmB
+mQLaEY2sPtRhayYIzpSyZX9huQvCXvCfClYn2ihNSCKCvy/KsUsU7YDmS2yozc8
LB2/WadSgmQdafnXhS1mX+5rQYR6AL7QLMcxuOzxIS9YEogsmWIf0rXZxlEc56Qy
jGWXe9XWhBEwMPxSFJwiKcu3JLtGBcNLwugFCvubCu4wyp+h6nZzs7El3plVhyZV
fBf+0mE5MoQ5tob4pk/xPLCnpMSiSVX4dQVZrrvL6VLeULcwvwi4f4lf7NZMTs2k
q/65QRfmwk3F1lY8lOt9veKcfs09SO6cJM+ePUoXrsRvKcPElwD66ArHeAUd7KvB
IPH2mAwI8JkHpkI7Vaxs4snYepTLrijkDoNaWUfQNeAfkJUQKagcp8FuXhjYwrBs
qQtsrckO2W5Yq+JIOE8taYqxVb38pRx3d1FRGF0U4Fi/BexXsh2HwllqVqb5dU8I
0wnxLvUSLINrLBurT3YCf3tU/IklsGyv9pkodLIUnWDjrWakR90gQM/J+URhdbu4
i//+PoVgQN0eSGswYO9zDEW5i3UkUXlar9FYhhZaSSrVro1s1tDkCXOCwPpLSR35
xspGMQZgMpY6fFt+uEbnLJF275umaayuLOHFHGUqm5LFfg05cJH3joklwMNYo8iT
LHYE606K8WD0IAQq7564jjJCtbQxIHPV6+cWGuhXqhVJWJewHX8zWjUCoMX06UC9
z73Z6vv6PofX717nHMW9r8driNVtSZQavXyppfIAQ0Lvm6xI00IcnTH4SCAn/P0E
TJ268Vfk7zcYG9ES+GaPgM3dQ77B10lQR5RqIfR2JZ0m0+Qx9mllWp8SEReYPWgu
C0iBW+neUSXVVLRPJ0OX2aCom0aHxl64ghyWxHiX0qVb795BV1aBkVI/Y34e+nki
JmwXY+F8KY/5lNvDpsmKVIIe92Fv6nJl9DMSqN25HqU/Mfe2m+Y9PQ5hk6s7UgxI
TU6RYkVfB9W+J+kmYZBt7WNY467BKZ7Cm2c8wH8uECw2G59FZXCgiyoaXtyzMrdZ
OZJDAo/HDqpy+wbsSpoZz0kRjGxJFAgp4OoUPjy7fRGQbcGj7viYNRZRti4s20YM
a20L07PWlFqUVo9zyQrc5wWkXSR0NmavFBvNG6+P8swJS3jhPMywGjChKFKS3ltw
rkaRSP5U4i0M4Au61Qlx68z+Hxu8dBn7qhQ6VRUj/cU4uYh+542F1nFungCkkJk3
iPzfhpbBUN2zFZRwWpav5Qe4Qi8sLWQ+8fKKfw+tjbDcTg4iqN2DwM81tH9UKIfU
CTY5VJ8/ADfWpgWtCn4XsoV1On0Z/NIYk/e+xjfhERUa9NAiX7sRsef9FyZp2azo
nUbKk+QFBKuM5FiAshzSPaoZ8c4Hqw0pxc4RxdriSKwQxQWfKiRNhLylIFTqUoUY
ICPvGppsppMTqtuMkv+MzsNtdNP5ZQZG6H1rg6lpWu7fTHvwdCbO5W4zrLM/Bo3/
T6ULpc8poOA4J5p5wQTrAyjbv/YR00xy5vbYd/gZiPQw9S6+lRgNmAICZWYsniht
cGzbBF5/aVAsp21aJWQsaZfrojvE5/DYg1SgsX9TbLhEEo5Op7R7qTmXlfDtigvd
vsaey8bmVS4HRosnkS39h60seIfX77ZCYVZfx2k7KR8t0oNf3q4xirAa9QmMDJfG
pVShkKlinsND8X5zkKuHSyfeTpqKZpObhS7JeGMcq1ZmPxFrvzLfzuuGA8PLZm1a
Wm45xw6plQfpBd15sEKBCg2QojIESi7mNB6Hmu75i1U0radBkklowPIu8xjzVsXA
46iGmuQypvm2ZHGOPZ3T3lKaj0xbWgrI2uKLdQ3+0s5fgNo7r4kJweVPFHkk1kdz
y99xONU3mHulhaLPlMvdQwyiwLWEWwih3WKckVse5tHjbRZOfNnRom4s1KnM8gKP
YDWfbKDvUst03iHYzw5652Elj3GrG1u40G+45W9HcHoKmyhNe1HUTQjfomuB4wn0
exmC7+l0XS/gi10l36qI5Bhkm3i1QGOBPVtIQ9IRh6fnVBIkzogSt/MYaUPyTGOP
Nfo6CtvdL9FWVKg8K7PkzMwc4i0NwEEBKkKG8SeRd/o8wiKRel5Cnz86rLFeqRWc
UUYWBYDJ+bE3wmxx/WUcPGTbcDKQFv9Aj8VfTuMu4sPkG3wAkaBgThn6xPioQDIg
b63JZKLmMVF66DCT5pzGLK2MOensnRSuXdgxrOaIzO/VaYQqMlPh9Qa/iXUHd3B5
F90zeIkjFvSbmWHd5X58vb84o+ZJjEqUNJnB7vPU8ZRd/i2O12vh8eEsXnE5a+12
0it6sZtxQpnNSTcU9p4Y0ymhE6aXh50TN6amdC4Efiwe26vVuIOqVv9HSNXyLuFG
fCkItaT4a/QiJW7lzuAJzGzftnFNkyteOiZ+W4NEoSJbLp8fLTbm7iYr3CToraIa
p2TtJ+6+nM0qB55khkkaLMxswCxUrK+BEIwkcRFtDFISBDftiE+yQ/GvqWJ2p1md
TBNZG0/rOu7fVhI0pCpWwuXAfge3C9yAoqmXFjGGkX51CyGWASEixCBN9WymMRRP
FpeKUVoo0hNv3a9ZbYolVRimsZJW9mkhQZY/tR6rbv5x5hSUXw3WUY0jBe0FUzpT
we1MLTJUAk9crwpPyI21UzY9UY6EkCCS4XFHfXmk6FB2gZ/PRKtjCUSyGmYYBkz+
lEKmA9loNjAqN5zsos+yw1N0gpek9nBaASMJbNHG4TAwbxzONti0aPX43cAqwSgN
rqvhqfqWjTz/Ue0yUiPOxjtpLdww2DYhD5SS86hwF4b3Fgyco0X+0kf9iAInFnnd
jHvQWT/CstG9fm0U3fIatR4BNS9+rRRQ524P4rvRb0b/LaYnWbOFtltEYUDad2uK
/mAvpSqkoB/W+QbYNPxps+ieRGAB70ENrcHf1bzP1NXDZO2R1vwrd6Vl3BDsei8Q
nhHfh4IpiQ4FKzzJ2gkJao5YJGymPndl45ctUckmZnfi38IbRotTOP2kk54xiznP
BVdeaahH3BjtXAwS+U+s9IKQfU1yfeyrK2exfIoafQ6RIgc/12KZmWVHWdNCXPsd
IwJlNz04UDn3WgX6Y8i2t6uj2NjyhxLmKB9viT6bDfkeb2E6K43lDgskLYRiCHHt
pfQpSLKCo5JpzbLpGayLQmKp3zaihXG4uemhAjojNCVymNLux+DMfO/VvAs4I5IX
+W/gN0hVmE1m6qKTRVAUi2x6J/pN1syeaQuJfIYfhF+P/Acds/dpnxgh36noR6IL
FwoVbuo7QgKkaKFw8DmDkduveCe8lE0vobP8/HOLb09Wzp//Zo2H23WJEDv7WIVV
5o+2ABd29aq5qgy3X/HRIpgZEVo6pIG0da8IF+ViP7iWdr10+i2pzZ6u72XDzgyh
mDICTyaKr2aHd1lh6c6SnWpZy6Iu7nibnz6VhbHSiv8fPiuxLa/uO6R37XH6FdwG
m0yYkbzyGfZEbTU9FEMqo2lVoLkJdz6EyWvATbkNlNFUQ6G3Qb7o5Kn2vgXJu9e7
gaTYwuJL8dp5vlSuegLPvz2EAzOh23Z46LNFdlAQYBLV98/PL2XI8s5lvmZcwvSz
KAechIFuD2mDXlzOusDoaAEIlYLp431KwgudN116n4yF2IWprFQq3xV/qRkw/ySm
JcH1d4x3/zCTWLUlFSEuMkaBxwEQSuRptWsC3f5uWJs203yVAvSKg8hrARAX19Lb
hLLrPB+y8WD7nmE8Mma3fuQZDqBflBL/DK+MiORP+1FayebvdQRG4qKhIxl/sN55
rW5ap/+cjxzDBfo9aYfpdmccapqCiNopq3bU/MOqUvKonera0/XCTYWqlELpbK2L
PMa4PQUIDkUgNOmD5WudL0kPL3ZoduC0LeJ2DBCxkcxHK5kkswK7+pbr4B04kvJe
tEy6sBjYu7LNjTJO6dbU54xNUFuEPd2p2vlq76IElzFT2ruI6PpSt00uWTMy3UIQ
nH2gE9ELYxErNFIXpGSRP+5u+IlPGGT+VTKvGJEMXbaGdhNxBIMC3aQRo+2zqEzL
90e8xWuljqid8EzSc/7CnKq87gowena8XK4AgUehjD+nG2dAHYULMc8hCXmzIkV0
XfL1yf/9pSK8fJTXUTRLN/jbYkGLAp5LfxXXQJFTDN8NjYeZ9hobWF4INAXZOJvY
Mm7aL9srsITPJ2gCVgIZX4SubBGb9XSyeJKnHGYpYGiwtULzmrddaUQo8sFb1IW8
59gxxuUhYgbPJO8+EBKJtc5Hqn7qyY2WbxYYata9aKWzTc5vQb2VXtuZFbDpLjps
XC38UKrFbZkxu0PbDDMg/aKp3wcQJNVnd3vQnZhKTZ+gyN2VrFsDH83DzczsT1HG
Vy/YilS5NkNozUZjmJ473H4ek4J2MbcGLi0sWs3vAJIUUQ8RuxnoClP9yFetKrN8
kAtYStWEs0UqA828NGFZNwM3qv3QTkxM3egFgiL2TKjaX9XeaNypA+DLl+uKs+43
Z4mEhr8uDoxuufBVM7qS3Brucm6pWq+BJooqvuPjOKpWk9iduqTGAmAPXj0PVma5
ayXiUkQU7/raGb+8jbP+lPXQUp2SvIOPvp93KKSMZ8t63rSw2ld+jxm8m5K02kEh
reifhl1G7cmXLVpsyjykAtPNMhCrhcrSly1rp7Pixw5ep9KIEF5GbXBX1eqHh6nM
NU1XVO7Gfs7oKzYA9fEA2w78ADjpiFkV9yc2XxaWytLmI1s02KDMsBhuBiEoM3Y3
7R2f+dTVBvWKWVnPVWm5HPY3tckwrXn4veSC/72dWZzhX8kLnwFZlhzx3b+zOmKH
XzUXnjYmg+nMrBKaZoU5SRdU5Kd/T6rgQpLbJmt/kAzpoMP34eMCSqp+MK8vC1RB
wo3Nlt6mWIGWU/A1gWyVaQ+MrwGEIKBykq+oCWkpKSoERgKmnXDApAZygiVE98zW
jjXjivSJ5LMU+2/vkzm9F0r08BYkZUxT767jEYg44k1wfZ/VVMw5+rP2jGR9fPHv
SyGMY9ugOS/6bZ5HKoHnEigwD/pWO6lL6oegSFNOoeC6ro+M6e0sZVb4Hjsst1CU
VOLIjwk49mJf657J5jBzO4POy0nfhpd6ZfSwDjtiJk23Ueji4qc81GDsvcqtVRF/
4y2ce7JRc725sF0EFwyfUdMkZXYR8eIgJ0+mUlQCnNpbt4zMm2kHi0veDgDeRROl
WedEYPJen2+Sw43QhEOSJ06xDtleb0Um3SQFsAH4TSBbaKdZvckSFYhyG2vRsJKm
9C9SQuOxJoKpvk4xiIuB+d+noixJg764TdSpDOnkk3MSX7A+cFHXCjQpc8rHRNWc
GIsqAv+aQmAnz2jDDJ3mta5BF2gbZ3059uw4BvJWsLrOVpwV52WNH0Xf0sacNrs0
IJeFU0ttDPkPCGMo6LwIxaDhOPQ3JR5I/61PrO/hLCpnEwEVwsTlRvu72gg+fDmN
SRCrADfUGVAI0/u6R4Fp1iA6k7BzByZhC4aTnTB7BEN83JaWExAkvHRaoTrVEwYr
2MNyiiiJenAgLxBayyh1faBSBKJw3R6E/YQ3MGFeBY0oIOdgJIMI/bSaZaHG7lWQ
/SoV268SVLcn789QZSov2y1Rk+ikxGEyPp+DcopmoW//iN4wG138cjhY7bhCTWyh
q+5pqd5W2IrDhoAhFNIizcGRfDy62AvNdfavujQ9TutJ/uin+1ZhGNgTmajQPPDy
JWfJVd1Ud4pF+V/NGZmqtzZ+jRJTliISHYqZ8MxaiBmmGeL+77k7xWsiXS+6BAeY
XsBZ4CuKDPaIhwTuGbV6Xkd+ruqubhSYf9T/Pl6Q1rMogJvSpkjeRBBFP9iVhXHL
QuUQ4G21sj4tw/7QKUxGIX6YvegS/NAOhVWYyM0F9rdMKa7ikiM5H+QG5I1/pOH9
uWSNMkVBt5bm9aK8/efTZI8V+iXfgezZNIfzDxPXbcJ7TCVY+nT2gjwb5ulPsFRa
vTL6pKBays9aH1Kx3/I3UkaMxOXQY46t5Fi/M0zYnToEX5qPrn/sk2LYvPQclB5B
t4pkzVQ1TC3RLHNGHcWdDp1opVZPCPjFrGA46UMf2a/c96XJAV8e0F71U1cS+NE6
7c85wIc6Tb0icH4YHfMvPyW+l8S6xUnPXQkOzse+p8KjOv6xxsqA+7ZcC1Xud6oF
17/WXeyoYd2ocvJojLYDHmcwNv5UBmx30pbAnKrZpyY7ROAv5Fy4bHFbDCWFqKu+
j789CoxUmwJgdpL2zcRCCB53D/350UazIgR5DhgPN3FQOkjweFsS9DXcWvskMFmv
aY1PGKzhas7f5OuO56iPUvYhurbL5ADpDr3Uf7/NyNzLU5htIZFgBGptZThvhp12
+R+hqYzJ6gIJScxnvwhDDdpz2sIkeDeyQmcFKp7kp/P6undjdET8hWQrs1RfXAGT
jg5I75rR5bJ9oXNXMLqG0fT7/8hRDWYKLZSic/fOUBWrHUUuTJZAS6eTp2VeBXaz
7u021zM/Xc/7tx0jnoMaGGAfoKGDjKcQ9mMcnlhWVH+IWaf6EISxEZtPq042mXwQ
USU0k48843s3UZjqPpAl8J+YUC4n9UHgZdoST1W0o64+r9jGQ4gjSajJB/NTDVNk
3Fn8QHbKy03WiWnX5kZ1jKOIYwNvGocLNdBJ9i05IAosMxIzzEs0xF5NbOnE0N6f
XZjt32ZXV4XJrz+6+yoa+iZYjpi5N6F3lvDZIpEjI1+n9aQ71mWYEd7BSM626+9N
hg3GcpcX7el+zNAHDdDIBdrpn32tf0BLUDJxFOLCsL1sU2b2dFEM9AACt5XBkZJu
a4KzrgVwt1nFlA2xNYhitvItqrtaQdwJcbdLzg+X0Y7BVfyhSQeEctrDKuy+s1F/
F5JgpyZFPhi98uyE1JHQfDbr34jk6/0xfVrSXT9qUUy5sTgwNWK0KkxCZRuWvbDv
RMOzsyM3o/U8Yrr8e0Beeczhi+Lay5GGN3XrwyMl9gT0txcYun54r7cHmcOqGy+4
sQ6/FgC1MgFRRfljYqkiJb9RN1uioXU6rJdUJhdH9BLLS5SVoVpRqTDrr5dOgW0X
WA+P1MUplTZctQ2MvUGSZ0kox643YO/NOPnSTjTVZsG9C2liAOcvXfLM6/nnyNqm
2uXVCKnVhJvRzdeIc4xAdqCrpyvSmpbfBhe34ClAjTu2ccA2bHUbaOvJk4cFYW2x
KPUFBz28II1fZsOXRv3Zj65z6vrdcIXPXdwXHGfjg9j0lYlVEuRCV4Zm1A64b5Gi
x6Z0nh/72M8GHmLFC3u3+LRGSYiNANdz0VdhvQAaNRQSRxpn2xU/NysJm0vMUuoR
JC9glQ5WW3s4YixXF7GF71NrkcwMYZf7sixeLFaV09DNuGU4+NkxErLLLbjZdPB6
Bt+el76qRLuDrWxH2mt15HP5NX520Ptdymy4g6yPdkednPwZykPJDj/VFHxokUqL
X16Nnhan90FGYtrsW2nYTjbn/2E+P7x7dtN/r4lr2j5xaF6McVsbwjfAQJq5yz4z
IRIV9Dr3GtjsqHRNHDApecuJ/oXpRC74NgvFs2FCg0wbcPIopdKIfz1DchGrlWCS
D/+ztnRJ546LrH/owNFmNymRAwiCr+0dwNPZJ38Cpjcu7+lwoBeIr8G9n4lCBlbg
qQKRScmsWvkkAAVKrz6w6gRLkuSicfyRRJGGCOHUMwu0riZ6ottaI9gWth9bM2OO
np+BHA7RK1R0VKU6mILZtzoKBuB9JxuZYDoKLB/FeRW5wBY5JZfE6XphYrAKB/TK
K4kj7Tvdi83GFwllO2slfGebfy7x7NpWFsrVYAsAOVxulGKxRn4P3eOwrzshjekK
9QlOrRQ8DGkNmPyKNDqTQiNgOu1lxajqUOoAKOMQBa559bzg1X8mzBF50NvfP6ik
485AgBJrKSScGSMXIuFB3bOCrvMmA6bGvyOiE++O8Y7c4Pzj9GbmWvy+nIg5p16I
SkFHAnG3RwfWPNnxEjra5Iu6YaE13YL7lwislf2A+fdD5Xugm7aCVU6jjV8ve1UI
PjskK/plgtkIc7aCi8tQ+zQJBflAzuwjdnnudmhb9RtxA91kholoRiFLW5Gv/S2+
nnVurJhqKo0rvV7WDPHwWcEBcLjxrROduZk7/ghGpD8CoswT1inZFOKkskwMLWKI
Okc++840R7a1f0jZwqHbmuSV4uiYDkiUIWTs9W//peDFYB3zF/qrqWtbSmuPU7uI
gxKZyS+8BqO1w5I/kwU2xch88Koz7WzxYIEAjlZYPLy1aKSUjYY9588INZttEdkA
an3D8/Ifyd9WPViNN4ZGxWAfFk6G49jh4q9OMrNMNrCmqIazkSumHkQBu7QK4hg3
Dunn4vVAMDPtDew8VX3YGpacYKnZiJZIkphhTXW6UXgYS8XAKwij7yn1YsbWIW4U
RurU3GnMUaC11XJUS9+ToyqACIMP2Le6Pgm5vamjf/lUkiDCEkJCkuSDsUUV0pPt
Coim8MNN4NUkDGqnovS5/VswnHAoZ26hYMNNROpPXodmpJqug1gUR4x8v8Rl0F5h
wNSL7AUk8FSNNpRKS4lDu8NBNTDD91CEpRypZ6OKprTqKoISj0okORsG1fwYSJ3o
ASOXxnXjLH614yVCox9C3DfFACQDzml4jRdAkJBej5uk4DqWAzg0IRwZaxzLiIlc
re4JKZV30IKCM+5CaMYy+XS2/ADPjFF2ZmlL6uEIThCykPrGdt8XjiFA6/19Cvb5
ncc1W9AyKv054Ba/rSXxR3jbb7E9M6A0M4zL/ICfJ7vl5oSAf4NHD7sjZ3qAXuxq
c7EqqLeYbNVe1oTB6XPKU61O2EQ/VzVGoQDf6sPeQw17aB5sZtzqXqZL8gEO0bX4
7nrv/9yIq3D9X2WJAy2OnLDMRfQ887YXv++hoOQ49L4=
`protect END_PROTECTED
