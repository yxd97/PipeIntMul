`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXuNy35EHuLA9WlgmLEaJ32iSRjE8OT57DpwLG6rosU5A5vjpbF0VYhpXJesxUE5
YEFwkkFX4fagtzDKsHhF5HmE58cncDr1gNk667X3c1/swp8pW03Fv75GmnGHDIV6
HOXgqKTuYIWHQd6BGr1QWUU0pf2Kjy93nMwPbj1NTjgtkEOdNpzZjzBaGbYM51VE
5bVTyu0uuyXaMXSebZsVpDzcdM9vduJJoHspsfIGbg9CjzFTPJ7p6eSUJnhdoZBF
0GCP8FPjlWg1VWkV2KIoPrm8oZcH7HtMoqh8hjDeKuRduKj/Tivw94F18oDWiRnP
stzwWvSLyEeWPNVPMSDfvXC5MX6a8Cm8Tp/MGK0G8nPZLh80OaYNu19AmA4VEDnR
GYIuHc0GNFKGc4EFZE1urAiT83e9tNU+L+Kh1uoRYVzT68j8/m2+533CYTiuHBVc
OPDgv0PY2KivI2sr6dWewQ1+iTP63bwJTLRsvRMLJ1o67TCX7m8QxYBR5OB40sMb
5VIdP8wgsgnpoq8HgkGLT1ZWwdxfEUepeSqmyGqsSjpxic529KvoB0lwAHMwyAd3
Cculvur5ADHowJMv0KzCs7kUaDNlGvP06BokV1q7P3DdyBi6h/x/buQlfT2Jr4lY
NAItxhyyLgjCTy3mU0jt71cVzeqtZuc6JM6zXGsk3d5S0zCVs5rnYIB5Ny3xosdn
7350vz5q32o0oW+jDT7RSNka2hb0uz0KyxLj5rPChchmhm+laBWk46Oi6yjxcb2/
XT6RzUFNoHA9v1Xu/+/qkI2N6FBcSIhbcUQLmZdXzolWjQV6YydMJcdt6vTVRWs9
a2Adv2JCJWIk2P1BMU4S20fvnfNfdtYFXBkOMO5d6+fwaywQhtz2RIfe/EuCvVFU
GghZgF9ld3UjvBMHP9VozowAgCkLch3UC8LZRpNk5jKcppitKPjs84RoBln2OKL6
mwS0snI2wFuXiC7fxB7ZfuFK8/wjf8oJXgvet6HIqZ+6JRAwwlPht5pntPhe63XB
xF/cMBuIe27qpMiSX/V4RTZrGs6y5p0uXiwht4xNqBewTGe+a54vaGmKRvQdrtdf
Zr0qO+aSTb6tLCPddG7TjnfIzv4AvZ2soZVTlsBf4olVX0mdENw6v//03c8aarqG
LmvRpd6MIOFzTq45tFSYUUWQplYQNXD1aFrLefEhlWtCwN2OEg15J8ySr2l+t8Of
A3Tx3sSJE0vYvQzOCgCSIb8r4mXpWdNqW7BTmDgW39/CDeLIFxXt6DAyL3mTvu8+
Ve4gi/TXhs3AqoIGIJEfTCLSLoTV9FrxSP2ZziZ31OH3lBtiFk9kfVA6L6/6s626
lVAL77iEFmzSA11i15cLA6r0jNzDAsLMdpA51eeu96e+eHsz/nMCIJxSZIdvI1HB
nSxd0bAW1P6wNe4zRFNGoSg5AovI+ikEFzwSCFsL8FGkTHuLK5epuPIMUuDzdAhj
aRxHBXvmhqqTuV6O5XC4ND5lrl6g+B8gcxinJ3GvroUloNX5DN7hnfPBb2V8JIFj
ftbB8X6HyVDqKhcG9grzVT6fvqgKFaFAFibeYu6j1Uc4eaPlxqrobWLgpz76dX/e
ljDMKC7idQPG1mJNfFS3jgRWUHTPg9f8ZTn9MinirGbjBFhztHxQytU/DH4YLOFD
9LFu60MkASxrylSKoaPrV/W/Us6fXrKqq4ptLKrPq15Ib7du6ycyM7+XxXb4leyo
4+Aqfnt87GGapF9EEeyqT+aefJuG6G3d7y4ehvgEYNeWTpr1vMXDx0gI/mtX+4yP
z+XYfymrLKR+/MZw8+8tZ8Qk0dSDvuIKK6VGVmEfVUNup27Im72DE0Z/4B06iyVn
TGueCDnWYeZi+/n7GmmXe2LHXGo5G3SP+G89LJBeplSv4T36cbP6HV1yiEd1nTcn
Yb7nRsh2PKWWlKT8M8lIi3X6RUbKqjUvrzZjcWEwSZNLC+1iTYavPgpyziakHVvw
tKQcx9DENkxhrBNBF2CPNZk4SEFskdGVwrmx0csZbMHmZcONpTiJ25t23tHaxTA4
MQI/+Cqt0eyNxuFVgOXgxyCpSfLwJBaLSAg3PQZRgKzc415H/3okW0lrPf+1ULL9
3OOthjPU2TzjNV0Bk3+S3kR3Ep4v2g3D/KETYd9/kraw1wRtykIYqCUdT1ZAG9yv
Cghc2/Q6dk8iixuh3llySA==
`protect END_PROTECTED
