`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rnmkD1V5DAwyFwsXvnDv0YLK3BANaiaVyWks+8jEV24+qGmOVGmjYUqbDQZ8VaQm
Ahxvpf7yRxSzy9VwaXQcMfC4uyZdnuzWptKGbbNjBVnEI2grIf142BObbWQD2Rb0
E1RKOJ0OBFDTNB9xtH3T0d1cFXHOR13qdUiq+RbP0F58Ba7weLD9g3Re5y5MBKan
UJ3e+5X/Jpn6nInN77HQoiUGyDuFdL6hWLQSJb1SmEUjkpQB911QGNzPOJyCB6fZ
bUsRL9GMLTvyyV7vp5RCBTcYNWmXVPXWoxFl3723f9VmGoP7NazDWqvnNFlZRaVJ
uWQY16IxCiBRSNLkkE4bN7lQ+AUlGlOJxiGVHCrhkf1SiphTkOffc24B1Rdqc4on
VtOkNnEYwMnUAQmY5jYnauoy2RZBkQneUNZU/LT4gYfRAkUkDzeTNqvqoqQJVFi7
ikrYo7gR0iWVMGb1E6gfJw==
`protect END_PROTECTED
