`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s1QbFL/VIiB9MxlkBxYRMmA+BrjUod8KJ/M9p2kk1UCGuNuGhOjS009etra8oOIS
BVo56DxSyPWfXD1CnfaqKy28Lun7C5TsVnE3pL96wxwhwnKMIfLPrUumG6FkZ9+m
RTevO8PW4+jNxKGjaB+W27zQpKY+uQ8A9nfWI2h4SZTSgpF1PVVS5J/PfghP7VSt
Eq/MisuzFZYOSwVdHiUc1Kzd/Gh579mx0B6YExlM6DPwdLwicdMfB+oCnoZQEwdT
hSYtzlzuvkxWQJ3MuporMpEoL8/iVPhujp7wo7f2DJrhCFj6Xt2WUq23e0SLpzjJ
Jcsg8nNXPGeTvLwxKYc2EjKhp5voxnj0+dH0RrEX5wyI2zLab435azJOkJukWfA2
`protect END_PROTECTED
