`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kYZQgN7SribnMOGrj1FqSyIaG5kZGytmqI9RBTs37c9+T8QGvXH2LlBwkEcAi8tL
tD+j18rIzUUiSM3Z5qjHGgrRV6HMyFC6G9PtlYYn/2g1oOt6Et7Cv+PSspeZC0TA
hnyWIgbjskQwBdFMfYEK31kC2tp0eOwfQfVzPHONpYhGwpcrwYgBbAJ5g1D5pb/S
TXcr2A01yLwQRz6RaseqtF6fn6pJqSpnFk7tLxglkB/3ztwXE6Jidn+HgcmhnhmT
koRozavU+cYfCvfqV3v9YsB3mHui1eqiIn61Jaf2LJ2NKPNIV3/DVI49kTPAOjuw
g9sD8bE8Y4u1z5Tfcmk8bZdlPMuaTY0F1GLln3rIfQXgpYDcxOWasufUHTR3pRgm
0yRAt/YZQ9mlyo2rrP8EJKoRn6FHLmzxrIrH0vCrWn4=
`protect END_PROTECTED
