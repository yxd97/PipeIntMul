`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2eAeEuuv+vdPYlgii0ZrYja/4welVz+Ujh6X4bEhhjocHr2UvJByM7O9vGlKFbK
zOhINFeLIYL/kpN6LTj8x+qxt6c9AWwKPlANqSfnXqxFgh7mBM78DW+GvJy7BgeY
tJH+f9LJjwbeDHVIZRI77U+5lWVbpr8gxOOGNsLrn8MJNpZ0ERP9haU7hzvWYMXY
ln150vRNVri0Vea7DRfQAtGiq40Kc1Dl4PCDe/0QsKiatKQpDmdPlyQG7z73pY+U
HK/tpQfqiiyq6P/Vnnj/cIvD+4QIF/WT5tDxVIlNhkUJrkEOWhiRjNqj6eHQvJSb
MDA7p9iPCLnnn7p8eky6fg==
`protect END_PROTECTED
