`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ghUJuDuu1t9tHRUdynsIfcm2Vh1WcErQ7MnsogIMOd3Ef8OnjkEGhmyi1cswtRV
YE43VZYLEPRkBfAw5xmYCQulhPPZAqrGRXuLss+LohLincqZpDcrkApBukyScfGD
MBFzffL+4hjrJFL386KDeQ5Jx/riH/nltGL4EchI+O82svOopNwhnlVSZfhFWzFG
Yd5fe2BSYfK3YsLFCa3rit3MxJsT27hiOaIsshYTWAWVsjsdzuw0Wg+Gm3HqjInz
YFf8SnCrc/l7Bl6LJd40ftRiYuKjFSRKgxEp9579vYvI/GsFRQd9SS+SIQi6IBrf
JN/qnCAF7umgacH9wMaA/8CwdluU98bou/8UI+WcBO0ex5ElVN8BK9SM2hY67lc1
j4TGEMczvc7pDQyYD9f3Jw9PbNIZSVpk5iA3iYiAxAC9pymmYck3W7jaRQn2O/Yk
JCowva6UePCeANuZhIgXH0vsutFZY3uogNmu0DsfW6MYE35NEULUxMOEAB03Fdfx
zu1z/378U5sHD2TFo30hYkpCH+ws30cUXa9IJ+BCKRedhvH1UG8+TxYBSgqP8Mfj
W0Y+Tfms0guL3WubsWu0A1ZAEJbnAK+ckbPoMI4Yn5u4dQlGF94uKzQeRRPdMGc7
59in391+FJZ388ZLfC9AQh76hWw1MjggRCIAARAg6RE=
`protect END_PROTECTED
