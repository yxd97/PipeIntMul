`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4mKiPuQr10E6GN1Fsj4MiRUDsRp5BtQU3SHCcJK3j8klY3zKDZkbouMkqQv3FXIk
n9JoryvQA6TwTLMogcKsOal4QMETPlSji3YdIbuDyvxZf8sAhuvWpNAgUoceNfIE
wGL2Et7iEAKU3QuMgN5F/f5qbFcsFKdp3Gf+ncwOj261Zmekxfj5MCwOCfobgHCG
rpaK8NEu/wDnwz7tFOB5Krsni0mJfCRnPM9yb7Ivz7HhrAG/WwyyN+8GrYPt54MB
epzSbxPxtY7FAZ4R1ZtDHjnCDM7yYr4Coz2BHqfB3XJg7agCs/BNsTCsjYrxCqOI
jlwsp1eUVcgdp/oNVc4ZOVa0+SjTfYDsUPgqfuoIgfXHU4yNRNl/J2Xurshcny/j
`protect END_PROTECTED
