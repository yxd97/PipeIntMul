`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/oSCTn2fdqghveTgz8CtGwnuWAkG79yItLwE7akYPl79eFDCpZq57YaohrneCmd
l1WHdrDZBb7wwz9bsbdcswZgly/digK1qhdzP2itHrsf3NF3WmmGs2tdsMG7/oOn
++S5WKxOiMMmg5DLd7fxkU97q9g00X5zG4IxtAgPGpF1uZqp1r/bxZzr2CMwm8wj
YFuhzFxFwCUfp1u861KewHEILGIe6ckg0DsCe73NSQImJX2rirVMIwCR4qpnbfbn
Wu9/fMH701wT8CzWTEIgco2RLhhZLve9MA7T/7CauBvLYe9E+ye6aKwrcW9h0PKX
JTOGhza1g1xHq2wJL84VBslKpBzyKIX7vA1ptj3EOgflZZV8c+mXdXvLGHk0jhuP
JQgX8l3MecleG2Y2LoNQyr1pS/eHTL75MPPcQ5Gdw6LYP3MetKjFPll+nyG/RnLX
d2vdHqhV1Mp7Em03tl33WVzkcvil2W/MGgui9T75I5PuOoJIQmh592USQjgqX3WL
N7PAYba5cNTlXr34XIAFcGjmJlPvkAf7zN42r9Z6DWc=
`protect END_PROTECTED
