`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iajA0Zs3IiJUtED32bE0UyAaawkckJ2gIbeNCi1HoJRRffH4CSw61iE2XbHmds5B
dsJ1ykCVBvdyoJEYtSgr0gtPcYrkSczTnXZEbk2YrL8dPqw+wmoQfMyOdHiO6enZ
hJb2oOlySOjJtqNXH54FuNnnSjeeEKJ81f4MbjY2EQjLdC0mU6pOoSbxeW3eP8fX
fJrx4VjxD6H/Jp4h4A0McaTiDm6gI4CIimpvcSTND5Ob3kyyfeLR2eaq32it3Dps
5MGaURsjdD0GIF7gCTrcpEWjLkZUWOWqbRmIP8sKdV1mjmZEmFePE7RlPv+GS36J
+J1fckAhq4V6xDKE3wXcpZfP99uFrvHiX09wB2bxzpGXRfyEUCFFk7g6SAGRLbWH
`protect END_PROTECTED
