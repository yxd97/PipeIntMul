`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8xxbT3bqOEiYIEvzEG4AUdK/Yammats+L4Nu0kTx6yNDFg29uAygbQEtGajqrJFi
rzAi1SO9vyLyDP6FWPWrQxFq6gGW/cHKyymalN2EW05lsEF5RM+rshJp+YLANcrQ
af6tL4+mzFt3rlNZuLSbUYReWkMYzytCoIbuQRdhklMMHPdB2EQQ/aB4wxiOhfa1
AhENO7nQEJxe227gZX+7vQbHhzz1SO14BmbXmsp/D7jnMLonM7R67QgEZSEe2wnd
X916dvOdYyJkXxQ061i86O+VYzVDyLvxvImwB0T1GlUP1pKdI6RCUNLwsyUC6A56
0/jk9Rlg8J14wgZxY0fezOOG6bs+jkgu3a7wDgWHeC6SD+3LyVNo9tqpS4fHI/iE
8GHt/bwxNzTbBCsjYL/7yQcZddYjyUI3CD7neFeaujhSSEyAjPPxdLfm2JtC73kY
QVUKyAudKx60rocujvQbKcyP46ckoSKCtZwdZoMC0/EsBZUcqkzMpX4q6O2ewogV
lC8a0JuYuUUdiaISJ7rx36EyVfrsLsQvXvyn4C/EEtlMEUKnKo/w2Xx2N0am4Iv0
eYaR54KxnrZHPrr41+xsCubrSyvuEjNF/b8FW+AdfP+pqzI7Z/F/36f4LYC6bM+C
zFoRy3gzhQYVQ2Tb39dhZBLUZsNGgjiuI6q9DtNyr6aIvurKnxBiV4lSK/swVaxB
6PulLnYcnwH567At5TEoHJvv03AzFqgexmcTVY6qtmLP7g7mMYLYof5cxxg2YKHR
KBi2tGW0QYB0y6UXmJ0HrlH+GycRA3q7vd+2Fnq9QV0peZQAMSOh+o2GoZ9atTgZ
k7nn94vvwjBEF0CpCyQtaD9Hy20UyalGyMPK0zt3s9k2iaMo35mC45vqNe+lpA60
P3ei7mr4LJiQjkXKQzW3JTEsH/bWIgI4ExThIX40G3dTI5kR7oIB3uMZXgyQ8pYb
`protect END_PROTECTED
