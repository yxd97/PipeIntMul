`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JxhIfz5TUyYVyPvxMnQE7ElXq3yUD7c/s1BMIZyhTbS+/41OPnFTphobROhUICoM
P49CDohimWEvsEHcnys4UxstOysYM9O3hlke6gEVghu0fJjJjCUFOy+8/0tySK5O
algPdKyc3ZaJAwTyp42NIEVpg+Yf29pAoqWnntfeEUX3ggZYt0ROSlXoiJ8Ecn5M
7U9VPccnotj2sEauOxEliFoiR2znUppJEGA0m7bQN8luQDF7Al0OgzUkX1RJcCZa
PwbRUcDZFX8P4Y4weOdJLz5lT+qsqc4QFIqHdb8C1DjnsmaIAxDMYDkKFMUI+9VO
CrL8JoZF1gvKFQJ+2wDQy7kDeyiUvb3PLfR+iRCb8MMoj8lYIcN9Rsgc404dNgLq
cFF8ODKRfvX+3yiylmGx6Y/anpvjCUpWp2U8LY9o3Ep4eW39814qj1J4sYSt/WUT
Ka2E7qPLrlG2sdinYhzNr3BGpe0zyvB52fhg9JmAFqUNCojoSg4HOaJbhbYBgLtl
/vL9QpcfKablYQUNYqA+Jjb9vz+69ZmNBWNd1Wksw/uhE6m7U+v3sgQ8UNZFCPnf
sFiWclxUHX11YlOveLB7/24sKJ14QeOKeuMtaNSfHNCFFJdapBQtDF+jBLWTJPLf
9RElA3La9wDP0fjDonV0tqCfTnz2kcwKBv6/z+idE2fBQHwFEzIszVSxKIvHH0qG
ZWXEFRdNlOL/J1+QnA/Nq7FuR/4IxLDKCmypC8NW+rhfUejzwOooNPbI1QCGzpyx
3zgYOK/C7uNA7keBCdRJ+UDo3lrV/1TOkany671svrr4EESwm5ghCf6PyS5e32Tg
xDA2GPx7r0/dTrlxgJk0iiTJBpbnUag02fgg5GYhAu0ShmTrSn97Gmnz11pXjYN0
0Db/R64hXt8WVQ54Z7ilW6I/zxT6910gmmAUezv/j0EvHIpTDjP/i2mBUJ11LcZa
IFGQZz8Nzg1kakLS46wAhPW/Iv4o0bVJaI8RXF8BbT4OymxJzN4eTa6A0gUA+P5b
fdlYnADECZscErKP2mu/U3fuqm47cKY+vFsSMiTEGNDSaZuQKwHlV2uSMiHAx5s7
ixXuiwGYdDOCjefbd8ZAA9WAtxlbiHGvyCcG4MNgDC1Zjwt6q5aQAVyNR875i8KC
dnIjb3mDIdcwvn9S7KpMaSsY3VvS5BKxguLPesTi0G4jzIOhQkX+ViqD2GuYWjfC
ijwzsm7NYmRN4DkjT3YYYqkEm+2d2bCKZBpEiNuQ5zCrNYNk83rb921wvSgwDGkt
STrONBpdWszCFMxrPgir+k7TpWZmRWe4MUqpl0WAWrghoixeIA/683pTnWIhdqZh
4jEoHSFJHOIISDi7azL8colKMbEQS1yAZ+NRGA0nOAraS1xNog9nVeuTZI5dFB//
YUbUDf1jnBEua1xnmlLVYxygB1eoUbu6YP9Cl8uVUPWWfYwzxVVaiGnU+H3+t7PP
WB/zlrt9Y/03Hc4ScG2JWztkYGqW3HyevgtCd65zr8No4HPnvSPBegmvncRKpki/
Vk5vTLwsbk8lJojaEmahIx2UX3I130HAyn3APHfWi7T6v5v6a9cdpDHYDNBN+63G
GZcu6+JU9/+taEcxWwOkLuhLMTWt9s1Mf+o33SpXhyudEzDUKK6Y/dCmjWRc3wh6
+TtbtoQcMnBeYBw31mTN2zbtgJ3OKFZxNxCpMnh0H64IJYKmTAKksei2/+gHO3CM
QbGt4pLdfOzc7kWLb1NbkkU6cZVV9nffXeJqlA0Rx1SZ4OeiUkFtSWAaaiTR3Av7
A7NF/29hjt+em/zKun7lPjt80LY0qFLj1uXOUgwQsKDgywwshbiEsZFJfZUPOPri
WbZFwaSqfgcGBOnMG+5dsw9LXoQjJ1TfkuC/CHi6WnjBbfc/HujMuKEADvY/dF3q
3A3/Uqjy18QluEclQHEzcpejoXHz5y3rb0QRvVnoaz+PtvrPr848fJOCQEUz48v6
jzaga0jVgBLqVzAkE1EEKxLoKMvCXUZvkeLcPycSqiROAwi7O5RiK0CC0ZFAI7NV
PFvD9My183Q+GfIVOcsxGXn8K7dDK2F6NDyPnL/lFoOZgB1KjEbZOBiMYN6PDoC9
`protect END_PROTECTED
