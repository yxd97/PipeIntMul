`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LUDdOjy8nfOQPGQ0brXEZVfjppJAgmqnKQI2eQIgZC1CnujiPvjeVDRRBNLr6vG8
Xr7wZ2AENvB8sTNrIP6EPhsPBcvjp/p/ozViZfVjx+73oCwVn1mgObBaAwdV3K0M
OM3+qQk8OF8EON/0F+7iR/jr4dQmlorHsJ3t4fiCjCpIuOSoqFGhn8/OWq7WhihX
DjgZrxtvcsQ8nIHSI1nBrZVYF4VhaOj6zuD1wd+bduRARg9VeitHDE64Z5XBpzMV
JAXCK2l+ScDYyEsqX0pz1Gs4jZODxyjMZwvjlHOCSt597INAgn1aDy/gAcpVUoeO
eTAoSWqCzVXhrxQTuVw6JzMsfqaBLv9Mg3d0qqvyJ+8VPG6xYAcYFHKrvbn7V8My
mLAxrHGh3oV6ICdVnh/1mWjhlPV6v5vDJwvc6W6DlQT+LCRRAqkxqwYuCON3cVp6
Ob49vqe/BrALGYFLbCKKZJWLdEonyHUdy+2NS3N3gKef2iLBYFj2vDsnOntwK0v9
84E3/19lPXMamd8XBmcG2UMbdOux4CBQLXTY2x+2I5zjad5PAtcjf37yOpwOnHGa
67XXrywEDbNQdlVX2EKcNnKrRAP1FBVtRjlt9OxbPbwI6Znw0kmFDlbJVWwaK8Lq
Xe4pxfj6JX0odEvk/nHz4c0KujZGIJuCW2/4iuNI5vLxi7LZogt1w7hZ7B2+lLSa
gT5vbinuZeqMLtQl7PbhcZhlQH5vlVmcBq9+dez6yfps2msZrLo8qG6oYrkpSUTS
0d/Xo9Rcpg0tmfv7+3xAugdBwzhAemXgcD+Cvv33YNBMUHqEYN0CLgZyJgWka8mK
Kk/QuD0beuqT1957BMIJz2CaQdH6+tmqptQid5SEmhSq//QBZIvRDqCybt4t015E
RnW3tRqHxHw+X1c4uFh8WOUixE6pUFxmZsZJQffbVKmp9aOgziHIRw+/bTccjnjO
HARl1ilJecGAAgCJjVvC0xeZl2lNmjxqKVc3fzqpK0TS0uRAQDhBBXtFw4WBfx8I
xzbppHFkd9eyNbk/I3nLKOnFh9FL2bxog45ovskoBmfU0lqoAKdXZnTLoXnmRzfW
xk18JHwRfqcrQVEt6FYSqmubr67Ciw8FL4VqljkpaCHMPWHCqBzwf7o2HjvyAad5
ySRbCWIQbeXRDl2ncxwKC0RKO1MubrTfFfEjXK+usLaY6FUI+RgtFAdVojgk9jbT
wASC23TIVMsm9ayxAhV3MLno2M0sJDihDFhJr6pYit09d9UF5D0XNQvltBKsbRfc
ptxtl6qAhds30mUiVRlJOGyYGw597oWzG8aWefbcEhKXiRnQES8p5jJ/diXtt1kW
w8RC0/m471RzvKCrfSLYpCs9sJE9lngdz9p3hEis9pUMioItgFLum7/HFcook6n/
87iNYBU0osVsVhDR/4C+cvOtPULjfdo2st0xgz0ql0P545RMtsnTssDpJ4FS5LwZ
ytt//iN7jm6SaNLvw7WkXIGqpd0DTODPOUEfWElXjwLLg8Zi27DK90KpgbHrux7P
TU8ff3MUsaivHzba/DPBBKXFHlerLMalvAyDPrOewkSxkjdxcFqj7UCcTJjUG8iA
zKTEkqtmnZhr/G1lt+DKxsdEJkLbTQfH3COHQR3UQc8u9Ds4dVWFT8NZ3OkY8DfL
GWujmBGo9rH4s0+hMh+3NPTi4kw3GHGW8XnCHKQ+kG2xnnKLd2hUeCU24HlgKXVP
uMJo/oMsOAC+Sy32RHPF0TgD4pTAgTdQ1e5c5yuUd6h0mRE7vbRzbTKLgBVyAX/+
SMpy4zGRZiiQ9TVza0uAXeltnWsetyipluM3OXNDbbn5cTUF7bT1Z84GTXjhmUa0
UaXe2HfzlvsFDqP3N+98WxPOg1S7od2tOJSFXlI/jhrSXH/Scpql0neLUq3Vt1Nq
0KXMKF7FCp/mhe1lRtOJh9a8mkmZYzjU+oYNLNi/yKdlHd4wDC2cHUiNc7iKt5la
ZsmjUymOU2tkmbGdbS0s1tJBbnUh0TcCKyUIZvhQrXdlwxBeuHc/LamIoa0DQz4u
g9YtvoTc7k9NUeTpU1XIG3QA0XMVq3gW0eTVYLFZBqJQXviI8a6nxEdXmwhyrHt1
IJvCTq0rqu6Wntm0UPFb9UZGOqYl1QWB9SfNCSijF91e62xuXEQVJgyyR5watHXO
q28Vk9Vy+O7VmgSUxIiAbbxtKqhfrUfVrIojRKjTrSUKHTdVPOBqgHQ2MvGNcY5S
qWdkQxbgdZQ5U3pSFXCxUkJueh07nU+32dShVePEx2qjKLPhDQfIFkH4NO2xZ78l
5ns84FbpcdSbRBeDZY7bT9Hm8zBu1k+1w/eVsN24fnZo/ZsUbgCAhvzOGsQ7gRSE
dL1TO7h2elDFE/jl2IdKvOhDddTrf3qLFd8IFJKX3UkNi4NOUCkk2zDbCHHh9raV
5pHmM3wn1FOgld3R+3/wT3GRur/hgiSO6AtV6Ic/MIqIgdWsiiDAafCPLK/sXkUU
TInPQJ3vhaXJ9bAEnHgAzIiz1MaGB9O60btvM9var/UVVbGwxRP/OMusF2gKBRNB
FHu7jkOdBmNRO0M7wMNajp/dZEMZYp3/5wrkROCcSqC/nXGhSNr7Kg9eOCkICVMS
RowWBdzfJd6WCJ0GuEo4uMkwAV/oBFeKcjmYga/p+bESAm03RwGtH5ksN7YTTZLv
fS3/PRNhNH4/H0Tq5H0JZE1i9WU5KCTMotEDoA//r7h/FXtbDRAVDELU8vevppxY
4GHZ8NXmZt5T6xNVWboswqh0h+2yNRgHV7VrxbHL8MKpHdrZYbjyb81I/UtJ+8zj
3S1Ix2EQh3wtnLunn8VjiQnaxiCOdES2L5lfmQyqrAbAOVL4nCPeh0r565NCP9cl
vkObuoy38inH9OxKMJjhGw59uHxzOxG7trNbbpupkc16xE1v8khdXaIwepiSxFiC
Ym9aM2nY1+aXFuoXcbC5DA==
`protect END_PROTECTED
