`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
js4A62AJHoceUjwf2ia5ghlx4c50bQscFLAqcdwEVXhCV9EfmRN55L8c8BvJrwqV
CAhCT+Upz5qb+EKBJN44+KpSfLtrJxKTf7+66WjhfOP/KGgWdQKDPZ2g1dx/TcME
Z8IXK0Sz6SqrwkeevyxU9eXparR+2zut8+TXxFgWWZ928iM4S4CF8s9Hn7uDwbC4
ZA+g2SLdmD/mj36oWvQumlF2e5fes7CNiJXJBwzewHyKaofZSTZFWmJM0IfEL6tH
M9rqQK7ZCh2e72J8LzliQgbS9JaI3vcMwlOu7cByMrHFKC0gTTI6tekSPVqbrZlA
5J2z7wuMzsLTY8RDNdEJYcr83YfYstugAr1FkDnBNr5J/qtGCyg0/3tyzF3+Uwl0
1GL5vxU3CJ4VTq3elnl2zphl6NyZsMNzgoXOqa+A3Hk4wC8SyvyOTz/7USkKixyK
BELORcYjrdz5jxRUmtJDGYVHgk6yoxqSMs9ZwP+F3wBgj9W1grC05sLdZVR+ckIV
DCoolbjM+fxYjQOnLUFDBkMcXweQ06kdRry4iIv2j0LjphKy4hjjAu5fPbjh5WZG
oIJZQdDhAAr0VK48EpsQ1W5f4HKP3o33KuIins74L6UevyhQ1PJGT9NpReHcVh1z
EBLuAHKedhTQXf7pt7FnGU4JlcKd9lybWhuVFRSzSzwIYDQO9rduB+qYNjMhdIJm
9g6EaWgJYtYNLIbdZVM7t3rGlyirdatl/tS4RH0WCnksuOM2Nx9Mqnnsa/icjQ+2
UfRD67EvQgU4eqRQ/sq5ALfOYqqV3haOQz9fNU6fQUDqQrzEZf4Gd4rzZCAUaDfV
I3SGsmsvG6Eaz+h8N7pE2ZosLscYV8IvjfJTe2KWlblaPFJaYSn5sk5sck1oo2o2
OaWmqNR4qk1UbjoWFPXE4yBRsjQPl7pr/eJVSRxz1im0oyvNH72oQetdh6/HXOxA
Ju8QAsHgXGBevzeYenLU2FUHF0ipiAWHbzkNwoZGJ3rRPbzulPIwBOpkyJt30kfV
ViUTazfJ92z54oZ3Z2giPgoI25IUd1BNXFskQEj5Uth8xW8AB4253gb4/p8mfow8
J4mShZsKTQHfyQy161kxO/Zu0+DXU1gFbqPzFPIbzAxpuYK4E9pl73xVGYkYD7pe
4QCukysXyiMTJiAvBu8KgBGy0FkcKlbHZJ3sCUmsvLPlg75XsFqn18J+lirOyBAQ
UI80fHXsMNdUwckyX/YiiFo1A7RXRfhvvNoFEmK4mVBNeDnrG5Qlp9QB/C54ye3j
VGBZQCyitKFmOlZGiITJwYag2uHVKFkXr4zesQFvsLCPW3cRbJBfugIlxbkUA80S
/R2HXyLP5EiFT7Xoy1pLzR+XBB2O86E4ERneAWekp6rZbyaAAdnT/CigdJDw2xnP
7wKGMCL5fyop/mglCd8PasnpGAHyWbyahaUtqJcCdk8AdFZZsRNMKBB7p5G+hdje
OlNpKa2x8y4PddTNOD4rp07tlf8Q8WF0hVdz1xsaV0atLWUpN6+r0dWgLiYQW1hf
N7MaYdtx9Wps390qd/fmz4CpgNAra8H2pu6IXjUdtvuFOeUCghCq3AR5SWsmsQGl
y93T1tLlgOjS/mi5+5y5A35tbOURc9QKCZtQcTISDzhgyqp54T869aNq9u0cZAkV
qU2YWkT1By/eEe95Qz9yO592gp8z/TIw7YcMaJd0aqMC1r/vLsShPCZaIyxER/6y
m1SWZTe72sv/g15ucXdd1xP40ErwS0ne2YNQiclsM2OCUEblHh5+sXLv7O2kgWGW
jYTP3DD6FXe0HrBbs3wcuF04aVDIXOuWSnngsOvTd4BuNthqPAfj4EPYhMuK0wEj
LZV55gICvndd2ND3kr5HvQ7jOoTLT6EqisIlhHqArxS/W24s8lJCMGuDzwsKEG8T
cOpop1exOjMwTnSTkTs1nkDlt2nreccgO1Q8g2oTNgSio+RgG24qXgUGTiNg057a
bZP49Qc4zj+tTeiEipfXgKeWeXBZOcn2RF4SFSVQMqrAtXujPe3ea1H4t7VdYXcC
X5ddVfrfUlaVSp5lBfnIrsrtb3bRNaDgrtuVfY9ibgzYLBqyEcXSPJR6274L4U4v
7z6X77jcnwgpTG+loRng0NIaynV/P+BLrQ6a3T8bW9aZmhTIswu7ArRaHftMWxFH
iCKCM2JLc9KQ36iID7FHVQVUoNAsDFKf+P6MowblB2xmQQ4xB6Ia65maauuJiw/K
5tlmr05uDAqKAa3JT41VwsaiYtgBZ0hgdLfg4LOWDPu57TO3IhzGfMhVSzXYwVny
4b0uc56lb97jXr2AqtyDEPJLR8VMOiYTLD07FAL3WxclrICorVc5BRGoLIjhdy3U
SoYtOZGzOT09tUMQ3t6kDgozamHs//4ISLaWQYRhOvRmm5cK87Z4PcmgKXLZGFjg
kePospEGjh1DJ2KdKqUv3GN7BHhm6fg7np7Nw32CU/s+VjxwpPyHd07Au2TtMuIq
XTrcJYyyEyD9lcK8aR3MzomzMi3iMqbbP7RAZtx5SZ6rtYozV6a18hulYDiOinqU
n9sG92Yrxekh2+4o9Sry/7O2TX3h9ngITjoshqjv2yy277K8gYXldO0e4uqnoWJ6
LmnS0TvySAQE4RUMMtZ57jf0+JD7fOcmvFzeTmAPjyqhZYw9sqVrUT7j55PqwezE
xfuzIsjQRWN35LD0pfTTO7EtmQezTUFH2xVrpQnbCtGy1aS87fcUpK/kEPxP3evz
h2HED5ypmFUTHuOobtT8ivVqblgBnpRMNqMDGFC37YfFGMCstCHcojZsznFSxyAB
C8hhuGSaKYFe171e+AbbBjlYpzR69VQEXmPb8fvUfaU/neNDQ83ak5cjc/h5jqfL
TqP/baWXRxU4SiRDQLSwSaIgKvbLIrgjTPzBbu/cLfC5qqq8RqO+T+Q6kduTsZA5
o29ED7ns1n+/H/BzkFpvrcyHZAU1+Jntn57EIZgvfWeKqZycPdmLNGcXMaKy6j3X
nzCRUMU9+s4+eSjXGvrlOOUbB7mUM00t0oixRRpRvj4LWueZ2NPHU/m42iE5uyPQ
fz+bYmpUiSKaK+NgRvBmxBK5h+F3fBRbn/a6wnAAcmIAG0rIhuc9+EtQJcFa1Cq0
KxkaWBx7leQKSUMQK2PvTZ06ClHYjDOHwfilvA2F5vhPZB99RY4KjdkPD3qjY8E+
vjBJgRxzNLTd/lYuYtSwLhkN0T3gK9Qjl7ike18nItZncnRsdYeNVyxItAjcp6NJ
zQkoAO9NN8Jv1sG2rz5yAVdY2O8/DHKD0+LYQVsWtk1X5nilCljQXkRF5sRWOy2E
7V9wqByuEIx+9DFJQcByHkgMFIrUSFc0cOlhn+9ohrmn423ohvIX5VlbkitkacxT
+BzyBhERVSTKeN+Z9lnwhYDx4b8rl+Mh7qArqo3AeaGNgijPGawjiqaFWduxH7Oj
0Ge/DvX9zqNQ8OSQBXthW0yUnEA7YYzFKX2jTOoKBphA0EYcrB+GRbxXb5MPF1iD
NvvfYDSu+uSYtiKJSV2EptgWMV4M3FdVyhl3pFQczCgQOJbCq9xQs71+vKTiJSmr
Yt8fRLa5eHEfEKITDH1JgK8uHz1vJTYm4plboTsvqrP17auMVrR8oM2oQp98kYTq
4M+viLYFsK+JsQMxFZAMAPKVwjTaX2IGjpDof1n/irynJcUIaZFl76L9HJCvP40v
WP8ja2GB5K5OtsDTShJO59R4ia7Okm38XVgV47ieDd5h0gAwPCQ8EkGZvhGgR04R
AYaQE/UGC4YoPGFGqQDbUxo1UQoj7bfSlsXmfpU/fgedms7dyFpxna1+t8Ms4XpO
pk6Xi0WVcSE9GDLjKNgrZF//78bqz5Dq1UAjo9hnBjLMlxMpFsBBccHnIcymAi2j
wjrJ3mF7TDNxxj/vEawq/Jljn+VpVqcm24h/NcPRYy2sAfMm/4a6lh/BVoYKKDmN
ujBfARRx0h+mj+gwWEFIzIRCJpykeNfQhxwXdLB1ues03hyUcewwsDPKu9OL1oZC
`protect END_PROTECTED
