`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EucZYZoc/MwvmBffnR/JWFmYHG15CW8FA58BvDp/bb2Ub6JXNL8thrVG8ic9H9+o
D70xkOJbdbc7AtLYxYEGObSWfKwNkpcY2Ew9zlnIhtzwJHuq0ieAsB5CPJ9lX40c
IgyV1d6XikFL2nt8sARM95YeLVaUlA/9uAelxb+ekrhZ65lI8Y28nXPg0BQZ5HF1
fETgvJ4w8vWFznw+RTwTHsg8D4P2zFiW4Lry0ijANs3MTUJDuBp3khnq7kjW5Vrj
GTKpIMQbG0UfI3/foiINvA==
`protect END_PROTECTED
