`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tz7MxkCGIwYW5TuEpWfn38UvEK9n09tY4aQQXSyYYGuQUWwcSsSvA4pjBDvQZAm3
u6DUwd09Fa8Kq0hV5tjD1GxB7TNwktojY54Tw6LY+vmpH9sjHCMPEbQ1BMGz1fiy
Qxma5oh7+At51BtJ6Hy9j8OGEbPfAj8Hoc72WrU+F1ep1+iKIi0njVF6knMkhh75
A6f/C+EE9ZdijXfsy9aCnonvm7/c7WTYtKPewHZ/pPmy7tjPAOZlFmHxmzCUooT8
P1Z4jNuoS3Bm0gNcd4Ps4EXuZoMgoW/VYt9DT4v9+liTwCkQ7toQcvLJ4tKFVQGM
fRXDyObX49F/6kC/UFYuhwWF0y2+b2X3k25PHAYwYpJQ73iGxTvMe4Aeh1XFBCwV
n3xsjte7fwq031T9TxHnmP6517fhkNrwMv8IKrLHGTV1XMehh/eQaxSuwUEcXEw6
4f1VpOOwhV3UxEqaE1qXs4PzOhiBmvJKvFyxmhWMd0xUektPO2a9ZnVEaoA6uw6H
z38pCCePtXTbSMTdQCpjhGhqPF2vl21adbitRLU7O1gc+eanXqb/ZdW1dJbMQGm2
p6qj6nh+ouus4ovwQ4bY3Xlrb5Qs2TUdhgtOPiwlte4GWpjNvU86Nqgg+yaWXOXk
Ny/bN4ubn6jqRh3DDecK+AI7qXRGhJwkTP0l3xknvL2z5qYykIJ+r71NLnffO/DL
He6TSnct1dAoj4rXIwsjtoaC0kou9gy3p0XohLXSOyPoP5ZKrFUv+ZsXr2YDAZk4
6rG3XpfXW/2zb/vKwxde1tGm7e1eotVC4dyQnQT9IMWYxXYqRskqndawT2TJPboD
Tt+DGiyLT7VkWzSAUlOAvra8aXZlMCmDhdZjXXZxC/kHkukEcMzVSjIN6KbmpAl8
6NRI2Hmu2+fguoenNmd88Y+c8VUw6K+MGs2D5OIODElRM1nPjMbyhPW0T4olmzQF
nwofKbMfs+WCcXLFjCdmfkeV1YLTNrM2uBKPwqBwtoAe7mrGFF0cl652oWP/n28K
G7Glifq1mGKisyJsZ/G3Sb2T+zgsOQvMXwrDuzSkl24x/nrYe3UzM6zQadUxyza9
wEKhSr+XrgBcNjepgHf/jZrRzcVuGfGNxAoX5AiJqHyMX5P3G7/dCzR+tP8gXyoR
9bnwFe9fwAnrvP82/AXy6Jpq20Ze0aen/7p3aT9y+OsefGm9ubewcRRfwMr5HSDW
rnJMtH8k9/IHZmE5kbaQyBo9Fpu5u5mmfGnV1ELEjgFYbgSabnP/2NS9Zz/2kDjt
Yl8MWWo/Y+j3/uVYkqiI+Qo9ycUZaYzpBXQzw7oZ47ODlnQRaNyKzCQKPOTTS4F0
SnnIpDroTFhPGG7bvPT8lMl85Fp21J5VwAl4qPFyTzx9WPel9DiNXUl5wMerKTtr
Z0L78jA2TM9lOXBAlL4ejMgX7LNQVQWIoSj/JGQhb1h2ilD/xRZATDZKjeMhSGKH
7KA5DRlnrOGCH714J8FSu+NjYeEsiFO+ua7OdX/fLXLxfTu5J+sUUUFFzOMIB1wf
8FwGzp34CqlV+qJKNWMiSrBeb9C1v5vYc/hVlZCMBQ+jpNqjXGoYo61HQVOm+nXm
pa0aPYrZuCG0n5Kjpf66DgL4Mft82AvIw+PNItUTFXaHYjXPkX51qy4Dz76gIQm1
l0HXhnICK8jwgu2jX/YsIOkMKxGWgl1j0qyfXlRZFyBvXEIdU3FXo/b8lYEqa5nA
06obxrBXYP+ZuiAFHq0hWv+LEWmFduK7tTgWJUQa/edttZP+X2w3Ad6m072LPfkH
3aNffZznhS5t/ZyZctUZkA==
`protect END_PROTECTED
