`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+Rrn+cdXbJuAYKRGJo5h2eel0y4UWDc0vWV6eF7dCtSjx6i+/8eNfBsrqBaRe6Y
zGLDUlyGRj2EnAxzddSkZjVd1IBHNwXp7ALTLU+D1vrv0ifFOG+PI8xsDvAc/6bK
CakwiM0h141pFzunk38sft4ZPisAIse4KaP+cUe9pXnFRpq/OSqoEhDygvWybeyQ
SeEFFmL4V3TSr54zWSbdoculCC6Uld9owm1Qam58mFtMzXl1KFssIjGkGyv+Ou6F
Ne9+lwsOFM9qHUrmexZlL9lIrDoimJjiBSyeHwQ3PxLt99rvW1Tr8CLz2RYJqrdr
W+iepElfL+B3iAaCWO6fuGmlNvqd4nasEotkUOl6g3m2/b7H0k4n/F6Bst3dra89
fZSIVbeFiDOxw4hQSKghZOAol2T/q2tI36S84BJKqDmCmMWFnHdGb0qYaD6M1b/V
sMvu8DfkwRDpo3av/pUDHmrHgwcTeQxAoWOl2Zfu9sZuWEVUEOx4RVjQykGDhHDA
AiqeGsbZnDkt4DjqNMx8pFls3osBJXS7rzzI5u4iD9m6eEg9koiUQ2TOnEKZbhCM
56SCCPF+pkgwmNpjJfTd9gSJRqo+MFuVsOKPpEt5DG9hHgeJFuUnsDXwTNBTjG7e
OQordUfmfr4bSy+hY2A2emvoDu8j7pWZULA/SJ+buDYugSOdrSJPbUyG2/x6Unog
hQ8pua5CfgQuvwkSrGBNPOUM7e8cudg22RDchFvF46qmuDAzUZUQ4hSX9eCj4+JF
+hIH7RGyQrmJ/+LJTlBZB+pqJp1ccn9g6syMZJiCHMdoqBF7KTF6YhhN/RAntFFJ
mR/7KppS/t6ZfEPYy+OLEthMEbClSooeg5hNfll7JyNc6oavlCIqZR6YVteVXEZX
xKqhTtasX2egsV7YgZsK5PXyu7Y4GRrD5dJAMfIDer8=
`protect END_PROTECTED
