`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQNDrOou0dc52POCrLCQc/7jEF7O94KIGvNPjBUHcbJWWLTwsctS7GKkDXFmC1lB
plK7VH/fB9HuQwRZXf7yEshyumj862ALfk/bCI6Ns4//MMdOcRDQQd2zexuvR2hz
npvzc8wS5FAbtu9Y+U3+dOdERklSBWhshYmvpKb1gb8fe5OuY1QBPluiGFYNP2W8
qvjrC4NxVF4YwnFP6S3fEyarHSkiqrmQim7rmy4VNDwsK6TQ5FLw7KVNrWOxRwTC
NJvSYUI3A2CsmtyUAxoXuT7hoFHsPpLE+mlZ/fkBWNoAgTfHG+feRPnYXu9LDVYx
Q8xh7V6/7UDqbkmaxDOa/Q==
`protect END_PROTECTED
