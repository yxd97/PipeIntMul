`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2JOJXOX8ZTlc38WWhwtT30J2yrF7qsOGzeyqbKRpQC+2YWA0CtZkAWnJCz4XATcT
DYOC+awlcDJeHGk3ZQY/HcCPee+P9UB9LAaVDF4UfnhC6H3qM/0HelUwPPJw7od0
oxJ6l1weOQSkUXVYp5Z/5KiTxcJ4b2/btN0f+Z1j+MwPlCIphfYZ0p7ZPKi6dTVr
3sjmjWDU8lAGCylj5DOoPiOV44+h0jfVLgQqy4Yb5xnZQSc8NLyWRy7WNbLTZY0P
isFElo8tgwu+JRiSpV5Kl4YBGE6u5Ad3LTU6WTAnpdZu3G10YZASekM3ZKXY3E3b
mzyPa77b2pN6dfubKzaK2wI84tnpM1cD5VadEp7W3RT5GPf1RCenCxxUw3j60cTo
auXWheaeFjL8zOVDGc+3mHKPwIJst6z834vvZ8UH4+S+hXAosWNxwfa+ikLZZPQa
BXlJFevwj16TZ696vbmlemmXdH8+XWKePd2POTjibsdaBZz9I0tHJFE20wPy0+HW
UL9on5cD7g/mIxqiXTg2p6D8osm21yZ7vMomOYaa7lL5DJGuP9hb6Mkb2VBFXMe3
mAUomvQkSlbcR5DKYNNmfCy9Sa09MdFlYzsrynMQj0aXQzB7qfLJZcWSGCO70iwD
uN2JtM2fJQJlUMWHSRC31CkAAKjbj8qc9YEUV084hjH9T+GChKf+qiDoBn7IQWeC
NTd3odg8DOV2kmLhhqUhP0P6g1GRnsqnBtlnEpCyL8j1ilg5jgcyYOGGSBCBgwvB
hg7rIkKeZ6axI7R0+qp14NcXuWQ4k/y09Cem4fCc1EaI9Ea0TzsYkmFLhnTvCrRl
Zz7Z5paFEEeCKoCs00EzDzBwJ5lQqFCdZzwbxYL5UJDW0/YJ44kFtRkwh53HmkHy
eeuS1jN6DDQftbUdVakozxIXdpPvfIbr5c88z6QI7kJN9kLe7isp29Df4iKRTYa4
3WaSuStSAZfok9xyCWtyHOkwbjOLgnDmnSiUyDsZswvsLj1p5Eyd0QtrQk8/cRyZ
4QldDemX842VyfRoq1xNiWpl4iINOA9YW3vDQKhkoyS7ZCEsWwCw58+q/v4RuOVO
SvYlH8rAaS8pFOCTZQx9FUfRn9AwPejqqInxRweU+T8uZFyTuyMDrD28MlQA+5i/
qRhX7Jxw3wsQQb6I0V824BwsLt7x23bvO1NLv4QPRN2ulZFXfsORez+rArW8Ay8j
Uad/ZAByTd+4EEBj2wl+ZsuKxmyp5v230BYo/NLTgy459GArgKSrO37fdPYoGGdp
qokAChcEQ945PeG7GQR1i+ltP6zvPilyHrQQl4U6tB9Hpjk/ECth96XjWNNMbWSZ
zieRFYJ9ixo2k+aiqlqGg11by6M4GYP6SIcUZ3MD9Zzm7iecGK1TlSt8rdnqh7oS
ZxNd87+7E0ZK6J969VSWHxBRiAE+7d6xyRVAq/fjBGVSRw3BoDwSmPU8No2poXr/
XBkAJ7FFCYUcAjtd6P00nogSviZ0aynslzOpZpyEa8LtP2B0W5VSaDZq+hcq67VM
oq8RsIfsY+uNhcv+lcb31OdGSp6Xt9qhw22BsMyeBUf309M5cWmavUU/01yCsewo
ZP2yI00yWmIVu0D2My3jqA95Af5q2mEA0OTHyfjUhLWqTkkxbrb7a2O3wKL8mStB
lBgKeYccAZMf9kyc4fI8b3nzakkCfTvMvMexr/WEgwdljr6iUUWdJHL28hZ/yxYJ
kXHc/RCGBla8lgnSalglGnUd8JjBDH+39VsRpNYHN62+zhGLGxXSa2DUjWuPmeGW
ZneQtinrhwyP5DId3PaA5lnpor0hDwfilK+NndxwXnI0d8O7IZvPZTjHz147LCKL
5T11cufWDkmAWpIC+wb9ffkEtvICX8uUYRf/Ky28MfqXQ1ASBFjTOBw5D4Jb6ada
I2BOo7tx8KANrfeHCK5xKylFQhRKPOUqQGi7Ao1VFJObm672S55rOF+rMScAyq3t
yqpV+GMOvafDpTGNIotEbA==
`protect END_PROTECTED
