`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N2aQyCSq9tbGPagaO0L671fQNE0UW55jqMGTEgBleFWo3gB1zPzdqS5OrgvfX/Ts
f51QhB+hfdlsgsXebS97QHYQFYYaintU/sdkVb19TFwPmR4NuGT0CRLOiPtRW5r8
jAyd2Q5Z8pmOKURIsaCZtDVeFPHMo5Jy6ibAtYxwVxcisNnvYri0lcOmjZUGrzE2
NADBD6OyNarCie9zK9NAc1XqmEcXIfUO4/pqX34oIr8QdNYfzMpLZhNTI17KpXft
GqhX9SE5IBNoQZ2Z7E7Emz7ZfNWK9Fj0G+dbSdBJWnFCdoZS0EybH0zmbzfvxIsO
T99K2k6//OBZ4V+WHTQEoSn10CTatcwIdHn7e4xfjy8Rn1OOHr65bbN5mIou+QLx
7f6bHcm/CYjJF2sRhlYwRqPm9tA65B1I+SjSeM55O5k=
`protect END_PROTECTED
