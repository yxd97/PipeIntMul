`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XU5wK/3xF+WpOCWBdsHRf+nr1G3wH16ZYmbvbFezRDVreuaKhS1XCtU0KDML+zm
ooUppS43ejQGaqJ+nKkG5vrpng7QFlrbf+4ydNbKZFlThkApDy51sniLNBbgbmTO
2fsA+TxxTRqJQqaNaD+jtauMm12dvNpp2LFFfVP867WhMP0le198t2k+br/M4r97
V/ouu17euMla0wM89c5i+3m5aXoOoDs9zAjN/VhRH2BK/dsarE9Dpx/HayceRbpd
fwI1Roiz9wBNLRs4S8QeVlA+VBr8pvuReQZm8RRZk1kKQkJ8tfrjEQEZbJS4Ijbe
UmiWKey+n20W861MH5uBVW1XxnS9aqhGFSFZnYm4U/r0G80VfAFhNdjuHvATtDe4
gUUjiWN6iCss5Rc8MBnvcVvO3wxTKOD6V6XQVGGkczTbuIPUhi/1i3fgC8eMBpUg
Jx2qiTl1ygmjNxqakoCHb6WfayhJfTuz9Rt+o8K/IZ4HWe6VH4/n1LHHXi0y6RD0
PwzXAw4c7+XHsvzsounoibCGH17UXyPyXjKsUuA2agVwJl7X/BJH/TqJ94hg21id
/uyelcq9CtpSDLHj1nX6i0D1YTpsHfcsUtuYSYZTWVDemZk5jBxeEcW43fiMI59K
PZk2hVhDtRfb8pgbC+eEr0krJcj26tmBPUaTd+/K/cY+QLP4e0wyvH6COds76sff
lIioZeME/Nhkzpa42xujw4wDjnctuqWQOpDajenLBqKV9jMBMIUBSCN840/MCNK5
BMpp3QvdGtF7CzEUAFvjl3I+fuf075wFQmvbW8GE0Px4Vr/JkjryuTcO50p2ZE52
z+6WbfkrJgjmdzJRK2lFHQ==
`protect END_PROTECTED
