`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zeHVFezqVH+MViAMZPSn356v84sFkgUM+0KrJtPf+Rmd5ZAXz69hjlMjjYUExGz
3LoLL0f6DMERGqyDM4yG4GW79SIxqwf6jyTfyHa4jDhsJ5TipHnYEJg/KxnsVPFJ
OdfTDRIUgxl9UlAHv9hnIqJbkKel/pA4YpkzWb1+FIqQCAhs2y6YKC6aJ8HuPjXU
zwr/L2FncGUcluldGuXBUj3hkOIIDw3lWAaBVeWgKY3vPEriH/iFsxP0AJy87VY1
JoM1uCRJhjjOOpy9geU9fmJDLiuzAuLxcz6AZ7uvU76zNDpV4dw6bnpI3xFhLJut
r5itQAMFsQTlbZgw7a8ijdU+P4hiUMpITRLCxY84meyw66Wn6A2EOo5nSVhNiYtq
gB413pWyk0pOYYymwSIkr6IUH+uzd1Aqo9KDlfXXMj2HjRX8iDYMl/wONUWsNYtE
7BWbsHTyCIHfXl1+vdSng+YRWW7+xZivSe/z1OajOskdJwewl7tQUufS7SdpRk7J
Ir4qZtpanqx4kX0KQslizS76+Wnw2LJ7++kLThY5r/95Ak2R2zsZwVipQX/S6mtf
1Wyp2uDqFp0zqF3YceXTKj7B6sssBWC2/RaPFu7rgNfIdAD46C1uT8GoT2l8XlsG
1pEu4tIg2Mr+h82NJhLpxpcxlWRCVvv/eFNtQOzs6gZDanuj0cLTfRdcTmL7PQFo
LLmldDm0uWgGO7ddS3apcJtHoUBy+ZVfa1ZP2385GTzu1hWvaYWS2gyITqPAMf1h
Sm470j//CRv4kRbiCBMFwUSuAhXPpw77qUuxdxBgZaQiOdO06CLtLDO5PJ0jfYf8
LTteiN1yXKZWVfbByN45e5GUe4Zaixbm+BpVk8iPrIskOOci88kyUXNqASOUTG8p
/VCPO8DyTso5W+LFYI6kfAB0nGCWymROfztbakszC44boV5lFReJRRY4cf4mHytW
D9yNBHwtDHG7HSHZC4YyAGjx5PKbuplR/l+ZedoC+9Y5ivqpl2hB/JdJN82IBRFS
u+hIbMTS8CY7uurs4JDDjS5bOdutNy6reohIimAqHlylhTbRSZQdHxLUvfhEdYPM
WxX9XUVFSDcytU26nehlkVZIEwwa+DGU9jxkoPlYRtGAiAARB4Srdso8/FVryXxk
1VhLUuBUDa2LT3KLgYxTiDh0vm9GlnTwhG5oVVxWeBQqMpXpKrngXXEEL4ifwzeu
bofpHyCNG7X/041H6AOBpo6vWddGP1pnwx+jEAw/F5AS0J+TEwgJpXU+Jkb8pZeR
ElgcRYOj41qsf0s3roLLqCj5FJCmJjpMRGp/HMdx6fozGZztS67lAsbPBybPnUUT
Q+UIthTUOoNJiGBl1hSUzM6zNtOtL6HA1HjxQvtbx9E=
`protect END_PROTECTED
