`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BL43LLjiEsJVELp+WN4wSKUQ+eQsfh4DJlMmEBrgMl1fbqI8kXyNSU757Su/OI0K
t2rXgqzD+vHqFjQYvVm7cqfSCgUeVcnw+ZElxzzsgJRdW8obBSXmOChU9/sRhJNO
FSaXISoXoGWQBrnTwULhyJjRXk4z8nELnh3koeRByRqs0pR86MT3RccwQgpQpzoB
quW8p3rn+BniErlnuLUcWnA3VIvbCGqBolCU7ixX50TncbABqmMT0C5/oMmBCfNh
1dnz1fyMGvJDVG0STOk5+iR0F9dlQuyLy+YwuHuMZE4u+R8pyShepl1n3o8dZU/I
CDu9FJ+It6qyM9FZkQFaCoQqZeZtAXmRbIztItfi08GG00OnA71YHB9lb2y+Zvhj
`protect END_PROTECTED
