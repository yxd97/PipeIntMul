`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ktAK34+cvnb+KSTD7cxemBV2w3uO1bFunrHXLoykModvJQNndew98ct8zXagQVV5
BU68PNQO0V9+SebQqUbnLcjDoorAJUPT8OVyABGnifpIVxMn8V9ZzPy1FXpbPO3v
KCxV3uMjvnruYRGaV3wUiIkFv6de3z5bJ1LM5VV3gbtUIx9KmVkJy2Cj0zpZB1i8
415MO+/QjZUzs5cKtvBEwlZAuFpKL7rwnASsHqYXvQaal37PjIYD2naGX5PMM630
noB0hTs1naA7ywEh/qKhIBxC+0F8xxrF+3MJ+CBTvTO4HdbSXpEs2gJJFy4D45Q5
EPRjudGjmfaWZ/FWsLdMs9oxvqfBrhEPhrNYA8jQ8pXO9kU15GzBrkteXTOWRgVb
wq5frd6gP2azJcMv0IoYDifa1mzufOAosuAEezCrnPg=
`protect END_PROTECTED
