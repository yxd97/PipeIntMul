`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WE5IXYvqy10KA5v0zgT3SznuKXyeamftCUiY4yfri1INMqMBIwCfhkvIgvyFIeN4
dF6dxehUtxVDiyNazJhOJCZvQOz6SJbCf0Ueo+jO5XmsszyBOboVaHUV4DSiY7Ki
bNUliIST51cFz5FVAms5Ji83hxIg3tzzbn8kkJhGl45U7QSbbBBNx5StgeTbj4Wo
e+qo6S/84U2QsxcnOaLieQ==
`protect END_PROTECTED
