`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bnuSP7nwlVrl944wBlLhXzG9xEvS+Vl9RgdUbd1r+KYsyzWH+Po7owlEUkOlUDi
W+jfyC4H/zEWwlaHzG0x03yKKIFp4+uRGEVFxEFNsJvSrEBwd2DXa0osVp2Meb8p
yJxd10ycLYYG4wbdMq7qgLkw2RFPTAjlNPnlk+19FqEeR5nTBTq/Vm+n9KmzHaGD
CRJscXDfQiKKfKA/zynvpCqXcBwyWpQmoxdIk2v/PGJlUWkISOfHmjGKOJU8g6do
DF4pb4gs5EfPgBPgK04Ix8g50vq7T690VDy8ntxmVPJZ2FDMftXX3OHUhAbDNt3t
`protect END_PROTECTED
