`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WQmjtDPo8aBVLHcWidhETgENNRlpF8tHdAfahF7cjRaAv+iMywDve2phJVi111Vz
97u0nAFsoSjI9IH4Ys5bohtEqpaf91yD7Ad2cTSecsUkKhTvl+zn04vjIzBdah/v
2SoulruMQwp5rMGps78g8CLesqRuOTvr61fsff1r2Aal/q8ZSiEqHrpPe4AFe8lm
PMiFH8VVmtXXWQ71nr97SJLYWiuKX1eN92nz5VIc3xoZWt1t5oOCB/wMx/T0PX46
6KMW8IPHyPDx3t/0LYoN5+NQNJMuxeC5Q+0xYBcyQGvOYkUH+TRvFwJGfqRM9UKB
R2kI6ADOGL1Ykvdm+hS8ZO2yojIyQ6camywYX5THAJPsXPawjtf8KEkq6jVNpnJH
BrxwEqg8Quf0/vQUIJEiMQ==
`protect END_PROTECTED
