`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1AqS45CrmViNrerAX8JtqczuiKt+Kgwjl4yfZOBl/19bQle1SN2IT/9K1uiUSwZ
whxLQB9x5R98beGlK7VOeVYZBEYrudyCV3aioq4uOUPDTkt88vU8gPDgIDVEUUgQ
t1FkTKkHHfm9a4GgdWil7iUbWsAEM9qOCCsvHdfIHeMBxCYrTzEoR5x8S57SNtxb
4WfWMFLmlIqneYGUvidEdC/FN4AqaXaJqjHOzBhnH/oJrrJ2ZdlAPQO0Libr6TKJ
sMhbm4DfE47ZvX6PjOetC5QUP2wvekZseUZuyJJhkEir4Jj3vV4YWuE3qOP87VRX
CFWBqGv2rSPWLAIbTI+zcoe7i7mG89JGqwc0FXrKpqhbZAQXDKMFZMvj5cukiUYM
HFNyGyzK8TgTY5fhdnFcXw==
`protect END_PROTECTED
