`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KYzInPWeuPeO0xTYyMRlgsCIGG9gUeOWW8S3ylV5ISBHMQzh39VWxKjlJSOX+jaE
gjQqAh33cyYKl1qh8SN5FpKYGOOcynsrra1PQnDrYwSjGnDx4lxi5biZC1iilxFp
pbg/YffAIMl10bsPmOyq+OCwRvVt+87hh7Vhf2Hdpf5TiAZAOaVTCkQVIAKcECVX
QVqNTTIw3GKvgAAMST8GF9IFmvf65BnYDlpinjse7J4wAhJDh3jg6AzXQKo3barG
2nieUS+ZQTcAxC3c1owoHZ5tVpIIcK1jtxa1Kn/TUogeO4v8SdN5J0xQ/gwNsd1J
zzaiymKXzNA0TZkRZRz7nfkm4xGp8C764zHT1bFWsXUKk4pmHPi8JGZ0km89yzs5
lUA6+FmZtBy9Musz5GHBKlUHhKtoFKu1kK/lGeFbVqy31NOWJu94dkepX5iNDwrv
jNIzdLqtXrv3tKxcwvc4oWP6XFsShcJACG1Cqu5G4Y4hzxMwT49LJrqsgJvkD17b
NlxgwbbppDGdRA2faW+HkoZeJjHra3/N/dyRURRXWhd/Dge0rdhuLA3WpBgrc0BU
4o0vwVWsuOohBeGpibW53lsqzcUvyy+pA7gvbrMnm+qzdQ6TPq634zpfgiimGCNm
I5lGjRE0q3YGTFLRINane9J/37AoH1hAms6CV3ZZ+hlxIS76WzOA9Egh8MYZ2DXF
4J8DZaw6WcY08zK2eVXDHulF00IggWIfqNTkN4VN9SfKJ8qOJ3XPVsIkQ1K6hers
mNTMoZNwY2WEvpqjTuCxg4H/HJo4PmaJwAHnDi3rs0d/RD1oEpAzFXYKay3hVmio
LaUYP3GS6Ky/LzIHtLVnS9SfmvcgBBjnHbnqVe7faqb89CSyBn+p8e4abOJhnJKs
S59QGwcAX4VNmcraFDfjcw==
`protect END_PROTECTED
