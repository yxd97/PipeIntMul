`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h3p0MIKW/hnWieDwZVn27Uy/IgJTsmsl9UBzTv1FrJSnKQVCSkpw2oAUfkVxx4ub
H7mLTnamOge5/05wYeN1we97wQzyL5bF/hKOLKUC5ykpT7Ee3COhzKb1I3ywg2VW
BF2fhwVqsziyxaxDclqcuYpuuc+a6Quj4rTpJgZ8Nr5j2MGQzwCaRD43PRvn4rCy
G4l+Ok6if+3v5Kc+wKuJJpYGnh6+JKsCGV/Ao7eYdE7ayBAI6bGeHCeXMBZABvcA
8P9KMDFNMxQX2rBD4WMlcAWaJWFmNVw694dldwiGAtCe1eb3X45o9GPbXjXf7EcW
sSEZuxVVpfNVxoBXcEA/EGI8DZpGisXvqSe7CcR2Zn0/0/nVbehIN1Oc7N2gXpnB
aqSA56Fe3IPKhw40mPJn6kds993/vZVKmvFYU10vdQuKDFidfJ6PRkLN7Bi2WiPJ
8+VdtwqjGeQB2fT9oVHKZmAj1fcT9M3KNm9YQq/MZgg2MwBbDoUcnNR8PzkTz5Ei
XBYmCg7EkZQB9lgbQDE1Xu+0ZVrJLS8qJmvIZZLPwqhaUsrGh9w8yhAprGBUpJT7
Ku5uuiNQRiOPSbGwru2k1ndQSHfjsnH7npd1+pg+/iZ7Lqr7/RTywDMQ++Oityl5
/KXut4sqpbQYJ7B10oRemSQRXW0v8+L92JGEPFhv87PzWC+vIWLYpl/L5vEid3TX
9SSAXihlkfui99tvRz97vfQWerJr6G+QWHTxb/lt+zCIwn6QDfVLyroCprMuJsWr
kO0VX5uLT49Lz464y7UFtxJ8n/R2xKvCeaYA+eV2wrPw6WvX9IiiVNn5yR4XGeqi
xl799Hx2zVU+xRZ0n0lXkCGlKOUHYPzRnt5pP1AOCU8LePkN3OGToQ6VedtvnLee
QiEJke3GUzf7Lz9E45ts5KyxHsosahky9tvnsN1OHhn8VCWGngRDJkAK/Flg6Gr/
PqctwBf5YkDWiI/jgCLJpSPIia5TJ7ZSe/F+Z0dfBm2S07+zRwkGxmHRAftU6rPI
GlxgOUeQcjO6XB2Ue67dbCFKSuwdXTC2JORMmpXBphhsdyiGiZN9EnVTPQm2NSAk
OBbUxpXVdXOJGiwKvdag/PyjHgam4JUQ5uPZrnVyr+i26guvFbV3z1BbED000BTN
FBRG4j7gePNZpvXz0TAHunXgDaRmfaiC/IQ/fWGp1l3OTHb83NN67S7hFbxFMY7U
aUlRlyZp3X4N/PADpYjJ7hn9/xljERFuLu1fmSssGRffFZ65D6L42OBoPcsAt/SH
GE/8J4PgllraYyiQhPofZTHWoYlRh2vXm6Nu4vQ0JMg=
`protect END_PROTECTED
