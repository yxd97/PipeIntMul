`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r6vMfIr+2wAoSmbUTf/mZkqFbvXJHmLX6dWGEVSUD5mlhgzY0Fg7JswQ4EFnJEJQ
QKCJAwvKuCrCIY8TbfeHDDPAm2QVlbOwb3qaK9urnjP+q1caBCjIvoUSKCNHMyK5
ur12T8jmzN7mZ0arxvkUHAtviWzxNiF2h2sBoHCnmcCOy1e1GlJOgYyk9Nao4Yup
rO2/Z6zGnWELzmTcz1XB880KnSVP3Ib+TAZPCTzusbu4aO9dcKO7d2AghLmyu8d9
YcmNgjxpcz2brPXn2E5Szw==
`protect END_PROTECTED
