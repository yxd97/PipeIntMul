`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ul1UdGxoE1a/Vim+FxghLBzvr9SNHVPg+OsMlEEUV21uTp7vSCRsSLRWuWSlkbqE
Jb5CqYIkXvJxW2KP397slWFlQlP27G+2XsXLpSMQYYe8f3GIqpd9crthUFpbspj+
H3AxtnZpoeIU/5qccpMUSs0LsUqkeYg53GCdx621dT60/CIWjax619e8BCNFt/Dr
QipVlgZuqr3ZgakFpceLVZHslxjD05ASdXZ/wrKAyZ/8xUjitVoQ5m2NUUL+33Ml
`protect END_PROTECTED
