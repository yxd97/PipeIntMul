`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRGbA3gabln0tBAaufmkO2UvHmFj1GTR/oqCPPMpbqOOgW0Y8uLJI+dLDxJk/l3O
dEMT6V1XNgmO4RXVxAumblRVXX1SlyJu/p2VTvwwwj0wUCt0v1uzhjV6esez6Gg5
JSZasTk6QVe0xlOSZ+5oyUPhfpUoWmVoLrVg6lS3iOhr1GF4S3S+2aJfD7P+g/Gm
zTHMSiFKUfs/h4WS/4Ljjx0ELyMqXMN/sNTLevD3q0paZ19WTWvwospck5VrCUhV
fjtSZhvXpCvyFiFj6HhDLUmlG05EC7/g1IGpnSuqYD4lDDGXmDAreB+0pIitUExu
9oTY2IxV3YCwlK/XBmkzmw==
`protect END_PROTECTED
