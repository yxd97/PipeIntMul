`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tLOUukD5X9g5noaCQoVE6YhT2ENTXh+vybUT4UX+jvIJNgpfqtnLGSEnBt5EIvGg
Ie17lPU6RUePMUfvMgFPWgyoDdvJA1ovzHv0kepIgjoTU8PrcIRCuqS+tJuF+KjB
89Zv8Rkki00MQ4pBljAxdPj/GOICLbGAP2KD480ThCfWjKGtbEQEQYr5brMxUzws
Gd8hUQOVhbcBK/LeFw/KLQ/blLXyji6wsRQ9K5QAQiZvPV2BNVRDGXntsOG4ttB3
ZPHjYwD2ChplXGENXoP9d9aQF1diyVFtKayCcOmGBExW2gA7d6Y/jAbbMO/9DTw9
UqeBfHraBlkGzbcXLwz3/QlKBmg0K/Qx6oBPSylbF1dboIwmw9uwfbERt7gYrqWM
NBARrtcNc8lev/RnFfIJMPix5qHhi3kZSz8QOoH04ayMmsWdgM9BSNV+ZSMSZWRr
406y+7mOgZ/Ob7FKp/FzIJCtaGGTKxsWhweKB41vF+sI/JbFO2Gg3NMSBnr5S8cA
Ti/Q5RKhP4Rgq5KfygGCfxIu9yBczytaurUyGnoPUbpn67HWe2QjogeCbwV8Ve65
WvmirWPBqLjMsw+edc+9NyPXq51MeMXUgrpzf5tA6Xb8CoSiR0lj6N6/uWZRfN2i
mnI9niITQEsjFjmKbaehzTuOVpa4nwdyQZR4ISpKFsPLl6CenSz8HZJmUHl92Eti
eU2HW5rJrNV4T5q2hsX35nipjoxxzJhdiPaNzLmM7iWbBXWvFxkorY0C+k1wmiu6
QkhOVi9oxFsuElmRnKEU1dGC2N1A5W7ZJUyRtwRVfX+++amSlEGWTZHcFHJYqehq
lXJonXZTlSyMCa1t0jZISp7q1jyCik69kd4N/YIWC5KKKntGbhCEBSxe375NDfDF
QbkMYn9MDIZi/IUPqkFSL3j+mqXToTsplZhH1rUZL8phoapYzKuGuGRvy11Lugfo
6ZT2+ijvVzlFIo7mQCs8dUVBQ613uu0ZZc5OmcSPGT2WpjoUQ2IRaGFp1KsfUDYn
ni0rkRphBk6Em0BbYqrKGMe1Rc8SD+wmIRImlOPf53BUzkPTSaxbrj6f8dFzFlQU
F4/8u2pMWFYfsdSs70VGjXpgk/z//QpaC2proY+5E+mtoy/K9avro8GGpwOGfPyw
AfT1macEyHG3aZaESdQdBnUKHPTo7AUpEc5gCuTJhCshytWdIz16Uk7HWtmvlQuz
t5B1dJwqcBaYij9m3yCOTYVW5QSC4/3Ez0jmG+6nQydYXKPk9fs2ScOw0Omv2b1m
z8PoW7r5BdPte/Dxxn8/7Wcj5A3i6i3OImpGUF84o2yRMvUkDqbYpRONNIdKwlwb
/qjvNRiNRRDDN4x3jki+LadysgSBIdE5h1syrCCxlJzlzw6mj4cLVrf+5xtWPLe7
As+B4/2hDBgly16YoXDYRVGQ7wpPudbkEPiHVnxYKRyHBbDS8rbTE/Fw9k2Jy2KV
V7NAW4CbRJDn2eJIUiSXhX7+JKIh1cd/hsV/RCkCgnJt1TvDJJnsIrgdmCbstjvD
EeQdN7IKMxFTvzAzY1zNT9XeUej+O/icTTIid4mAxGQhd049FlpaPqsJkZe6F8Ci
CvzZ0LBOYxKYQBCmVna2CJsiD6bJS617go05TFSmD6FArWiLOGjdCUVnTT97U29i
qfapUwOSZd9Fm15h7XzxrltRz6WX4FFi5bBGk+xWMa9GYQ+1VTNgpuaSGrIUT4U/
fBmjpAckVteT3pkRXTXaQrJv3H/XkPF3pTG4sS142zabdh7vlLDUv9UKj/EmKBSO
+XiV2XhN/fEp2u4OSvdJFuhUWGOmuVjL8F01vTVG7U7y1O+LqPCj6B92y38op+kS
fUq6xkmKKeW4Q8xFaK3xrNp/ZrRvAxQgbSvSCWj3ANl3quVgbipTKW90ra0dSM31
zqaY8cg/pkJMg/W2dtoGVG43KXcik55dDfBZqKtilMvlim3BPSseOgkH32s/GStB
ZpGOTi4jPgMjj2UfuIW2UAeyxtqahKSMYjqtBtcUdSH7DUth/Qqw5P0MXQo3cjdS
eKgpRuVpd5zOB8YgEXEB3vinH7wI07Z+GyGB1oyWvkqGf+j8P7M7uQmu07OuEoR+
NCDQVMNis5vxRMj/1q2zkjIZK1Glm+Mgz2rFNAvknvCy2koCnqPyehZAgWak7GK1
sTD4hM61cGg8DzJ712tjrqcrHLVFokGZhvyJSLlJKu8CmBGYQOd6gjh/+jwEF3Lm
qB99tk7j+LuHVxQrI1VJviAVkN9jxpJQiI7u04pHSoU0QveQG+7yfssPjqZp66pP
E5tBdNYvNtWZlFT9FICCk860fDTN/3AbdmaVIddlXPViWqZaVQBYQW8nEl05vVeI
MGlONyxwAmQ0vY3sztkKxgTLIDAAiyu3h0e3ryfSLWJ6cocNRePfxqdBagz3tpir
9bGtyIhwoirgfq1NXbX/CDuDMNq0zvtX5aoQsh+oN7TrOiOq5Wf6dFPqwSCIxc22
pOJ2YwJppth5mW4dNrICjszbskYpBEwxS81jyil+ML+ncou14OdnvF4m9SKc3B5s
OaTAqzTOywra13OKNrUgqD2+9BFRR9glEBudQC+QzEQG3cGMxnwBytGXviJTjcAo
xqjWvCK+GGjsey7umKGNweG2G3JLzrfznaI7y26ISeSSwABttspi4QZwwGJjSXWp
I5pVcBe9DmSyQU53vjyk15aPX6o99Q+zmPwRdPE+bCaipW1iNVtlrqA30EZGUun8
OGq+HEaax9cvnAJ1+mvW0qOLkkRPkuEJO3YJq6RysT6ZFXJgx7uLhpjzzQXmLEpt
hroUF+mcd8HU3Cvem/JngszqKFnAm8oYpw7tTZkBb4zqszVU+kXzFeVMgaYPNpu3
06AJVWwWy4pO2LOmQpqFGJHqeiqU5uR10nhzL5TbPvIeK6MX8kT6Lg2x2dReo7at
rTNJLKJ5vlZS4BfEHgCTYA==
`protect END_PROTECTED
