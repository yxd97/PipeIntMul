`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6v4tOL1uoICcyZxqXefwCFUEmbMBWH5WvuCsR35PKhTJFOOTXuzYOgnS5mVkf3a9
r7vfNfyCdTTW9JInnsxEo8w2ustq9rqQjYSKjW5z3JmCO5bH8Clun2L4qGXEKUxv
37ykoLNoA89cFJ5WzNwJ3h4+a9/GT9go+AgPVtLKQpGRDWc6nGsoBhJm+olm2xvM
1n/d1JDIeJOMNRNL/chHrUbz5Hp29lgdAe6LxygPvxBwAB5TvIVnNiddBO27XUd5
4BLdDxYiPL+KHwFUq/HCB+jsl1QAXsPOdlvozGSig05xHDYV46mS8FPFg9YA/S2K
gapc3b9f0gi8r/ze+MB0yuA3KlYKsADaKEkSQqBwT/sQ4kYNXITE2HdKnOZA121c
S/ze9CgRI/i2rYenRScaxRqGMSSXgh6VXV+Ew2MmfTFUSYrz07nJwM+J2mCbobQf
kEWNy1d0jQpbMJ5tCxQ/eK8hvaNIYJsmPkjHkNzrBSoo+FuhqjjUhaegixh7hqbb
1aUlrf+ISEj5Xc6z9rn/jzbrnRT1cVnnaUGjJneqlBJuFIBlhnUwnN/ueuUdmUP9
kg8+T5SgzJeRAbNJlwBga5zYwgSos3Yr0LII/TygFa0kMyKGvcglLEwz4dcsAc2A
CtnlddCzCoa3p4uGkuzE094I5jGPYrkYfdoBzl1I2zlh+86/1Gnoqebu/ffVyuKD
8QtCBwd2pQJ3mwp2iOplmjoy1f2mmdr6wC/L5QrfwNeNtiMEaJ/17mf6cqYdORCJ
EQmjlTxPXUYnonZswiwwQWMHu2C1P7773UnQ+DF84zbFDsewwKmj7P2PlCH12ld9
BXTMf6v4SbQobkGsIMw7bTHhGfQ4Iasw0LnCPLZYbwk24gArxHnebECmudlrcqRP
NOJRr3Yt5HjWNqpJtOv4N0TxzNkUwUhVf9zm/9YymGZqoAykDR/8bZH7hfc+vTuR
qRlG62BCCcS/jSQcRkxR3O+aAOYDouKHZoLN60tEWYR+gJ8oVKCqoksOf6AA+8yr
enyHkjbtdQ+I7QOW7djEmPfoy+42VBp9ftLFzBXsy+adPfhaRTA/wdZ54Pttb7dr
GImArUqXjkY1zdsKNbx1iBN9QJ9vXHKMwTMs5hI0WMa1zFIasA006BPoaWeTN2eg
l7HGdP9Lb059ziPwbwMRHTS3OzLPzpfNtXtqXOo1tiXmYHLH/mTFJaumHucpTiFG
EYsAzdQC5qvNYO6RXD5cFt7BEfhkUZHHAqXOBGKHIOjlAOvbEtS124ad+m1tQIgz
dDuBr7OzeafKtGPMN3bYoLKkpXoLnOlmODT3W9/712rUXioTnsyVHKXlCg94eVH4
Eb3n+i2Ke7a3CkWKZ9O3OrZ/TLcEqTSzbqkvebyNEG84blPeGqj5b+MUU0FGszwc
Qvs6Mwo1idiKt4gp1XEpYveS++D78PKWj4Q6+2d++SkgAkOmDN/8NxsHjMf1pPjj
BZRTUFNyIupIp280tw3Rz4WhAjNUwzXKKUq72iWgRtDXYW2zrM9s5hd116tte4DF
auDkVPQcu2J+AvVc1l7lFXTwzMFUhHXxcvGFgmeXovjx7Slabt0YEPa4Bfy7gPe2
o51Sq00JykEbx6LHgkelvylkQWPAEs3SfSuuylfEuZJf3vJihH2hQFm6pTEgvqGt
Zynb6Q/jk1nChGzSjba4ai+M1P2mpt3itU2cADYybhXzWhWvfsyIFed3mvi4XfNS
VAriGbtTDS2zzDwtfD2UGvrGBIQEEhZqTIIkZ/WowvP386o+8aJbrRcFof6RcF8e
zuuAOZf7KzYTfIT5eMPqvXTPntyWt6WlK5+B/g1A0vqyJtIYg7Lfp5OmxzCPYEmu
wFsq7DNonQ521dmiFnZPOAsSQgIUZITtAYdz2ZLcjIqc1E/2O4n49UdspEgC/9lL
p2cOpDCRNnyxppL9n6x3SdwSMo3TSawtUgh4WE+Xjkn5oNokeVKL+wn8mYXF5d0z
WoyEz4/+59MVomEZsIOE2G/I8J8ECj+d6z3cPcnabNYVtVohgm0dYwtLIH0IR2D/
B6DDbzX5MtR2hT6lnDXCXYCsARj2TWwPCD+3pu8xhbr1p/vl47YMtRlP8jz+fztP
Ac4S2t+5TmVxXYyN0rFFowtvfYhQWtARqg702QNCUdSGdTqu8T0wMrlJ6DRO7Max
+INbzkRZPYviKhXVRB14rWuP/5kBdZgx9Otob1WrmGOjaoTKQqIgfbDBHemIWjLt
uDqpKrfJkxB+xbik+Su32JF74B3Es+X2LBS9NkbqI49/o48zSlx8TexTteqZrNMe
3z8+GEXB5iwY/1dQSaWyt8uSlzjr16QP1ayA9kOVFnZ5EYSrz2bQTS9p5eVn8NRf
mVPeIf/mf8VFbGVuHGC0Ws6gm3UlSFWXzXnYv4OZf8paM1/I0D80WqINROaMuN92
slBj8x96f5BcaXbKqq65YsN1K5UFr8ZVSnksxOgmQnvIJar7NuKKSHJ0P9Xb2TJe
5HA5P6d4bKvNxVcaywZ+l9ECbKI0iw3prrtYB/LvUtwvFt3yTY6dHUEKe8o6Neh5
or39yUCg24PUAeIwALs5WoDw/e/pkLgWudjhY+6PZfIiqcrHSc37GqX2V8/Z3+10
KYLlXa3eYCTfk3BGGzhJL6YdnsDkYl1mq84a79mXjrlCHHd6nHdiNd3ABD6SSLwV
Ll4duFbt6cFGvnKvnpAlPjrJD3sApctELmauNx92U4wuIjEqzCwqGXwOK8hkpmA3
VffVSPyWFkrWGmXFjuqwbQq8IepqbwMUuhVHwscpUlb5xUGTREFBzcnLwfiY5Bf7
fVtadH6sAgDio+1CeSLtUh7amXXPqPcjs4DwibYj4wJAUY6zt0dPbE/PPguQnCHs
BByCma6g5ZNDD8XZWRJT+d1A9nFu2WZiIMt6lWDaUSvJgZ8jcCMfWwhmroCB/rcv
d3V0GpRFAaM8yTS0MpN5J2XmhicCsInlkdjSZw72MbEMcIg4d+MGXMQV+PE2w3G4
G/Nad3U9q3aRiSUrAhPWl0x2/ahU35VxmiRok4GIJwINSb/+dOXeDHM0JMVBzjqu
k5yS9OYgfJO2K6jHjhbButsGhRWItbjHuXorh/gDNazKOastmIC6pUM3PUSr5p+a
wMNmOTPytscwdoob/x/SOyZ7d5F3X/SbuG4ckg2z42sYrBOUQ3nuQK33kpNiVTQQ
1v2l7GljXBnmkb/YPSJ/o1Bzsf21FXU3c8uv8tohA+/YTajBh3dqAU6f00hEeC0u
nSAVeEWIksjVF8pSMpBP6dfAs03n194IMPy8sd0D7b3O+6XrT4ggeF5F7GKJsNPi
Gc5QRXtTMnuhK8wSpA9NaEkpEapVSBPpPZe7rVNSCiawXrVW8Lb8/n3VNpwKmZDV
3pBVlTvb32sjf6PUIJ3looLuTJ1O+LF3Pjb9VA7Vfz/7S8maNQMawrPSaSU5P7sR
kFPv6BMv752hc7bwDIW4znBJxOddRdnONQ35bH3iYYCjrVk/KkAhYnJ75EvdeG1h
n/peg/bpsPtFbG8Q25lm8v38C1CajOXGuZZoQtInEK9Pb0tF6OjB1fehOWl1/Uky
Xwf8oUqJ00Y1kqEYAbcbGzoKzI7A1iL3OZ7/PBukmqTQ2ZAwu6S1oDbNeKpT+OlK
kdJYCsADJg9PN9SrbJdRV4NRpRz7kOqPyVp0arzG0LFfcfpvSro8Z+v3GxynzXAt
ctMM4oBB1kUmRu2m/czc3/TrEG2O2ODFfJPCp6ne6t9jzPB5RE4AYGcgdzm1yroL
+6UzpBVY33ZeUWHB7BdP44CvMGaT4kQ8n9TSdoIV6ak197swpmKWg0Pp16jHXWxn
UgAEDO9fT3JsJ1/9pAXRoqQV+T5OEpGf/PZQAPNsRQnCps6gVjRhNL2FKXsX+kZ8
aAVUyGyU5mbgYH+vdx3Iw+dmOaDn/zLwPXFfFsfUI9jSs2LVIkLGMDFup5fBaBOX
lfWdb0/jBcawkh6lXa+IDx3L1LWhXVnZCQnuzX3acXNlCAitPGokQVeEgFfixnIf
m9xA9fsFRj1eylfKPxvdLKUUvZa3EvtZ1yjqJAEbyx+r04isWZN2hJxHglGWOJdQ
ySkBUTuucYgZeRQ3C3qHBJaWWgjhgz5IzRUjoT/52uR8oZK+2yBpdvEH02YBlija
VCFnPA8MjyxXQVThGsn0eKIngYF4nyJWg5vGr1KNgn6iuS0hahQ6Sg2TTYPt26IE
KZomnxmcZKqo8Aj7zgKdgGzjC5A2iGMRJmwWCiIIpGsg9lz0jDwcNQNbcPF7QhJa
J2LPKrNhs7ngsyQNeMTVE2I6RIek1VNTfJsSBNPWg2JZfEXXDJxZLlaF7d4Rq/eo
jeMESp7TyCTs7mc0kJE6eNtKbRr5Fm2GBUEO2KPJ86s8E0e2Y7svKDvDNaZsBVlD
JRA7AcsRzj+L/qNgWyZ5Ovk/VKUyn70d2YUtYGzXjDZGMNtzU3w4169DLOBSM1eQ
1ajL3UWOzZ7Zuf849rEjcdPwebJF1AjYlai+6xn/as0DltsecgcMptoqHInuFurb
Lik26sndCyxx3KMOM88YdN135ZnvS0JR4wl50DswNW0nHq8Bkn9loag05aVkCP3G
oNUJcdiyIVqzJvns+fF25VjSVjjv/UMuDjPyzZNxE2fZhhUwAdtv9KK+3EcEQB2v
96f+zbAsIWjf/56Xuuio6VoORzHyasEViAbHiI1goQyqhIARn1MAwt+6ivYTqlrr
5jyofpJ12Le6GBNIdJ16cWfE5lwLo4F9mqtQaWckuMTQ9yKCrwh6v2g69cYFZCgP
Ge85Gxbcs8YQFb32co4znPEP6ahGQ1/CkQXztpbSw4P+3HiDSesa9C/mPOY8+io3
xkvQHJk88uxZ3oQoQ/B3XBFaUmYlvgD7o78uCqJJwZ6mIS7lHgua6bNMR8nM0+29
7q0OePd1IIqYzBdcnwmUiGzxryxc2aToK2CTm7GuYM8Us7EKCwqTOigSI1oXIqAd
drRa9hb9vPEEYp9rM2UFB9xR4PwQc64Y1VOxyJTYkvzapFAhJVPS/eR0NgNhXrfd
GO6mVlEiu61qg2qEwmsk2O5Rm5leePU9xFnxAbfGXhH77eOnRZGPAHmk4jUdC5lX
vEZTKqtsz4Et25x5MWeazPs3Cky0wlmk7D/dWt/3TD6ozbbbLc1AhofLR0G67vIU
cn9L8fFHnvjYNmIw+WPpwtZmetl7+tHkFtP244YQiIWObSrUJakCndsQRmgzzMUT
vjiQ4LTueSWEcXh5re1RRd/5c/F9WJPRe3YLnyj+Ph6fOYIHZX9a68q3CW1GnDED
OWAzP0OljCGLWZbJkmfqSk3zP9EXACydGIdAlvD0AB/SdtORkVESJvaLTbTXbVQd
/+QSuCERAYW3M+yIcZuSIYBzjblMxDL3RWTDUDd/ad24Pn996xDxIu1DJaJXdM4C
pxnke2XMYDZouemdiqSgz6f2gPrjoCD7hCqBgiitEil54IUuxU0ZhnTp1+x++88m
UfwZh1jRKhQD0n6xDHKg1mVzNGWnYM5GeQio8/xtY/QeIPh0SlNUni9bxuKAG3kq
ACp8tuoY1g5Ruq8lh5Qikp2qEeioRu20d6OOZe0K+oj5xyNXFkpP2c5CttFIHujk
BZGkYS6ufkpDI0Kq2CTu/jsw+NZyeSr/CXq2PXzAHSCMG7fWX2gvd84+BStx/7nn
`protect END_PROTECTED
