`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6OvFSZrve4opNI2ZudQ5/I2NUYYZqJxHhea4nsXnJUFjMLJTlUqstkhlfy9P+iC
2UzZ1Lpo9niu2sf+GLQP+yS1PyXhDsMIL9S6BnmHiuuBM6jziY3OTbsxruM2Wcs/
unOpITGXgsKuC0gdiOZcEJPkZsmEknFA+5hHolwIDhZCSGYngN1VWcYioqSJBUWj
tk5xoltTEPMF0yKOciW/Mt2y85tK6dtL+0tz+BITdxcKNLOepd4ngJICirTUFJfS
JNevX5sI/j/t0+Wrdvw9CiY49TBTEv17o0LL1d+SFxB08QBc5yxNfSr1iyntXTb6
x2oHHw0OF9AbQKhdifB7LICgvyA63aAWOcdg1fO7oKYOpS3pQzit0o+c2HH403CC
CvXp0KtW2ExBD6T3sBUmhrkvJplppUXaIrf0mHbLtin4HxG1rIDs04+ybk+AuDQ8
j2VXxqTQCr3cAXbUVk+cLbw3sYOV6Ia+EyxG/AWBnP/8uWyhNelEY7GANmlVH1OG
EKBC+RDnbZfrmdm49gJi/iQ64lHQTZS4t/yCRIi7pTuJsKquw3++Fbd1JHc16mGP
YPZ/G3qM5DXfely2NSWE3i3Xb33/ZBPqx/7iFV+nJp2RnaABceMau2+w8np+8irS
lqQ6IEEb2HlIkEZe786xLC8jLERMAzg0OIvyQn4tyId7mfyC2wnx5eDrwpXdAuet
wIp4YeOylHDapoG1lnCwoGNdoiya9BlVfH+RrEWsNEf+FZslM+O0Zi53lOxLClax
SoVpgbvQk8AA2dWM1kTaz6CM3Sg+5vNiXf//tRqAwlzJYZQyKXJ2A6AzGmzH8WLC
3+Ufre80H4UbKItrmlDqjqUjM0BK71owkL07q1f1w6ZIVCLlPAiibjEnmSmE7iF/
Ad7q5E9FsR02zkDqaDklQ+S7wttYuhzT33JzpBCW6z/gV5SW4I16tZmK1hPxrPMm
BX+rPZUzyNUMZzHFTNnZz20kOy2Oo5/Y4Qjqh2IKN8GXHSG4rovHeyirSHRAN6I7
5+QWvCOmKVPxkClQjPYoxHFTd1JRfiJj2DIzlkQ++8iLC6575EnF4bo7dkqrr9t/
vc/Q6cfZYo4a1U0AjpUk4Jqcz6g//YcpnflX6kDbmX3ekSdSecPeh4q2XXlUis7f
+masF3V0mqWrqRmh6Fj8VdAnxZeONl8fNR0VOW1YEng2OOGsldiPfWdFhJIlAaYX
GbtXscplyMqC/PfdssU/eUd+j3c6Tv18FwmWQnELxhiKE8XoaoGHik2z552RLo71
LSvoix8ugrw5FlRQNEKK2V8XG5JyxfxMOLhs/CrLFjROipoaF++lNQkEw+OoMJNS
QPU6ZTyquFqhFpxICG/YlQZ3uIIWqPxueblCqDoqHhV8Wj5XcDDrdqWLweb/olgl
V8aZF9zdvgtdnDnAZDpC2cFbD16lTZOmLUGR2LVfDk+TyYb5BLDTkoITepXKQxXt
5B1OVEx5RMT8ZePkF3d5DcUWfPmUXek7MQB8oudVuk9TXRymmN35sp9taJ1gjTkv
LsKlLXut+0f2eqEBHOS448bqNSmiwQRlZfFE0rt99p7CjXgiJuaIBN0UNtM81zyB
E25GIecBLjfm8j2UnxItlenRNWs6Fasev34cbno2nOlr6m0udCa7l+7H3f/a159O
QgVKGHpn8SLz7YHec6W7cT1gFVAYaEASD9W4cvvptSrUyoZ/huDYL10kcPrRzrCy
OEcHBuGRLnnxJw7SLX8c1PAO2/Ks8Ko+GlqriFQw+ty0D1vRIwNsH/MR3XWS88RZ
e06AYK+oy5jiBi6OC4bvjCg9jhb9ojn+uWPehY5BM1ibimP9YiUB4HsjoZuaJJwT
DVXAppAxkJFu1l5ry+FG8QyG+VrJGvUilBUqyoUJOnsvY1xfD4XA6bgI5pjv6T7K
1JuQ5nRPdbSV9/8w44bCDMbHQhngkw4vQVwAKFm/wUtsTYhDmVvYEoTMV8/3Ntgw
EXEDOfm1J1NgoNey7FUnNcfNaQx9P/s7CNLn3sgYQedDwasqj0exV/IcDI7kqp+C
B/WzgkvEqlkqzz29hu/O4nSm7Ws2XyZzYvo84QtBGVZYVva/Y5OKhAxHXqvJ/Q1T
f5x5SBTQM3GcH9Wt6wTFGA==
`protect END_PROTECTED
