`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkIj+oSdBzRSaoyPIjV9ZioktoXEWvQjt+hJ2Bfq6Q3Ryb5akD056/tPZ7BxKpw8
td9cGqvKUxWPt1HxswSXpzuDtagGfQTAEXVq6QOAOzLL5Mgv8b+q8ioa87t1aX6m
trEfk5+kiXEWWyywT2ZLYyT93CLIQ4O7i5/gEzL4k6nPrQPQY5DEWdZeM4B/51XQ
LBELZVFbbK+1ARt3VK9HcbgAVMsZ2pP9A0R5JOnhJIUjfikyCzZh7G/p3QbfcUjW
5sFK8fS/grG18ytR4LSr/azh80wLi6irw4h90rHPJsBwK0blwo7rsbRcppKOpG/U
JXPpeV1XiK7HmHOyFn7r/vdg4Nu2kPfAiRk8IKQBczAv9ImuQxo2GJG/UXXrQ465
DK+AlonHDkkOUtmCRAR+xsD2vKPIZOFiLVSEuDdIU9OnJG3UQv2m1NSrFE3TFvnu
90mGv+Vp4M09EvGU3AH8BkNET3D4rtxxNpZ3kKxo1BbDgQnwFQWA3W8jMgENT1J5
SCLD4IfCFam11cL7nQWEVW27LuOxdtUllPejBHehfp4=
`protect END_PROTECTED
