`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMJhmxh8gNWBeVAm+OamOX8BrR/gaKjQvBVCZtT3HthAAaQS4Y68dn3Knycqf6Yr
txdK+DYAl+n4FEN6jbAf125CecwaKFv7Z0FNb4ynqHYDV1NlkjvaNoV2g+pJcqRd
Td/l8hhDfFV7YdgIQnXDcJFpWc1AI+k3sHPhknBraeqiqQXcv/S+WmNyJi3QMKHG
lfrPZclKiL0sU0cUs4l9mHJD8GBm08+ZfSsH1FHvyLeykykgkeTk0xP2HSaJ7bwu
aj3JFtMHIfdJVLPu02Ej6SSdfmnImo2QOA9qO/1G9Me9YMNJdQlKFCpFnfQGG4n1
v63Kc9o0b49xA7gwLGxD4UjMkY1FlF5YMzM9ZesUv828gh1C9OnrUfTNnfpQn4Hl
k8RHGfVfOX2tZTGNoJxZJGpj1FHctP3uG3J8WaV6igBFcJZebWUZteASjdXFLDAw
M+FKKD3BqczEz5YZkfoacgKKvW7eL3fopH0jXtL83lkpEMz28bd6z/Y5McTUYycp
UeUXVgfvKGRow8+014Q3Q9wXtsiz4NhbKfDzGOEGuqTTrcFDMDFLDBh2m1rB7HJV
SNjyq4uqKqZwR+al3fGwoR25YUUwP7h8wTjk88Xxq9Q=
`protect END_PROTECTED
