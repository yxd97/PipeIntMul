`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24moi+yAW0ivzQEcfZK+JAwn1Pca6W9JLkXQ+zG6Zg/D4MK4+vcv7rUKJqK/nc4i
nsQIj2ijdnNTpDSCNMn7DOcX/bYyUXHxXyiF9CmD4+Dj9hGe5CEd+7p9OEMw27Xg
s2xcQPRC/0Czn1tXpPdw6mH73HqANAVmuibSyISLXMcQBWqm/GHSKc/3nmRm/zNe
qZ3U0LV8FdvAEqX3m/vGgYCQFbBzQJz/v34bkbJJwWWjYDyxrmr6/JRXCyGJ/qE8
0GkV14Ty1hUaJcydsfj7NC/Jcvj1MdoPvsO44/fmvcCl3R1wP+eIe1tp6UW9TO1j
zR67iLtgCxQ68ADxlbYPxR4Yrp/m/nHRyDVPTYkfqDkN/4mQYsLU0XR4C+AhXXmX
tJ4HGxyEnRQ/sZPMocUDD+UTjYdu3jpZs3kAM1Sj0KKQIXBQbzQK6RRpE5gTR/6z
7OGnnbYz8BcaLzNLUVPsgiqVo6IuoLHvrM0EAX25gij9v8KEp37qjxxF1kF+PQds
l5szDYEg16gGqBOfwAwpKkW1jeyJ4FSxPnb+3mlvDUbBUAfFXc5bHTh89g6rO3Or
iSN4xCZclCSI9roKB+3Nb5N51TrQz/wKF6a4MO7DeD0=
`protect END_PROTECTED
