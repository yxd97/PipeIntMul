`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqCl5UA5y2q/yMsOEVZAW/PId8dqQPMK08vsBC7w+c+3YtuAcoDXCDVhErbZuwJZ
wTRc6qTZlm0PTU2O49GSho52XZVPzC2L5jMGjeJRe9lxzDp+3ntpfaIKdRb4U7uh
HOkigQQLFrfnAfvJQ0i0WQCxWG13535zoYa3D5+uSOywlPiy4MJrntyGzhIAsJXX
63VlC2C8fjMWJJkRcs//g+FiRjeckOLX4Pe2vvqzu/UE6ub4sKhcbUhn1h3oJjrq
J2LoW9swttapuvnzjsynUa3BQMYyTkkMzTLmkQRwVIkVa4srxdDu5sUSgB6KfQIB
yZjDzkKBfjTRx/iiqjJ6WlgGxg4DkNCb13bBLz1C8ZMKOvHVxulHQN0GNnMEDmmg
NE2nYn/eROLSmlzAXU6NMgsAxH6PQ6b634RAaaWGaIjZaEbfthWhUfId3HYV5npZ
Hff4L4hJEEclqcFy7XvAVJC2wLSUWloX3QHjWXj9fdDwijxIeFM4WSQCArOZT/X4
dbXuIf8suq6HqrMTy9ipfgBz9oMyxyKA6xMsOhPsVeR1uaxyP+CIHrnj6BS92FhF
LMLDHmJZcYY8P+96prwFAg==
`protect END_PROTECTED
