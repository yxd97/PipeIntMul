`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKNuiXI/9zdWMaZ7XPAhrJd1CAC0K29v25jPzT5I8z21EVfDZxjICfEu2S07OIyl
UdFVliHJctaXT88wzh5wNdDAzPaVIUFEFJexy1S0avLkyL5zR/3Mojt14qri8sOn
gl++QBcIExqtZXWytx4vhqcXZmQx0d3OcKNBGPEyVfF6rVj2Ik7YU8+gIgz/6r49
SiEGKn7YiCu3a5BmBz7j+IrHAMApb0tJgSr1JkBVaMzFo/W+LtE55LLPYB3JhtjZ
WAiuSc3OgRnkirIj70XdssmW8M4IIUO5b2JUDfxz3jjWjrPJidbnSk4mJXfJqRef
32++DUht7hww2FrkC7Wl7EEc25SeAK+NDP3UdH+tPY7OQYtC7SN2D89jiJnjsUdj
b3hheio964qiI7hsEMNK9AEien1w/0ZVBUJ3fLtDMgKTjlzBHONaBcqsbxpI0H3N
M+GzI4JonVxjEyQUcuiDCEpO9ciLnQ+8bLk2onQPwX5Y2nk4axLTClpwZfWmilZt
ZI1HHfKfaaFvzt1r4wsW6w==
`protect END_PROTECTED
