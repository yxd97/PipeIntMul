`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMGr6+Q6R7/fCjxJzU5HWV+PRriWPgaCELG+N4eWmq4M3h1V8jVDL4yrl8SUnXwM
tgzdNMvSVXr3mXp4SX/qsyzBIXZgov/yfycLgZl300r8qSZn+qpyZ4VRIJcevbUC
zLvqIQsW4ai9gEjyrbzntiWhS8nHZDyGEVdpzywooep5Bmt38hlrDQU4FHdsZJ1h
9IiPTiuT6Ybh4/NcqsO7SwbLZh/KiiTU/q3P4eCRh70+h7WXuGBGspE9MSImhfJv
SEDzEZQnncNY0PEIqCrtrL8WSrW0WRSrexFVRCTbU5IP35xlgOMUIDyUUURwU53U
fzIMBvDUA6JW0YCFrsq352Bg8grPjPY2zHa/vjukt2awscHUTxuhcXlzyyyGEPgw
7N5A9pXOXDvJSxSmp8WhFwXxg2YMav90MefNEpbcbah4wlLJQ2gb4Bg2FnNFuCFu
nBV4oEbmRz5bovys7Y50ziG2wgfRB7SesUIflFPMxt37ec+AvBa4oiBTv+edHnnv
kZ4pZX6aJ9W9WfJPvVEF9QTpEPvvwYRPWzCRDuOOGRz8W+haTqoJpcifmtxde9Ed
BbL62vS5OQK6MJryX+2qUSbLiEVFP6JQ54JKD4uUw2ENCzzeXm73cEzjzyAfNd/u
s3ZSBkBd1zoKmi6BNmwj6ucqqT8RGZodTkrJvS/lKbWpdL5wB1l5ss6E9HqzDedk
lCzgQctq4Po6MRrpvLHVFn6Y7a43PfWPUJT+J200zlkW4ydrJJ7Ns8hs0XHAUmqg
bw1HnX1Qlu9JWNdXtJG39S7HbIad24Gguz1gm247NFG5xXsO0gEAUyNbp6RHhLTM
rPY2iU+ht+l7NzxrHEprzF028DgPuadO4MNhTtHPDwE+jL/GkExxZ9CcNqCaCRbF
uy4PiyF81pHfQk53bM/slEuuOT6tvRcfI2QQ3EQDRp56QntiFAAlilj1FGp/BHUs
7nHt/bCelu0BIVKrdoiV5zLhgT4iHsrtLDQkCvD/v0wz1nhoQT0A2VZO96YnuKgl
HW3vwBb9uU82v16Ftlzs5Sk0zxWs1TrlnGznvVjvqP0kY5uRpLpjeOs9ZPG8ArNg
/CUNRCAM/14YalB9P1lErdvbnpvl52kzAq+QyvfdO7hgDWI4LTXdkBvr8q6cUrOg
mPKImietAPq7hbs1c+Xlc/tRns2nViUiBNE1EL93Rsxf8XwwmsMk4TSzCGLDZgn2
eVKIpUBSikFi6ipLzhZRK7vikQMa6MXbsEJVOjPSlJ2nu7Kls7rUUtDatcbUc60d
eTy2gRv8i2rIjqics4Eztzjs6JJSnXuFkT6xNqLUGxYKmIuMpT+oEtxOpthOpxEc
3vd4TrXi3JuFkcZflKH3JdpVRvW5aclC0l3WPExdJyuF5FXiydk1E5iHoSzCC6hZ
ny+sDyvEQvCHf067LP7rNY9qhnGJJUfLFCz3KaS84hvP1wEuKCViin+aFAbfEgw2
3/N0hQWybOICee8edIvdVdPpCBkHG/lgAIDk4dK0mSMZaHLx16gi1fhJPxlFHxv+
0/xB6OBRKSrMGrvUpa7ZL3al7MtpqnTbQJH9UMjpVtJWeZoXIf/J/OMFJcTMyOLw
uWCjO/JUWJpjEmAM7VeA3IlUhNAZ90+W4vqxBX1rH14h/KtO/kUgMpGCJnmLlRpQ
mAqvDk1kGJw+TostHd8IDbA+OaDqL14ZPs171umf460k8mPTKfvgTnJkPYKsUXZi
y+7VMKDRv+mD6+ekwZu3Ag==
`protect END_PROTECTED
