`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1vxz3WTWIt3GE7/mlyevxfMtTjI0eVdw+ZQmktMsGUN5oRTYFOjZLi2YgipZfhw
OpJJY8m6QXGzTqqAHgTgZt7kmRlmydHNtf9f0rpf48NpE97ANCX9z51RMISVLIYo
vHwIvGyFA52yq/b1E9AVGXHsGv0rGs9ge9f6uAchjaW8qHek6wI+sbBGxqPM1MHM
VSXfpTA510BZfPXtu8Q8zhlhobZpvCF38UbBuGn5tNQHkXuIRuWeiZ4BUYOES+yM
ogClnRR38N4QCS57TkoVC18yOunLB6x/SFNxUyvBgAOaCaFyHHc1sggqAM6SokWK
M38vWlHjUwVmmk4FMB9CEXkqQrEGxnKk3oa+uu3Q7X3QuLA6dj+o8Suj/05NTB/Q
wJddoAfqgi4bfnN5GdaHKRDCx4AFHH39xPTJintF69Oq7snVZr5VAhTr32zRyx7N
Pret9FIMYgupDgpcstxHxGC5HcB16FHf9S/0601dZMOFv9fQw5FMLxZKeSTlBN2T
sNTCMl4MUwfn/1YPinvqjJYPhSYZFZ4BDLx7jHlrWMJVwKuQmFUGItesv4dTv9Ms
/1zy+E4l7euJPEEWO7Ru40a+50Z1vb1Ob055K+ABgBLK5XDxeymirhDBBiDTiHSe
kXt3pbPAmeG/qTSfPbN9PudEyvubBNDzdcxR/lcTs2ZHQ3ouh2DB/rAiDudbsNZS
JyhSPdbov4/H5s/+P8Jc2A4r60bQUdl0R3lEVkkAk3tB0DOP9xBSysWmqxog3b92
gdmy65UslaXpaIXN8yPjjOg4K5oLRb7eP18x1bi9G3Htaiw7ExZRoTr/IcgNWuOQ
YgyyEvydox0FjxKcSGI2cd45Ia3vq3RYLJ1fQ7FEwkj8f/TbHfAGmXlvjv5MJmBu
URgG1BkuZ6E+Qew0JFX0X5GUc63iq8Hw+tH9XbGrS2uIkMCDhebdD5e8aZuxh3/d
DrU1bHIaLSusr2eRpaUuDmsGj3T5rFpUWrlNmaTvv506AYXAZiPammhHjL1KqU0b
sihF0GgaowrL646OcBw7M/OWkDzhsiduxWfXwjZ4HiruQz5KxKMo9X9+z1QfOBMB
hW3/CpmMsgDJo6LvmkV6n38vZ4Tb+KhKbpHK1dpKM9lYqPmjyKAWHQVyHARvPoSQ
7sDIwCkIND7LwTqAN3B0w18Dr5fzS8TTkT5dWcq2oVWFi0NYe345kS6tW93YStR6
UcUCsGthks1ChywhE6E6LlPyw7iswCkKpHcJPTaWk9MeJ+Tgul0lP13NAZg9rtGa
l5BJC44kUsCH+dArEisy5IsKhxyQVzuZOo3KxLOvGcNxeV0tlBZUMLBQb4CHTkwh
L0cHesA4pss2fAJyVvlJ3Xr7avqZwdo0rIiCJSDA8m7hh5nlV964JbgP4HKiK5e2
BKywndrsGgJxk8XERmZpSKZMgN++lWMuOERLV3Uv5v1GvuamfnAzFFlsJCleVzN0
ASpVHVAad4LFUvNb8irxaTrpjQk3Ij8UKEw/3UJo/PFugC/n/eQ8SEoyN1e+jC21
IEi4CF5fYnIgoC/bW1nOOmrnioFqxhasDZ0U/kd63s9Jpvvvw149gqV7j1+auAfP
dca8Iqc+U2i2GFSr7hWHP6WznUEz8/OiOYsCZsUoYpn6TuVXdq/WvRbSJ5THpE+f
gCjBMMbZHlYdv/y0lhfknw4QfejUnaY2Y/r3XhWH1ai4HqgmznhlNoOYyB3YmH5+
5J3piNH0agVadpy0Ojgv+DBJXeA0g9AD7nKVYm5s54VNV9ghPQIMuwWgpQTD/7dJ
16O33cK6rntB3mf/X6MmsrO5oB/epS66mZkMgVE3btXL88qzqXZYXe11TvKT/xn7
mDkXIGqXPWOzAwl1hscqfbTcOQb1Y6vCPQRsY/j2gRpGSj9ycS5WD1jOWla1KqJM
Sjl7h6S5uBdsXxGUw0hqBpD0dmMxwvf7LzXfEXxOw+oZedq0XiLLkoUxxiur8Fuf
jmsyJVU5do6NBdNavKmCiiyOHHdX3y+xldQ5PS4Xkqrd2aaS2R3kI9xQDSfxFrPs
wYp5HGfuLuz/roYHj9FEOuV/3yDFTHVS+nlCKkOqizZfFuyDaxZodsG+8dGGo3O4
8/M4U5U86svtA35GrUYuFSfsYCkUhiHZ4n+A2AOdlT8FkfnpWZkjNDdtYxVjvjYR
XxSiLIgZA++xDyCsOQ6MZs/7Snezkn0S5CNFzKE3p+6n4awKIwt7SiLlmejYBP19
xuCrHh113H6eyRvEj/UivKA+r7EZHuSj/UganqyciSxdpcN2531hq1kAQUC5U7C9
Gs31XuPhAHuwjkq0uvBRoRFdbx1nPZG+50VYPi3z7ZADuI1x6QXNWpyje/LdiRx+
Jhe2up4n450S7RZlDGHYapgEKt7GRg8eIy7MvSB7nTTbimRpmRqcAPt73VMApDQH
hnxF6N9e/7tDpUwv1RCdvS9bt1PMUrNLWmFetPqcGE+Fb0zysJJDX0oGyZ3wAr3O
6pvlmNpbCKZWRz0t1cQRWcjJB+58toLJLeqv8z8uGmGd/gNGHgGTBdvrXkI+GGCx
z9ksgU1bpZhAbCtTJEyMV5SGn42nF320AC8VF+k5lol3ZSyK86aq51T2IqD3A+0B
8Wdz6uv16NqErW8ZJw2XL8LSnasmeASiYmSKSZy6KH0474SEQi0e3sfq38wz8mGf
N/DtOHU0zMZE4yc5pW7wo1erqFTExGjvLocxwi5nYRevLV4ukmfIOCibp8R24/IV
5RHF44TJJSZ/LxOcQBoUF4QQ9icN0WyXKfEcH4QTbDkDKV2Zha4UZXFfmTsw11n7
2eVWFjHX6uR+eZYs3aDWUh5wSz/xAxtnqPgjQW95MqhSqcDtw7acLo30LPh7Fiy7
3oF6JHoZTE0hDpdGe2wtYPaeFTDSIQK03ID52tH+EcqdjBu9ERyMDRO/P0P78NKk
e3YMmj512mxI+P/ZxsGDd5oRkFVOOgtJavPu+FOXC1+quM5XZkM0xGbA36vJFqTQ
OrPlp4dQjz7b19VXH7rTyY1u2MlIxiU6XjNwW3IZcYaHfDO2VC22lzTbaceqxRT1
46XmCAh2e2K9rSOOF+41RK27DxgWALEB1gwvsb378RT0KJ+Y/Nz+r/VwJ3gBQcnt
nreiRdIgsNK1OViBxrLRoZ5o1iIMQZuWY39g5N2NzZpCW8CujjYg/zXzJk/P3kHO
psmMRCVKd8WwOcf89jW3TU6H7gLUUKKzUKp5oML6sD/TESa3Rt9/VFE96w4jqO6a
uEqCvPZCiA4QQbjl6PPeijw85LdtRvIe4VdWJw29shOKhCVRmibe/UNvGLcDCNv5
NHh6bWJURaGr1/18GDRYBsGgeCI0MNMEvdjcZTsj5p9kb7a+FWCkBWqZllWMGavJ
D+gtM6DNvegjwkdJHTafo4KnCXVpR0X7c1M16irlsYU/a6ykgLUtSV97XpDNzodU
Os7uQ2vcz91hCkUaiPTRvHDSfvtJv4mXJkUjKx0+NRr+wC5o7OTS4ATP5h3sPXkE
xxjtyQkm74il9Dy0IrEFGtF7vEDY7v5FOjpghy+jtbZVyA+TB5pWKT/OcTworOWN
+yJa1jETmUN27x2hQNNBx8rvtGE6BY2DPzMYuiWiE7xUvpbiClsFx+BCVyasqOlW
r9ipSxQvLgwk+bZnc7l8Jh6MJTXEJcFPqKBYoBo60NveFkwndQZbZ3LCYNfvLnfN
PwjYURqsuH8nMiK692skkdpo3KDSa1PvHA0DAOP/fCRtplZOHrGECpS02dSnaqt0
rFADPFmbLP2CzCvbqyawDPJampQJpABES8luZ5DW9eyYmWFf9V8ok6YBOPT8MdU+
bEiGpTH0IO3jy22RKAIXjbl25ul5rhzgkEQvOPA/oVoP414zEWddXdAYTUTJj2HK
XSd4OcMZSJ5WsJkEkWwrrOOUMmXLj7ZBykDI7yYBi68hnqAwKht3DufcESP0itVw
XlB6+cEqXtBzEtVM7dljRXACDejPj1C/cvwXfEkW8oi9yM9Lt/gyUTqGGQP2+TDV
rT9jfjvFulO/E2Qac6oG60TWcmhu6pCLslMtWTTlMA1yqQXV/fgyeZo4YlceN7uq
E1WFNcoa0BzoSzX32sbVyrVnE4AR+4kGohESMasgSu0Uuffk2o/ZkrGxI56H7MjC
MzoQos/Brvoh8tZWqEpMd6EwtqkGhXndOz9XUeA5JtXs0F1tg4Pw1AQbRFVP2K//
001W6v3GXeaj1Bcc4e2RxA9IdGnx4ixVZZ/hJ9RzLB6coC9S9M+vb4Zqzw3fOX7e
2wEAthnBSgJ024/Hl8oO5nD+a6BkEiUVh6JbovKgpM3r6xudTVdBv/w2ERFl+Z+1
EzCxT/9o2l2/5r0DgOuOFlDcVmLQy/YOHY4fcuR2xiltdQVXHTWHe/G4yCwdL/b8
QnOUJK6T9R73OFva8PJM1APt6RzJy09CejZaz9RaaG1k6fcHPcbBdg0jGPSRBnBl
QdrQ6cxLxp7neaHguwyzu5QTiQN1JJh+8T5b83Z+dWMSzQoU3u3UxR4kfgqXe6HB
SaXSM1cdYBmW1q3+xx279UwNJTEvzSZwARRCT98Vn5EzC4uiM+0uacOIXiTeIjGT
b8iIIfV7ZPkre2UAtZw9SGK4IFO8yqV9y2g3Aw/0NVYuqEajA9kSvEPEZbTp0Os+
74CvAyd+bseUy6TZ9b2HmK9tK7bTw6IrfKFi+gY5SjzGDkoc3Ddypo8rx8OqnWue
Al7MUz0E0D44EDBYGp/dJeXX/ni0znjg/Y7AaOXBC+oaEnYiIRFUua1YArAq7kJn
u922Hp+9oUSgA4YPcHXTcF/IBA6i2SaqOXQcEFll6KD26v5TEa3ZjUk+s1fd0z6g
EHCuD51QJbVQWBWl8z+b+vliud4IjlaKlBz1vSLPTlnAHvJh0bYywBe4gKDZxTRA
j8AaQfb22k+rMjk2Vn8tdbqJAebhyP8idVNavovmKu+75R+NejpiZmsxyK+xtvtA
XMqi7KX+74PDGujy13ejmGvZyh3s8aKwk8uuf6+URLFVDYcq3QehxaBWLS64oZF7
RSSiyM40l2eRdhKoFUTKvU1M1y6ZX6wt/ayp0Ky1GMF+1OxMK7uEhmmkzCx6Qpfm
KIO4bNt+t10PlRPIq5/eIE2sYomyJsFdf/2imluscAWbYmVB2UnvA3suxSl1n35C
GiCYSgR7GhZzregBp0LEtzWcH0TIFSVEHWjXdWR2ZWvDASXnd1Xb1mOX0LtNCi+V
yIiFv0SD6PCfLVVxwxXry9qekpzop4syYOQBxy0Y+p0wvoZopME45vFTv3NT6uFJ
bt/ZyKEN62h33/WF+SewBGyLpVo5ra5QgG66RAU09nSxZNN8da1WDft7ieowfd8e
APuU77DiKtqHvQdz1kADa17qcAq+bK+lhEtfGDqEQbj1TBEZ0Qtlr+CRQH3PqP3M
uOP31uam6tb/26U0ptsaKnxeXghqMvRbig8w0sQZDvOsvIavt7uKoVl/4Ev7q8fh
y9E1flIMP1avfti+OkuetLETlwZwwKBoJl7NuBwbI2tmHn3QY4MsqddqfHUGyVaJ
kO/r/q1Z9dGLD0pFZJqDRpJFytsDa76ptGMup5ezYdZiwoVhejNyNyU5g5OGwndU
snnPmbTwrat2sbbSl1UCMW0hmPCpRjnlyj7HQM4RlDsgS+iaIqRI1qJIjYKpOxc0
auDsYSP3M0FmGu9axPs3W6LY4TjtBrPMNR5m8HHTQjrE0o0rzCh9a5lhDl9vh3E+
GlRQS+Gc7taBw2exzVuAM1q9BzVE5ILT7FTbJKk+yB3U59vuyudKWT2CJ9YODfsU
QZeYhW8TX8Nb/Wggt7q1kE7de/61dYvIuahXzDa57VM9wEGs24A/duqRyxtmB1Tu
O78CZnXrG4YxBj9H5x7MidoOTIa6zII1pZsCiiUZlPS4430iNikXCtvVX1FRYDdj
gy1XyQ0nDUXmggn0LxzmaRn+M1/elompY47PdRqmuuTU1WisTG7eI3dflUHBMWSk
NCDMCuYQFwTUnUqow91zVkvq/V5z8QQ//wPBAdpz75kkBtbboI8KvzYknVMgdx4b
Tpc2XRhx5kFG7gqOKr3GaZBxFdGV80v+wfq8dg9TEianaSu1C049qtiui2RwiRJn
JMzawDBZzhzau4pSkIy6kDMXPQnES5xzHkyUHrQ3ycEwgrwHIrS83EGvAldPgo0s
ijkjI+CRT59D3+pJeCh6m/W+RWhgNLLI5V15Y9IKwQ0noyRsNoV8rQhzc+ENBBK/
sUCoi5L9KjAeqKdak2nZJ8gj5av5qDshkJyrLeQQT2tP4clMBk+rM/itHJuwnqiB
fIauKPYYor1iSt+joeSh2Y8uRuFGRWwQAcxP0qN8xwrSqBws8BXXL/QIT4Q41sph
Ys4ABRncnUxAUQNxCSItcSXUi8i8DQ2iwTmPAJZJ7j6mYCVzl3CDNwCvTgFo+UxO
37uEzXohLUrnCa8njHvaviJvPsB3uiMRDq23Dv/0yG9jxXTqbBWcIInOWITUOckS
rK1MKCYLKVu6E/8K2wCk0H4tdv6OcF9K0eN3ralHjhGheQYBJvqRLtFz0QFH6GF3
zVK6P77vn2o4u4tpmWlNFa7qDDj82Kd1Y6p7r+34x3Hq7hFD4bIzKxmRILdj5/I9
k/x5jW2enrZFkl5J80wj22xVG2NO0ZvCjQavqm47aOsf6noSAVpR6X/beElN7BgF
FkXzx40Q9bDLllkZUiy0zdznjw55KFThu556BTDyMScxpMWQRAKccfyCjdXzdRg1
z21TTkJa8o9pa/d54/5ygIxcJowUU6QbTu5k3+A6HDuF+q+BoI8Io6/DhtxnaH4I
PNfQ8XwJR0omz4gZAefOsafmnk6gUqU91wkvbnkCou4yd1uTMJD4xzwprXJdaFH0
pTIeWK1yNblrGbLYFCEslNPRa2b0Nc9pZsK0DYXtNahRV41Z4lcfOV6tteiMamOm
vCG7OoWc6+SpugSvNBxEnAiWcwTkY+V9yXDSZBm1glbUYrZHOQKr5cNiWRTFQ38W
jf3ExYxDx+E42CPs2M7uEEdYm5+4zJ2m4nu9OqU6C1VEcN+le8JSOqXsbLxofjyE
cwwucQUhzyuZVr0msUEJYhv6+/QR0onCCB4s/YcNxFD8R1x2RMeiJdGGo/N41C4f
8J9WHugHzn3NMT41p4RAjHuX7ok07RCt9oTQFf6S12XQY6mE47LjzQas9qJTN2a2
Aupwm9NDl0ivHj8+9mHK3jhe3sHr8JH0ZGQQQZptXLRn43pjXE3+a9KwQFe4mmoY
ecQ6JiuZ5Te01bkI+8eB88WbltvUxXU4XQyAao+evv2/iAv7qjjcCXLBu67wGIRt
mMfrsNq5/HCItET9YtE7U0Jx5LSVYcogwLJP52eK9ZuFwxEU/LxOvt/CtNdZYKS9
i5X7uUu9cGI/F6fHRhiA8nx/zuKrJP2NmGc9KBPnuOevueJu9HdTnmf74lrzRkgD
z56b0jwPxqEG2Yge+PXeHmN58lSUXyE+KJIRv5eG6PyzCxIH8Ki81iY94EgMLdUT
3LCZvy0tbrB5O0ywEKP7iE1HMt+deQwuDsSfv/kpLAWr0078J+wZqaB3XxmQdm0r
6c5BQQC7jhPtNxoI6Smf5QoVdUBBfU2cVs45k+n1uYG7IPdHnuCB2oBjjFTo2JOZ
kneTwYw4PrcFE32P5qoD5SVdIYL58OgTtdD40gwjmRdTwMsWTa1YS9qYZF7er9YE
o4eAQT2Nz9BQBbI281iXGApbNsCZL8vWZ4vDuPBFB91dLVK0/Bp/T7uILr5n120/
YFiFq79xgOj62/JBQsm5ePdccLELanoEtw1i9jH31LBESXd6rXr+wGGJKeyYF9b8
CPlTn2+8iRLxc3gDkz+dKLTsYItibJFzHyal32pStvaM8asnHzyDJepo4oGK619K
f8teskxpD/n22Q/y8wdHw20tZm2y1Lo6sMO2L1yHkoAOOVOnyeB6ZeKsy/I9IuKU
Yvw4FIUzuv5qati/N8ql5t/nvnxUdcDirww8+ItgVk8mxakF+YZga/YFa51OKBSE
SkQMLxdgHmhM96QIuGgXjDYukpVfXrwHJhHmOvas0+fDADKogBEiKU7EpIt/yM8K
6P+Y93AAijXy2IZhsB9XJv+iZRKKO9wLymeLE2oWEH7LJ8YcQSFnqSLhDFwiDRdN
pQLUw9iIB21nqFqN4kXa7l5ZoU23laCsQh/GtECizxIQMKzvL25BdDRHSmq5Uuvt
IZZ4xd8BiWm6fi3ZgHxF6dvhznozadkXKJZWukwbN8GTKc0ZpZdrYQqwBG3MNWKe
gjgL8QxNiDPBe2s5MO+8FfQNN0WLJRYr47PJxVc2+E/H/FeAwTfKGoE1CJxXXqnx
ioDe2GXjheFUDGv4Zge+wVvQZE5Cq1lIEQYnWL9WZAx9VLNuf4jGX4UsjbGFNG2o
Xm0I8WD7FqGMDfqMsCqt+ttaPCRzCTonWg1bYRk7WwH+Etzwcvr7tSpmeckc6WPR
BbuJWbJpFuae7u4EXwlNjAPslwgLxAbKdesSz+zvJn+kKRkSOeEURcFGI/gI2SAS
ljoJ+KFRVTeBjTlKJICdbSGup3s/xXMJfaK44xT8N6WdUyqGUhygXI7aCgOFtLog
0HMPq/1R3rg0FNVZu2tAevJyynhiU653v7lwqpquGAyCiAIytEDZKcjffMDR3m2X
28iTY+Jk3zgX+yuipCRLgXI99xOGPGinHHfBPpCmX9XPzYoaJPnzFCKP3tCwsb0Q
UEHu1hXpSwrZ0Ux3GWT4Mcgx7GdzNGANAHTrJVyC+p+Hwczygww5cQhBpwtQoWq7
qGhe53HCjFk8Hw4/nnTJ/SzwwzJ0AGTeC+SeQ/X7Tf4kI97IKyiGQuzoI9kpese9
lXD5k/OkO+KIhw8syz/6EjgSoacyTgbsEjZwNo0kxWNxjJ8VTM9QR0Ll8Itp+nxY
7QbDI1zGzsbZDIgb3DrDAjhZJT6TufB7GfZw0fWG86QspcN0oSrJFFqx9Iu4Mstq
yEXzOKgC4tPY4G6j5l4KNHPt76kWaRxAkaMbaqqEQgusItYASip4a8tOD+mVbRV5
cmffUeHFwoFMKDXJAt/CeDFsDCFDVmsLk/2Rgt8zGauWP61t4YgVocCrlTCbdK+s
cyZUuh0AVXQ9pQuYsXlIiT95KgwHvRfW8mb33zUO57guuh+QRSePGmkgZ8fTMZF3
0SWKS5+42H2TlKWXofZyefRPTHlPZ6QjUpK+fPpQcVIjSUqCP9briEQTojJzm8IL
PiVP/Uo/vT9az08qM04cPdBZ8Y7LaQiskmklGUCQJ9J6BwFbU7fZIEL4eZahjxky
leEaA9o2wwOWwABbF7EMBLVbeHJXfPsiz2E6l9JHArWzyPAmsFs0HgoZNZS0+SVI
Vhp3PRtsmbPoZWGes7yzxoauOFpKhAUZjrqYY+4I7hCzGrpRdgdEke9uSKF8V2WR
7s6WLt/vz3LKDsYQPkSg3aGG9nrG3czzzA7/XHx1Rs+QXvSX/GYe1BTVJ5be+slG
kja7vgdwCLCKHSV1ddGUTs9oCq8eJ7E7VZE42tOdgLit/DXkz27YDh1rNByPtXWC
WC2Dk5vWioAwrZEmPQEjrth6X+SIpwK7WV6TaMRNzAerJDuRq9ge+ZUp23/ZMhjZ
++w0T2xfCkcwf7kEVIkwKG2CbB4PcH2s2XZw6+DTwJEGQzt23/DekofeZnfzKPje
nhg6OggamSCwCofiOMYaLEpsICeA+ADuZizdkhu/RulIJrz2usx4lAR4U5b+R4KV
vBF3/niWDe8ET3C/dc80fBxBokVKhrlM6f6z/C3cD5SC4bLkomYJ2A8+4dXA/K0v
yywGF7Z7ESw7leEcrgkAXUtTddI+LinSkOCtsqrWPZ6SpJRnq1Iz8yDYydYG276a
JBBVnDOTE3Pbcgm0n0DleFaPaT3iUwKXCE8pqSGFCBBxJWLmYNM4riTQiVxpSBTW
3sKf5SnHu1r0nCZ7WUoma0itC3bFLFZm3Aau8xkLT5GNkvMjfgMGybbnafbLjVLx
UHX7mSoXxOiWVG15uMxmqEvNLXJauTheclOacsOmSWypXoKNRa9xpYS0jNgTZFfi
8aeRBGTvbbfeDzfZQUYf6gvAHu6aqkCAdfjqw/hHSeC6F3pjGcte/LqhGqmtgsS8
lqNYaJt4JFcGl4hIERaszupqgXT580rw/UKi7N2mXN/5MFKITSrr3XlnXjyfxD5u
/61IRWCRrA9FXp6tqNmUvQVZT1lKJCJx6Ey3uLMyLsVgOu2Dc6h5kXfWQN9QRfTg
tGRPE9Qn3oMKjV3ls0kSUR9gHkKMfEoogn28IXEerL7FVStWy6mYGTQaa+HiUhiN
vbOSHUQqiLTxN/OWxynYKUl6e2rbiTJ0QRSl/s9ujHKL/+AiqNtgFe5Xk9yv/hLB
cCWWtBj2huBpYRCoPpfN8PdkK1gj+5Cbpx8VuHUd9DnzNF3ZXaVEN/0yOZ4jQEeD
5oJP01mt8FPWFA1M6go0LwOjaFclpwmha1bJSGi+XWps6BENwUae+fAutAMtOIi9
OS+jhyLHdCitgQqd0j0Y8x+jiG7F0A+B/9v7qK/H700o5pqTQUB49hiRls4DE0m0
tfihfq6rLyoYZacy0tkauJ2I/+0vt21H82cmP2HRHNJ0+5Mrfc0dxlxElHVD3Xgj
AUkDtjOANWxpMroD+J+tEFZEgv/vwx0nm78Lz5QMo8m6PKGoIGDMWMRoZksIYCdx
qiGx0NEztWjLfv2gRz8RzHvNv4AjvGpkaxpyX54ZLp6gJffMx+FVv5M+aGLmXdzZ
PQazaknPaz41Up7mcVTcUGbmvfVam2kwt7s4KRfHlxFr7U8cpRnOxKxQ1hJIkopb
7vzapcEIxEU0cmZKhhge4vQkRTx/QUo7aiZZVLGZXhFdo0NC3hMRPmP8LqU8nqNT
FAJH1I7l2nQCKHLxpyrpioxYwGCqQNRrw9k/PrHXGWYY+PMy2nd5zMrc9lFKbj4Q
BNSxzhLShPT/W47svuwziui8FxPse/XMjpVcO7//uVWeb3VOgWjx6G+sme2ylZON
RqhilhiNYnUwkdWmWkc7OzZufQwJVo4fusXdQOmmkxj9wsdmp/FLs3R0yBKx9BeL
T9x1id61oItL+gyIyHNR5IfkIJd7yNnzlOXaZZf3ui9kKQPEIokmtvlD+ReewCWD
7jKCUlbaMBZqyEsYvR22DDRfDW+0VHPaz8AI1UVouqNfL4tM7bh3qEUy5tLtD0zU
8ibkzfn8yPstVsH6fJ3aoVJdLHNHr9Ywt1wUB+HG5iasjcM/FohIJ3jEJ8E8XG9O
aRrHbYLfv42zXdOt46k0vbLCVUqsirLDAQESetLnefEaxYpYJ63btih8b8HODCXN
9dsKN8AwKXqBID8+xi8kwwR3I8zVDDWfBTMMccw6qjRULgYlEy2W5wQ0sQ/jSnuF
qFhQ1cuCkX8wnQ9o5HZYF0mVuhyfgc7XVlgvEUzfFVW47eCN6nXfXuKHeti98TGT
Fl3h2ftkW+dYF7ezCQFMdNacKxhYH1BDIOIUE+49fn0+rnCLcAKwCasIex2wF1WA
kDdj8LBPQQ+fgrlnCv1C/BDvDjxFkXRprFW3Fmm+h6GdHa6B2LevstdO3tyesDGN
sXsI32C9FPThgpR+BdjRuydV4+Z00LKX2DCeBr2D9hwb3m8Moot+B1QFlhavSzMT
/NBQntIExgyOz5UedgJiMPPDdyBeRCYdYsdvyo5FgRR7ridCF//q7CPQoE8sQZO1
J5DImbYAYaeQmx3mkZd7gu3f+PjpajGi7rkFp2KxujXH3W/MClJxPC8ulKOF+i2x
48zDOUIIgTBkxH9bqRQeKu9i0PFUeNhJ8oEAHx3d8EIvd0iQOBSc3oG0Rk28M5Ro
1kD7DaLeU779tlRxm7UiZpFoEilnfgkYVLqJxz1TS9czgpajLrNawDlGJu6gcC2N
hU5tTmgyZewhXlZpUDrrJsqzPoYZAoY4i5sjB+PTzEOE7QPPz7FgCnZRjqRoH96M
m+hakRGs/u73MqKEX69tzERKDsjEEiZCxNSo7cSNajKvbdRHkTtgWtgP6oSDBPi8
puebNa/guVXrH9K1QAO6Ugs4YrrKRvBJwV3qyqeX9fjCOKURoqXG5QX+IpYK/v6+
E8b/yJCcuHbhRRPMuuX1vlC78+AlIvq0g1H8lxA3cMiyMiNMvIJIBjXEUUIGmAI9
GZ19VbqPKMgYMklIcKskprFMQPqa9nyfZpcGEGPpufmw6U+22UidVp5WG2SEkPMx
z+LJmn34eccd87VOIeKm4thhMfZjsEQNmIbrkCgAsUyz0bF5l/U9j1NYaoYzKcoq
Ls7c0ZeYO7goYZiwMB4hZdnvtUMNTJCBHst09PqhUDIC3BPX8ssc53MW7UQEZtW+
5gNPYIn0Lay7ErKfHFTKM2JJRhVP47/kgDjmGpIvslvgj/cZ5DCFuPaHEqyExmwQ
7fRE0RlK09aj6eTQWKJxPe08pyPx/IAP9UeV7PHxV4n9p0+JWfuu7/p/wgPHyb2s
KBWHr4dq5YjadCfd2nm6nUgRcr8vX3oO2OTFGWMTD9KbTiNkUFPX3XLcwcX3eUzu
I91ryJUWQYANJX9/m87dS7fzzql1kqpIOfYpT69FlQjZ0gZKKNR3y2F2aw8b3501
n43HDkPlKRlvmETdlfkfh5NBQf88nk2BPVRR7xEFz9X/xN68cEFr3Rghp4zRd23E
Km4Ul2IGvtnK+oSEtY4bRsw73y0sTKBxDkoNDR1ua2w7Zyjow4YO8vY9amWsVGNw
jhtIDjnFzjDytGbspYGklPEGYcgWVvgAcN9JscuyfsM27/f2lah9MS1IGIXPK9ld
MPmYDTK1Y576k9X7uOkuyBOqBdlCyRVeZV8Q0jw9CH4QBpE3K6FeECa4bgbPrhBo
J/g+JY2d+VRIswRo+b/HyGLr1pNSgiSDs//+YN5J2y/Vl1reeGP6+h4QDk5fb8Rm
cYMITeo+Tps2PajtMoM7d6VLKOJil1Vjgvwzw6MZF2LthlJjgdLyaeovXSyD0m0f
r2QMIXnKMKclf/7px4MJrV0zm3ZMH7F+wgkWyZ8QAYrqEYpoGq+DEMO0Ebi1YfWV
P2AdOFz7Xzj96PbwxuCSLjJtGLr0fFsqU4uXma+fATYkdUvGGC5q8MBLmq9tdrTg
3PdRYbBBz93zzbhjDnq1Yh750isSDL8M046uW1f2Kdhj7iYN9nIbEBYt2pPTfRMJ
VHGQp3YINCGwem8AW03WWW6441z684nDji3MQfwWMJA4oYTISvy4/1mzZlsTQPJ+
tbSCeF6fHlPP2g5SmmQrwZMUSIRNh9DbGQnpskwoxHJb5MDQbBymJgOOdaPeca59
tqs71ODmDZy1WUA5zouWIUy7aXUMpCjoZNyaeh2T2kM45jp+Ab+IDIqXfY8HfvW1
P8BepIEH+TWdLDIdA5e/ljqQr/b9j5hKMeL+lpla1Ouz3n6iTpU+Z3fS0Rn/upyu
7CIkbC9vOyHXEfgHs9F/rLD3+aqXepHQEzBvE78kynqrdAA0zUi441lW5Jc8skhl
Ys40f2wJjfCyNdetDuQHDftYhvYhdVFgVbXtEBUoc59zXEz1xQQeEH4oX1gTlzfi
+BJhekOT3jTFndjLuzapZ5y+tKSfi14MqAUAGcnrNINrCOXs9d5Ez4ucVrrshJQY
GNRKUl9iQmZrAs8L5ESdhrubPXZlwI8Zzjn5nJr9B20UrwE5c4wt3L7jNq7Gxlfu
XcHlUeTHuNOAL4Ehbl4l/oaF1B4M6HofOFG7NueNJAqKcLvoc9YFuLxjQYFdJhnE
fFmESnHOwK+OPszWwg2b7Cy8Z8GiKf08L3cLnd3bxU7HMgANXwLkfB9zfNAb+xAI
NexOnoWnU/cKlZlzHfrLCiYcScngdNAwbRE2ZSZq8m3LvQ+yMwLm6Ee3g3txWhba
3ONgl0p8uy/PtI1k4w3oMckwEkrj5TBnR0JahIbgWHQWvndL3oc6MlKeIs3oT/5T
X92xdZB9IejtnVffdAt7e6O4abVwJNo5U+UR2QgPFK89OOGFAROy30Ghfn1IPhKK
feZ2yQew65HnfxcO8/POIL6GlnMpXeZ3UXSI6XNh7hmr8msCT4OlP1bOpCJrMydY
nYDiQ7GXx3Ck37zuTYQk6ffvz+y+3kUsXKk7+9xPpGwSLdLYkgF44cgiEHIAP3uC
fCCr4yQCch54bSiwv53EvuujZgiCcFSvMSHxEtR/MxDKf3DZdDvQRqSDEZiuWo1i
anZO20e5g5mKUAxGU1+m8Yu/g6XJS+vUy/LLJpgo9AUhpAK0LrtHI67/qaY/STRj
ameddhdSN+QEdz7DaUjnEk16WrZjzfS1Fd1/acPjoyQUJdFnllaDjAUA6nmHmgpt
ptJ1nnw6sCcyCvXxHiSkCzg9kvdQMjJB66biLEh8wdYA1KNkLBBhiuB9E5ZpRqWG
PgivR2l3+4tNDP56K7GovGnQsx9Y5RXnOVUdYVohxjuNZqKLVeZax/XJIzrqNY6G
EPjZ0xUdjaJKGxe4OuuTXnwa1jvFYz7gBOYQ6XmXhuFwqyiSYe6OOb9NLgkq3+SS
6wZEJm62c8WhZSpnYMj5hb4h+nobzp5lM9BRKSywyvpJX5z3SXEuH87EF9t9QPAG
sM9CZCDjzXhZAm+3q7HkyrDV6pXAlJ9GsDI36eydKRgfb4eXZU+b4J0I3g5Nk4is
9i4fgqN93/x6cepbAbxFmUnFch/M8PHWh4z3eQu60RezuleOm9Y/E/jHtElAqQ/E
YDXF5KS0WZLonU9t29ez5Tse+rRmfqGx9K8CAaz7m/QJBQSucgFCtAHTS3QSByhp
hjRxdwcikFor4zEWH0ao7WNScaJnekwCK6TGIHmDRh+uWAyAT9/mH6eF/63Qn5um
gSgUR9O1UMJr4ehftFFMIrDQ6rf5XTjIVEAxX7zgtcP+JEaM626w1P/pmTR/M41e
2SfE13g/7jCzgg2mF4pSUPWxxe8vGudfJDbBb/84dzY0+9F7VWwilcKIDN49VpBx
gbhKXs4pcwKUPy+83OgVB1/dT2hP8eOnVLdNVtVbfDSvqL7dzYJovswqRND2dDXF
NENb7sEM4vt1KFZP9LgdmlD1wRBmqkir0CAyQMURV3ZJLVOv6ULsRmvKWjUnwuXB
fAYHskJ55n6lsHBmEwY/EvSECZEyFs86DHYZqksdQrHXCxgGrEytFyOFtxpQMg5D
883ftCR2UMHl4kcXkdIAVLTBQtiUC+6ZEn/GS1CxH+Nv0NXzcmitH7S8mSAmxZ2p
KPCNgtXjqUwx0XK4YHlKvdlo7Q9OM94diP2q6certXKTPCJTG7HpDRVFU+mMD8Gj
WldFZIV2QNIQliGrjw2B2pkdW9r593Ip0UxWAUS1r33VrsXXQIxVsJMfY+pHMTAV
AGP/7mgoHVJ/dfoOE3jVQUrIus+gLRFSRqDuJ3GQNgqZTVkl2GupdD2gEQWsEMue
ZR1buALyq1f1M2W3jOtyBAdQmvsIlWPOopOZZ7KUP7OoXnwCJY9z0y9ZEfffTEE3
fs6iK+UH/M2hTPOKcWcM3qVdZyB+Ue/M6oHMP3/XDdSOeJQkeATzxZ9FCWE1B5WX
BstUfChTNj+4FqRVo3s7FT3REaNc2DTdLufb4NM7QJ9a4VQ8GuMtWLbIG67zoqth
pUos6Yka4ezQOaQZAxJHMWaq9O1QPlKNr8ZknJAt5uiyMQCDjhr791wsjLmngGe7
fThoDcz8/NllNFAaZ49w+6zs12JO+407VHRs/r0sbYgAXpVXteMp4agCOJlZl+tC
3v9MojXd9Y6jQyCsT5BQQ8UeW5FIrlMfnYkjAAvMJrLJiouW4PcGlhKYU9RdF2Yk
Ms6xPpsyWQGhpJ5wp5jG2TYozAvVxbbhsuF14hiScRWJikRyZAhKijBH+VYsX+Th
1fndIr5D/wfRp39tIw4Xva3P6lDR4kbjoO6z7RMEQU+snkIJJaq4GD2U0d58XZSe
stbnxsXr4mmLHxW/mzTOleDp6rNEm2XkSJS7Osih4YJQxuNv4skPG9YFWKEBYwxo
9IykICcNTYVPjUL3TmMOzefSyfSvn7BqWntWP3q2C88Lh+GxPhIYE7LbUVISvCs/
Bc79DNJPrFts+sG3JYfYBLMY7T8fpnRthjxErinPaX100aKmaPc60+nFSw0GxKWl
BuvLLGQaFVNU5alXqQm3Gq6YFUjJSisb7yTgpu2nOJIYRfQBI1wwoRqfsexQ+Ubw
8nFUoUro+EO+HyOK5I8Bkb+RImmaR3bsd3uiUrCsSc0C2bW0rmLW8lOpQdiI5kJX
wLUXCqxzlLaw/MuTYP31x6L1kw0FtpCOSOs2xK+vOhdW0pB26ovGqvltRDrakfyW
CL2c0tLpNaoPqqZwedTANiYROkAGbneqRuFRfZBpvC7NGPv3anC5UkOwYz2gxQ4K
uoRbOXl5PJ4zz5r7hCjMacskMc1XrTqy6zHVGmo6GZbQ7HzLHFeD/IhfZxzIUqDv
+wi6aNDJ1wFkQZrFyOEP9edrBZ/AL40AxVjLkjg1nU7Puat84Ukt1uHmOkfvUQfw
Em/oCHYVCmGNLC2toe1BRMg6hxWEaQoTLN9ru1cOPT9AfaqKE43O7a1RVybqe8qV
9oq3F1VJauY0bU/l24zgEbPsHQ/xIr8GsBRYA2GkNWcRe1OsDewhWtSQ/chcew56
oMYjpzlFx3U1mqVCj6tCCuCudhy+/8lVbeiQFTTtQK6q749wmnXiGe37NnqrgF53
E0iiptn4GOgExyC+xf/Vl1jOwvG+qYxeoXM+cHSHpTCLHJFpjzjvZG8LnuThl03M
rr3HeL6jPFUG69lk5rMf2ZEpDvQuG6lilJASfpMQb/Y6tAIvpe1sIZWYXcIn8QWL
ytq5KhKvdI7Xf2Vmzgn3dxI5mIQtmt8gou6lj4ykusnMhqIEU2VAxSnUrWHi23Z4
weNTydmQt8yRLocyxuB/HThk6c6JCWnBucemZFF5we6OKea15E/5tsQzHINQzRS+
buloi1zoZtb3IMeOzR31IjEPaXWVSWQZbx2p3zevqie78nGvLTD/nX0okz/seraT
O7wXtBXawJ2wH6NZi8oeGTWtiJHh05Mweof65WyIauTU7PdsFfafj8074+BrcwYn
zfHGYADyqY3bqtNwd/e2Wi0AdimS3CQkMLnyrZ97RvapPIrbGg4+miuebBq558Wd
U4yn+DXgcLyfsGp/Z34sDb8uaz1bCl5z149lrbihJ71lOeLz8Rbj/a6LPVIE/3RF
y57m1svETPVibc76b0MVa2UVSOoyUfe6W9mQfgw5Gej8LWF7no6fEx6f/GKSVyfH
B4IOjF6n/jyilHTwktueVsiDJQQyr2dxigDlSa+Y84BagNuNAnE6SDsnt5G6Huab
f0nROe8HPJQBJt9OA5SdUb1TmShl52ExW+iWxNqN+hDK9J2/DS1/sOXTETSlnZfw
r6fvFl6k9u80ueuccipBBDYq9xFYD7aJ5YKC+zl84ckwnjXwGY/UiYSvIE2rN88f
kqmyWVEA+KoyKb4KJi3V14cPWwDKKyDrob54SQzxBRUAjEMsfSlK4NzNsV3MBLbX
vKuoqJv6x0VarR5kHZFxWQ+0kU+p2eXv6C2yHY1HMOTUsWl3di0/VH9PRGKFJlVK
7KKS90P0stKGIhmOH+I2ZnOxIB5j5hgOHJjPOsYgvjo7uQLYo9WyrvsLOsJvECSQ
vFVdqLxrm0XhAH9cFZZYOF6naNihYNo0W//cs6rk0+NBuDBRD7Xm8s8XqNJK4+9l
I/JW6C59sXggoPy/cfp4ap/glJGVxXqwWtgnIt+znXTiT1KdYVkpmGvqKFCIVGWM
ScU+i3PhuV6QECstcf2RlI1faLMG9/8aRLmLPeIjyS+aAaOOZf++igfiTsqw/pUf
76DOLsenusHlAjWVgaihDIskUTtjad6iVRUHVZPk8MGXxNd8taR0Er52zmjMQuGw
QOyrmx2onxtCT2i0ZPnWNlGrB83DcsglPr80UJG7bvJVROksgkSXN0Vtx2Woy2BU
U29ZysazzDTbmBfWFEqvxJ6ML8zmqh8KKwm1WC2Ps2OKdRxOfMt2+5gLP/4zX+xr
xl5GPcOIE95AZCmu+cVsm7RnWM6JOZ9steq5Dgm4Wn4ytXnF9O2jFri6zsBclmqg
3qYEzOu8L1G/amYCBz9pfPa6LjYSSgaKqEhL3dPJX5s0GLOObMg48AwRZEeahPnf
QRDDzuXFhbDUARztvQxOQvJTFEzorxoIzjOhuJV/Gf2VnxqfAQThOhFsI6iK2HWh
bjJGxLdqAKAjq9aqEWkOZhv8krh6y0vNEUqE1E2Y6pFKUr9K4pvnu+TOi3nFrl9r
PgTfcL/UiLpTmlIMwbvAcTcpf0i3jboMc4v5tozjmAtR9OymFNt9DUhybXuxHyeL
rgl2GWrEIgRDQiWzQVutub5sKpzJGjp7AIRilhJP1haxtT2wXE6tBhF5184+95yd
Tvc+++y5uvM2CvrMXu10o82loeMvwjUIcrV4s7gVmWwxd9P6teRgW05ExSiRoKqg
ot5doethSn5ScwFuPFObm588L3SjZwwuxKvdPqmMlcTsgLtfjAlvmp53VnnqlreQ
prv7GhuZZC/c5YnG2Zd+NmhP/9AaSAW+tcKj/LobekAXS0OwKCOh+PCNa6ziD0i+
wAgBlVW+yIj/vtrUL5+9KaDZJKop2c6yC1AMmTSdP6aTn+t1zN5elDubsIgHeM1e
qMa3oGlx20DDIsojpjjKKdZ73ciEbmSglG/nKcscIjxiD1bcvidr+RhURdZdT93O
k+Z+2n8oszHhlxG+yiOZlORD2xKAYUMjBvDtt8KnXq8cxdGttxPwGqv3xc5H4gwu
OzZ73s1RBY5M9nHUaRVITNbhrmFZoS4AWFV/W1/pm+lzeS32Rr5ofIWQLVy+63Pv
jfq5n++p3UWw8Fbt9RXXPT3rw1nttCYWdgtwdk4uTh8o1aCInRtqmYjUID5O7EAf
tgLzgD63FszUEc7dZxMMSnzcjifvRdWZoBUIpY7VOWVdDIzA6mBuDMHYzE68+Bo+
qCIeG95sphKwbU4psBEetIsjL/nP+xgM5EsCfSus+eltD5ioxP/6u8UCV6/qxTEA
0IXj2MRRuDFPJlURG1ZB+b8A312cqMHlxTCmBUeKE/M8BRmCNOsHgCaP8Rz6bam/
qQ25lOZ6u3JPprg+0JuKHBJl1cD3CdOVjDOsFLOGtNI9byshl5wAst4p5zYF0XfX
E5aAfMYwVX+r06hyNAN/402tP2FxsaxTtDvlKPMdHsQHtmqTtHgcuVPEIFAhsi2x
aXCHrpx9hCmWYwViNX3x6GFCLDMKnITnSa5PHI7BBkaOhYTK82EOfyo/HjJPAguQ
4Y4fDunJgLt5oYhGuJyshkLsYw3BMcCyPn14vykXUcH18/bqUQyVsdoftmIXISyf
iLQqQAQ0A86MoMZMkElKzTn5RVfoeXga+Gu5bMqypT2Qfkph9TCHS6+Qx1mYglth
yXF5uPqccsqhYMSmiL8pjPms4KvfQDQ3h664zVhgIHgCig3J5zSsDmb58ITHe9HC
+A7igtjBDMje31XEvBTD9BaydvpOOdil60vod0jKRMQOhSAUUn7zck0/4chzFNJz
sF6Wo2Ms7YKk8hKgSkQ2YQ==
`protect END_PROTECTED
