`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVaIZ6Vtmu62fL0IUKiG/73ioTOKw2bn7xbTQ0yVWAHX0glMJ635M5MPFHlEn4Zy
ET9szbMbWPCt2uiIfFFvcFr+pC6km+uNtoaCYpmuKYE5jBXiXrvDMAmO4ToSyaX9
szx7ZZN3Hv5lzi6JGZnpaqZN8kzNMIZTGPu3llEhQykxt4dF6Tm2vdJe6N7SyKWG
fsAVjJA7FkTbOFsvh2HtG9G/RpjSgV2/27K7ZMY7CDA9YrXOQtn5RAV4FUs3Emxq
8JwtVESdGaDPN8T+edERcDRd32WL4Cvorc4hpD+mOijo4I+wkS0VdjtEFTmxn79F
DsswxZ6S7wIcJlrD6NhtATnCDluK12Pd+fGoWtcGGrv106ogqZdBIYvLtU8XqI8h
0L6f3pp+YgN+kuJ1vTOE4wyLdeem4oTkoTz0P+gmNvbj05Cfk2z6p9zMHRXvB0M0
7j1fVXVRkXGAV/1CvPsP1QnVvSzLK/nUm8j6YHdAuv14BpbFrFoRkg1w1oLpp9u2
j52Dh5NOqWnPhscTcvLWr3JKm6pU7+T4dQQktd8OG8fzg00+bb/XSpbSkLBmnSlB
cwf9jbotb6inzjASPNpXqz1hWPDneTCaqe+PSRJ/9MtRCvXmG3Z3hhf2kpxinIoN
0uCmq0V9KV55tX5Fs+pLblgSiOgNvsMTd5jQ6CS6SMMNiXtULc29lR9DOnGQzhsi
NsRmyiVrdhJd4vCUl1+3Uw==
`protect END_PROTECTED
