`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OXAttdxAIOrqW9Kr6gBNOJcMMS2eVCDkCeEKc+pnU7O4JqrjVSLrOXzCvaNebEBG
8ZDlK0nQF6Q6E1BFXKezLpXFY0zCM8hG2SgmFNi0qxHInVuFUmcmPp/BDWoELCwc
V3HbQD1vjXkaQuSs2tq/OreTTSp0dOADsChfRpYbvrlt0UeVq8QWlM5zroAZx0wC
s1I/dzcq9cCmpYrDpMJdcSRzXUwONjV8BcduG3XGUDMjVf9Tyfwa42tdGYVQluag
bdibg7NtwEPIf/Y5UsJc4xE82or6hLtcGof4oS8jLHJQ0aATU2+pRHnkLtZd5EnV
At1ykrTyXLm+ZUQsdsyQnbO9DDVD/r9uALGp5RG+jgIliNY11kiLBb3kYRsIBrAx
4udkmnjhboiZt8OLHfiUyP/9pPXR0qDxoi8TYvQpmUfGTaCTgQSII4H22GbZCMnR
xSuBI6Zr4vnXBf1fNDoNCv16P7rDyihr8wOVhLUGus+f1diU9RlRZtianMPoNOgB
Xi2MV8kyh7cGRtyDyYWvwldKS6KcgvZ2jN+fJKzI+iqpr2ZE/25YqXe4Jqrtf2LC
9qpqlAxRk6CBXGrnsHJruECly5b8L8E9+UvuXG80JKsYYJSeJ6oAuOpENa4i1Rix
VKNeUjTJlDhaJTy/g/3LbViM23a76/G8k77+4+/E+xrUUYJSWPmyJveETmDj2KgP
Ajlurq8/k933CJhvfnUlidJsi4VwLg6CaP31GuylM+BEIcKaODnUelTikR4kGfSL
+x9IQqbxVkIzyoPfcgytO11pS2xfoi0CEKuWX3P2ixP4hGKZZRDL13tAq03obnO3
mpL4IuF0tgLwTmcrPRxora17Xt4HFBMOfogfirnoWh2PN2vj9mGWUL55EhCT4AQ5
AUCQLNIBvYn5xkR+dnoV4raoBgOBQABrdjqK+p0Js7pXr+6oXBFfaTmdcFJxfq6O
HbAfg9ii9Fgpg96qo7eupNehK9k3G2uScTMWUZelte0=
`protect END_PROTECTED
