`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5vnlpzQDtSby94eL+Ysmx/GhC5DpABCAzyGpcyMezZDsyeivGDThpiCLmIz1/MM
HLs9LilPg0k5xjcRKfrYKQbri8WG7MLsiHSiIZvYduRx5a9ZZv9qpgIOX80ZKOqL
hoTVPBbK3pzWClBtF5TA4lvhRDdrS9d3+i4I8wi8xx3v3YTP16+RIzban1vi7xUN
31y3HppeeivjNKLA2IyEEB8UBhH0Rfgr2BXUynWmKxaAK/JlM0Iv5xEra6XIFnrQ
Vgrqv9OphAamCh8/02X9FVfAM7m75zv52KqJyN5b33Wk6fGLEHEdy/v2ZiBP+jxA
ZukXUqrMttam5zDgmWGCxRhR/oeRHgE2TR3pC680P93wyyWO/NJfK6qxySLkSeBH
TNPFWFtWujjGt4C38e9Tci4zGZ+Owe2ccSLuA4IenD5n9WTmogoWbo4kZFqpdNGH
JMByM6/sDeFEqNkVbicsSroaiUev18juwLDfDGjB1IOFaADbVzS44SGY+irNznUG
Gm3YWDzsyN4/fL808WnmYj86mt7nRblTHa/vSrEqP9IeSiXqJSOO5x8NeLUlZ7O3
`protect END_PROTECTED
