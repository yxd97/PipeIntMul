`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFZtp/CyYtNW5GCfDJHNGsK6XnH7sDu+nUSzhmINHbHyMCu6CnMafzqSsCv09aiI
qiQ+XXsgvH6DGnODfREJwe66U46QkP6efPn6HqOzJGxjMADs/cAB/lQVHFbuQItD
wjWgYX4c73cOSLQn4Lj4hIewvVOzUTjq0mwK0Lb8fvFxKNfWx0XeTblIqB76wqjW
4+Rqn2V9D1z6yp46sPols9fBFoN3zi1vL8fM3qx6vvXmw5cLQwOiQzAnr/XcNJab
5HUcMrl4x2p+NUAnAHl+Bmaq6lCg3VV2B38Wl9svNYr+b1tRjwWE/H/DHD/633rh
M8hz6wKnyqWcEVXDmQXX3e+tRxJUnrxUHXWwcAvdcp8gKsjpPEYsyUs7/Xq8NumE
p5Hg5cqnHUc5HlsmnXfCuPQu8cK2yWQSqwslBUL9gacomlHb6L+fIj2Az8OEk6jP
A3xbFFxQ4b5RFCeE/PZ3qE47ykObxzwJXzy8u9WKpFO/8XTv9We1XGSHmGaSJjtt
6YD7Mp/uFfcbr9tsp+LD/+/YDhHexre4Cpu3E1FVOuY6cez8LPcMbjm+OoMLoMSU
tQYaTlXv0axnIpahmaYexKVYMSaXyf4lEbuy5OdrlbypZ6phrbWTRpd6esAd9Vtx
7vzS/2g8iCvxRCrdW3eFNwzV0jNQ7OIH6m/kNBkt/U4zeBcQlfbj//yQgiOrAP7r
qcozIXcotXAt785TkU/K3RJxgD+T9CzYA//qHgX65ZMD6mjMTvCWnOOj1ZUvvWCG
Ago147qjAI24pr03LQRkxdPdJ/o2ymwmewMvoOv9ZmKLyfL8Hc+vm4E7t1Tf2pRt
M29d0Tv25SuENPHFEo39RoHFMx3tvVGCJTyKYnAzW6EpZ0k9EUhZKyehW7wAWZpV
LfVWKNLgT6amdsEWBjf6ogAXDf+hokrgDTiOWpF5jUNl2AVxes0Ln6WuGB1atq2V
X0dVge9ViLcdWIvfJgJfDLLyK7xBHZbroTpR9aALXebmvjJEfzO8D1v2iS1hv+Sg
jgFFFK4HAMTN6K+YgSZbDrfOeyMg7FzDWdvompi+hqCb/97y6oP3T3aGIJ1QmSao
pTX7wjvtUZssIj5f2agPhU61Qd3k/Pfx07wDV4wTBRTkBN61Gbsnm+/SzD1j5cPp
FmlpUc8fOD6h81a3qDp6jD4B0ttv8Fy6FWLqmXNpXcY0BZvPzkqwVZYk3ZMM6rWj
BPnXE98NUWriBhuLUOHkDSgWIHjGsuqz48Nl7q49atclgLPqWsTRPPPX8ABd/l+A
lLGyuhv9GlRn0uNMmA2Nh4D7WmcgylEOh2QPgLXuNjd/hnjsoymKB4XPiLsgySAD
N5aU5mK+vgNL8pDeDrUlzlpdC24K34GMeKiuCUaiAHR/9cHyYMlO8Ib4GBJE+gqV
dZXSC0P3Bf7+t51tehXN9iQuljGj5gSrtJ7WRA0RV87rIdJ6f0dAx9nRsCDKkhc4
nBWQeImaXta1/IKat9dV0lQjcIV05KBVFSZZsDQjJQRVuqZVophINSTvlwjSxfD1
O2eOAvCY6IW0ihySjJ6zJ0MLnE7fnJcZdYHc12Awp5UhOvG0+9HMXo3NJVJ87GvL
F6YKs8Y2yJqe47jB0IHKE7UfMcM3rgdggyLPldcqJc645zNE6+BulDRBpOW0+9q9
uLGaMGl5VcQcqcYgcYbHHcbb8+D/tyDxy1064Uuw6ev+ewS3HYU0qr4++DpJQZeP
pa1qNDOEOzi2BtBLRgDGDMoJ0Wla3re60+3YNltMqtIOfsIMT5T7BHUAd8Itwdob
+BC4NKUaFPkfRVmXfVNkmCu/eKdTi7nv8yzdNNR2PBUqe0xT0FVUiHDRlZ42xgAq
ZRrsAPBk/DYqB7cu4D0JRzRYRw9YSInnMF62lJZAnJeNiFUWfk0qwL4WaY21NJSh
q49Rkiw8guveTBQEHnL+jxc1p/NysaKYNTqGYXXiNUf7zrrwyBjPusgiuiQtUftg
WszPUsthFCguVO6Zs3SZVim02mrOJVfSF0P/aiKZER3jcA+wY4daiUDVKgamt9TH
Cf3YNZU+zD0vV0VA9s3r6aBi3o1BFZg+Lg/tHiZFw5j8Oz9n1vub9fa9xOBwu4zy
/SKNewIk11CMp0FbLF03bS2C2dFUVew9qT91jo4JyWLsMgCrFwvSv7WeKmICBwhI
Q7toDn2owgqd+a/T8iG44P/3oA5Y20wJzbwYx3qmGYP9XEisBptdJ3MHOIogJwnW
3+AW9tant/ciWJfXU/Nx5XcOj35Z7b5Qnn8xKpciFcdXmZA96c9qIQC5K2MB5Gtj
UJtT51FeJXCsVuC/AoUTpDmqyW1U350/FZwQeN7CabbpvpI97roo4mZKfbMYup4u
Onzn3kB/KQf8SscwfEvxIL3WHdq3B7G6gdiuAsc5KRexFPyiXiA4oYCVwXRRB39x
hzRUFxyHRTP/CcykPvXnFYXeAVqn5z4Hu+3WmY0+Kamxws/LKJ41EpzPzcokVaec
NwL7vHW5JIgUB/pZEze9MOEEh2jC+UdkqqARlGrikP8bHJBhcdYrKhjYtvUpBVBB
UoSubFqp2cP1UdIqzpsmJT0X0Epk3jnyu0C9xF5Rm0ofj5vhk28t/m/BtuTaAffD
dKUb369M72WF+rh9Vn+8kJrqsTUlj7eqRnjbAn+3mfnkfY8G2JJVNEQzBo8/chji
lAkGsG3LjNgP910X44NQU87AyG66kkNS33Dne1SxtyuLAJwHBnzqAU5/YrhByuUK
kur+2SAVyzD7i5DIZDb00HhYuZghNpWIvULOTPvNAOb2UYUAZc571n34IN9NeePz
JQ7KM2M4hwvER52p+r+gLDY4Jzrt8iHE389AtY/hmoMrq5qKgRgL5J5Qutwu8bgD
3/XOUndd5FRyqML6AK0siGCwuxVPYB3a0x7DHY5Lc6f8ZoT3gi9QOQh0mni+TA6g
HA393PiI/92HCzItP7We5NKB8Szmk6m9tQDX2Z413I58vb6UrCIwZ1cgdA70iL3B
sK5CE3Br+RL6AkG6O8JylUSNTs/7Wxe4bQonFjV25l6TNvAP0qzGF5Lsnw16I1uw
rfrtu7QJLiu1XdaSPJT/aGJq5FSGeHC8bCKR1ng5BTcXATagsk8EQzvzYiMFj0tZ
EHRaGuCDnJ4o3eTaHkcnUSiy0zUKUaJAgiQNj9O7hlepDABT8xwSrfLLohfmRBc1
3vz6q7ScpnKKFPCRnXDxtc3Q8IiH6WxKkNy6zYX+En8OKz4mDD8mLBsRwjjwhGcd
Zdl5yX7SDvYLWSp83r359Hrkcp9Es338HAir9uMqPvsV7xsS5x+zaiAY5fbeYmio
Rh0tQbopRVsxYs1JWTscfUQx3CyXftErfSpw+7v2sxBrqTPzUK54JuO8FUnLsxPB
qJu9aTdqy90OIy7Y00N7uz1uGEBUJLaio8ODlFBQdueboLEe0TDa7HZA5MyDgHQO
jlB5OAluwtTF9dD5KfEpnyK4SsPxGktziRcVzYbDDA07BhGT79lgdkFNjxZ1lqQS
2CpmpVe/DxiPnz9oYy1ddMumiCHerLtkF07bH1fH6iT/ZslZKtLDoXcwkZn5tauw
RBY5+NZ09wbwIWt/lETsSeAlI05DfAtu5CKv48evnslHZFo5nU0JZtW1ZOvGi9DL
bMiW0W7mGzwYAZVPjuMdSEDu9trixf45tr63ovDMtdxImZL39uDysGpWaSfWofuW
fl+bmMW2XvqTVAm1Gc4ufnPb8SPgx0q+sywNklvR638lm+GJ7OQbtsVd8+P7qfRM
UUafcyVMrFDx7z4QsTywzzTvvMW357SWwtRVUHMeGN320qG7UNofWbnhY2pfc0ma
+kUiEe1tBDPrffSCBvb1kqAWzc+ytU/f0XixxYDVFENva0zEFgXUmcypv8wIwaXK
VfsFpUKv2OJNfOtSuO8P5TLEzdwZCmFWdFg+eN2OYFg4U4QUlYGElko8m+bhN2Ev
sWG3j+4WDtYHa59kdbzZZvQ3bF+BARqNl7z01gGeBPABhsGYdq9yis36sG/UPy0n
KKO83tDE4p8KEBXxnNEYTqbdrVHUKIQEJCJYdslsUIXEqBl+mG+BGzgm2waznrKq
PK0MNo3pd3bPYcfypmK+8SYWxcwrQFVIcIJvuRKsQY7+hTHgt9fpuftRp5E9Q+7K
9y5kekVGH8ak2Ly5d/5Ja+kUlIgBzLJC2MeJ3F1covCcABjKH5P2rlJxfX8gbG2c
QRbzjaA5MqDJlBBDbBp9elmOQwdLjqp8MqvmM5RYPH8ilD4Qcd2MF+v8Gb9QU328
2DWCmsRnDoQzdrBq9tJYpJ5HjuAI5U8pzFHhSsRa9/P1uoazcDUj7FkVNj3KiQXO
vQ8YfTToH1UdloE3c1Bvm/Ejkq/nSt1ToWe3BJg0P/SG+zEbYLOgkOkImEuZLWgX
voMn4Wt1Q3NN1+lnOApciUTGAkE9T0ya47Bjf0bjIlULVZQCNSYvZvAbNWc8FrPc
9jWPV19nJy2s/cAYesf9U04htrIJqqjxk7dmrgGysirmSjYds5BuBqj/kaGtAJAB
kMelLfn7acnSQqQltrn31iawLd+vFAeGc/Vafx+th0aovwEGhePLI9yuK+/u83aA
mxCr7mTUuvq8wP4cLEyD9XttUDYWHkHOcqTGuVmoVcwCQAc9GMPmv3DAmBM6dvuW
kcAafrQxO4S1nuKZ2Z/QGILJuuHUZF6jkky6etQdUjJk4q4g67CIyviNi8IkLGJ+
A8eR2oRR5txzYGEpWVZ+op0e+8wGixzo8sQzS01Qf2rQVL63cCuiYtq1p36/Zc/D
00d0aCUHZOt/qIg61Zo8JzAv2EQC5i7X8guDHRUOvMzQ2B+aTeBarbBpj30Erp+U
KiTiKS/hIIdZAe1pwJu1vXnIfyc0Dq1ECBlMpSPtYRaGqU7mvDYjGCjCS6No7G43
p3mRBBZGQlvkW+rY/iKEtdQAzxQSTTRCQNYqNMsm2gQLM4uUJ4HHaGp7+DDdh4ej
5zkkzhJ7FcDO6W8g9L0yZiIQyz7agO2z8WSASTueu8OA3G/1J4WFuWnmqARuZuDQ
jXd+Wg95Hgt2fTWnz+D7FkgXVEubjPdZ/Lfi5E2zDfp5PjOPqDNa5WZusoWuc5bs
DV7bZU2ni3cVi9yKihgb1jAkqO0eeuj19tmSqvxlNp6RPbTOuYKqbGjIyWf1exe0
2vZ8I38vvpljGY6loPhWe5tzHihO0Tny1CFgw9KmsmRkKLMn/GDb4h+YzAI253Gw
wCSgFpHPbHERrXjLBVK+d+qrA0P0DypKXViGVfIqJ+U3+TfWB/FrKkmebjjkdvbE
wVigDSO4/D7cNqfKQ0LdS4884PCIWB1k1N9BY6obr3ElOSVUDDQvbEh7ZrOlHWxk
WYVYr2IzHeaESKjaGFU7sNOGG5y3dqiOhZwXTcg6PGcqwW2JBkEK7aHSeMYI2Mz7
qKPZtzM58ZBHtLmd/bTa/0kprAYCrfWureCtasfGvB/Zb00teh+Y5dxvPzdKSu3v
rglHEt+/wkk6l2Dzfukf6iLlqlqaSD9YZjglzhlzvT4L+50mUE7ST+jfbydADKh4
XF51hMU00l37BfDePeYbfyQJp85p10Me3ikR40NTumxgprg+vdeCfkDDhxupV3qR
TLUm3a1Lp3cFR5jN9Tq3PWg9/0HlQ158vh7qAoVYcuHAbMDh+bdhabO0QW+5AQ/b
dU0eWunECmSE6gO/cNKYNYdQ24v0+Cmvmi+EFhT4p5nUo46QvxBb8Hg1nEcYq6EF
eHmFF7bqtn9/dcNqpTWQG11r6lGeA53ZUGVOu0iGGfyS+I76yX77HnzBG6qe5N0+
H0rag9ZZg3gAdi3NMhzKVC5tMvC7HN+vnofmLZQiGOo4SADjaKHGB3iybJ3DIzHY
fHgosic+WDABweQRX5bEKiBiS7tOZ+b0ur9CQq/hmuzlLvJVkMJirTq1ThqbzIRQ
F60yxYxHvrANaj3CE1UgPYyp2kjLKhtH0pW/6jEENn+uY9ITSUHVkbz3DNRmpzQ7
iJmvC97LvZrzzVHkHzZOPbOQirJeZUAImkNE0nKPWVrEspLzEQL7O/pUJZ+Nd3KI
3hW6lVSEDNRqn4oGzFjcfEdvGWnUUBPvYHl695BWE5RVblf1Em6hvok4htIt/Zby
akwtc3Lm9HW3iMe9lWu3yYP6Bt6XSwCTUlvP+aO7JmXsbtemkB6HyTQ9dclOjm5r
8NL1ocbUr/6t5ajgW3QgeObILg8/2mkLPB7LFML+uIpusfVz9CDWwLcECGVQ7iaU
EwXwvgmMYql5gTNiB2Hs01WBqsFm8SUjh7wTFgcO4Brj+kooUJZrJrVEtsSD+/Z3
PpUG2gybdEepU36JlHKoa+ag2KnjntrVt4AAHPh8T9G+chAHfhSi/r6Z6o4sKH4r
RO5Yu/OJx58/DXVAy38DJhJu297RpwtozUrd8KJsvEBdbbnyYl2FJTrPQPvvLdXE
wjKLs/7sMkAlDbW2zHXauo6Tx3Bt1mcuwrO6N4xHp2aIJXKd6VFlTy6c3M+N9YiI
kpKg/KA+flWjYfF5MPEEl/Oo/JjWJhtN1Z5mQ1QJiOV4NlDtDIjT3iXLxKnwcSG0
3UEn+2JR9Oy5M8EHRlcjIXZ1orFfjzpfRPYB9DIl0n+Q0INNfKg/9L40jCmM87fo
fHE7SJzyKIU+5dV5zFifVUTPUhUvZ5jhgBWmypnvVUudnlIT5N0tjfqWdV082Ad/
ZMEG/PBBiPAQ2r5WRaJFMiusNd1xXUvKNPDk6Cx+eWEqEv2LOAn692znLOPepJ3Q
nCXGo7uDcy8xgDgq2FI5ckviRcvMw/TJJoZScXanLHvmVTbF8xhteQxOng27z2jE
W0gHSsvwo+q8qIiYKIkLYHqkSlnBmlcKog8mZPBOYmxAHuRT5RpqtbkJRt/6xluj
LTLvWfn870t/BzzNL+PU9EOkO4dH9Cp/dIESDdHxNmZ8GZrAMv09KporJA9gd+T9
rWC3tjLEDBnALMCjinHRY9PcKafe36rV6fGE7PirzRDAvAe6ZG6HXMUE+6LlT/ux
6DgGTLcPpApYpAlpc6Wf+OtI4yE5GDnj61EPBpvJVnG6tnQA2CtzDCqPYCInUQUX
tmWbHyFgYDrRSUjVru7uax8ghRVszHNj7hZaZ4vRvDmitESFDcYW2MFD1sD8mqWY
eDvmtd1MR24hJ9cvVsBPrCyi/v2hVv/8eZ5qZNVxpLPi9c007ptHeu6xniupuGkn
wxPptJhLl7aIXIPNT/UaK9rCKWurpDpwL+t+f6xwRCmCB2w4mxtsyymBLqBNMQQ5
H7jMPIxkQ3L7oARMWUGmtxQfoTPrvBbzaP5XsqXvbGkHcTi6zUrux25xKwZ4rtP4
e07fIaTZ7NHFUO7gx3TY5hsDXzyaEcmI+CrPt54IP93ugF3/FS8Us7UvvNwnI3xS
vCOlLUQxZdZ7/o9UebKrO9s728ItGuGjmLgezWtTHvLsO+JyzWYbfcKGSAi1nmD7
yBS82RLmAFo8BDfhYRvsLq49mJNHHGKiF8AAvrBgAJTL3C3WHmwYBgrVimInWmHs
+R6mGCo9f6WvdkqTRIu+4x/ej3jZn0a94dIBkPY+r7ZplemlEPNmvTGnMg+5UhKr
pYxwHjex3IgWWzIPKb0tFr8KmpGRntHpuOCS0jtFLyLbICj9WlXMUxOyAy8kzBTN
nWbF4go84FPq57Ri9h6xI/pl6Yw0NSM5mwUCP+gaMVgziCbUQIId5pnSKBbkB1QP
7O6XAEJFdAllSZij/ZgGjeHbVRRtHG6vG0wplaz02qy8vnodj8edvpn+L85vvU4v
wLmMnO4p/TYkE2peZkqqsF3qHPKloJZZq4NdKH2/nqDhyxhgFRI2oODAjEVAQFaz
41FkqMPCB4xCZGp+/W+ZttXQssBSLy2XfNaNEDH6FsssGSKz6AjlfYQPiV+lf2+V
5o32ZfwgoumrWNQB4I+Dtvp5U05LsJp94h8+lSpmI8Re9XVKuRun7mJxG3RhtLm2
61Nn7l3/oEZ90yR+Y8MPMgkAvYXUwXIuwSw2fttlXxbP717d4alvBrxj18E2J2pw
Et4jnUUf9+VFawzphrpWghGaG6/a154hkIhih3oLplY1k5Go4HWNpiRzj0viEBKc
U2XQwpvh3y2akytBDIRtVyzslJ91ml/aiIqkw6/UnePwedcvH51RM5paHUm6HFas
Opd+9mQn61SQBM4Q/Z3D9B2YHw7uqYdtjA0p5lwKuXw3WdHcIScWSP5G093uD9CR
beJesCgLaLr/Aqj+5LjrdB6lKeu1m5uThnpr5rwc174JJb19ZgvfRXG7b2KXtiHC
pzd6Ry3RXcSzCUrQ3K0/Do9iSHBPozAf1eLd744l9it7qJw9fb1dwAVbOCHeI/3Y
UOFWvSs2XyDdk7MagKqD+N810MhcwnxOuus1NOrzwHeGZ4koiIGSWydDIZHfoHVf
LYrbOlRD4vbB7AJPehdo1h5zZMlC0KkgB9omqPBU39NUEtJ7++NnPirpM4loRHx6
yQZB5DnpQjER1g2pqC+HSIy67Uj9NMjy7mRUQiSC0kqTSvruLzOBKKebsqiipYYS
HgyL/DPkM2TvJS7m9NYKMSpBvhxIjkYgzXWDtJDPN3ty1zenh2CJrwf9yFH8YWKR
CPDohASuu5twy9IdExPsKjdnzBXjlwxjlZoL5Ew0XUyGcRN/j5fkIYHi47i7oIe1
47j1dYJbrjq3xOsw8Ak9ReNBm5701R6548EZNGnMIoHuXwpXLEuNjwazqCBBdWXx
VePObsJs5eerzLM3DYnBqkTRq02hsYa9BfIE/Dht5T9NuX2casWjYClIgaQsilVb
gElMLY1uanbDxbtVmMQ149zCk8AZhK/pR6ASXcsXSrdmjiRz0KLGzTqDs61VQP/c
PPUgmoCyVuSBc21ti24BN1awsR/hO0YGNakNMb2Mc3SFnL1sj135uzWJuTNAV+0r
CV0bzcDMWwIRYtXM3Ql1j1mBLAFHhuWhtQ4A6T0hVV4Gqhjdz+u0sgPJ6Sq2nGT9
BPeI3cIaE4r4Zk5ys441f/J8oVkRc1CNjcznjCi+KcrwgQiG7w+gS88JXlNBr1LU
zuzxVTfTo4SmTn0eLJrp8kwqtCIUkbfMAN3KmjhsRFx4EywKwTbirchL8mQDMXCx
n0HxtjGiTbi4NoRhKA+rZh896x0SXANmTGViEfFSY1e0ucK+M37oaL2qwq3X26Zp
BegsBoRtmICG5TwzI8W/S6YS6/DiiNo1NHFau0WQnIfvJ5ynNe+PoRt/GL/QrRfd
rYoFPLOGgY6p+iUq0kqDYP0iZmdDrYkFORbf80WRXTsUXD2yRS93tTkIXOvNGd44
vMu8edktim/SSZNNeRgrxX2mB+17NaYJQSJFbTezufl3YpQaYWTGm5sjXvHr5UuI
J21LnyryGWYzsM2D/O93pw++4TCXX/Cv4QsnJJ4Yppi4QRsxd+cDjlr06raoFpdT
fjIoTU1O4cgB4kjQBuJTwqKdvZp4ZgYBvR7DbLnk6ksynHyFipeMywBkPeWbbCkL
LZdc5EQQoPpy2oNnvjasWSVKjRYlwoIYpoqaXDyJSe2kmot75Ea35jn0xjqFIdCt
hNB8VnRMlPchnKy5sQ3x4RD9V6NW0tyK68xyWFhPHN+E1+xVlqZggTKa+CqYhwbD
tdrmDGCrHvR0rZZm52Sj8aw46YWzRqImk8KC0z5xXtr+GWaevHvDmHOIIIN5tHMJ
imzGnw2AOV3777YBWcpPyD1GK0CNCP+NCD9s/yREie/lg2FsHgG9h5AUZRNTdfaQ
NUVlo53q0LTp0UMFG5Qw9d3SXVL+TT6OS0wEzMsripI3DTBnbDKX2nw+lZ7asnrA
K8xbJkV89ihOK/b8bPeYB/Qqg7FTpEN3VFodjEAJZyjPhuQjnUlzcdqDdq9PHmi7
QQ16AANA2K1dgWlyXoyZUHwjffG2wnFWgyKy55+uDMND9X2xqh4vTsVRPYAJ1fEH
YPFGCFejG1lY8OjBym+aDYYb6DvkxnBWIClKZFVWzPt5rB/VzJYzJlZK8B3Lfu58
JHmEXmvd794EFzggfBYkah5C5UTWt73TPof8TVvrEBchQNxYZRkKqdlpjr94DWq5
68pOuhoKq04BRgR3CcWxDmO48Ew+OW0nDIbqYxdrS/GmIj+o0pjE4S+RE+70eAAh
y841ST0eDc0PDtLEvWA3APpp41hxuHu+dv2vZHOFj0bNo46B1Fd2aP6ZKSmqeLKr
um4Pidu0Jz1wORZUMXmkXzkSGwp+SMSX3SCejxpPhSwPSu5LiENoFQ7xnV7zZsLh
e6uolV0UsLMfS8t0VLsm4ey9fFqImuapm83rCzDcLz7AoZIuvimt91C7HZX6M9hW
3Xx/7Jjz/voaytfCIxbVm/gF69wisXpKhaeOwaHH+pTmRNdyobq94pEC1wkAqtpB
inGrf8fIQG378x81WfFNv5tYRgDPIBL2YUF9BC4zK1+Bt/mcB/O1NoOUbOmMcVIC
574ZiI0iOyk1Tu4EThScIpO0xwJNMFvIbLF478DUCIS3erqaL7JtuONcF3Nw2+l5
Nb2tdIjIx6Eu6dTiEdxdZzBZqtKcIsjvecf4Z7vTXMjO159AT4j9ACNuFdXT0XxO
w655lPbEWjzESe/x6nGs5f8BNRxnwUn+juidO5zEX+pnHkvivRgkwsNJDgseptta
DAD+5Okt5ANDooNjKZWSFjmREvf1sgM2ULcNGvs/Lt0Bt0JBqpvG+Vo4c4ytg5sg
J1VGjI9G9nTBoRA6Lf086Mh4bvrblEPZdwVCNpdEfDS6zquUf7LOtQb6AYyq2iJs
APKg3Q3dBMQbin2uX0ELbe96/qXcDbpW3fpogHWwS3zFEksMmrMETq+4NdZdko0X
PsRrzAoQ4KPO3EbqZ2sunLvrYG+8U4aw2NJQyfDsIkXajtRWk1lKnqoE84jrwxc+
9o6Dhm9MBujJ08PA7hi9G2ZJcf1pFGmTlh5PYWXOH1XfZUpJsSZtj/zTmasvGWPR
0hB2JifVDKUG8J+y589FHb6BFmcdhSlqgegVPWSvSFJODvdXhgErtp0HJsUrGizp
GRl2v+hRxuECtfy2hrVRGeO16Hl6r+slNOzy9UftwatN/cfuvm4g8PuIlQsI5Qlx
z8+xjkE8A/I6PZ9lvOGbsGEA0KTmIDBW5ZDjIMUxB92GoZlqBypEdTlubYIJGnK0
GESLa+J2VCCgIDdB+Aihrzm5TdSoDEoJobiAd+LzbPZoLsxxhijSfWRt8UTcU+/M
Y7/nJVV3WywC/XThqOKi5orDDk8Pr/2z+BG3EMSyoUNnAs4o5rCxpvLu+tMVroFu
rmtuXflkggHyRbFHqYgTdaEUBpkx01vjq2MoDuLaQ2JdxBAt5R2nptiIUNXa/8FX
NawJiRApaL64mh746c+3Z1hDN1VN+hnNQl5WzddYLeVS+i/8W+xZqrTroHv6loAe
vQ6eE6ydZsPFCbgjnSOjDj22M5t1C3BSQTnYzKgQ8uylDerHXCRmY+zRQaNu23St
c8Vq3RCpKCVj24cUB59lL3NBZVZmRMZ+zRJEEThUSGLBmxTTNoIul9K6aGRfH3Ju
rQpzYIlNpVwLH70L7N93n2nOKPMh57neKAf+BlzTVq7j275XVbeAncGjQ7aYorsS
K0GEbZVDwgKLqwvOU8i+n4S1E64CnGqkYpQz61wxoGIOxnn0zwYj6WLqQTvYUgOq
22RsNLPSWty21Wx9Svytu61p1H5Jcr4gh6EuXqVA5IYuRt2YfFHxcOuL60LP+Ko5
jsZcp5RC/0ec1uS5VsLh9pS/CJbchKavojzi0ay/rAFJb6cynlXDXd1XwnE6c3xc
/YvoRSq6lXTzPP6AD9hXq5UkbLwIvVoZUtK0f2sUEYFDW4QOfadv2ki+HX2Irese
BmWwRGSvtZdvor6XFgDAZ5/D+ASYF4l/UiTVS+QoKjh7yv6Q5DTpxER30Apuw/vk
b6ISG+L9ciQnOkj/t17ca9TGqbeboV1OatODI1qBulEckhVLXKurb6nTm3Rgct90
XarRIbe5/9SQ6LeeQ3NFA5+ET0yRjS2rf3cgK0soGRZH8vKrF5WxLb/R+zmhRy3D
8OpaZ3mBbhQE/eJW/s0PSXgMonpEWH+EWVsDBHiGT7FAwZ1eSa55fx3iG56avXW5
bemAZlOgTMedU0KTJDfnHX4XzKtXGFyZ9s8zbHIc0rsAf4KLPNOBMU05ocnG2wfP
XNLp3KrZfRheF82+079vYVikrePdG+Zs829M1RD59WUdoOf3NQStn2n1wiqJFnRU
G7BEGb4TXhWiGiY7aXGaxY/yVPRAoNPg1fKRlF541C7awOYz6jP0fXesUXuo/rA8
sPuwp37SWXun7A/8/zmUDKA4A/N4jjjewqt4D19FFloYSTUzQ/G3l1T/icHLUPOh
fX/0sSq21cTkS7Bsjmy3T6Nmc+pd8Mjy7jzH5Ej43IVtrNuE6mNXQS36aE7AmMwD
6ki06xUlAMFByhVFlgr80K95E6l/KQiIU9J0ixEn6PeeQwqoQJ0p+iCkQLF3unMf
n9DN/nod5bouhsZhubDLgquCCvkg58KXZvvODqwqvc3ZDlPOUARyfYvAwvXLXwx4
EL5kXZgTHJz9Ip7mdsS7kUnxmjye07WQJZ3Jzac20kJzLjFVZf/wv4tDO4dEcoS/
qwCvLYGJkVU7y381dhedbVDwvs6ovH1D/Cp6fwwTER2XrjQZ6B9+An2U8JLAH7gv
MvsPtSXbBtOAjsLiT9ueb0e430TCCG+Oc0bPqZ1ymHuqFfFvk9djhQQHjGgSCcTe
Y45NqAZ6vmaM5JLJl0A6MUKXGq8RlfREOzMbUrBfjRp9JDKSwALdxYspC+Wt95Cu
449o/Ji4iO64M5SV6gRNTZykagDttTN3X9I8xZTSl03Ji/3ENqYxu28Yy6t6xJlY
SXA+QYXnlc87hqgsHpOmU8P0X6L/q2Zh2LlWijbzoy7yJXTMrH8H4/qUJ/EX5gQl
1HRkpJBFROEuXJC7iD8nvacjxd+3kxY0ChpzwYk4/c8VIVqwvv05flxJwoRPRtHF
5v+FAVvFnA20Tz8cLgDjLQOfxPeHAjnEvLDdLauCcdAuuZ5dyDFUmYScR/VWXOGp
G3a+w7byUqSi3VHBLacfHzKpNMEFqReIkXVoNCJZMYvj2/1rUYlGicqtpU9VBku6
ls7ET64Do01Pl7hZglm4huUE0WMZELAxsamF6hEgqG9y6D9ukQT/qPu269OCNxox
UTace76SpwTLtO94DtJIYgNUPYmnwb6+wr9I/tZb+OBZ2J01UBB+ZNr4q5PAgCHx
A8/JtoMWjFTNBYv2/ZT77ITFjqo4rxHuuguqtw/JEJlYYjkyH8QERwv9JMGixCni
oeiDfJuPi8vhyRsfWsTpAAk4MxQCURWtAgeeOrAsvbj2HgUx9u91Ufp+jMeIf/tE
6DckbP3smnlhf6lcHuvnfkFhM6irmGkMYAhORfyAr/K3LwCBrgnn/P4UJPDy1mFL
lv4eVI+qzqIDFGIzDxm/H+u8rMm433ajieH0VuHCqSnxpudhln2l20SA+IOsd5Jy
DEtHvntr+TQGHrjjmtKoLCzJPX03uqewM85gq6gNk2D/jc5xqgEw3ZjKTUTd4d3F
srW1dXjKS3x47Q9t1X0Oe/xQjIAl6s8BSxiMFMu8NXSwXB8BBejuCcjiLh6mTTfD
5KjvIYtvRRhFWzMPezdzsThefyNov0q6ss9UBEorQg8C3r40iDUpQ3y77E3LZbYy
KnqJFvDv5cyopC9+WAZpCVvagufPcFhnvWz1FHFO3nJo0qS8ecFVeFbu2alCRwq8
TVbLoE6kNb/b36wJb4h0jo2flAyvmdbP8WLVMvaRuUnXQNqFOFIQq+g+C7je3I2C
TcE+yfmHTMfKXsWxJAODj4D2MDHF+De3xzPl34bBBDCgOvTBeOeK5qCOzlWkINmv
5cJv3wkJind8ONe3k43NZJFoKPIErTw3M6d04EbwjfzaNQ84xuZpF+8jPS2Fcezt
ceotZjBd54//bil1CPyO3fvhcZwRhGDUA9jHilS8/vwGWHitBJiXM0BReo6CND3U
w7IizI50qFLwVF7MrtD1yOlytitMlqlkmwbH7woB1nvz4Y+RwXS9MrVh6gUoHkcl
OZrk70mM24xeYJWA9FQDjcadT2rNsNDjLy2zSIzFUtGGZjZQWeC8bSA/Wt5aS7Xr
gC1G5cpGEBDuf1rGNT3ESZV4JM9nGwA4G0uAszEhZvK8uf6fqilBubZKBfFdnQP4
DZVvmZC5F+loDvYRfsQs1oSJr8GQ+hs1lf6UdLxZVFxBJUm2P7J5dsv8zQ5SmFvR
qQQhicLfFDhV2VtAhgDufr4PFCygkwJ99ZWo/w5Gx//hgzv82ufG+bAOe2xOpgMW
ceY6sjC5f3SNcoXhi82ARKUaKrdxBFdvfovaOAN03yUO6D2rlIOZUSmPpbjR1/o+
jUzsA64hmQCq8SpuLYqRuL6Mhzg0K7HIFNR5c2PENhGWvMrYWVaHR3dKqVHiYsdJ
CSIG9V0K87UTez61qA3WItnknDhRKCvbtjoiLFnp5EZWSRiXBFnwod5GD3q5w/vF
JexROKn3sABqKW2V8ADByFVewR9HNrUvXFwhGtmkj27bLmiT6NuGPTUY56MHzBu8
ZI7R6EXe9hpEkKuw4H1uZPC2k2REJeNuKC80rbrS/HZYaWFJrS4B2inFnAb8Vjbo
PWaPVHyHeoXF94A1x1buxwhsehILxtA6Ex0TNCtfIbmuk3oOeteJLpErF31Ph36R
45CWXl2Qin45IOIjeh/rHocopWUReSfE6IAkg8JqTRjEC6txh7DFySLYmY01pIlb
xywDFejtjr1E0SI4U8avK2Cn8svYn9Ut4PH0nskPsNKCyQ3600B5+a+lJd1rHyoN
6v33MouhbNnMQRqrt9DHe8RWuY3Mw2l2JnTCrRGRLA3zcdN7GD/9RyvYSGq+UbxE
x5Y5As3oRzsw+fpwAqtx4OayEC8ETe3UwoAYZNlxID8f0Ik2fJfE+ADdeS+6LjZa
0rQ/UITwYdI0VJcBC082pJvxpHdrn03dGqADzxafMN0m3KZbRNb3H/tAhstHtfsZ
+qTnBNWe5c2iUOKRJm+sj2c/6o7x6PVY+aZC8a77GX2E71o2a03ukdUwE+K35/MQ
RB7O1oTrzLvqDW+TeSHx5z91G/2CHQsMLi23cA6cpYbjpT9+7+d9gDSqLb/X7pCe
d0LwF5v1C1AFmagtmEQVwz4nXn19aKbgebIFZ3am9zl7uTMBaMk6Muagv8NZ8mn2
dvuGodyVCMgjTWxyo5KmVElLbFQnZdrB3xRcmww53HDb/9prO5MdSrMyrfpZN1en
jSBEJ5sTdv/JFV+VDW4NXY0E+HBhAhscFhVodRE1fYnk+0y7Al91sUXP4I0dgE/s
Y7gPRIdUvGRpmPrHb8ThHoeV/kCF3+g9npZw2q/67OtrD9mSRPcEwPsTgm212a2n
TcJCWpVUwU8d+uuEZX65tGc8L6yL8s/H+EEgXfeTd1TCQc5ydilbIe0xT9MtBRig
vnloSZB0+Qu3SV7+10n3JcREYFineXN6fPWxjzMPjmscrli8NQ3egQxhUA6MT+MU
MrnRD96I+8EvCSs2Oeh37OADn/tHnqGOIqV9MIv6aXmwA8qa6y4/5mqIsYv4sD/t
lb8QGl2DXnRWjgnXFxo7ikYY4KfNwOcmYPA8cunMmUubFI0yUc3QSpfymNx0VSiH
9ZIEeGpzKigGBixPlK3ba0d5RsLrEjqmjiZQWYTyb+KSzSBA6WgMayoneCBgWOa5
L/qWKs5Ia3+aKIko43dCwEmSkvCCMAo7BpDFnZxCQaVczqEIr8MmUlnSEBWMUn4t
frx7kmVEViHYY18oXKVf1Z4vnNGB54eNCaSjxZp67RgMGHo4PKDusgALpni76/b+
ywEkc1jUK84QxthPFzeuL5opbQo9EW2X5vOa5l2Iv4FmS314F+RTJBL0ZVViE5Za
o9/M4elwrUMKNfpyy90v5mcAj2M5Mam64kQl8wJnAr3IFpa7iaZ7iSdW3UYsHltx
RRmvIYpl5fgZ1PWghNADqnMycgibxcL5f6zYlWgVTAvdbiCjKn1k8o6l2zYxvbRY
jJb/y4iCZvPQ+iPvShqVT9YS8hbwiQqizZzi+F2Our1QR1axEdYCJ+dz6NwpkQWY
GGuFEy7UszrgYXF0gNZhl190Q3R9k1TKGCkdwMN4FLDLdI8vc7ADBbau2MAkHp2J
oU61db1+eYKggM4ZzuMdE0vYos0mVKJ+1PF2iv+JMO7huQfE/ldVvkc1v3YGGSHK
MQr0LVCGYN6FbHDKY+QOts+r4KodpoVHVrweu2Xdfs+m07QeOxtIHq0EDhLDp3LA
ZgjlUS2RH14ck+AfFaCfASd+GkVLRxyxO4sgcVjtnjuiAAYdU0AZMuyw3PH3r4OI
enSEwwKx6XLVjQzMsC2qupi4Tslx9jouC2CpCyHkYdObZsM1cwGm7OwQPZ9Lg9C8
CdhAVta0pE13wtDo56vVPrpzchwIQGGZsxOin00nSO/KUiyHclMtYrK/o2WppfRI
3VUP3GUHaAuEi48QtWNVVEPrItPR/TKDPYapAYaPND4plWRPTGKe6hM4XH/e2fBg
FegCrZ4wbj5+qp9PkhaHqwNVHeuzzEZt9EoLdjhbTE8rXlLvfT5xuwJkX0Bbt38A
qN4CJbVy0f6QaAP9/C1tVsgbTtxsAbcgmlq7d0jW5GW/fleE4VNUo7iE/qQQ3p6n
pFI4ylv4DaerHK5pDBHTr7OQ07jwDPCl0nhYB/3aQV1xqRrbrpA90/b3XJnS3b1J
ZQQYdn0PuIOZPp4CsjJyHZbIs0nWufDZUGY+Ea0AO6S/zCi2dLg/yWJkzopw7rQr
hf11FJfevOSrTajo3C5X6Mz7k2wYAFZFlCeHSCacjSicij7egSZsUsGaXGBotzvO
OwbFpzNrw/LhW5PyoftIbwDV72VfTGqytaqSZ6/AJ2hROlt5X4rM0DdxNmTsX79q
qa8drcSSpWvlvRM4syM1RQ5rXUUoYzFYKw6u5qycJaYUafXEI7QB/ZG5Sz66JWzq
RqDU9ZUhuWAeImZxDsZkLLsrk+f9jeB3+unW+9/l3wjjEJZnDUtWQyCDGnLluKsn
ItktO3G5GLEdDShUWnYOfFBI1KYTq3nnJXOgljxXSMz4gYhTIqR3YpJVf6uK//Wd
AdJvesNQTUjzR+G0zN/kBArsz6+ZIcCqNaLq/tEEKXYV1Vc7dLyIQdVF6JarTisu
MelYiwH8Q9UJHwA7VixVvc3yB2keXP49Ff9B8rBmZrK//jm+JECj83DOB3GWppw+
uJ84w9FP9k1x83fD0kd3qXT2tZohgYx+9PIFwCnjFRQDwJErFwH7JK1K4RYeMlM3
CjkCG/mR9axb+sQs3H0bm4c7RRwrblAg1pXvzMiKmdKApLaAypF+ZfHxO1f/L5Ci
7ohMuA0ob8zH+qsN41hKa2qt4IW9Wrc/QwncXk6Pyd3HxfXNufZSHgi/ClUyENMN
l0rkFzREkUeCukcwO36sZlcQhBoIN+tmBUygNGsg7DBlTeIjcEpWNszCdgo9Sm1J
F9Zy373sOg8FF5o5hR2YywXFr+kVRv0VgaNBzFgIrsT/7HWqHkZ+yTqSntXlruk7
GR21XWIkWJcBilYMS58GgwFmozyU17bg9yh6VrJdbbz4FvfPlSYV30EDs9pgv4Tm
OgEtdRLneAGfzlrOjLu8ljE4yzZOFeaKCrdt90t2wWjCdtesEnrjJT8biCar7Fm7
yF7lf9rfwIRIBuDL2iDhS7xUHZ2njPGb/bVKEM+LKlsQZ2OIJ8Z0OKsg7L5/J4MV
znqwkZE5vCwPXyRlSOb/OspWcZPsXVGAdgOQa7KUOwcp88EIJuRy4XP9bP1bupdr
AKGBMmnbsrAQh1VIvkC+svd13yBSkoGP8QPxs7Tr6yHmJ8WVbrQXWtIdtSb4Sce6
P/PqJ+DSHC+TWqO9liZv0KAAjrpiQPJPrzbfQrGIG+7+jOCU/+E5LUbeuSt9oCyI
UolFFmYJpK7vtQubBl1EW/kmjcjU7dvLRan4x19F0FHlBW1k82kt4DFwfucvMfCl
0qfoQKJ63sN5LSwLlUc1udErFimYVXDHiPj9NoxwOilFshSXeuW+QqowKSGlrYpX
itLtHfocfNvAynGOEvib9A2iDIDFRki/iFy95uWqCVc8PNmImVcIOrDdB+3irfYy
tjzrDf47W70TUVWAE8ZlTuKgUKJda5r1RLuhymJ2fINBjN5OdETyi2cKiQfSSqhg
XosTV2X7lPhsgwqfydQ76G8fYzmNXkc91jaCof/9b/YYiin3Q4otjkb6jSg9zaT3
7af9o7DCtX1wswQHUxBLXfTD4cDbfI+GYQLnBEDnwcnAZ0wlzUpR6Hb7P3pDxAnZ
7ug09FERIJDTzSLvdyKCekTzer9Gs9HfhUvt95SkRivvsGjYzk3hjFLkcRP8Ql4n
lft65cfdbAfC6XPhS33Gu7apmyZgA7gI1DH1v+xTr+6N9ELbND0Vu8XiiiIkKbA8
UpPoDeDOxRrAPBoKc9/vAw7E6JX6tJBKeo0QRxO8vMAkooCZm3sYMhi6YL6EFZpG
sI0b0+UyEk2vfQ88vRUBD7IqjmdGvy2evOUDvW2x+Gpx3vDiSpSlfrZLb8tP8SNk
lKxzDfJG+CXaL4fBfEC9jq1+THePjB+gTxs4HbQWEVYhJeeTCA+Fgo/7tQ6Ni46j
hCCZaNg70m3ESkvUpOt9v/eofhU3VWkz7ASpD4f+zdOyWF5nDNeCO8o1u7a+t3Iv
bXATjovGj0p37oPPqch/OlFH42ftLmlRxrb5Kjzl13Fi+l5EOaiLwV/avvWFbMUY
Y5hdiwDukJB6MaNZ4sB063FfZr4983PfLFtTqxLVvjBMFuxTUnLcKq4COCf5Dv7O
7OgjqO4LnlAml2WihOKMEVcvF/D9VKYo8FVtq974OFkz184E6J/KOzbw7Yf4NV+A
1uSerxm+jBPYICaulqnD6Rsk/TfvCKMb9Oj1lSq4wktrFkzsNFJ7YU24r1wooWKQ
LjxmUTCFhiDtPExHh/4Ce2dWeczqRd2rGu4CeOLlv4CVDjaowINZpJUFRwY63lyE
eSWdjZ5YYSiEY8j7HF2bgYF2/rGv/Ub6wKzwaLZvq8T8J/Nzm/S4rfwCTwwB6i+e
PNkvVp3zVqTKVJDOnSaFu/2u5SfGnQ9al1e0CJiS8YNoGU7y3tqv7fpGoUjiIm4n
mDXVlDEJThNV3huKQUznLafk4qiBxgC2AcewNJAUriaV/FFvALv+5i+pPbI5cPkV
qvwLkRMLZKDNB+DduuBoyaUnncd65tm4Rqdt6ubQHiL4SWKh32mtjgQdClBbbBcA
4HZTwPPOi2JueUzA+JZOBKJHvbQK3QA17EgW1yQitbtqt63T9XnzWgYrLvvtU1a/
tp2Brx1+ZSIQmus24w91SqFhZglDpJN6XSOBa3n3rg9BJBP7+/M2S4U+Va0tM+e8
oqRbdyGuAyUndSuYPQcwzLllq1/O/KDFXNdrG56dsqyEANqBxBx7mriTVcp9Xmvy
1uZ/hRTY7iErdYPLUvFWt8ye7iG7hlSEp3sTZzTLf65uwhYr1D0XWB/0GLfzJVUc
BrkmZjhhmXuuptckCC5+23WuNGVttk2bEi6YmQ9q2fdu7VE/mxJxziD5CLn8xYu5
psXpdMh02+CxrXsGjbh88+axW468eVzEphb/KYHbYJhktYWD451JZhxm/pxeRrdu
NnjSl10EUk2go5BL1NhQnCOsJjag7dfOKsO//8dJCPGEY+RaPhWDiuPCNkgwfvLD
TA5+v3Lu3ffMeHyoDw6nZTBsQWNmRRkdqHYplWXjeTczPIgYVhiVEKGYqVcSOwGH
D6i/jKVVriPnPNzhiCdxZFhV+8duFCC/gUIcIouOeLos5dHSAnvInNOF7eNuloBa
7pRI8nUGcJQm5iFEOFIorUxb7c+gXVyn0Y0eBsj2r0SlgjdfQCOi01Xa9w9bZIq4
y2NJOMyxBecrZZiY6CB4BUObv0LGCkvz3spt/ljTRkwe6ODTnPUns7dush5Zt1oy
6oItcpbXG5xI7z81CNNGtxs3HnG0nrQFO4tZ97u8WEaQmkTIiZbBNq/frxLk+n2W
NuLR/mXvPNAVyTAENnagO3/fc11vIOWElJAGPE5dJXeaPAY5BzPXJVW/TginSxSc
hui+kOVsSH3Il0V3Unzox1Dhy8Lfqm/mznRv2VkMaGn8QW5t75nSc2bk0+N2EnJw
CkyCcPWkqrEhDvCSUSnI9SBmqjYvKx39LhiJSGb2M8u3twiFofVugO1GYZmNhmPv
R32NvBFsNEaudu+rNkS2N0sYrMjJbbEhKPdKNZHDSlyU0IABO+xb5XZr4RG4nGVI
6+knRqPRJwEwvV+f/6FsU6iJ43p3iAvfWS1609Pjo99xiGBvHBjILwCY5y4JjGfR
ADVhVzHwmQWVfenB4pK0u30FdO7tnewLnsJ8Iz44rx8ST0ThNkIlUI9Fvmws89AC
GObPRjeWRYA20YaSdcujHbi0S+JQcLVJKUQtqkqGTT3DB32LfjvGDKj5o/8AGjHH
a7KM8khhfXARmat9V7yyFgeS+0OHaE4NtMS+Kzcs98r1cm4CjXO3zfSBWxyXZQxo
s9mbjN1zSvoLaR/kLZ5yT7ZdtK2HX41foQUBYEHG4qo8ZvJi9HFVcNUaeveR9Gz7
dZonPrPdZ+y9ojvqxmiFAbQfCY0rwp+OW74Po/DQrG8ICmxJL8s0XLESPdMS6TkM
kDy7HOTqHfafZdw1aabG2+0Wk09FN/Tv6n9NcFBTIk+O0nC0yFkm1BP6KODHIC3M
cfUxCXDr66dpgQSqX/UkNDT/CcYSeYb6seGNftlajUPhtVjq5DbN71VHMcrB6kDP
vyilqa30umUSjqCmBCqoPszxP5MK1loMjo8hNOeav8m7MccOJGgkOUZ8DW6FFKij
d+ANYnY/aBz5+VFkzXDxXNR1anZUyWTfPFvYtJEwSc62dIT3enVfr3cpkrauAyxM
jx9wd6yheQN5OgMH5YwvaKxeh783x7GuqHzQM25aoQ7lUL+n0Zmk01ySNIBFPhOw
5MjLDMcMjR3tzqe8GuZShQFOGldpFcSFGEr3hbYMnHlM63iWWVgvy0pei0+AaHP/
PtA9hy9brvrHtPpcOGSM0CXaD5ji8z7SmWEnLYj07uO1Vw67WJ/Yb+Z7Ty+gx+tB
FPiCfY556rD559ARznb1Jy/cg1WaqGEaI8QHlQjedEKdV3UCmUQ3VHBnAPOGcMpS
FWz9265gtecVZ14gD29hilOPmy1mxy+3ww9+MQ4/sTjSxSuyC8Em/7/6ZLojWbGR
sgN9Ze0kPvSxkieZ8cZ/meXQmu9J8tBUIHIocHCpUvQICqzPvAednSdPjfqjnr7m
3+XfHl8rfDF4GvprPYNaKncn2sjI/gN5BFO+muPh7eXw+1CSgJ60gekqD6RH0ww1
Zb7fBn8R6uLOdXBQ5EDa9lDbmNPSPhxq2Ly+ecxrNruH3CEKtLNBdQMBYNNtmRdC
sJGkHGsOZroe6e3MxmI+Z6/n6kuZ2yQGmPbhyLWzXzxr1v0Xxy3T4zbBevNgzlrZ
CCGwYzsbRKuMwnmY7Bd8ztnxc0fxaCP0W7oyWuKpFREfRwZl2Yfn6OYx4y1wlCz9
NHdRzM4BrQBooq8XsYsvClBccaeMNus6tMJGRX7U8BJJvtNmWpAg8bOouucRNapo
suNYFC8RpMXPnQbAwRGSw2yaU5vcNJOMRVkNBdqaLDR3CEPcIfala/wxqjFjKWDx
mFdwgzcKUXK4FlcepPDo1LgKfZ6wO4DolP3ZG6LfYut2fBtBMohqdcEmPxmXKr4v
CwfBSoggPjgek4KKp6+/wJ5LxbyiwCxp51UagMm+85BDlbAsf5yZqRcDofnwKyDQ
PNG5c3cCsx0kEPbWEapSJrb4fHdM8R/VXq3M2x51fOBR96awldjoAalHcsqIxTsm
887AAGgPnQVvI7bdIxQd7tHAQElrHCUF4eTlOhKBPSWPbvMS0FhI6WiA7+EK5fe3
/8cn8mG5X3DvRzchvnTYTVEwlxLqEkuOZFNdnYav/ldt8T5lknaGaQT7wRljpZZa
SYYxrkypa091TYmyKkc/P2M+oWGFIwlwHH3JanzJnn0MX/OagoPjFEahZou+04je
vpIDzC/9hHBF8/rkpxJkgYaZ2m60pM7w4UVJzWRn+j7jBS6YeFiY9kJq2kzxalat
swrBJIxpLD1tDUcIGz8cNkLt+PQh4vOb5oFIwELMm7nJlpX+CORu21/ieYmq7AJt
fJn1KMgJgiXFH11qfaBVa5iHHEy9EW72i8lveQX6qImDDdWVccTXNxB3/hfsRVta
QWFJc8HtO8r8qdpxVMpZU6hxqGoTl9P2WW5xaYANkm66uW7OQnwu3yxI2gHrSEoY
1ZNpoxcwPxWaCvcHHhC1sQtQRYXO5IQV7zFauCKdEkziyI9JkqjuAY8vmvZJY0HR
3KxESJQT1xr+FbV69JDnbqvVBZYGZwEe4EswZvi7up5MfoEatUNYFSC/11KbpO71
YuQrDd9RyBqvEXP8JbJNfOaFYhHbZSpA3Ont5EvGpQMF8RmcUsiL8XpidmJVZexH
29wIDHV8k2ZoWgyCakwGrb6OmzErescFxAFGVR92mZzJ349AM0Hj4ULKVQnnGKNw
AFUN4KgImUid5mKxsD6sk4zWesfO2UVfvsG21Is5EIUh8o9y/wUdoFWVt+xLe1/x
Oh78w5uw2cbVZUGZ6Vy1Pormkrf2Br4E21cfC+L5JziYMaLk2h9ugSv7ykhA/cSq
xjEV25mIUpF27NnIZ8lNmS5jwpK940Ztk5eTADvFESNER52PiZqXZL/ydX27JmEB
Tb6y/Ir9UmDLHIsDxubzrD62hG5Io893YspgaThL9qT5OVVWswcOe88z1G8RSiSj
uSTl/h9QAJaDLH3OT6NbNegkrYcJM/1CfUh4rqu6ivxTjg8d0jlUZboGNF/SP3ob
vdyTKiuUKLGCp3LIWbNquKzRPfvZyC7qMcg35jIun/D1vUAP2/e8cJqpOJwYBoWg
W0Bmy54+W6KqmDsJkCo8PoFrZz+YgCpXIIWj5PrGaKV6CPqpnWQrlKZo8M8A98IA
W6G1DvsSjVWpOB9VY0v/oaWYJBAy+g7fGi7pCTmtg5lBfCeEfEl9IVhwtF97RT2n
TiO6eDq+hJzfpZzqSd08hb4IUkwULPUEu5F37MsFoUcoFopeFqcaucd90oKJbvpq
VHvsxEzOe5SKlCAOUT1dn+oRo+FTpjjnTBKxEt3BkLx2Qys+oTdNOdkvYwBdwlT1
6Z1WaXWU46fzx2KmCpR0nZgN4L74BT/K/brFc73wkl+Dwuf/VfKnnEbx2xVznvYC
DNnxX56bevmqt/JHBq+LNZRbSYNPLG4Ya+LlhGrjiw3Rvn2MYJMEtxoEcSHTleae
1IZ8Ds/OkyFzo4mRbuZ8fqMWm+WxDS4aUJzOStDUxhkTKJiNwW8Cx9T30jMuJYxc
7nIJDUS7zOBXTWQT6rA1hA9kxjAPfYjx0MilCZC+v/fL98SUCtoSwOpchJfLeeXq
0HLmLdIOb1lJwun0loda63lxpGKZQVVWemQbE0iZQOmBWuZp/L/hQFetYrrYSYYi
s1aozu2SZ4JNNBjN9WezCQ==
`protect END_PROTECTED
