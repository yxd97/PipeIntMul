`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y19l76AvlRDm09tNB20d2Qbya6DSl0PU+hT36Wh8DpNyhb5J+p+qFsQC1tDNx/2V
JLWpuNKdsqWL6NBOwuvJ0B1UVA0vtp5sknKDq9SOw3DFHAz/8oqVX1Gyhgcq0fTX
hxeNQ+640n24aMQ+8O6X7UfeFLpYvgWyTs7BVYuAfrjR3eKudy3yoeahOkwAh6BK
EBvhSKorl9CKSrU1EX5AEvrri8XLQ94r4F7xqK0fIbTc7q5/aNP/eS/5LcyaGhRR
tyUn8SY5M4kG1tq5oFzKpecR0aikldkZKV7cGCwoL8suhhIBardLogvFGS0cMD4q
l+Ywkw+iDZe33QMzIOiOrrJPN6BMH9lD3Nqnsoy7bQMcYmXfRl54cjfZxI6/rp4P
OhYyYCOT3oq+cHlS0QoWZuJXtKXy7SPTJrIEzraWydvos/lxAXDVoAtZhsi7zuXP
`protect END_PROTECTED
