`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqJ6jgWbZWx8wczUlEZ7owWjVkTPGtsq7LWV1US/QfzeuR2H6peu/sHrvMTEo6E7
SRkxM79jUOkPdWdhpooZVlzsKXAI7zNH3UYkN8x79Ef8hVohJG8qjYB6ddo6dLNo
SpTwM5wfg+hQhCAoph0RTL/by79Z2Pq5ZpQn8UZWuXCjOmOkOqnkWY94Zy19QQCK
nLi4HjtHxWKEWa2wvYEE9zYLNqhxysi9PQy/sImDAqb3nirYXP8tmbdgzlLX1rUw
pSoHEDmQqSGjwABOS56ZY4wOIfWMYms0z4FY/9Rm1jG/uVL8qt72rGRb6I2dS/7i
RFq4FXuNbQMt0jtSq2RwVUFN5r8hI4Q/5GkRkwu4uLyf8WxaA5krMxgKTB31xK/m
ntCMioDrXWvGYQ9BSB6VcFFQzi+BGcpCJ748xYwl6qBCzFu0SWoqaPlMnF4aF/lA
lZv8HRcEZon3BJUjyIeR4qN6RMir7VomheeWDCCRXgueCrAAIN00c6TRjjKiO/BO
2e0tpU9Xjh3haQY4S/CtMNHLMrKHPsWBqNj5Q8xtxnN/WXFU0u9GyVH5uXVAz+ps
kDOYlI7Fh0nOT2klGq6wjQ==
`protect END_PROTECTED
