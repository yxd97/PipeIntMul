`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mVP5dV5ZwlvoAnBTMgxmTzdH/1OSRIBoTKEmqWcJUF5nAo6NgYzLBORrZpKc3xX
jopXLmfeVYsBE66+2AC+hBpqTwVbO/4T2cvMXxkB5GbW4LhxmB/XdpIvyRew48ut
122UDSFISwF9iPK21SBRMxgBMj0rlfC66ZLTKS3rX0lCxm08L1+XmvtMymEFcZ/8
xzPllNjCa4B8OyIkd2oFtmrvOXR4W+ZS9chkEROb6vSx1eZnfOvMXwXXkYmfmQE9
sVTUT21fMXoCrCHwyxiYWQ==
`protect END_PROTECTED
