`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WvcbDL/RvVb7rsoovzFxEwKSaJbqQOWHx+w0VtaVXuds6kq+l4oi/nfJSTKRr/f4
tqBoGpez2SwrqIY0kT0bQZ0s0tsRMu1hmvU+Oc9odeFGtBVxxe50LXLX5wHw/oTH
H5RxhVbCEDA5KhxF+TWQlhjEJFXfuKR4I25BEPX3uw+ySk0pCo63Ez3YtGztEWVY
0bYh8j8KcQFGCifG7KdRn4p8/51LC/nofcE9hWLLLKmsXJsNllccvl9FujundLfS
PtB0DKPSTGq8lbi6udAArh+4FIDsTtNkmpzptSuSTPAnObdiebB+zcbPMAzjWVYY
dtuXfYkpl7HguacGTlGKv58jEivOwwzZ/+XwdIjTMsCw3Yr/o2PRfKJ98vvczp/d
L/ZDKxcSa9WsUQM/cc/WXdYUUBrxghogfOWzQJ12/s3RokB/LwJcytseqrwpt/Th
+7GqFj4EegloqrqMWW6eg5ISwT8zqr6+XUfXVPxYZgVJmVs0laNJPrGanaru0MJi
z9FmFbx2o97yfAfxnPhy/UqbLdBr4rXgH9HATheeYwDMUC5RwwM5jT7x+Z905WXi
+lj/5x/s9/RYj93YIoBYcf/pt+eCEpHug0//jnEFho4PKZPcnIdFQ5gBU4MfXPD4
PZx5gDNDwBV3vu4teY+UFSG6hcFWgiVUCb2nl7L57ut5X5Po56uZFsUD84wntLKO
ZUm09L3hIews8vncTTumF9knedYD7bqWAQEHTkjn/H5CZSOCe6UGBLGS++XzY+hV
ixJZJ8odvJWuxNu/Y1PT9Q==
`protect END_PROTECTED
