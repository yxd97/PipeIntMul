`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e0d9Wdx8TsYtE/Uno/Ll8FFZJPdEVRWhGyZ1j+Ym1y4gAuUaXZSVrGilhKeL+xDw
qRvR6SiYSEhSBzo6N3TV9UQ8r8XpU77ZOg+GFgE270tZuTNEZosOOIVVlKt6AO//
6kYQwu4mlcx5O2IkujWrKXKANuLCForJpsSktVOX6TTyhaJt6I+dtQrS6VoHMXUQ
p1Qh7rorRn//5PPnpR70j146z5yapXNdiKu3/Bce7GOrQXGqQH0C80jpHnCcT+TE
x0mqbL+nwfx8aG+Gx4R9+HLZQAo0aOPOdRMKzDAcJDT5NVt2SsQC+ohJJ+r/AaI2
6NB6q8MBu4JylPOYhzgoQA==
`protect END_PROTECTED
