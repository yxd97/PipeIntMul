`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2QKsWmyZwv3Nhu8JEauIu9YhEgjKyPf8o8Ibe/AKWoUxCyXTXbLGbyOs1GOAm9f
bv8jBO88/Q7Exn2ATnjK/mdaxjRTfQPtatGGagyfv/Nl+KgGRvjITeO8bEu+d3t8
6JRthIzzuK17L2gPOciH7yXR9p2DeUEp9XFOk8NZfTiomH9yH3hF7OtUJ0n6wTJ2
IgIEU6QX5Vapz1G3WqUTfBRIhfimN8BkstBWXV6sfhm9/moYwrwBMBnmlIeIs7uL
2TDCspTvcok0tDaepEGZIxmXb/HzC8SQgTkUzwFY17KvgRdpPrnK2T1Q7z04aF/E
DiitBO+lwd6eMMDKIyfy8Gz4lLBFj6ABAMm8JiOW+SzvY62C3jeVF2tLM1Y2qfN/
ekRRASvrDdgAkcY3GDbCIh7lRlhOgWPdtFV52aRWXdSKd8BCkvilydKE+hkKh+fo
ZpqOwgjuuLm8tN8sEi0GR3aUODBT3y8r1VH6jwbhcG+2nWSuJ0IhU0fnQrjYsETN
tAg8fGZ1OqzDacgfYg0+wdot7y8Fo7wiq8DYggSPNOej4wGo+wXR6qBn+7VSZKNR
G/ES0p5y7VcPdV4GLPek6w==
`protect END_PROTECTED
