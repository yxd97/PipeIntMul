`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pUFHgvoeIuGX+3gQLZAXjWy/UthO1TZ/Q6mKZ2lihSPEAdSHL3maM9Wt21/GWNBB
+0dqtTFidO+gl2aS2jfH9+bQ0GULGSsQ3Ahn/i2WgG1s+LP4/7Wri460x8ZQBG5O
3OAcSujxQ2AcntP/70n9OIw34t8zMZT88EzhbcDanKZMIiJnWDLQzGqHwfMrIdq+
sdSf7EpoZIfGcR9QMxqi50LleatKkhXPlt0d34UE0Ijpnqb5bUtDiSDYGtkAWT2P
B0y9RXN+ON+Zl4pD5fs/9oWmCiKHHDepvoAAPvHw69gPounLG4J6tt9niLNEPEH/
SC50isk/NoqPmValETvVMc3nD5vYKe8sYiReeZkad7Ksg3baSrS6iQ3v5eBab1jB
uD3xvtzDaUPxQD6IcGJmPWLTxmGnh7BiIyDQo3cCtTvpaQzYPGW3zyyv04kX0WC9
h9MQMQX5tLJ6oP/36JzucDsjAUFv5sk0bZnA1ytqjGzEhvz5hpOuRQzvkeDiGYY0
`protect END_PROTECTED
