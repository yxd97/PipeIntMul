`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4emtC/oWE6Oiv68DKu3oSYK7ZwxS91EnOu1IgMpoRQyRuXn4lNpqwOquL6rD9U7V
/OodDh0krva2uec33bbrxJ4WcyLb9VmJXLHamVHjizKPGwH47QjFUi4YhRmq3XHZ
ANdnRqZ4jVOtxbspiD+zfbHBfmoXZ9b7/6gZShrCtAr6r3jXfrc8KNKjsEAieUTR
81iV4C7wWD7VKnKfaCAl3nDMJUDHFQNnXNTk8Ny8fwPl8giMOCLFDLWoFpadsF3B
eMuZq1e267iNrfD7xsJJL85zvn5E1b7gtnaXsUG7UukUie9265pf3zSHLj60g4D3
panRjnlODTwxf9qzg0xu8Zb4YP5IxuX/FkoBIAfFfYwMTO8UFbqLjYSGBUqfCvqG
MRIXSRqQvXfxD/BtQ3tlMbvFeZD6wXu2EJNcZlh/MZRbkAuqXBGZ/1oEfLJVVErS
G3OfGwrZHMZJdL17msECVazY2zEbcQcSLqZ8Ir506Bt9ssTgSVSEevp5w8j8CMw3
`protect END_PROTECTED
