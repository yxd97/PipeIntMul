`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Z8upMKhZms80XPwokYkHsdYcFaQC1ULReco255N+xCREsAU9QOjKDDa7+90oCkm
KO0tDnGVmoasQ5xRr83avQBsj9I2a/6aeuwg0IMXKbMfBLvRlzA3abCszChloDRO
j+JaaxvyoZGM2WcBQNhpXwG7WgBWmSHySpfKpb1VjL+ukx5lnj8mdr3xn6Q/p1wt
0LV2Uy9McW60fsW6Mj/eVhlylcFrUCypD1tzZH9GCV07RKowNxILQJf7CU/x9F7k
3BtObtJxhMM9wgNNgOlU/Ce5/Gnut1x0MN3vYLPCg0Ko7l3HJtCY1nPJxYk8ZW1+
PIbNOx4K7NsM0h08wQNq2tdtWRPQMFj6SaB68M6w2Hg3Rer5FyYkSDupnnL/Jk2G
nDvYmVe+HtAa+A2SeIQKcMPh+oiercqbbpBKmsf0O7oTS7b+WZolM1+/IqaxXz9M
xfeTOuaeX6fLDhN2PJxcjSlT1ZW2XyUnClX9Xo0eGT6+sMsvTW7DYxpLg38hG0lJ
AEd93ePTYefCJTU0cdhE8coaVT03uhgvIEbi4OFzzP0MQIOoA97zJ/sbOxrj1tYA
`protect END_PROTECTED
