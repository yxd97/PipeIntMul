`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFNEv8gEDShg9rQPeH2z6PQfYaEKw46Ok4bXZKalgZwswlHVRQLx7wanjAMIUhv3
yXrGLlMXhbZixwMSZNQYtLvFdsuAYhgOCb6uDkMfenOplqWqdKOpS54xTprALkl1
7OI8zPEbor9tqIhhoMUY4YvghieUBm1kPw0hgGhNhBHXBCdHQbZhNvf8UWLhBRsO
AEF/LWEGBTZd2UPu6d3GGaK83jfB2v9id0bI4Y0GI1trif8jXo5lOFIRjIs09jMY
13Qg6W0r/YdsUazu3/nK0/L4oRx+I9r4ErIhK50DwsS0fIBEYmKivIPMFd7QDurZ
`protect END_PROTECTED
