`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2j7sn2wjdmQu4kXG0gl4tukFmwYp8u/xPz9lZAjA7nbmTPa081RCkAXToIf7Wue3
0xR5DaqJy5213NNOWJAejpIdTU0eu4gU0LWAHGK5l4orrit+yEKcMGNo8mUwVc9z
FhyLM7RwnFuhd9KVJvUguyGEEiIYulF88vvAaELpAJRNIxUju9phgSB8VpqTU6sP
E350+s46xPJoKrHtnC0tQquBGOr1malWHManRtx/jInCcapbGjJwNtJW/6lq1pmH
GajtAs31tclPqLLKLjvykurWwZQw1/xb/DBc3kMHucRhlW+DuqNjBkmmXaeomCAz
rrNsnuMisDHQvZSrZ8MM9MJA5+sWIZw+gpFgzVmNELMW2F8cY2dy6oKyyhZR0klX
mYiBQOHk51YCJ5Xa2Rz5wAfG9YgXWX9x06QbvdNj5xEfqLm2d2cLb2eXPOKb90hF
yQCWjFJPw0tDghkExL7jKqds+TqNahuWFMrHxESXlC1POzywZjjZhSZe1/5KVS2J
JLBzqPmEZCNzHEmzfgEvN1t/yHNuSu/OgUKD995EkyhkRQjWoJJTE7VsMSbTrmEV
JkEKOLTrMzD6Y8G9LbzQKDNiIPO2MoR6i2yMIsubDe7FjSQj2v8bz9HIzRnO4lq7
kpmAMrQ2Jrbmxfw7RXYpgT1HMPEXxUxNSJySYAyGdU837YxGgZ5UbmUk3kpgCyKE
lPnSQF/H27bPkxnoA7m4zaa+dNn3BTfJnkxn8ULUTclQUBinWx752WHH1aJHa49p
DXLcdsauj7Vp+D8hg09tUOK3hhOnRAaQPObjtqqugZhAOBc1nnU5qFCXtgw8Xg0k
v0p15JC/Dz4vs5WbdiGyHbJYVDLlp1BZz0xsboY+RUxP4K2+YvEGEtrxdvufiw1z
1byBjHkchwt7x+f6aRN2ebM707/vhDPPflggeRnHNlpYuzzq77SNaLbJX7MIOGoM
wNJITNPSB8zZADzUAwZESTgUeLG8mJTlZQXnzmPaNWjmrR8PZ98yIEcNgYmjxyMG
7DO0Z5DmHhFPzmyF1nmLUQydckU6QSKK1P3knoDSsdX/FIcgAjgAqvYBQs8S0SW2
hU3wumb4wjCNt0+2UltPkOZQkUcADtXw1rARbRrsCPwmumpNOsqByZsijG5eJlMw
Ci2tn6+Sldn/x04UAW8ZcFtWn4BZObwJqNkTgX6xgwDN0a+77n9Dc/pEhgquYKfc
OCE8Vhc9tP6WN87U48bwqxfdai4KwMQjZvyewf6oPVXkLjUyp4eGU4orCeO7PxSm
IHDpRHOASK1N+gfGyJJt0R03CK1M9ZUbN3Zq9k+BS1y9vx9fzOHgkBjlKvpJoAX2
4YsAhZEgP/D7Egby0wFN7rvvtWuKLe/TkXG+pfXGInHu9oepsoFo2GGYNcMMTSSL
4TR8Kuz3oXdVa2NfqS0yv/NXYweBgN/qHsvOb+0Osu4I8YcJ2oxlRT4j5DUmdfLP
Khm7AAXUaxXG+4MkwRTmP5MU64dxJa3g9I3WtF7wSjm4v0ooNdq2rm+bGez5oBvo
CeDqkpkNq5PCLfKCUbPMv2+1rJosTEiEfR65VlolvLpxqAp2lkEKg0zW6/PXJXZ9
MLQjisRzKtpJRn8G6wcpyGXQp0cy8iQnitnqtNGS8p7bMPcVdegDVH+KUqQ1ljyl
9cqMok8m1ML6xMCFyLX5hTjtUlVREnoSf47qbBTIF2hgjLEhAc5jO9wWUXzvGyf3
hTS5vvsB5D1wFeQtJY0QPB54pqZJuMjcm34jSFlUcFuNOMcfAQa+6hfm9MowUm/u
Us8jVAdrAc+7UtKu4IQ/46NSXwtnoqRBgmbk0qLZuJtcbt5uNB4dFeAhGDCROD16
3tOxnRFtbbu7eXZUiDfVzsRu59USaMvSumvS3StLYroUd8JDSJ5gxpPoS9qqcpmK
DtcWG3LhmOJm9oSBdSlMqS8B7dEIkIfOceAWwHWWUCGMSOoYr1dn6N9kqGSO+DZZ
DE1x5LI+wrZSVKtYg6VNA9m8lp/YVKLu8W39kuXkRk0HPYoIYecC/wJuy6TsdWE5
seDX8O1N/6DcRPpUICXGn1qbNjg+tIKnNvNh84tEcvJV8KxRn3WqouVKfo3UQzKU
J1EVVgKbsNBiVlNagnOPH+38RzZcm3p/ixE/VNTAC7zw5vCsh6sJC2T8oQPASkH5
dlivg3FEpHK2LeIDILV19UfXbNG+ieiWfQ1gaNS26w78ENUzT/Mj0l1al+Cbdg/V
Hh3G5DVAHji7HDRnLdB9DF1BEXl+jDICQsjfRf1GXwIdVZ5wsjFOxUf+rmcVn/LQ
7RyisK9B38iPhVHAU0cjFeTFRSzO0+jzF3qmTL7Cg9KIM80DQ1dKN6rN8cox/IMM
2achjetNFBuQQuZLE5ThK8YkgPi+X8YBXL0/Ouqjla1fUHkCcvBxQ7IxeHIvgP8q
0GopxhyuGRLWe3jFM8El3tkqDXr8QRXEpdiQqEU9X/jEEkQaW3A87rGX1SXn6xs6
fncipZ4rGK1MUKsw1TQFT/TO1MiO5EAMBo8nBuE1OXh/gXelcBDE2XwKLhLKKboD
Ea5Ia6hRe7fUZPEHiQ//R41PIIu8mQFB1ofE4SKbfqCv8Z3/MvsA2SKIqZa2KZNh
5EYnfIl5IbstzJrybDHwAOF3jitP5grhMng6F538QeLh6YRWxwXqASTK+F9NXZYm
xvqJwwAcfmy7Y0JrKioDnr5FyVbh8Vawa37BKVRKOSJHxwkEgCZUxP8NqpVo6fq7
qKfTMczR5ycnKeiN7Xxwl3FL3krEupbtxbadZFDDY5s/nUfemP1E3hQuTduuz50a
1HfrOLw7O/yXNiC6msMODRnulm3l1nimS+OsqA8q91PVmvhRZYlRXiUS2WqB5kWW
9f1cPT8gGWRxBXIgabf/LLXy0O+pY30pbFxBodIqc+VMMI0VlWE8fk/d2zd/WA1j
8IC7XP74YhixB5hIFyQcdSwtJN15e7BdFyfvDod0dYHAeGu01d4YnirObZfj4jDr
k+iXx4IduGN/Q8UrVUqOnQ1rYphU7Vh8T7SiYlV3nVpWR/HIBW4PM2tsidIGw9ks
NZ7j3pXPH5qwc53zwrtzQ/J5n9juChFL7uzq5ekTInzjRYU/EXaRF6+4unxN3ojg
u0E5BlF/N+qh6daBl1oJ63hnJ2YARkU2HtCuF3Zra0tY4feqytxTC4R3g6tIpmVV
j2FnjSv2Qpm74EuFQgkI+w0a0Qd2Ep9eeDaV2lXEqWyd9/0KM81ZVULoMroKGHTL
qFbeS+ufPYLumDl1BCBS/XD7W8ZTmxR4+zo3kD7T7IHOlI7hsO5pIphcTif++vDD
E656s2/5mP9jZrK23sydxqCZN1iMqJVPC1G1NmW0iSwiazwpkJXstTgVTUawy444
C0YFQkDcXui+0BbMzkCWEUZunKOGrcKMsW/KkqYSa4P8boVob80sjRRvBiC5yzH1
fROs90sXKdhVWeFJ8oAS7W34BJ1iAlO5iKbgFPRPIWeABt17DDuI4Kww+7XLasZe
S4wtQ2Nr1Pgaqc0mR70fyZPiyU7YBK+U56buU9YJGNq6zknBpxrPAfgqbSz33mfc
UkIVjoqAHd19016dXSf70YUMd+hpOCK51dQAsKyPeYd24pipddBCnVMX++Mm8QhU
W5EDOeC7yVyk2piqLAM6Hhiim3e0o/yVQHzIEVLS2wt04Vcd5fX9CftkPJJfhOUT
CYH+o/53weneYv5C/7/HEUbRScu66lCCCj+3EYNJ+NI2DXsDGI7eIEVQfcTKcdvV
N3TdUgmY38vF1VE2J9UJ8NaOzgPnPr5ycd5wy8e6N8r9GYWXqf5YTt8EwHfTyKLr
EFmeq5/naOfImiLx9oDpEaiFr2MOPHNXfnaGllHAstYmyQbK0EHpRClZdZq9kN/Z
nfd44QZ2ELeTVxvO11PRVOKWGQ/nRpkGz4PklFtGFR79Wd2UPRaF/uuH7jG8TfD/
5Dmm06nxXuXPs9PDZ8DOhn9XnWyy2r5I17Snad4cpFVZBWV91maSSGpiOnCCTfC1
4kkjpUDmApebSjYBOzqMgFedzeR6+DgtMl0mvqbqL0wVQS54/pMocYvqTOhVVhn1
3+xH8FjHN6/He776dlS49qP3vI/tkwrMovovzJ2bzuAnuxEJvg6NY3GdI18Y7G9s
jRgDV8tgoWnawfseHndXOQlILWOaNQ3+fB91RahRQ2Nao0qpoPDU6ueKbmXrjzLg
oHAU/ppnKDwdc453BuZ4VVpDtgBHn5o/HoHAJnTo6ZVMwTB/ahjXOAXRYxAo+3lY
teTgUluYk3vX1RgofROvcLWXWP1gzqILDBVRxB/oe+1eC05OwHC72u+KtQdQwRDj
lZdJcOeh670tRm2EXqvmPY32yIPvkuzfBTGb1pt1VRe6TSop/ZTYGKuYoL/b8qpF
npqgdWoxCeG3xPmgQ/EwlIj5u1jchV1wOW+L5aMByjSpoe0Uc1z4YDiLtBTaIpuw
LMHGGs4hmNRd12QVVI21yNFLzDEk2tBNjltq4qlFIrLb3QUuaS0v7ZAQie4vbdfr
Km+RtvHkQ34cH35oU5PuG+tPN18ZCB9H8h6GcVTXqI5IbZV46JLtgjysMCFySw9K
jjhy3uM1Gpsgbibn7pzQfAKcr7xwdR83zPFlwMOg36jeq8o1t3UHuuZF3+mngP7R
Feevtc0SDQ5QYPBQkTmQOR/OupVCWfCOroSBsarHs/1m0bqpfpqIKjQHa3HBubmv
oNyfJQecCzYx74/SfwgcUXUubHO8yYnB5JI1QfdJ8bnKoNU10E6xuOwGMkXp7vF6
6CNwcwa1bHakKAQTEZDGSD0ChmkeRfQKvMk/MmQyP4CC916UA4ZKQk6apLuSa7oZ
PlCHeGgc5HGFTxOniAPdGbkU/L3X17QZFssXHGeU7VU4fkdEz9BnUKcfZZPCzqoO
3WeQ66bOm6GDWfEW+1aU8Wmspmy8ovZyMLnITwUnL1OslWYBNY9J12UAMDfXLsE8
1oIA6vG7QOxWfcNSES/AVa4DRP6UQbsydk2UIspZCYe7sjJJMeccLCqzsB6fZClO
lSMD2cS69R9Jx4zMY67TQl9wzdMTdFPB92EHFD8UnV2mee8SNQ8zSHZjDc/Xk8GZ
UJxSUPiqLZTfL7I4cgQ4dPAlU9yqSOhPOdfHdT8ll18kbXHhHCJL0mP1cMHRWszw
ZRwxRqKjaQrHekAPFXRSeseDdU+MvtMxopDcjjYP/GRcOZ5pNFngsctpr29O1Z5m
e/Jzy33gY42fHwIRthWoI5zE7z6nD/OdKM+1tHPoJBzmbWber9ZSAS/1nrmNc6gk
VYZYYAXuK4RWYO2YpLoEp5Ih82QDVpZzRe95qnqMNlW1v9Jc6Mk/ZFSOWeQXOHPy
Xnah5JXmgfRHqWMgRqXukGCkjNeqBrWcfn+SW9TT5WQQubsET4vFl2QGfMnqf+On
EDJJb6qwo4QoGoB1upeW5iCeKplK6Wj6qQpVOJvj/Xm5tBQvwTZ69qwCgmO79KZF
wTZgKZXu5z9UGNabFcX3MG6p7rtzrzms3YVj/LelUfX3vzsxtY31zlKpG0J9DXq8
ks5lHIv+vk3+vP3OIH+XBZ3IEdwfswSdqzYhQLYYNcicXgHIYUD68JKfD6wM2kpF
MOkx9U80IZu+j2sJ0dBdI8/DUkrV3dIkpFCu0cxxr9yiWgAPLPfIGkOsy1KRhfkY
DjtVDbWVEGcnhNIk1sIZCz+u9tQmRAQxJUbZiz9nmVA6/oyS52+nZ/4MYVbf5lHx
HIN8+D4NX8nyLkOm+wC3t2ShQfrW6cNjFpd6dVxsVgIw/9r+pxgMUY1Gsw0oZllK
HXp/rg8WZcrM7h8HMd+VXyC3pI+OZNlaBlpKzZ1YJDsOca23LFDTzz5D+M0rIPAu
db2veNGtasmcIUym+duUrhbUnr24pMBkdByTsx0cTOLHyZ19FX89uFDq5uyw5wMe
F/nM7+hj+ZWXkSr3rMJ1PByUDR1fyQ8IjB8OMnXH3AvCJfhyG2HE3X4fAfb3qRaV
KKHaEu8ZqeYQGHJGw9RW5ZP7MO2Ub4h83IM+MK32BdcBB2jB6tF5RCufxONGRFBs
lvPpBB6eG55qUF4Oy6KjllpWgWTmQnvXrBFgbxf2JWdhBhhdzp6AWABxh7eBFbgk
Ie/5Rux5uHphT1Uixs+XxhtM/31/YKBC1brRwyiz4hgEM3nC9G65NErdnP/30eOT
xHhgm1yxpu/17RUWWqhe/hqEq3Y7KtE0/9f+E4/r7UpY6M0L9XsE+SSZB7hHSJwC
+9yYGQ8VLoNrAXMwNEKpEjVQ+BVn+TXAIMYgfXxkZ/LopSgvfuSbZBxAroixteR/
QP0GF6RfWFruL+OaZ65o6cievM9si5Yr6UoPS1utWcG3ZvtaUGdMzekbjbB8k/A+
/aQmG+floPLgIkOOBv2si11PHyBCjxe+d8d/CS+x9uJkO4LaYuTEJgMWEDH6U+eB
DFk0tVDDVuWdokgnIoV81Lej6LZmU3DLcPmcqwrK9xv/Xg80EQmSAL9ASQOxxgXH
F9j77f13+LfxzWFoi2lGKWE13G3F4hKNeFLJqqO/M/QG48FONT3f4oKdrzX/HNR+
WveLHYlwudxsNjLkYh9N6w9zPZoHzabvvzWKOr5haLnZqyVUmPIU6Be2oxvWTh6W
rIcj4jyoaF4pYQpUiYs7acAZUjSshuP63oTKqiyKXV7VXGaMb4UeQpS0uS5y0OHv
8d1S02ceXDJ6fIIfGsVL9yMzGMMmrXPJ/uqZsfN7GgfCpr3xtPg/O3NOEt0eT3dB
1AbQUaav8u5D4vhOL7eoeMruAnuPkRUEEKDSuWetGuIas/WHK+A8M1AKmPEFAUb2
oykwGnjTIHPAf46UUhTNotzzf7a6Rj7X6n8XOpQIkU9ot6etVfxiovZTztQAdWcG
lCTOIM/pZzI2TOvnBchw/ux7qFMkVbPCM5DAZbaSDNH8XR4l4i12Hj6GQ0rv3Gns
tFgF0YQcCWWEQGrDrf10SDBr2MR1iFSFC1c3dQYy0G4u0QxZa0rba7R6HMxdJSPF
6Mu0E4rAPLapZIaXTCQVVeB2bCTbTvkYwU3ZuEZCtBYIu/FUAyiSW3TtKtFoHxF2
2TqXxfVfZgwIZrxNmHcAgaE3fSx/xUQjsv3eKs1XUnGwdudSnaQ4Lh0KmCgKMat4
DizcEThT3/hnYk8BcGNPs8vnF1A/Tt179dqFyLMafYmL7gE5k6VFPbErpk0aUOPV
1noO2LtsOgUCToY8jU/5kqFcaVwcBYFHJxnaV/Eghzkm+lD7zY5X0wWCw8ZqcV6Z
Z0bFSBilrUvc8Jf3uZho2bF6HJbhd/kU0qpFzNd1WQ/DG7iX2aRgeFunUxHj9mBf
sBYTeavK9lCEOFw6NUU/YHNo+iACUwmhHwsJelIrDh7YNMv/QhAOEiVlUyjHuF+j
mNjwoT6Paun+1VVUV+D0Ftabzx5QmM/n4HAwE2yOKVWgxF939GZ0v093pX0TU0Ko
BwmnaScX9dCjwJ9Py/ZJYzV59WrjTLp1pYvZHAtM/wi+rFKCb3JPTf50yTJTjwMa
E4r7lXvcdqsbkClhwCywygqQ5AWrzjFd1k38L85h/BWF/EKOm8OCxsyU5aWGJNdH
9c5tt9oNlXssjbjhKZ1Lec7pKVpDLH7f9KZ2TMqFR/f9+Xou3hs7DURxYLQGGjS/
alB0XvJcs+nAYUdWa7AbLWlx9CSbKOOHc0yMDbQ7KD+vxOON8Yabt089PSycpqar
tc0Jrj7mcl5bZQQc4zfLRP3dSW9h6LZbyLhyGHHCBywgNk4/rWhphlTYqwybDNh8
6j5Yt5cf2oTVYFOphHAfA35VPR8d4qP7msnzJ0gDb5r7V+4igD4VlGe0D8OPypjy
rkn+jIqNocYyHalhg+JC1QhsLJLGV+tR1CMyMb29nbl3rKyqxrnD8vstb5e0j/am
PlOpgMWM6IfaKfwx0VIgwfjNEWaO3GpGBM6ryvb9N0pp0GOLib9UDoKx0F/U/vvo
FmnnJ7vbiZp24mbrwLwdfrElluQk1SO4X4IPTasibQk8zz1ILeWDOLktwfCd6797
G+Sv+A0mpzVH3a4bvCTjYUVdnabk2U9gBHg5AQaV+RoPiQSEXQ0XZw6kaTWkKtzF
aLcsQZ0RqJ0fS16UI0N7flgRKvSKuOWFa2lp1zkhq5jEifdmFvBsL/FvInZ/Uto1
dGsXdEabgc+oUGinUx3NvLhnq022LccRHqvIftfigCU4FuY5xSBz27gh8b3vbHp+
fN1X/uoMFE0x3I7iTOS7mfnDW1SP0qXGnbwl1i3G9OjeSLU4ScHICR6jJFqMUE2e
nBMToWXKossra6i7W0jwcP9EyNr748vNjr1ktMmLIVevR09Pwi4fBhcAOg/oBng1
bwMm/hSHQGQX66i1MKuq4cFUQZRtyoBRcwh6VcWN7gqFexuyE//LF9k/DKof9RxK
CVdPnKWoeSo53M1SkhpwegL0+4DAii5sa2r5k6Key2NckHKxOoEn4m/AlXTrjMat
6PDG0tBQr2jgHXFaFXAFLMxqcDmrAWqRVX8L5VR3PRH1WZDxF6/qjn8qz3ipoH1W
dRxkWSo5Cun2Ijqh8ddL4nWjqqanY8KkG0aWPxF2dPMF/OWXfRLChqk6vNT7cLma
TyVWQQl0Yx2QPAwO5kc3slX6cxyOJ7nGRYx43DWFvxaWJUGHuU48vvlazfQVov+M
f57nC/5A0jEDoeiF2aI1eyC2qb8uhVvKIXNxa7sSXos4LsdwgBSSE48AOjHpnF/M
dPb9XFn8VdUQRNlgQliMlTCh1DHZ/Kdi7NTAS2hhbnD0EiEVbeNLHfv83TV5402f
xHpYgprD1kdG3o2tfN6eWAu84cKPMksON0LEtGvTSQMoU8YIEUw0p5HADs6QFmwt
ZEUy6WFP7GvT992Ty51Bpwae5qHTCVKlOPKfNoL9GgL8rdLYCx6u43+taFA1XDnZ
MRaUml3eIef09FaJS5y6pEXT6HY7/xwAEOWPW1cbM3gvBqVbNt6SqlHgPM0Hn7Xu
4/4f3/qXEA7LzOUuwqFceZJUhM0o+/Iael3aZ3Zh65G4uuU3aLaUdovoizDfyOaN
d1Hce1nh1gkFud8p+BkEFpZL12o3NsSNpuF0GlRFU8BLtCRBIhYTNc7HRu/IHHfq
67TtxzcnFXkxLUuVlKYAGUUKxLmR40t4z+RVDN3ya0wv0ktu+KhrhVmTPqNiS/U8
EPRyAGQ5N8wredWxQs2r5y69Ybg9NzyD9DfWrpyZsz4j+x4aiufPxSdJrdTRjN6r
t/KOwmmpMlAXFgk1GUjiXo1ZzNcEqjghL1qgrQySo3hle0tW/6Ebrr9DH5q9gvuK
YxaNM3PdMZ8/+CVKjWZfew37VNKUcExM41MEeTanYaZMBDAlXv3YPkvQMMk9djNR
0ZFtdAAQHRTRaFtn4MnDXoIbH6ENxVNAeU8OTPsWCrbdpgRznYv4BCePqbgPqpvD
OdPHpDlMf11kxRr+pqqVTBfKqLO60JIFxkwq9mbmOUbRpCsYw/5tVfg3/rKgr/A2
zQyOfgQjhUIDLk20i7YBGpg5dByb/D+DA1kHjdcfQsOZmW8iehAk8/hcoe9oZgC1
Uqnqdu/+TVXpYCeHQOUVj8ZJYEghdiA1Gd1wjbn1WaUx9nyWXZWmmZQwSWuAiB67
bUII154CyPTNebNzP4zeZeFP32ZqkoXdQnLgB7y2YGQaS7xz7+xXAnel3167y3lB
qwXR/R98mGhQPixyWBAS+1QnH/kHnCOPK9udl3VfkZ0/4wHPEXs2WxXkgTHVJTWP
KFkH9bTMCYNkYhIwOUtWvtwtxN6uXy/QkkPnMBoP5hgo4PfM6DGqYP/P36NpYgzu
aEXfNrLh2UignE4eC78j3WVSHTzjb0rW2r/5752t8L0I9ed0LGITnZuR449vihe5
Sc6CkQp5FA89zMHD0bjpMjzrsk09JsasSNMtV9AsvqlRL90KQu+8EHxCVYUgddG9
N6/MVAbeuBoRdaxAO6KNwfSbMMmV7YIReU+eIURcyCrMBU3BM9mLAAxAlFxLE/jk
5rjgFvV0vhfJ9/sT5vGjmtY2vqi7myB6kvfzB+gK9kVpMI/wP9K4Ai+wFtcorfxW
j7Ot7jo9Z/46YNVp1CBxOhdQW4Gq328SZJK2fI4BOkDuSh3kVQrsGfoq9f2MwIen
iOYUua3huDuaERz5FFPxxlAr1UOZtogopG7XTZrp3B+zBBZ9q1hC2c2onIhIBk0E
N0itkSOZ87OUyFjFSUmkvaSfbzVNe52HyEBApNybo36pmEC+IqWSc58N5DsOs12b
u3L+eQMr7U/ZcrLHvjjs/xS8JpwQ+4OMTrwA70y9B/Udy6lVgEptv9pTLDQNF+sg
KeMHgJ2k3nVzN/i50+pqueGR+voa3sJ9Sg3RrOwv3NalQsQ8gor2/n1LzFr9pJ4l
eEKY8q8cYY2V8JXVYTIzDqYtNtdS9jLGEk/mWFyrftRsZKitQwG57jLR5URvb7tI
xP3XtHzFnFmCop1McElB+dPm4+46vdKyxGSA8H1s+vevynMR+V0yC3Bp9vGjwEBM
70j5fVXMvfoTAwbqT6OqPSCCL6xzHhonzcqMidou5fMYVrmyk9hqrq+vIZcZmpD0
enndergS2a+Q4ZJkLPNFCpchvGam9ojP5VQzlDKgG3lhDYNO9W+gfpGIlH5E9lQd
hME1YMEDEIUK1i53dNGA5r3BCmohkUvE1AEphw4rVJ1Itx+hGFf8ZjqWghOeP1tA
DvcN8I7iUtyVkLX/pMLwnWA+Z5w1EMx0rROvJxBBCbrmeZBCnPJbScXOQBFSFtNx
WyxoZRKxV53zzl7+GtbFfe4d7Wo+rM2IqF+tS7af5hTrKvZu47DT2B29F9Dl8VEQ
x214HdGvb83nVQepDhafwtfICm0s/ZgfNaVagBZRG1fqsEkVTW4uIKIobfcybFWZ
ymBIcz4lKzj7pENMaFZLzWY3RI6W/z7bFmmlIOYUaFzH2IwzmHVWhdRF4tfI/mv4
h27KNzUeUm3V6AodInQD0owcCjT+elOiGV10YAwtfZSBzT6ZMhQOECftGJbabcjx
ybKLUObT2yxpoToX4fPVnRA8RZSNcxrIt2WDYn9PWDDPtHhBma/RzZx19AKInfh8
b3dELqmaXBbU2aNv5bLvlyekWRHmMM9nQIehDUZLjOWrUXBRlXxCUylivWX/RJd/
5kSSo3jctGD+SMJoQuoe6NMCNG6eoj3lxAF9yVqIoNUSN1MUkpdylLML6ROh4VAg
LdUI/AZiYJ2RbEZ/qnHA2PJYBiRIMManuIqOw5YHjWdqr2MLGuDx/ko6YRsgu5wN
i/mlz9SQxnL6Chu/xg14+afGJJCnXxNDUKbAopDeTbEoZdFr6T4qwsXptxngHNgy
DFogOgjFFejqo+W6/WqJI+tcXUm+F6pHkdvw7S2aqDOdN2/JyOLwmcTDafX8wix1
NeARsomSIvGIIGxMWncxFIWTlVcR3Bi6YLm1vRgo/3KdJnyO4Du3ohHYBuvChrww
hEOGnnN2wHvVcv541gQVAtD1iMhTgi64ewGxB1qBLff49iiORjRW3Vv7qXl6QTvL
gf+lPVd8B5lhSiHlozV3+dixU95fh3rd1AyYjW2lRzQ6/iP/W82W97QY8D3IW6Mm
V3axJiSPJuGGTTKJl+vMI8Q7sLr/u1DHmTL97uX9BWmb6Lrs09dNWYdEXH7ep5Z+
96mO9o1hecncJ/Xjvbzk6ey40Dg27PCokNTzdNppWXH2CLEMltm7JJjI+k106kDT
isxkjfyXEZX/W2UGkc68BMY/KnZ12CwbjDRNu3wzFgBglZF7TJRyYNHKayTy7AQk
vsigTODjzovuc/L9CEXHq9sqC2k9+CB1+OpKJ6hdO+JZIXI5wMPN5EoVMH3BlCtg
ZW0o89IgSdGJ9d6et7pMHCa7B7nMN5XSKfKMWcnSV9ypDnKc7jdRKtIBDctXKG3C
F/4dikbdjJj+z0voJ6bmR4V1B4oiHjH/ewQxnkuP01bDsQeb+rcZYFbpkKMBuAhS
S6+IZ/PwzxZ6hsHwQvd+B+u/J2PxCRE8svA6kxPt2tBOVrLommzCBsEdtBLhkjE5
UKFzRBvc5Rg/EbUAnDgRBpOuwcUivu6AnWqkNbb/7GcaN8GYHicfLyHDB5HIEoGU
ygIwt+dkCQOTMVTcS8ZwFusd7Gp4oUf0t65u/eJ45rIqO8ub9EW2N5oOhgDEqhxz
7ACk5DdXqrqbW64bYizcqCvG7fsId0o/MhzCs5eP4c3k8EDzvbUzXL+XQ3iFk5v1
Py+tp1RQROHCGD3y6iFRqxi8qRQIoTrKPrf9X4weUwGf3N5NNKRq7UMhuYUZZs76
iCt6njaisjEv7droD/vAqta+m39J2Y0BtmOSsmOqRCkT27Q7PTYFFshHtEWTOUh7
Dhyy1uLVGZDr1fj9EQ19JucVR75KjDvSD20h+OV/rVwni5lugYGiT1c026jIVjt2
P/JL9q07O6nf2epBiBzFAZGMNbP3yiDPnJLuodTmUPCQdheC2Y/YqGC8gC51rFUa
ARhjfneNUz3X/mSaLGWu9LCB+z6iCLxrgBtUHGai7UcCIDlUdZYb8Ujc1Z9YymU+
d82dOAxNyF1x1kclMRHdSLc29tGX2DD8f7F36L4P4OiwBqWkt5yz6hQ/x/gVc3Ig
syLsQRMZmQTOIX99FdwbX2TcqQDUGw6ecNvioOKrtJEoXkaHdCjzjZtxGaMnJpoP
oLTv5gpMYVYt5TqHCO+QsAfQV66oUg3j5WLbejIVRtbhs6Z8yQzD0ilMG3pw02k5
xiJg/Ir12v9k2yQqWsbpVUhZxTxsdXoAlX36vy6ZR5vlF6SdtQ7LjtxH72ZHTBTA
L5ZtFeylJDHa/LTID7nxgY7zyQ26I+qS7Xahxlb6ofWxQaeBpq6l6juPMy5+O7k3
dsG/3tuECz3IdhmmYiBqo96HlgQ3naHoV94aHh7N47oG/RW26XTsOILsM9ib0lgN
Ltb2kS/PWPqeS+FAM/Li6XoJ3uS2FRvJYpkV53JtkhM0GqwN3Oatvf984IOH7S+n
gflasuLjSBVMWKGa+hNQvyTQVXjVdG+C9CtmlLS6JrZYuRQtC/GhdhghG3f8/S6q
2SV8BcyHFsuq0+RQ2wcmS1kN5lvpdCH6AG4VjexXXTZWelfiXEsdSNB1uxInGB2o
jaHflQUd5vtLhJdAvjIUcnusTFJS93E1Olp/PapherhDOtbpqaUwYh050u9iHs1o
SnVxPgl6GKN6xYbFsxeRKRQ/tAdK8ji2CwVATbSAJ/L0DxkQ92GacY782BOhF0ck
s5dpU4Hr79nNDuT61EoyVVaiTpAh6/hNYm679aRI/zA1utQ7RmQibsRu+Kz6Puu7
T08Y7RihcKP11/zcYgDr2p1IswuyU0WR4UV+LeFdGcWmc7NslMhUg2UkXwYQccjF
bmo4yhfU28HFEyYjlz5Fj2CslflSoT7uXJ89u6D493SreU9qOre+IrMzxdiPZ54m
uEzt6DMx0h14SKawadyeWQxqeS9e0komLH5FDbPlCrWAO26C7/d1mh4+AsFSoyyZ
PBfDjjlbqZVJZ7YGCzIET8+dKLjvUKT6M+uKyXP7oH8CL9NzKZ7IU/bc+ttrxp4P
F/S0bI/weTikmF8rVsnYsmDFFcrJNbhZNDMYDYXr+gypUvmM9ggLH0sW7hZhs8ct
+QWjfFB/o5Z6qaH/i5ouKBDGOwKProvgVcKywTV1m6sY2WffS/VYnc5n1tGinDyE
3FVZqQSDLO9yNq/oYHXueJG//ab3BZX5vVZRoK2rK3N7kklAuHfSEleYxPxk1zQX
UyxXsCMQh1sSbUAEmHAwSvS28CWCL3pKlxAhF80sP7RQqk/2KXhOOYmgkE7KCLP0
Q9MF2vwg9nezmbt/pu1gVdbbP+UbbhiUMuTzJj+ouoTVdEqKGONyC9rwnFaGj50u
w96fluRBrBa9TAj404y1lrl77MqAnPS6rn5G03910/B00Gzbp3qYP9oQE/ZYK8yb
PQG5o+Ljbxx7v8p2os2cdhDO6HszNHQ/lhKQNjBjfE9gfBmG5w9RsdVQP/M1Iovu
WLYLs6Hx3/GqihtVlaVz2x4PUwfz32Uo1kNKD8leMOZHsfqSEJO8oUQUViRFrVzH
el/nUmpu4vDeK1lC43EDz6ofqIERdnwtdIcCDrjQMYSjb1Ba+D8UYZoD750wVq8h
jQ1vRhvYp6z8IxYXzelbebNPyPJgbrVTDF1N/ja5bNZMG78pdMC+6mkZH1hVJDw+
vVG2hp2YsFlHQYidam/FsxhOmXdnoIXJNJ6tIKiZ+eKDmftpLrORD5rsoSSFugg+
JFJhc89y1TAYDgqTv0SFLwXUp43fURK1LDyecvQ77rENggaYimO2fY/FiKEy8Pf3
X81AQW00ltTfyCs1yW5SZyRGlXVLJ49cX01Q9gJ+kgLU5LPw7d7XwzrjbanGFDlM
Ni5IOCLB/HZjpRjITpiNS2Zau7CrfP6eiYznw1UNinqzuHqdnl6/73NVlx2985eP
g1wtXD3nbKF5JgtjO/xGFworO8hzGP4kiFEibVaGb8GFw37e97Vz/xcZHhY0LPgo
MSLxF7a0c011LqLosj1Yb1H8knB6RGAU0jE9JxheHn7SiMlinZEbFa/ku0D2r9nd
FTd0IYlOt0Kw8Gj/Qv4ZBj03Bsfvd5tVTACRTsCuOSPrp9hgeVZAOE5Ei2jSpjXk
80syPe37C5klPTtlAo40l9GOinoQRPSZoo+vDVTYPJbK5wIz3koKA9WLw9ctdRLQ
33ui7BkAjFqlBnoGzjJ0orLa28uTSfeOTuVT1dHaYWuEXbR9Z3sYG+NgRPxtw81k
2G88WlWnNTQJt2Kr47JLCmTeaBXnr0f8/4k3Jtix5ML22aYQ7tTQhbYfSPGhwp5s
R4b8PSXg6SySdZLYhSMclepUdK0gJIh3D3HExqx3R+ZUG6plerMAccqtQYuMMF0t
XxmNDg6OPxTfA51ENu3zO4+HSNe5NG56AlEcWMb1xykIwcK1C280RpSPk0IWracc
N9+UEZ/1GsPP1Dly1s5WdvqWOM3Z0BNjQdpxkEgSzZ/+FIYI7jq8j7or1roEtJEq
zt2e0k1ofUw9y0qEXU0vt6XR3mwn1PC52MrL4BV5a1xPQBRG/oBMGLIuZZ/TwuEr
9PBLw8AGtFKMmiNY4CeCQwJsVCGeZqZnDj6wpZ82GNBLHe7bDqoPheTJOWcimfla
jP1IOWykBIirPoGCVBowNziJ7mmf9Bxf+eBjuIlFUsMGtL77+5+ylIVH9OkEdbjg
hDx42JSQ2RnyxAtvmc69BP1NKbm4QEpY44wXMDM7HdwM1uryqeQWkAvGovrIdc2X
IqFYJnUPK0TaWlkL6ejctGJ15Fem2jo5b1Pn0yeO09atVz0A8vSUTXBB7Lxt8JPD
L1OMgiza7UoYsvXGey9gN4e89JnMHh0IrjQdotA9rtmecfgQqZGm8iaWNarsbTk+
NiPL6+FwWKSHu8RdfXAr2ULhr8Gxo06wJbjWA7IzHFW2cbvM8UJaJB5T6df02Nzk
wj4E7CZIID044Z36WB809whxqFnaufEp0iGwkV//3rZ8XWIoDANc4aokFyP34kb1
KzSbupW3LpLYHR8t+0WeN7avp1RFllWgjOsKw2HYoWhSZ4WFszKI6SMENPiIPcw5
cikm9y37NORF+tqyUX8eT84+wFn6JW0GPoP5xhLeaoRvBOWCvEsnrfwJeFkEal4D
kTDoMjC6XcIYbJ5YCzS/G9umOF9KUBWxNn9sUPIiI88MWPx/NeCoOczYzOO4ziPu
yh7qN2X0BHjd9hAN714B9d2tm+L9zKSxJ8aOd9qvpNmkKLyKXnxrpJmtDs+X1YyI
FYhveJYUc3a/KmiUQgzaQNKeOrIdnOM8JQqJzMsjd3Ma6WhsZmND23ZAIDIVwseb
T9L8LSh4VRqdwRgiTgULZA==
`protect END_PROTECTED
