`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/0vl9PAz5MjHNK0pq7ku4qNtifVfqHy4DIBE2pSoLk4JO4Gk2xba/l8AGOczYow
2z60BJlPMF1jcXzdwXGHSHaz4OOTuD3qs9Ao7+lx1AlHjgYJGfRBOeV21taRY6Sa
vyZf7pjC0cGA1Vi7Jm75duT1bQFPJ5Vr588NeaG77CCaXzBX4RCLfgYGBAt1z/wV
kGIBmntW0u/SQX8AeMye10x9e98Po1NbmeeL3Mpzxw5qz28/BMGTsnrSxZ8IdS38
2LaSg2Pa7/F/sQTx5jswyhiKeGAhdOdMU5vsvvKLjwR86Hpz+7zqldGYG42b8f6y
MMDSZ7ERuJa+aN7teXxv1YR+dir1ivJ7j3+o6hXhluW1nA1lwfW3xXaR3bIvNzhL
UVIuuHEinUga+ekhv8Vlwt4y1lNOvFMOwcOr7Nfnwnzwa/vR7Z8u6TyQvxFpsfWc
JgZU7xqPqU/L941RHKfHlYpYhgLEihRZajoknA9E42Y=
`protect END_PROTECTED
