`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6nAz70YwVn2s02OZR4UA8t8rYFcLPppplJHyk0XWPLHE8r0xH5PoLcNwBwbwq/s
5dF+8A7fcmviGMv/QukS+MUWIUCqJpfVaBggqQ/e4/Z7+JlagMOgjvQBfhNICDVG
Ht5HfjK6Zp4J4v+0F6CpQrEpAqKmLcN5VHd8fovp8uMyCSxdbcCoDWFZ6JGx+BLi
QeK3Ji8igy7H/xYvncbGVKC4UAqCwOievOAbI7g6Fj4cwpICuMNoJ0SCmcjiDl+K
ZuoufvTSzuok9Ilf6hGAkkVLmPsd/sO7kevMhUX+JUODA6ijelww4QK2E+ieYf+j
j1AZNzvrB6I58mkdTNNOu1tbxDz8o1RZvFiKWKRU78rm4NrgWOv8+kyZ013rYJJb
dw+VXx/260qyA1GRTyjAobN/5QgCgVvOFpj/gCDHCIKz6CwaraTmjF++vWEjXi2G
sm1s5kqCyovJfr4SwE3TnPyvB6KQrswoBmYeYAo5hiA1jd9nATSqm4fJ/lZiiWYr
+g8Rlk2XsiamAPXZlSF29EqOMAZePTBawRqXQzO/BMIuu8LVy/mOxrJpm/QyIZvg
78vewldjAhaho6MBnt0UXJQhBSxM3T/OJITEWI+bPkhOzrgnAhIYeR1TIXc8xgT/
feYzbS8kMfrZ2BIcbcEWWDsBGW82OXQeVxzooUGXOHmWXL1TGaZav/iVgkep5hME
M3doQZExMSBluB4Gxpm9gadG1n8niAEg+ov/CfGH++CNIh8K4+SZT/BpfTJHNPpA
z9KDg8lm4qXokxrER/NeG9l5jceaod5l4tA/b/Qq6qw3e84HvASlzXTdZ9U+u/us
WaQJ7+cK3NaZkBuEnpGxWyoWuS6JQySHexDvXQBbfF/V4KcFF4RtLPK2lJiGVvlS
SyZJzYXpoKCU4iGkcAAsWykPT+4xsdq5iK7jd8bnF8U1hS+WlhiJ0qDRA5qymnRq
ssT1LQRK+wm72c6aEXtx4ogGj406P/K6AJ+L0bKOKUfTq3RHa8+siM7C0RxDxcrc
T5KdUhwzGTMDmmO+t960Ub3nLuZd+k0j6HRgS1z7zMyoti6bnKFNVL0iv8Vj8sxU
qFla1E5i4QbO2B9YQxp3fdWtMJS4JXz/Y8tADCIyHTQAfZoGsRKfTTEVfJgvSJpP
ZKSzUKTVo4PKswXDZI32eYqcYxWN00+i2/Kg4y0rPlMH+Azm9JQNMpsfvOSoZKR2
TwysYkXi6wH5uxhLrk7KvB4SZvnMrMMiotKz7tx5vzR65jPHBi/Zc34P+q70OOIk
HQiJPK7N+ZD4hWlDkeKTp9Ze1WY/HSaFQFdZb3TW1SvWlXbV3d8d0p0LBEoDkZUY
sUOFcyQEs/XD8/v/tgGYKuKYPUEBsh7I2gSpbFe1QXEGYKW/F5mroWbBopc6/4rT
ExYtcbWPaijL1UkRz3GqQ2xDC1Zb6nC2pgV0MedIMdie2pohaaH/K6XTWPDxyLQo
pisRk00+8zSd3QZ8/6ABxTSbntlGCQ9SETgl0crBy5QosAL1vk3EiZ7KbKJ9nuHp
2zsAz3WIN4CeqC+dTCHk3uhw1HR1FJtHa0/g0Qc1mltA4hyHZtyD9Y0xLet2eM/N
5X9Q4f+duRQYNc+otw4VxioLFldrn5lgfH9HgHrtSLkY+NKXI2MGDPDRz6oSdizC
DhYzXH6r+VmwE4sZEQF25fJmZlhFmwOfZ8mEGv+cGrpeZzvkeell17MHC8WLWC6A
DP9K7oukIl9q0q8dqpYqCg==
`protect END_PROTECTED
