`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swoaqcT1YK6dB6P/hyVWoHu049zC7tGhDwPwdwJW82WQZQGzGvK5g6r90VHUPCDK
m1A3YiiKOf1VJExdAFrmESWMJYQ4DAMH8eXZuHxgExvD7A/T4PjbUaBqgi+5WILg
aJ6Du3VyW/raZah8b8GJE0no73gbLCaWyWmxhp4yIUEt+OYenUgXE3asrDxH89W/
dep3V+XYTAP3l9Ul4z9vp6V+4f0aEWuF9EypWLnGLZI7oORCVCNR+KpS5pvSr4rO
1ixYpmcCbk8Gvng36WpOTkZhK2i4nF/evL853t6WBZ3+7pKqt5JDuBBFbPF2f19D
Uj5krJUA/pqxAiooMjSMPD50GWh5l25IGKWxOL9hbJAgMqUtg7slQgRFsw1/LtGt
c9QTUM8LYPxC/FZ8Kp/rCFg7Ze7x757Ro+IKVlbi1WI9RzRwpWDU2I9OJZvWGCWa
KF+0+hyuZpyBn7BxcA83HpS//XwRXOrrk0Z58M8C3iG9YmuUOxGQvlWGQJrdBHu+
+VqE72LcdfGWlRMMndGjLyR8896UiIEyxtis0eNdb1XQRd8FkHa38zhBu4g0uOxw
`protect END_PROTECTED
