`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6S3gZ2UK3Cy3myvDhd5L0UytbHbXhZv6JIR04WMtz+FkKNv5JD811FzSaI4fkQvL
opEyr4YTsw0p2ePtZj4XZgCAMwL0b7g4rvBE6mAC/LX5m28kkukP4Ksqo1b4JF5g
tNuZj9SBM7bvRgSHWU56mGLfcMcW2NzLeZ65xaVLjBR47tzwvu5hNSGLgwHZbMOi
sU8yPl6ye4KMSpjWbQdsaL+FbaG+PedFVMdFnXSUeqErQdqKK1e3qgzN4jD1sbZm
LrY/DzD4X76rqdRRcDvgUkbPNXDWn0rJ0y4UXd4hi1544u+gJbaLRTVlEOrP5FDZ
HrLNMXcbeYeajOGIyIxjNQ==
`protect END_PROTECTED
