`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhqj5Jf4v401PsU1rR3rkk8ZpxRamDWmiDvOKCrAM8OeWUnDtpRUsdXc2+xhnh9T
IOZYai06WsXMsz9br6eOtg/gM5L8DkISuulYWI961fHncFyOhByCX0msZYNRTg0t
Nw7pzh+f0vjIKwo3YhKYVUrFpCAr0i1zx8pISX3DNaN/if1Y0ackQh2GAGJiVJYe
MLhUmvvqc7WytJcHaSEmB5Ccn8UYdiDpqa3XALLhd8OL9TuYLKHDp5F2gyJ5VTol
MKcYBUwHG4zoxbZTaRSs155MuU/QdedTkrY3hwsGOAMdV81n5RZ+zVb1OvVKfKgy
4M9pWq7cjRtH9XdWuBeMua8TnbZt30++zXvmDMY2oigP8JrJDJAoYgDsTV/cNSD7
Oancsq9KnZ3DrlvebdfdGsst6upUDDFIfOwRo4GAOJVzjRG6dGCe+wnN/6sopHYJ
LKPfRsOS7CFkL3hacrJVXSgl+3heb+fOTPetsFFJDNqQph45p48QfD5JgSt+blNm
naxpokrg/PA9Nwvkr5xxLoTo8AOPJ/7J14d3Cw4hVLVaWgH2vMSBcXWc2pxaKR35
wc/RnOgQ4y7qcraRoTZuwUmGyqw8Q4mxUj3Tt2DjenDVxkgnZlVymyAqFRTGobyN
3ZCh5mivBZ7Obf4Ae4QQpMfvWZ6aQEFbXuCjzhj5ZmXnrQ1ujf+6UVhhdM0aYjxc
b682Kdaj0AlMYRI6NLMar3EChULOs4OOPVyX5nIK2BPOX8BIGuwYJ3LG8tQxZg4S
+5tenEowxFmtLR7w/kM9vj0od446DZk0zD+SVSCT/MnHnBZV6DzPyyCXTmk6zTJM
OEUMe8Ra0ijhlMclAODOpHzZoek5empE3yo91Z+1exUmFfgDKjdpzdYixGl2Xb+4
zsZxAD0Hq80m9QlzXjoILZLAsSMPbQFm/mETBUbvsj+3MHpc5S6VgfPRoSfLxrwk
3TwAT11uYTTpqfF4V6evX3euCRlK1YLJATIgXyoCq3JxDY5QbDL2N3x8A8mQhbP8
eFX7vFktwzQ+4EVEYWjNW8YRPvXwefhdeq5eCJ5MrwUk3ay/pPW0sD2chbL1/eTF
OlVIkrufZePauJB7XaKM0Eg9hJOxiFWHGjn8zgVEccAavk5hvDwY2vROu/agTUZG
dY/th278IVYVgLxXFyIvS+OV3D751JvHBJ0CyYB7DJcXurSbfC18Ks31fuK/YEpD
qpFg0s7/oEvue1rkP8wxiOuOyodYX9JL57W/5fixNvoLl/+fGdZlGdKftMWRCeyT
+2Ev9iAPMvoJzv4znJMBhP7JYMaMio8mC4mIrI7ddxv9wS8Pmip3fV5AuNzAP3dS
Q18KfE3fBmpMppSMoDESSK7Bd/3h10NKWieT0k3bwYj2ZwDNbKNlVs2pl0PAAITX
qhsbPGoR27UaSp9rFFoPTrDkx6aYQw1mZLF9F7QLO6X9H6+yvvi/OYRLzsV4tRSv
kUOrVjeP4tGp9n7VQZDxa6B10EpqF6kzO4TQMXDf4NgQODhcrmh7pNzlXQp78fAx
Oe8B/hrDTzkz0Lq6kDSq3rKheDqpkOHLnDnOKzr4pHcSmK1gdkxPBFEKJrj8JpZN
gAK31vZxyf90DCidlxl2RSCjTthHm6nYGYNtv0skDrRc/qEIi9rjdp34rLXog+ae
IwxW0KNb2cDtJZK8UrnN0r/M/rVvuLg+3APqLgO44AfBNTTvPt5yavq3tx2T64sO
XQ+5yIlgcUFwqg6J2pwn3Y1sAk7mOccDOnN2RSNzdYKpp3PCVRCsCRiWB353EcwY
yGEEzKM45y7U9kcP1qXNSCDnTNeRENdMteJ0sVqazUlbIjnJ1kHOhM2j+7gnhnoT
KMoTuzR9ntRN2LOEseU6NAP4hiyhC1QYyCJ7lO0FH2TUEvTkUSzYRxkYKiir8t3W
R5Ot4K32+d0dp0x8+n+T+7dgERSSrgUqR697b6FNbw71msq3kkGcP1Zvh+wozlBH
G8zJb8kFeVlNE3yz62lFo1K5vbeWWoola49imOSOGyo5iNpXzDfYv7LVQWx8Be5z
L5FC2poMtEibvlxLmFVwbEG+xzKoydqBMTHFNGkhdjI=
`protect END_PROTECTED
