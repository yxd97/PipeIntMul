`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ow2E4SndzaTDoFeokR8bSLr7ljYczoQBBq74gpnQuPrXlur/ZkB1E7+JiYwOaRBc
+G12iwp7aLeVyaVzL3xjyt9GAoAshXs0wBU1hXX5nqGn7lB4saAQ3M8vWVhQGSdd
OCVTgwbXB9+I2L8MXgTu9iAkAm8V1UvDMM+HY/supIuBDc5qohxuNrEDqyM1qiN0
FK81Omb9IPYs22lWRyDh9T5Op8gFmTinkPM0MkaurT0I2ofZsUs9DHg89QWzQcHI
K8uyTYpfvxe+I6ZXynsKVYvWZEOLN90S8CZ4IaS/Nanclaxgp+J+CjAOIqMe/xmt
Jmr83kqKezVowNJ7tTUS2itN0pmZlqpcOGwvDdWl997LtaA2M9HR+SdAWcq9w7TF
/pnamKyQYoIVDEPuMQZ7UblE9Pl2KngejrRQfoyzHEI=
`protect END_PROTECTED
