`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ynX3le/r8QElTCyS+c8X6Vyy1/tmRvRSe3+cWFO54zLKniQ/um4f7FQwEySWvyPd
3DnilEF9Te4jMxEfQaZoj91UqrerkTo4iNFUQkLLrsmm5Y7s9GLs83imTymB5mhz
0HTmCkc4O4bsl6KmBe2JoZKSedXa72hxAFqHPBKsr7IRrr4F8drsHnhgtADn78+O
GESgAlhKw9cB5JHsPvC5pZbD7R+Clqk17ycodl3fwA/5R/cghjjEidAHQFphL0lC
QlxRaMkRYHvbTflJA5aMM+42X5r5TfdhNRardvvYxoiqiBsA3GGOM3FKTzjWAC01
EGbMFAOOt1AJK/SNt0cBC3Pig9dorMXhnKMsymWghxwbNpuvssU2jbS/IirQ08Ua
KwAOMdTdBy49NAN0OWEJU6CoCqlA+w1Qqw0OwtdkKpoyesDfMlde2xmHrfBc6mQR
wKgT3cc6eQWxqEV1DEEO2osuFHYUHSq4nf30EcpQkTImrPsGtuHWfvyI93GNZjNL
M5uHIXB61vN2ZahQfPEKm0s5wuLk7kTv6DBDonJLah53ENhEt4GgVvtJJk/UNGPF
lBXXbsb/htzniljPYGF0cfFKL/SCgjcLl+OI+9mjWPl9kKh+RS540g19ZKNNejtY
2WCeqXu8j+pkBB4xb9p14yUJafYpAjKFc7a4vBqciIbMSofM6A+pOmiRZreUsY2B
dSr34U+lGHd9aCAfzXWrA+qa3gAqQbPqXu0ADZabpHVJSkKJDrE0WBjnDv4aouxV
FBsa4BNVV0+tfuEUezfTpZsMrVpTwmr/TFdd3xx5FGo0lzD/QcOl7PDOTs6/eWyp
BHMRjVPgBcVYvPO8pfKU3vcvqsiR8RB1gpEh8CeElfsJLZnSM8Dq4NxECSxoRfmH
cVVJjyvqGxhmBNGHduudLQBVahpvW9u+IUYgmb/9GPrVKE6/UjXDAyfl0b0recEm
BAlDVNVIpCp8cwLxkBrMPqonZGgit55J2vR1A9wtfzo94a9oVs6c/aIf/kvepclO
Qapid0+8gKflhOMVk21klYt6Y9JxjeWcw1E+ZjdCbQxe3Hs2jXXaRkG5HHKSrHzZ
P1iGLgwPC3pq+FkZ0VoD1lJVpIFBmAfzsEeb/+z7uxy/2HWB3DbvudoeWvzfISQV
u4hxV1D1gT/5KsCApLxyGkneXu9udtJV05dRcVthXhO4ZkkEtT41d92fbn22M9rg
HJcpvE2HhrdCerMLJjmkHCj+r6T6kc3a1454sUFw4ysCP20aBJMaagTcZo1KGnS8
bdOasLi4Of0TxFlaLqiGZxqt3nO30EVALRYdo2OrRZ1yJZBA8NkIMsgoEUXfGsFO
CJLDO4QR9I+ceFf1yV+Iu7LJHWsQMCS2ROiFHvBe59rwa5fpuisWhu9HwtBC451S
igfPsbBPZDp+cYTsqdaosWHxcCx3hBosLSVFUFzNbkQ=
`protect END_PROTECTED
