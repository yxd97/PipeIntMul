`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LnrSnw0HI7p1EWGLxVW0P3asianEPnf5SJM7wtNW9g6qwqGNrXN38MEW9OeqDoPD
NyvCs+I92K+cz3/X6MPC9ZS+xh+vUsc/65TxC2/OvDc4k7Iz30b1WCDzVfN8ZZcz
PhW//cwcHuDeG7BbJBf9/NbBreZrLK9hOwbrNlwGD6P4QZoBv86n47IGLDts96rK
d7HNXjYVO9vf+wLn9w4eVI1TBN4zzL6yTOa4V8a5IGuN9RWt5VCtzbjLeOb3Vjmk
s6M29u5+An5U3eTpNY+LzX3s4mtA5g94HOb/a3lY4icn7X7C0pVI8mzKdoeo/F9D
Y1i1fPJeUqjg37BZpczNxAtAfhd2QFPX1xsZ8ki8khVn4fY84pjE4TxcMltP4kWQ
VDAPIx9Ul6hPKiG/usK/C5MxqceQ3KBlJ/w4BWlyJXk=
`protect END_PROTECTED
