`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/1RMZ5DJU3f5Uu9c/9JOYMITmDU4Gk5msk2ZcTODHDB9CF7YBT4NgGKVznTFYfF
PnIHgxD6z4pLgrAY9oP4gUTUZNkLKRYUJP8BtJ+GyRUzT7Hg5Py8OLKFuzgmdzk/
1djESmxL5h2riUdioCRREcudTqnmW2MybehisMjVXlY9SEeM7Rz4SxcoQx7vcEPc
dtlHlg/Rj4AcBJnmJzrBZYsBb96lQv1IqmIig/uKxrNDzPFzEjxYTKulJ4VXW4U9
oD/55kuxEFsNVX6M7lHJv3SjRiMdqlz8KNbz5bkrtFE5wxzOzPfEMzJzEEq0ad2a
S3AeeCH2CkfY2WJwcVIV98HOCMejT4hznf6LUfVp7JT+XqA4ABuEOhICmnhnuPcP
yaZ0ekl7Qw9O95ZZJvB18TKwSzyT9M3QYnC6BSQBp9k=
`protect END_PROTECTED
