`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pxRa3dIjH2sSIPp/Bk94HuG9XKiRGymmo3SqSfWTviTU07ne+IPHjK6x+uNPpT0k
G+kLVskG8rzhBpe1uqz+KqKzTNZd2FeFZQVTBSUDmCKnMSi36QWLb5pYodp58sx7
X0aZDz0w/Go13pmUraW6W+VWcaaHuEICwkqePWHFQrbdaKEt2RepEScJuyM000h7
lTVRICvAwRzLHKJPgIh6F59X+YesOhKZCjE2e/d9Ph7JKb69R+6bFSQJpUaFTsmQ
MaM2sfzFIW8gbxZ8SSl2zouLlvnGycJJGIMjc1u9RON48JJ/F+774u8YIxO1tC8I
GB4JmIAynJ20DkZLyJjFjCmuxsi2kqHZfnuZHhGq8HHKTnlMaU+bd4nbSGeUOm6y
`protect END_PROTECTED
