`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
prM8oERKpq0nxyerv+ahjDy/0MpCzN4AlZlQhkgN/iLItQg3yyuQJdsVAuGoXImh
Tb/lIx3IbvZW8VFEreEVYQgmp5YSwej5/CabC4adGym2/oOuIIGedaTdKx1U1HFH
VG1NrDj7IEmwYfdNeq6qbDqdj3NJM13ocuk8QF57gZTHwHkXp/Sdampr1YWWH4vE
wp8eyI4bsjk/D5bxC4gKJi1z8aNWtzLYL/4h3e3KQVYzvWbWtBG7EaHhDxLYk1mL
nSDqMaqgFmC4cZMzRe1fK9MF5z9AKUomSjmQwFo4nnmMhxJP4+Ey7t2f11Wo/K2G
9VL4GnmhqM6SMC0hq34vB/Te4eMnkR0sd3HPw9p69ySz2LX78iWwQZDH7orF8HNE
jOtgoekHij03MC2isZ9CF9z6Puht/RXCwTWCmr7ZV5XKqBzH5ZFjPAI1RDYBBQpD
uuNKg04tPxPckMRkDIAhsg8jKeBKTYkNB8X9sirgqVMVPlxYZVYeYw2l2QJY6mil
hF3PqlA61x1twEC7pXczxBjmKu3fObwdAzIQHNC7j4GVEAr+NzLmZSpIWbWs79mA
b8gbJZkazxCvSl37VlAFLhlTAXj1IEkkIEIIi+lZmmPHiusFZ/+Ojv17ndFeBRHk
HL9zagRTZ8r7wPPldNqBFD+fl7w0n2X3LhBBR/wal5ZYYa7Ybvnk8nrpunWy/vne
5Xbtz8WN/jIyyfxNqO/AeHhuBhjc6HSTQgqcwLDlV7U=
`protect END_PROTECTED
