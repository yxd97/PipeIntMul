`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pyjHbHU3zroooK8ePxRRbCkd98d1iWaP/hw/BNlTbO4EoS4GKoDTJMPQLFOd4KbR
C8ILi9wUYOe1ETl90bJvWjmEQ4998i5nr93YYCdeRSdHOM4W6vtuNCRAaAGf/odD
CKy8JORDN3Lubl0Qi0k6pcDnr7NqxugoRAMNJgHTGZcaYI/1ogno6Te171jRf+4e
nO4iPU2wC97lJ5kyNaTNjFiNY0gRvbSVVjfXDk/lYWS5lLcfMDgUSVNbVvBN1OKW
KAxFJydxlkk2wbdSFYRM3h8FaeBT7OCuS/mmMNANvTTuRQS9rGHAuoZpCseKf9sR
GRXxWWovy1+tn5DRIo+z1XNs5f6srn4fccUMyyw9Q/yerQaHL/xyz3+6d0StpNlc
x6FFyKGK09Z6gHyUmS7uGmwioJZbGNm/QVZ1OdlgRgfijaBkBE0AaxRv6XQKzImS
2GwtOhjptwvn+gzbsq4hXjwhF/rEEMaAFSN/6CMXLd11h32rCYqzf56Jue9uU2be
WslLM22SGPR5DiV++SsBRbLVsD4f55LrWRmq2TI4yPhbdobiWyPT34v7aYP7j+vK
Yfcz5edZrm7uT1dWqqhsIFJbkiXGymjhI8miRblz2M9vU9Fr5FzXpocAmwUEsnKb
WU5H0QHB24yHaPI/LSG030n5RbIpEqMAtwq5Wb0g8Ap06ceSOk8NKyBP9jvyBCO1
41WvFxyrNsYq4wED/UgncnwYEM3jFtyhSVPb19/vIYMXrWMxEOZ6G3Gz6dMUaEXr
LxDntFFF0rUoHYE5VwXfAaKkrMABZ0Diya+XfikZsGBDvS5tmSEoxYmqeo1aqrB9
9HSyxcSwl49lgAoq1pRc1mAo4RKdx4KcEX9h9roxGmbWXzTOV274tvGpYn6Y2dwQ
6AVD3l1bcSnPFkmNkw3nFGPDqKTbeC5YjRde+fPnse51S8FmlOHt5OHXVgIOPJhY
i8F+1aihVxAcZ1e3dCIE47Cw7X3OJ9o52dQxJuc7kyySdRU4+WadeEAfKEFbHeOv
CO1iHDWCU6O/PgsuAagPB7Jj8xn2d9g8fFj4V7CjkgqReFw57c1blSep/R4eoNna
u+cSGfjxNgrPqfm4l+eovSvQVR/jcaw28tklWTvEJQ+BR1olDcncI2HmbeGhpdIB
FQEfHacc3f8FeYyGk0MrvE0+4HbZ+8vOM2HAy0ospTQzGstClUwv8znIj2m1gx41
V3f/i8bND233ThUUelpusxuwFCKtIHI40c1cIhyaVQRhT+CFLayZoa+fkrB3Jssh
bFlze6OQ0hmjjLf0G1suKvj62UVT025ZsR6QVDtYKl6aCUk1u4CAeUhM+iKBSChn
fJESi70NOOWmVRUg96BPG7V1DZWgulYxjdvEfp4kt0PryfwO2n+gsT3R6jIYtfhq
7BYpB9R8fQ3us5ah6Q9FbfwZ8NoHjTwY0eK9Nl9wLEOD7rd6gMhaHE8PEL0M7n39
R0KIOOqmZNQS329/CruZ6tuTJGLBpB2ibf8y1b3oJeER9TuPLS56B+UgNpTKEjzh
BMdx2w2njEHeSYgExUUYGzoulio0CYLMMTSzWmn1+QJtdF0cBFMAtHgOuXz8dYu6
PCsyIa2MHBaZ/xaiFclo7ThFrIGzr0NYTM/Xcg2RLENy9LPoxLhOZpYoVzwfGqJ/
pb4m2EauqwCOjrDQInM3hzZo/1glIVcBdVY4BeSbB3duSKddsUuFGSPqhgg5GIgU
3z57VP9Dv5p3WXU7THGHAXYPXMKZJTi1kp5cGU16dJ1G24L/MZT9+ZOoASIEFs5b
OmTpQWsdYnn57WgPlX1PT6Fi0KKcYnnY03DML1zZAAZvZyeScoo4SSNwpkM5EstT
R8Qryw3aKF2PbM964j1twDkajRg72256AzzVimCMFS9kJdWqs4y6Yey/wuFQILvR
hkjrQDV6yygOYGPHXclo9jBplLqtGlwGZ2VqYAA+cEiZ+BymzDnBpR3qdRNTiK+7
t8iRE/XR21reRp7EE1shNioK96a5tYnHhALR4uAJ48CAh6g1JjTp7yQSiBl2k7Ab
XhcBOK3rKDy++aM+wECEH7FQks2p6Id0kIjZD97HMif5/mvoZ1jwFk7avT0tRWS4
9zNFzjH2JO/dDI8fpyb9lgeZfB11Bt1IHMB2DvMlCTxYpz1xznpTt2CkK54EWgSt
ophOqB5N1tfUCwyZmkaPnKDnBR/nU8ri9UlWDxQEjIrZEaVct6tACTx3l5VJSKqk
ErpNnqDNLGAZGaXXddXQmaCm5eJGVyQfQelh4ldkoYqXa6lDBOwEWN9ZtgK0KkSy
0o4oZvu2njTFZLDfy+RWVCDr99WudRbjpWsDS3yw273KGir3W+ownWMcBWnLjs5P
r2gp1qwo2ablabhvv1ql3Ei29CwirKE7y5xu2ljtOuUtRSfs6A+AhnLJ4sRrOVJw
VnVGlSOre3bYXRG2F/bzHdKzMqPEYka03sNZDVfTxoMoBM0jveFnqGdd4BW3NbDJ
x4cIZFkcXwNALydNEPMLdI06M4QGlCRHMjlZL0+02yDnPTnBEUJFq3uYGhPpJlb5
s2x+io//nXVdeATQmz1pjBm77Lp3JicCVpBAYTJLUPO4BVonQeY6NEYgrF3c7ARL
8D3D5LTlyNUV3PcqZj/rgxo0eHtS1zw6a2vkvyr/PHIS+8yNhY+xpO2+VQ3gfTZC
v6Bv2ng1SKmPGpDFYZfokCCoaubcg2tJzxTDcwG4bYdGbVX/HgAd5NK00uZpVmRq
lKBSJTFaSeEye9teg4aG0mR7d2VRZBFRz8tWSKDf9G/cs9w1sKhMBzQan9pjbOVM
3A/PfxMr3WlieWO7zhHTEwhQ0X7nKc2UkTX6WzxEKCunw17ZHhgCqSdyZRDGVnLK
HY1lok5oV5bO+7SIX2/tyr6mbKp8ZYdTws0JJaVlDgyidkl/6OrOcKuszSKCF7Jk
iiE1LGsB4xukz1QwDtEOndFnq+Qxl9UYzl+RJeSd7/ZpoSS0QETFiAtKsYDqqKuN
awKbZxfNCg8vOjcVi4518Nbq/zHC7QFwsBBtA3GJbWTXckffugrH5nj7GCvEl33F
xtMeQO6y9LFzLtu0Rc2/m1G7zuxQl28eWQcX6FkTh75qk58yyBsDoI2eXQ1Vfgv2
6iYFotFVTJ2JYoiT9w4FWPjSvHqckjwDn1PCUPofj8s10QGLGTqGVaIgqbaKb47o
vOV86LitgO4MQATnFI+6u4fCJNXAWgctyf4hfJmbRBC59kqE7T/eQ69e6zUnASnE
sOC1phUAwvzPBhn8sQoi2BWFVvYy9VYVjs4iYQfYlDR6x2IDz5/dneG+WryGnURb
HS4Z5ROI478+m3n+6tW0XitkRZVC0aZih9cSZloxgbN5aWo3LmlJmhVzNJslxIXT
kBbeVavfyWvgoCT4p8yDVBBMgIaGITFP+fO6HMqoy9YdGGp0koGFjLB4tX7flSTP
uLTLyTfz3MH2Cv39KnIAgfPnSG4SuvZZqMP7kXTWxfSY393oP3wRutxLvErZJ4Kn
5PHmTwF3dv7QmLWv4mRN7ogFPYslhGpeP1W3wD06sB9nB9WYcYpjMzzdzI2LycDV
0JMig5wYdxH6EyBck1dcSzhi3sjrkgRYaklcyUkyZjcVLBEMI6I+k+NbjEchq/rz
ZC2lSLI+akW1SQ0vYTstBLktqz44rf/MmEGWNtwF+ovkYgsuWSCtUoXgDnCF2GcG
jIpqTLxVdT5Xrkn5CPo2bUx2LLYBnnXE0esnBox4h1XgB7j6/5fEwBXOgWoYhZWJ
XFCAQO4nC4gQw/uGSa5WdM9Yr9Yb1VXFeIyMD7r1jybR6OZZOLQrc2S9QRxsnSTw
z9H2acBc8uNVvCI9AIZ14qTRrPT281tz6BBAa1pDs30EHiWf/WqobVK6eJTlujlW
nD+fwISiTtQwoMeAmHPxpUXks+hS+KOFhmVWQtby+m1eE+VUGrIaMKeP81PFLBV7
kvsw8mC5suiNHmNdSiJCeoqmZLIH1APH5nkhnJTpVS0sVHpkEzNOZchONUho+RMy
TqHrxSLBK6kACEVd7ZGrK9XaQtLWagpWbuHwQEa8WCbeBHu96Ht32f4Is+YwmgNQ
XRm80OAJaq8WeqNxI6J/pNsm9A8OFOfsq7gybV8EgxGuIsgntVbrv4gylO4gvDge
Ug4cXNZwajTwSYyBxyXFmEST8EwwBNHpADB9ynPtdE4CBQzSLguDS1ujOu4EgaHn
2LXhNLuFhT1E1L/gRJIBZknuk6er9z1lcfiPewhTXsSWiuykLENI8pnfPV6sYMev
iF3iHTMtzOHhRITkQIf6rIt3StivuwiNwMXnYeilC/jbqzlFZ0GocpJI8TwuRPtV
4n6j3JObw5feB+9nJumfsFpwgqvXwnnNxSAc8Mtb9hx0sDXoStYY2gD8ykZtJbR3
c+Y8B1E073mUpXu0AymDeQMdc2GO3oFfeDufb4E+T5oVhGsTYApblcUtt0Zu3qir
nJjJfkGVEESqMOkNJsJbHB0dFTkq+Pizc2xIPWiNWdduUz6I7xJnGi3PemHKwERd
J6JyP5SrXARg8TZjW0z4OCvA6iv7ggF7veohtcJZaQOa4MF2StaB0Az4Q5DyrGLS
Vimo2yQi75AcuWyd0dy5Sto5Vn1FKbannsGcPDdUklBym8F+ByxFAcMutFXJhzAX
BKhGH3CobPfVFaZBNwp2vHrYzYQA23ziIMQL9lKyOl580D9RLdNiN7yzwzk4Uo8D
NZO9OBKvt5yETKgcnsWQs3bek/1lDhEJZPPi5UxbQQ3QIAAAkLj/jeVvBIKcBRDB
X0kicdQsWqoH8s+k7dsDHgeRVhO/wIsomqNDQVqPkN6kcRZ0F55SjEvG17ixRvMM
VJBEIhPcKMznKjdWFNuQXzQ46EP1kd0tQ2AdtEcVGRLrO5kp6owuzS+fM6sl9dUA
1ilP12D/GjVnk7NYBZuFYl3HS1w/cUpTNmkid7x2BUuve0McPpTrIKmeqR9gkYFq
pr8W/Im+VEiY+1OMOfx0gxdFXcFlcjIlFPJG0pixR94ds+BGp99ps+Rs/k8QyQ10
mkvIWz5l/stBVBAxpW+Dh8Lj9u+/NNsoMKHwQRFoXjXB1sg5IkO3Ocf9Av6Cjvxy
zUwQ2vZjUOWOahbqusf6wKh0r9XId5PN31rsHBMgzEWWGzGgUpubDAEWztFwHoC1
J/nH6xdv1dK9xah8W1hl0c/lnnip4ROTIa3VJlNvJ9WKI8vUIoavGQ2wPKpWwXv9
BCTjMSM7d5kp7XR5v7MExhuIGK0v0GZUrqVSfmR3ZHPDabHtoPJ8ccbZ6LUSQnNy
mC2OItKlttg/G7wt6nltDHts4Lmnn827TBv6EnHaGfiT7BnKcwbQ3HsmlN4UiCKV
PrM/Av7J+DgVyTO8PXEi+rCqL2pVj/QuNpHxvS3JCb8RvSfxCdJxs/woC2rWRWBG
B+XKye01RtjpIlRVt2jlAxRWz4NtZaY0YtR3EaTf4413+Op8M3xx8uo+VYg/Hssm
JU8LN/ZBZKpLBUHCaLVCZ8KIbWIAADFanllacV11VIUSxgJAAeLY7k9HoL9TqG7C
gscqzp7bQIty48OUArLc0T+DyO45lqKCvTCQ/v6hbya5o/iORJn97dVQXAWGtOXt
na/xoXX9edsQWjNe2+6BHw==
`protect END_PROTECTED
