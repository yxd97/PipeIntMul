`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ZbqdJFps8MTFsDTxwQJgxgRBqAWcIgFn7mL7Jww75c60CCurBgXBxxbvJypG2Fs
Co9l2TGfjr7gx/vsR4r3amgH10TuP9/MVDVv1nOrOgFGL2Z5SdusA6UM06fmJ+gU
aQwpPMMgSduLlfMTIo02fGLuLRMCi4zLLu7uIQJgGXfQWDO4Q/o8nHYoF7XOEw6Y
iw0beYPOHPXE1CU3GRFyt8Y3+M19b7zeVxtz51WDJSbWiNenhBZd1UUREjzrbzLq
PNVZ40tFGi8+O3Z8WaBmx+DDpVPwajZWtNlkqar6B4o7n505zjaoWM+i2dG6liZx
LbIrdxzGlfF1RhRb6DwqhJHJXKYsC7bjoPpQa30txVFPAT3l33lYcKwEHN1iYN0p
tH/o7BAYy+aTyG3ixh9hgSCg1tPKtPd0vhcIBIhdQJuZPOzIs9Zp/xNevO0Y0qkx
cT5d8dwM8i+5Ls8kKdYRi8ZC44SQ0qcj5/xYTzkoSOSFjS5SH5I97DM/A4BJBRNl
A/Yk98ssH5kSqpThEel2q/sRY/7ifdZkK/NM2tKqRvo/WT4FtK5fQAxgDSx8xmKp
0RdM2ldJD9GlukShokOOhci+TtilljnBqaWk8FxQ7hI1dzr/Sz7rdkVcdRuQHi33
eoSGsNgg/9bbsdqGi4XcZPgHv5Vxm+kTN0XEXArmyO9RGoNhakMjyP4szRZHLvXE
s4o56j6tvHpIlsuv8Kg3yd2YQgBYT+OPgrnCeyRaBMuEomBTFRdR8nYuCAfX750r
POG7rmWZrW37IR8DGdNOKvIDbmMZWVuzx34c18q3uTHLDf/ru3/F2MpFaoREg9OF
NX1pFOJ+SitJcLfufHf04qaBHoAR+8ZYY20NsNCSKKolPH0A2aQlAfhaK5Dh3IVe
ygabRR+8X9xdHZD3G8xOH9/PkBvADRtJu/Dn2gVNIHiEbp727KP/y3ykF+NMbMka
n5steNbAR/d2Jgw8W1h+opJf9NtERsQuQyNmYSWNF+OxCLn62Kh4x4qHlC38a0mA
RM4P/g7+jmIXXnlcgtHsEYFcGzFJv6DAQea2tl2LC8a8v+20L+XoCcExYNYYV3IW
k6v+ptPXAo4LAWOOkg9LFcAYHMvwec4D/zzQB+QfwbQj6QQwGEcl7TrtyUQUQEPZ
3Lr11STfqIhmS5fOd9LSLj2adC92e7X+TgkdpkCLnQDh3Wi9BsafUhRTZK0wbDNm
2HvTQFwoqcIqqebBkMhzsilWWcW0PczFklPBLvnS3OPT0in6Myqd5SJttGjLkb8v
ZkEcHpRAjfbTkwXp1F3mBgcNhcAqwDytWlMkRaz01g4By/K8VQXfVHn+dHBHkF+V
Jm/g0oMQJk13ZFy6h3uutXLEbzSm7bPPsV7tdRaqWLWW/2qpsOo4i/buCudakoKG
NGO6l7J/chk+6FmW3idIclFHqCgcNLdiiPdNKA7PCkcoUrxr3RUlcZq1oI3qP7Vl
kfA0JClBPBWmcOqJAX9qHUxe3BWvm8hEZrqQeKd9w66uMWPC81I2c4YUYxaUGznU
M8Dw/MndjMMonB6SJNQWKyC5jsUYq2LmPC0s33cKmBnZAN4heMomU/iSJKZHCVPK
TzFiaP3RoJhmkGy+0mJ/c8CiJQfGgS2qSDzaSq31NuWxwl8n60rb06tN2M8TXjeq
2MO7hRxVvZF3Una1DZ00IkZ0MjWjDs1tVQ9xhyDfkxVjsA55e9rPKA8jAGHYZ/vS
cgWP7baBFwaLIKCSDSAArFy0NM/l2/4TQwaOKRyOqGMK3Ohso2XQ+mmZerl2Icq6
ivtWR94EmjB91+xPyDXuTzZmB2Ax8LhPeTTL5Ip82/cDVjn1pvlAOmUhBZ4fWaLy
apR1jbhj6O/yb5lIJk45ZLa/dpPcrHwOKNd7KUsyRtLsNu13KH/xZjXIJYEymy+5
OX/aF+4LLdY9zXh8+kZs2U8ZRgbWm+mhzGfWzuXSNhwMsWN3dxELPReznw/i6vxB
u4H8M+3yBK6Q41LwuZa/K2zbQ8B8HoCQkqQ8EnYFKfBPMByO4diLHNuAfZycmT1y
cn/ysz8lLDLadafvUSm9Pw==
`protect END_PROTECTED
