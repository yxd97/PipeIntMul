`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZTsL99b8aeELeAE7+NjXrPqwwZeojXcPown7XcizYyvMttMP3qgtxzduywXHCzo
2jMv1djaNt1OI/cG0woL5r2Ok07fjihWuTNUMf++g4LBuIMXoBunxPBqOr3RyNdS
8Va+0w0iX694o/MjQA3xmasIKTlUOucngPfgqI1BEpLWyNvogDxRcrEJ+Ems7UdN
oF/YWm+8+GekxuvQznGnqjoLBLqBf/69EQpKZaiKpO+wFiHuvf/F2AxB6p4iAiMK
05LovX/cYSefNh4R/AqqGJAEWUGagzDC1AzKwOLHE+mFP+enqAHf7/CAhczPZtRe
fIR9ha1cLuZHFz+tx+k55k28QQBygX1/ljH4GW8cvTZ+ipPoHhW6GWHYGSIIsUrn
XuekMFkbOWXkiIcBEB+NCu1jjEtuxZPoCACA8BZfDX2DfOflgQTTSUZLlB286cEw
`protect END_PROTECTED
