`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GKZJUPAqNrDFec28Qse2AUHPjMZ9DQUbwwpuNb6TzKNCJkhCmNwylzOfCoZErUEq
RSrUBCR7m2aT1+Of5p4EOq0YBpoyLwQtJwK8S9i8LYE1mA4tUKNQ3hHscnWjZloI
muIU19+yd0C5inB4Ey0FPq8OyBgaK8F5lkydUx5TkftebJvYQajrPIMe1yIf2P+7
GU8vAqkmeUwacAKxTkm3KcyuyvlN1FOm/UDZ0CnT4+m1GDd/zpoT9VKBmhwVlAes
6z6F2HxZaFOcDJuqugZZCfb3GbraqzS9OzCRn/ADTeg+vFLUuLv0k9v86Ua8QMUt
GWzLXcFPWMF9muTILodXiEhctmogM7Pu1g8z5tB8Cr8wpY/qZxSAzKRFbfUyQyrC
GFwOB7cVnN+iF0wzN/kq7vj7j3fbp/bw0ZVccPF5iL7XuDupXkoVh03RJkrfNNiL
3RVeDzLDVPKhLXgWuPvqXpv20+4wJeDcCO201eJGvz6EKLpjdnDEBqQHo+d1MDUH
9HAK1eWSFhhAtJJCb1e7YqKVlT4SiuKKDsFzTSFsVLfTHdc1+GjE6QwtTNLjRYSh
tCSmyqKD8wZKNhqQMLyp4VChn2NXJ6zBdzVmbMAABe+eMfMwrlZVc8OevkHfspoD
Ph2r2c6udDJYpO9ORf5fnyvDK3QtjvMOWno/ecqMUwLvBWvkRXld35D6k+4rxr3j
Ar8acAcG/rZI7o+FsKkawyIeHJtk8YMerhiQMfMFT/NIrc7/UNBbcE8ADXlv/ADp
YcT9pjSKv6nTcMdHv/WX54YUdmdTCb9jw4fbBLwswtFW3ZW4zthmhFRRX9ZMWLYS
3ipm+eB28CeS0e0A/WEL7R8vSfL9HF9SASp1Nw0IUPMOuZiDHzblUuyMMko8Mxk8
QEKD9dNBkrffj10elVALupcR1mO5sHBqv6xRIKZSy7o++Ai4M0zzRWrI05dY2V1G
hL1RXUXvk6xj/iFAyfL06nYLTza/ghr43Iwa1o4jID/a1hdnKMsvKHp7/MMRhSuj
m/elY6QGO6QASjOpOC3t6mkmvuRHGFd9RbBMllvrN0VLMTUHZrMrbyBuuc2TRTBC
V15aTDGVN9+r7+TQ30TL/ieVlkFNNBnnD8AvfOdYbC8fOhHGmhSRV2G07BdP/03D
QOFsRfOO5zRwej+xjotrrS5NpguAtKiK13RgcFJayykVN/x1E10RRFeUcztF1DtE
IBnsv1DTU0jKAuZQ+D2XDQgBfyVhbuwrne1lkSH0COfk9KD3m2pYYUV6B3BseRc8
l6flrWhtVOv00/JlWntbLQDz08vqFjvVi3RO86ebETLBs7CRKxI22owJajPXtPDD
XOfQIioaEg29rrZ76zIGLGHjXiOhWz9dvNiFPR0YxpDhpFkCp24ltc+tVhILFlLL
HsOTK23dn6XHOl5KZJHPo+FG3ghArwURjYB6bGP4Jy37MVpTWvuMp+hqVvak+9iD
Yk7D5/Gl72xR2Fi1P5Fii23YDJ5mZE/IZ6GavE+7YJjhYtsjWw1SzRbLL16zn6X9
AaKcMzrGI76CLfaSyzTLUc/aA/Eo8HBUDlUjaZ4iZb1kpwYpIqAn7BgPt1wCZ6du
1fKO+I9iBPGKkY8GZY2cJPVrOh2QemwkFIvj547A5EWrid/ecREG8bnQE0oBHheB
ZfJ+/dL0K+TKqO6Pg/6A9cZpb62Y0gQz4bia68XrwozWQsyickpFOr/su5/9w8K2
cn2tXbyfRUehGoX4xJnRTloRBWt18/S7I6dB1+40f7PwupGdMXR+j3YS/DdZc6Sv
oLwYHokCYAlPsgjis+r/o68TkdPio9w8gbk1KvgeiHRXXb5siJNeZoI1tAukG1MS
sbWRzLz/+bM7oY0POOvSIPgPbUbac50TejWc6Vgjxxq4mgb5FrKGzeWpkmackNn6
`protect END_PROTECTED
