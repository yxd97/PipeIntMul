`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/sGgMaZ1YkNfE349zJVtosafiUYe2KaNTRIxwS/C/4WfowWdS3DSTk5L/xnRLSRX
3GJNqPoAFwyniB3NmiGba7jliNcnd20Ydc9/Gg4f0oUG5t8UA36znvwqwiw3Cji2
40hlo9s8QM6+MBAfp4MTNRLpwh8tq0bdEzOmpI/hrYTHnbzwHVyhPVnjZ8rvRRzk
2++xP5lirhsBckosfABLdXBhdUJlLRqcSkFWoGr3spYmTHkWHMUi7a1OQT9pJ7wx
PQQ7gZL6bwHtzhy9P3WllEdDGbyD8+Efag0ULm30uV6EsBbis8Eh3mGNljbYWtW1
5SQ8QPiQf+QFra0cWDfVnnabL1DpHA2IyjCmcnZ33uMWqQ8K8xAEvU8MGoJNejh2
opLtSzXm2XP1Mj7JDmGSVbVv1Azxv+zg/BxodFoGWI9JoNQc7Ekhc4RwKxI42RCi
7yMGvaFtW2GqrNI8Pxu1zFTmnSjfHsI26WiGh6laQC81oTml7bte1Q1IulJdH4I7
/i8jmTIcnCkjarcZimxzkwdNPeosG7gmpjPXLY+erb8rcTUef7XMSpmmFvpac5JF
Fa2TMtwosMCBSgcGVaslTPkKQzA9u00SSr0BYkEEG4SAKX5c92yPZoWseGid1tbc
uXOZXn2U9klDx59j9SYOfRQo832YsRZyFraVvFWpIceg1gBvpIW73ZtfI4T318Ys
IwiWEAdX4Cy0am1Bx9T/GaxlFkPw9laLPVclv4h3SiA=
`protect END_PROTECTED
