`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EB2vL/BMZJjmFJzjinNPuBZFqf8WUpoi60kRvQ1yock19wLjQsbUZaaWCUZXiI8W
MQdxEq8hE6kWF5fvq2palamfSpg15Nz+gqQukPyde5RZ9iPOMsTRbGI+07PQVf8B
eQyCiCbwEADU4Q9blXYcIR0ncrUGJNS/HctavahgjFjTYV6WoGL9vTZDzKp1jxG8
3D0pzYo2bLdp/GAahAccKeht+tbPutExyvljwmBawPkhSZtHJQCMDLej1QTmj9Kt
bN6ED4bqaEFtTd+lHuazusbw2/1620z1wVmAiVD6hYLhXnmv3OFUPI4BuUidvz4a
F/ypo0pEv69Ek9GHeE6zs1tm1qbmMDO8PkgtRtTb5exiQz3D5PfnadgzEEHdwlPk
W6l1XpC0feXymqqk+ySwp75TrsWhhUWG6FVsVcH3Qi6rSJa2hJ5jLrodwk/xG638
DwSyPenabPhTpxmzYBinRDikvqL0Cu1vZsVcFEAmIod+QVQJ/lfemBE+/CbK8vYM
rBkjCQGlxukRfrUCRdR8WNNTtI94EZrk5RqAfd0qGKCO/WHLSVG0vfk2n6sMBE/a
/nKpcGAfaMBCtvbhWtqhC5DPRkqWH6rvRADwwXwaUy2D1+ODx6DaJ4ofy1LeM6u0
6/Syc52QsO5ccmJNMudX4+9oqenmHOAl4ipypg7j7ygOE9Wbo6TTp8RsWccjuZIk
uxISsJxXcP5TY0Kv1bA5PmV2MKbiNZ5fID99MbSnWbXCpviNQFjJtveJBBDMnGLd
fpiLUmy+suuNygRL8FriUYGldlvsavl8pneETw7Ofqx8i7j8npKE/kvQI1P54m5a
46gtcmQlpgyP4CM9bhOLiqG6s6ifvhkb233+aDgct7woNEsZrr0tEKDsJWEmAswD
F743fULGOpvKwxN0LQxh+5qKMo7VNP7hMEJb0J0q6Sd5tvIZonQNi1+6iun6N8VR
tzHKKDtwM8Cy0NLj86cvgG7iHA8TFzzHwn/brHDTlInoOh9wik8YdfqqDaPkczet
f0Yh7jQCP299gn1BeJ/aIWpIpCQ4CDe4H2rHh5z3yImRMtlleHrW+Fq25VwGM4Ay
R2RaqhvnHYlKpykS2Y5xSif1oNSrji6vRjvtDElv0BIiMiul5Uk7b1Ih4Yq93Qgs
7eDjjaa/j46zbWLo92aURI1rqAP/NTNUsmRULfb60SecmlUbYgUfJbyOnVFZPEsG
3wWFGx/Ubv9O2BazHtjgEVq6c5sJAuZ9LN8GDd+biweqJsNsAZiCib64cetFA3Kv
YM1VPxvkkDMy7L71f4vBfsnfn9zTyERpgskcI0RtSslSMEsSeh8tqrgpfHzROug6
63mNsAPgmA1QMXp3pMCIQihAIB9/9HRgTGrYlHyDkSW0iPE+B6eOoRRYJvQkDDCb
zBPnVoXOm7Fie0WTxFNxEg==
`protect END_PROTECTED
