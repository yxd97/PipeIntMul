`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YfYjnDFVPT0aoDZLvMRcJ5a2KActnzQLUO+o5yrTuZbhQgzHaiG9nF6ti8H8coWG
7P11tC23NNu/i0TOkP5CjQr1CZ5gt/8heC0J2bWMlTy1XgosrQOGoQG+vbnPPYRv
8pwmsF4Curfy1PxKNIpTKUvLtba7hCKqPe9r960FaJhXNAYvgOKCxmR449eEn3OT
EJTh+KNze+ff0/LN3gPIfxnyNQ5lWjEu468b6URKh9ipaKLEyjjI+9U+Q3uQJwtH
3GDXIszwwHysp//F5fMG5Gz/HfXn/uaNx2g5JDFMcLH7Wesz8mN4UEcHk3r/bG6z
+EjtygypkO4M+QPSxKG/SHlNjSggnOAFTWUI0l5xTbIUfvOkwToNS+iVkb7xeUoP
+H3iBG+uuIqJ5JEYFn+4tA==
`protect END_PROTECTED
