`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufuuAYAwnDoWk7uqv4tt4XjufpQ/q3a1QeUvFLrst/P1Hv4cGtuU+mQ4krwdarN7
2o3lKpJjRjek9EvFua6jGsTsaWxB2YxfDybBPRsYXYlovSw5FnPX6kOoJJ3HL6Dl
IX/UEhWtLRrmgX+V42g7kKj13XX2+fG+enk0/SNmyXX/CK68e+XErZvPktCR5p6v
Xt/aRC7dGpd+TGe1mpYOezaBLxyLKzh11HcZasznrhqpF/c3YRRDn6Y6E4PPLw+Z
Av19WYMibxCc9hvqZI/O39aOXtSAFFS1Z3bVjgloboDv5UYnrLyWhHuNDQY/FdpK
SUzFnP45DakzxuqnorlP6c+sY85uHQSgjD14HlZ8OY1sGKYBuaPbEFgHkRrdrsZE
O0n0jloMrq0QeFEVeEJ/gmWyfG085dUYzw+qduBdx1NO1fjRfx5wSQO0aoFV0dkH
eLlSiWpycujo5Gc8KXiYDJKW5DmRVNPPWcCvXA6Jbb6W2jHMVKzKmGUGSNMzFXkJ
AwiUkiW5hjzGAZQmxurFXegCxwzDOxrhuK/l6XGxfVF0iYIUawovCkdO88TZDvaB
LTj1VE+P4sLa8OOWfRwOoNZ0GyDYJ70/cTO8Ly5SThoAL3POhV8BBdf/AtTYbrQp
tpTUWSt6jvtqxEsoCxqSneJ6uy1MVGIWbs0uci3/LrJocbGObXEUHMTCAIv/p1du
06V1/x4bPUs2eSZ2WOPkZITvZO/oGNT6+aauZCRHbFkskUwuBe5po3CrndV4Vysz
diNSuQKopdiyDkPVT07+9s7hcTcdWILcSxmQT0U4oj/iglYeHmawgc8ZAtRpVuWl
I10nBHhLMYqX6PpqsJbbtqG4oCv2v7Oyad8yhS7jX0FrkOM7jzEA6jMISzDyNjLC
pfWrDxVKOfBk2OOmhaTaUVpohtXATdSInIrDJXAPfqmn5qKiaoqjxKjUMOG26/Td
ZdN/ADyH+f+dP4YJKOD2Fjz9FvqfrnaXFMGPAovq/qiJ/MnMzYmC/xZChnZ7shrt
HNa/szQu7xQAFlwlBrR6KTuVVTOfV1awx883uUpypspi8S5C/W2hfovsFXilHmDn
aCWcX1T8Y+vyAQF5ba2BpziowK/fz068edsu+Kf1JfDOnY8nfdvzWXT/bE5XufYM
o3LT2MWqxyNokkJlghzfUZ+Y/nWzZYuX+oRB+4rmJKTq1Y8dowKHfPV7x33Mx3zm
Og7rWv7yxqON3RgJy+IzW+tP0IeUAolR0DPrKKhnyytKoEfcze2PqRNFU6jOO3qF
dZicEThQ7hvjaAAgXwxCOsysleb5Pl7xjmGBGOX12USJHBVbOe8Uz/aUtWZEHWUH
d8AGmcjAvFTn8pXuFRN0UD0SIUOODn/L5pMUuJdgcCXAwDvQkd/AYsq78RVyHszR
/Vddssb7cyWz1hJ4SJVvxPppGSIq0wkiZGE6oVOii86DVZhMwIpt1Kf74NHDMnGS
c1MnvdxG0ud0lovl7cFOcQ==
`protect END_PROTECTED
