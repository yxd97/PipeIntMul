`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vDEtoi9juYb6jUTrNXmI2B48qg2UgJ6I4o1qmeHSrMM6oj/Vke9qpWi9oxTGiBj
+MqtyXGNEHQTkgZNR+8KBSQEgIN7STr/4joXi97bwghrRACxHo2ZWTLlAP9Gwca3
ZobIirwFqNvM3WV3JW83iNW1++tAJc1h94c8adHiNfPHr49gS3qYkdWInOCprGSw
/kPFGg2DKeZlLzq3hz0MktZVGUgA/Ave4wTBwzDOduU1X7Zqfa59AaHwB+ejHPX1
aprMhUaW9FEgfTfnxT7xFfmHa/6g0sjfIf+7aWTHNJnf224T6n8ydnr+9gwvEctt
RJvtgK0+0hKxx0RI/+aZUNoj3d5QJFlWgU0M1wjsT+W0l0oGfZ3lPLtkYAr32hq4
14olDNHvP00NH/iFKeizTRFqKl4XX2u19rqgM+l4OWRrZjZCdB5xWEmx1Thphs4e
e13iHVyhQjEBoUXBQcN4QZlkfKGMcO3LOwFZKHz3AF7js3yxSGfTQsJaztHw/Oub
rzAB/DZBAj4NQCUmvul8EvGV2qzm4F0xVBal3sc8VowZs5lPxXhQGXKMns6jhW3e
kDlXds+a8OsIGHX3IHFieHHSyA50AN9xFsTkBYNswPL8+YZPFwNh3SV8zEB5TxoQ
0s9rNY9I4HcbaywDP4T66ZABYzGbJ3xhLvzfZ1cIQWE=
`protect END_PROTECTED
