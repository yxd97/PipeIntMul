`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5IZ2nAYtOizR8eECmJrWF9lkIGKdauHeYif5zeA35Sv1Xcy3TUUqkwKnLaz25rLK
SigwWTlS4OW4FZ9otJ2M24YlwP863b2ys82J/oFMj3H4ASJTzFX7cQWaXHRe9fdh
Z8UKZec9hqTTzOqxLxEvYrim0LniCQqYjzZbc2XAu8eLN6iGG34d7rfNvVhWJJ8L
W9aK0WLARwJe4GW6NOL4dj8+lR1Ssna3Pj5BUTnZE+JJynDspTUrXJzn31xT+Ako
+kbHbYv+B0kKz3FkImIaIOgFzPp9Z06FWkdEaQhWFCt2tOp/U7TrT5jhaWz3YASv
GNvNIm2FDj1rNjCaCUQrBO5K+F1Zi+2X91ChuyD2S7LPZBXKlUASdxALDyqqd+Fs
`protect END_PROTECTED
