`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m56177eB/vnwmF0n7Rsrkn/WCBblRqfiB+iJq8ednpw5qQsVw4w9md9dBZjlq7re
HKWpLJSDuveMbck8iZbUhdbiSFW0kGgxLYF7zqRWOsdN8Y3wfLeSBA0BVSw3JcVE
yxmWfeTT2CZcvHtoTiSuH4FIpk/e5xZzdejuuO8mwEvZF8ZBbHPxoH6p7IPIeTQ3
cVexiVwDfZxp7udQyBbQR5kpcpcqSDjVlaP0Tp74vuWwnNO7Pv2xIStF4wFuUoI8
QSrLPhKI/FX6S5a+EFehdkKWbtuXhQorQhW8UCWnt4E52NeMB9nGmLba+N8wePG4
d35uS0uxcXQVxJHJuA9tHw==
`protect END_PROTECTED
