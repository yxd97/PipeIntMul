library verilog;
use verilog.vl_types.all;
entity FMAP is
    port(
        I1              : in     vl_logic;
        I2              : in     vl_logic;
        I3              : in     vl_logic;
        I4              : in     vl_logic;
        O               : in     vl_logic
    );
end FMAP;
