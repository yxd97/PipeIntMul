`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AzXOnmVFb6YXw4C/MPzR3VGYOmhR29P7FgYIhZDlAtIZf8FHSqwtJlS8SoF5xOZK
rkwO8lbFClzSfkQV9BsfbAx3FjXVclkjmcgmuPV9QPHf5SipmkhBZf28OJwrdqtc
bwMEQT2fuaEpqbYihIxFXeukhnsxW1bddOasKDGfdFGJoDIw437Sl7FJCwJ9bR+j
C1Z5arS+6Ih72iPQw2KOVUnjmIAm7UHEUe+vhjsqtGs7P4Ve4DQUTKYAX/YOyQiq
TUie4niPn9OJRV9kx2RKh4gL/A/WLbJTaNwgVZSxGcFakd585hqQaiipNMJMDaOS
mJHVtb1E5uD7QNjdeQPYubj15QKR75H76hVterA1Fc9qFlFgoaTFqudlXNjk8KQ9
hfBsbZP2wKM3E2bY+KHLN7YZSEwxxm1pElSegK8HGZhSqjKgnws2IUDfMSyy3Dyt
3bO43HFmVReGtxvFfWTomfCPs4X9SJFAg6cW0Ws6VMRKnw4X5DGhCO9A6h5fKBaN
`protect END_PROTECTED
