`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNkAkoqAinjhtEe+Jotk93HV4BxgRH/gvL433R8FVJqoiu0OmyNvhxMxTtzktN9s
czts1LQHm7hGAVBBhGUEm5gSWUyY6wyxfxCdkjvDD+uS8WkWulSXS74Llg6GVPjr
TM26RDDBhMWwQC51n3hbprxGIAJxCSoBQFFIkzP50dvBQ4h7mvwRLCj/Q+DR60rQ
OxMJee8H/iUrR0vtGaXQglxSzzX1m54G8mACQlL6wmLuJi1LTwzhtiPeeiq7Wn3b
2X/ALXcbPKUQtiZ+YV8ugQ==
`protect END_PROTECTED
