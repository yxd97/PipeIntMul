`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l8VHYtLq50qG3dtgpNWu2TUhC6GBWrphiJI9PWaGpCUM5rqsjrxncCi7bX9wJmy7
AivlEsKxLEC0viNk5t6ztj1o2uga7GbempzbV1Prz9HE0g5fd7nUIrywqnPy5XlJ
pOhK//kxIgbSUncJErGerygzy6pVlw+gfFX2ZjEZF4TJZJXcbISpt80tsa8QUdkr
nWa0sqd4DStX6nBpsl9gCs/DxsNGte9HWSak58ovtUGH6+/j5/DxVfH6KPKPqbtF
PRYI+sqfofBRTvWHqDrvye8LJAJHOkjY018YJiV5Ic/Ng5BXEXYaSv3ow/ifW59E
b+xVP69fXrPEPZoDjtk8FkVZ3p+g52aEjnOE5CB8VICcG0sT9rBHZmak5eoMaNz3
V9yDnfp9S9qiVOLVUkthySBo5nPh6NvOzwqoI1WwV3E7VWVePGo+xNTSCc7xqY5v
AHkC9ccuJrU0WhmHYadNpKHmRkfgB6AYueVHIvM5XoIgJMZ+ZqTQ7ZtVdIa3d1tk
FiLUUtcfJkIs4xZAhN9Kvjd2RQTW9l/pDdFcXE/bNUISW5sR4mQnj30VC9+YXxXO
ySgjs9YYfr6McuXciXbWrMJQpK3INn33W64gT5fBCgHtEuFHcUT9BlHEH/UoJO/Y
+vQg8kwt7dmXGaqpkf5vX9I9Ufy7tS9buPFETr02yJAb/FA/h83rlf3pSIjgb0Gp
B9vSOVPc1O6G6Kwe5kxtXGIYyoyM7BrV6SCfQDU6BPM=
`protect END_PROTECTED
