`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4G8/HEkwKP5yoL0WA5fEQp7uEI0tYXmg+alq0oHF6IFTcE+miYPFho5OSgeQTyR
JTWAQ8375M494AYG2mt0wEHu/UMvaCcHD2nATjt5XVslJ7cY7yiBr7bFdDqT/Vzt
mkIXZ37cZhLgy08GT6HK41qLvMtZ77/cHB63+nxjM0MuvOlDzXheyjfGwapXlSzv
iRy1ICaB4sRINvNuqI6RosGP/cLpBM/m7TyjWmNOmTRt9RLif6I+JfScXLGe6wg6
O3FsEIk1xArmNZQ7VYncBodSoLczhsdCWrr3LqlzBOiaVn04jPyDh4miyNiEXXQZ
Z4KYZm96d/L3xV7TFDdM9tuMzzZEuqsG20N62XRQGUqVRHY/lvp5CZZvOzVd4lcL
CFrwr5A9fO8NhpIglxi1RnqsNeA52//3Yqb+Bochw5OJir2iFCSMnrpHfwkKb4/L
Lpn02CT8+3QNM+Kh8BXEAOC4W+BYrLyhTtmCdjSNt5XDJOJ2Ls4oMrTaiRdFm0hc
FOY+MuXYRcQTCaTqBfcaNH/nFg6ISyAVNjf0QdhPAxE/rM2S2zM06kR6bBwTyBi3
`protect END_PROTECTED
