`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I95lirU79L5Gsuvud2Lhm6nEqXg4URCTeY9ywJKPkDRk+Yd84Mv7LfK98Eh5R7Ws
ps1PvtdlxnBGI9zPn+MsukBEUA39ykgQ3B2l3uGyZCaWqkbG+07sajJbujxKzccJ
pG2f7PLzYawXCju4J/UjwrDIUMQpqyO8uDuayVyhDVj3o9XrqkOewxFhjlBz2gwe
yloLhOMxJgqliWR7prKFsslGcYWia3BHokc96siIzVXxC4+ab8q4IeRiqJHBsR1Y
V2H6cbrwgx9XNLR/PSiZ1iZ2pG2toe/ov9UJ+E/IZfStdGkz4U+Pc+bSVspgPL+h
99Wb+DRBjfLv3IEf7id9ALrIN7hNUTlWvBv+VIfLhG9ycSGoZLK+Uws5KHDCfIar
QWcvh3lbW6jMEucGWAiL07+hjloe8rsnFffbTy8OtPFTcEbkJomDLym+NhpYi7jc
`protect END_PROTECTED
