`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SX3ZuJvanohEsxCDmB2YUjJ3zKAwGnIJsaKNPrcDAFdRKlEEcNhtc8Ypi1Kae/41
rMGWD3HGuMW7dPrPk4eyEseu9IFxupZ8iUJzCihLLQAjxgm0a6H3wvSZCQJ+Z57b
EqzEU7ggRUWiW76iLhIdjURkrowXg+RxfFn4KFPFNpzuLmi9D+6aK9ka/eLAIwLV
cmZKY4UBxRiUlCaQgapiL2yJTeccEmFLsGFgRV/3eYE9cWcNgcQoM1lGR2j/pCEI
2wKdbFBwbCu4Vq44R7tLih0AT3PfUMw9EVKf5Sk/Ko6y7hiD9buHqgRiD7tWRECW
WrHGI2OiRxcaePqGHOniFQwNhImZBfzzqVhkHtXigZ5J4owlM10n+anOVuWUCgtB
O1cqLMK27daku/EGXmqBkyo3XYbek9bVioignK2JD5ovKvyFDA1wg5Kd+EjpoSLw
eaP0I1BNL9iD906D2PkpuLazhRSUTm4J4IUGJUQ3wg4gV18JKaP6WS2v0FfPyn6q
j8PR92KAJCXZ34BVnquMGvGepAi2V64JPjDEAtiD2NiVUCCnUCH9Q2gHkxYggXhR
pckejgMUDJdfe0SKYdoF3tW8+XS00z5FuphPa8C4yEs=
`protect END_PROTECTED
