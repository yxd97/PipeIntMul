`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4jt7dc+VvvwxW84IW0niZ4T9zyC1LyRv64Rsr3VXGQHmUybMrbFr0NZkIBogSDG/
HRGHm8d/Xyh+JHRkm3YJkFSblWjvbmS3T6D/kIVDpFwZLbGkP0goQjadNKNAZz8W
b7LGYWuzoz5UyWMqrhKmnlGJGU8wC5F7RCMfHCe5o9BU5u3XGjZnFsDEOYmiM81V
96HGrJY2pwhT5SvPqmM/7QHIT9d3t87m0pND5vYTfLk2bXaybYNasan8rwe8nhPs
xHqsyXQtgO0wyG78vNmZODc7NefeqSO+3H0iIsca4a7rwaCQcukOBu4ucEEg3gJV
c35XbjEu7kdNFCeV0zorjR8n2KIjwWYMmehmPCenNt0llcFUr+aht7JS8gvOL3i3
elCNIzXd6tsX//DRV+y59hs2kHB00m/Lf/XO3lJUGdXS9ob1WMhoxWNSnfyeT7JW
L2vY+JaMihJo4GMsojNpxUL7bZFlR/b+msmgHd7pMDTIgcVkGrTEzHq6KduGztVA
0fl3W8OqwxJZVoz4k7tPSjvZX67CYYVUOffz32tqXMLfLIb/054ZhOT99mXiBdG9
DWOOWAiVt+mNEpOfOIQ2d6dM4BvFiYWr6gNFVwJ/IsdTIiQ4Z+pEzZ1SBDt84kS2
UtC0ZdN/ae4gdk/3hvgOTT34X/wB7G4DIX/R/J0/M6ylzv7M1dGBiqAe8jBwSItA
hD06DfSvIhedDevWMMnEJEp0MFX2rnotS0Zl2pwPDvQ1gf7aqR5tiS5XHXGqKv0K
VvdVWDDJ6F6opmbEp/tIS0c097Ny13o+vaHIJSnktgTEj1HdTaeNhzv1a2NhiRPw
qGuIbG9psrHGrhvfV5qBsbYM2jI7rV2jz6JzPY3ffbyy6VouSdlUjbK9sBjSqVzQ
IvVmcollU005FJNNpPQ0XNuFq6PuQWpVgEf0DReWEeyqlwW/Hfu0TqtKlDUAkfzh
`protect END_PROTECTED
