`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t6crU7X/HOCTxp60NYgQY1FthiBsYl2uHOLxutaeT+xphx31LK2rYyqWPUK+nSP5
1ZPov6OJuo6FQiG/QIUju4cSzxiQao+FWHL3nG3PX5Oj7Z+7YTPQFeFLzObsdE88
uIzhChJTIOacAA+TfbV8PZIPhVlpTBPJTDfELroEUX0y4q3v5didPBSsK28a7Fwu
Nro4+pm1dNKDUEEyAfhh2aGTgDzZh3gOSSYLRv+Rbl2pzehPrWE+RaRbFIsMw8u+
tqkmabqxJOodVvmf9qWdtxn9ETNLaeBnU61JLcTa7wuv03pG/jdx0VDRLxXXcCJ+
EUTal23ahhCowPr9HGnR+LBpwnWiA4zLfY0/z1WGmmaaONR6/nX4yQb8Txv1t+FE
Iu4xpZ+Ses/BPsWRdDdHwA==
`protect END_PROTECTED
