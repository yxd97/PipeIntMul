`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fIgD0VRA5ljXHxG8xTtB2EmKvjdPU8hYq0oxpCKjVhO+BZQnPkdNd40G2Mknz9o4
O29xPdyZjVWfXsgIcfk9rr4mTRmAOCekQK2iDje6aVm2b4TG7tm3Wv9ymhqxkTM9
yK/oPwAEb5PVUpIcMhXKXZtL8oAfVB5ORmjnDOAOct3ZC0ItfdrVMC6twDNHQ5OS
EV8tIx1M+jhzOdL1a1eZJ9jnPJv7hPHIe3GnQHd3SBPBFchbmTnpmwhxCP8BX+Hb
4+zlmg031RB04b9bCoZLf5SlqUrxYt5Rk8szNA7RVZ/IXsj1iNBsA7PSP0HIk4a7
y/Rafgc7oSpMmxxLJ2xi2U10Ex2nQnls8psQQAyW9jm5FqLr651kTNJo7Y5zYNtb
enpNQ3LbMHFzoSij0IGU4MYFQfgYuYLKrWXL8l364lscbxVHA9LBmScB/UbE1v6d
DW7R5A7UMII+3oj2mzHqcZyBGcF7g8AaBzVqFTQ3s+oRvei6q3kRSjIlDQf0ozvv
p9pkfs+g6fYMdjIwXZdMNTmSdv7p7szSm1qDdQjVm/bkQUBypnZs8VUcn62gnV3v
bbZriZAA2ycQNUJcqM6InaRQXp+I0bR1gm9ACCQ9DPowQhFNYCd1TXF/KSjhMhd8
igatVw/WvKDE6HgFZgQC8LM5p1XwDkOWyMGo02oJx+rs7ZHQAnVA216n9D0Mnrcr
+hpMi3nl4wKUA8mDc4BhXcMFBIk40me/RI+VNGC4I2E=
`protect END_PROTECTED
