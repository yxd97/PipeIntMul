`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFrJG3GGsr2zHVHvvWuRvUTHsLr73t3ZkK036PYA4Zw5fLTCTa9Rg0W5wtJTOZ++
rah4pcMJdaYz4PpK9ey6o19e4m5RHEcbsc3qDmX3kgeDmvVcdbY2VAjQwKiTWOH9
5UFMoUzugQJom21GjCHy787DOewEATA5XVEzWLoOFkkQZ+EzSh6+PTqYNz9JBI0O
XkqDCU246zkm1SeIYBSZ7dvIlpCa5Qxf+drpj0Zw1/UXnhy8pO+U/GWZTVebgVgN
0FbIBqkPzEGI1d+HnKtDHIq3EJoOZZX7vtOMnOXaJceBNcNEBoWTM+D5N5+qxr8X
viv8A23lo/Eeynnx2A2yDWQlOEW9URhEZoQ5zIkfFyBTI9vGrlu3Bag0yNbbfuZk
bzqizfqFB2h7vFdlYSVwXplwdD5yTK2xI9mRUCiePztA8CacBQgIorAWi52DOKa5
dmdiK7ri0mSk1HXK04byiUcoVUS1sFNCqd36Gmck4lj3TLXy9RtOpV8yEGLo807l
Kdi70PceG+OUo1XhU1w7MzrAzByTYa2xK88K4P5e28MGeMtP0hOvn7Fj17iEomc4
Vz/hnuJ6fWkhYVJYTCFOwPQwaxymq76+0q8svOvX+m6pNGdSo1tnSy5TDuzkUamN
CBUMw421pq5o4j1ARbnBRRzOY+TrM+hmRIlPL/qbIApqQrnf2EWIEXQaMGqfv5/t
xunJk/H6BfIbhgvLPiKiI5FJ3fkrhAeCos7bnK+NhTSIiYmxTf8yHW7lrgDqtEES
+hyDlPwFRT3mbmpMy8pbiVhLX+UG4+iSPSVVeYxBoLnpBPI1QJwvbJ+lfE/GsuJA
/1fWxl6p7S0AECJ6fgMvaQ==
`protect END_PROTECTED
