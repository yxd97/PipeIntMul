`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JGt/ob/6xfE9vuplv/vQBvi4iKXkqtRaiXyeMzJCeoWmtvDdIuya+SzN6dK5iBtY
U+MK+Ua5xkGmZuGs3t0qg8qAkzKGMOMNTdVx8iACJJ6ONDj+0o7k8sG4YF+2nf5m
yRjvD+WAvcxO6lCFuVznfS57NyfnZ7G0QdMB7fg86v6AJFhs0HJnn+bp6BLV5G3r
UYHAGMSdmJfalk/1EZ1ywv1x47bmbAudAuyUxLw3ZUUAYZtMYpurtvX/Ijcs1lUE
SkiMHDzq7pmb+xhLC8WE+RSkMyCAjQB8ry0bFZzVnPElzB1Vq3xIbh/JR8BE2Dl9
3WSPC+joTStBlKKxX8OotsYJbcMSQd8oTDQXt4fcCk1xmbnmrtrc0Bx42KzZcXX8
XNkamOCwyE2WtGq7lZvUWFqmxdAaWW4cbPkbEajiQVfMb9vGGwUsW8d0xqgPaBZx
x7/DSCjsVCO5h4eSPedvsjpCump8mM1Iq8D+ji+xe90=
`protect END_PROTECTED
