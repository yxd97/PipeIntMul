`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYQQ/cGygne+eAR/7TKKdy/J7Unk7IyiXPa3mgpBVGaoWjPUI5IOB/dpt/WQRXP1
d/fXvKzs29Rsk8yYuHd5JgRRXjAepYgeJV6M6jTN4j2MzbjBPE+UYEh/30aSoMHl
YEorh4RiP+knfvnDnaqfcwbBVy6dH4S+NItz1/l5ZfwoDHtOdBrGEF4DlawtiDT6
CfMbe2r8V2CRkli87th+KUKnjR0qBr5s2u+avzLJAo6ctArGa+03Low2Ls7DCyw9
aaNT7vSeyUuDq3YikXLIJCKHD8EPr3PH+hH84ISSbRRPF2jyczPf9H3AYAOOtWaT
4G3AO8zQJEXWT2J9h3ygoxzSeKLAiaX3H3kmVhtN/P19X3q20orcvBW/Qc0AI0As
OAnbOCvia/WgIN4Pr2FnxQ==
`protect END_PROTECTED
