`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8k7DnbKDzaTUlToi/IXv3apfiv9Wn/6q7y6bBul7ZhRmqO+AqXIutQv91h7OHJJ
zCY2+53rb9xfP0sdmDhvKUu+rEhOV4Ztrh/BV9G/U7Egg/LvIoDgIGQBbP7dqZJV
qD0GfEgSMkM8RragaRAtioRnkFOpDHFGdry4JABaHOKDWANFX66TJSwbW42Go30q
dnVvHMgy66LmXNj3YToxy4Bo7M3ujDgLpRhhp7TErAZ82bYvYK4Psaj8kFr/swqj
lZcir54cyay6O5OPYhapmGeSgO4PCih589/e5T4cApU6rQquEquro94Itvd8gbPh
5CKN0Vp+XS6zaTexKe2RnnG3IjjTDxK+HlI7CABhz+xwdReSRG88p2HXLLQ7Tflu
GypGcO/mL0ySRXzVXMaUrQMLizTC0k4wX4T9SZPD+icC9SIPclFEgCq36iW3Bet5
WKmf/T0U8+kcC9h16nAHuhTaCLmdd50hOBrFCAq6rzMTB5PcSTP2pMIhGrJeJraD
GNpQHBz0jt7nT9IEQs0Gby20hOBok9Mh651v4oEUYDaQjx+pq0ZFvnylA8We50G3
SdcX/3G9z6MlxVXbTZGB3NX2p2R+bZXdsipTI4MV10AjX3oejkLg1zcPsg2bJogA
ZTzdTHLgIq9b0b6wzQsVG/RTObNWW7OCtc4vwncaQwrwL/V9jIwWrMt283pUsq+S
mj0EMu4wemMeDLTqbpT53r0OEEKpNwjtEgNx4/E5vpsnjqD0NkmBzzOCRl/PDIvs
GvUIepDrHS9QJtwcFR33uInzxm2dMguhuPYILR+eeFSxqdaqnbFj3nJ2K6NOm25D
5gpdYbKXqvJSssIHcecm2jLcgBDzlvrBV7Uo4GWNh0jzYuX3z1DE2f/3G3g4oolP
RJGmgf7ufsSyqShlJn5NRGo2bQZuvWJ4zj3n0WiBI2exCiKfV5WTbuJ7xUbNPvRl
j/RimOvp98RxoufHMliY6WPN8sHjIzYDX/fYu0/cL2DAaHv6hZhoFrbVc7a4wgix
7P8yF4n2VC207KpFf/nPW+9cLv+QuvLHWLL1Xi0lkOGloO9baJDhVDc6OWeeWoiD
WohDrcDU6ELNvj9C56l3ES9NQLLl5iQtJRW8FvxEp1gmHpgQa/uDq1uxrtXvrx2R
`protect END_PROTECTED
