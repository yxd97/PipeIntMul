`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A7uLu0XNFF1cFtjLnvyQ28eNhfeg66eXHnNk0TRQqjUrk+LxVFAqdL6T+uVlltId
27UA36CAVD3F0dDf0ql69DhO9+TaGrnVECTMLUZ9/CfZV68oj0Fiihqfq6nXWYt5
mYgnXW4pqaccoW/+tfMte1800NUBwctMxn2WoXhkg/w8DpluzdCOLwl+XF1oGUfZ
Ga4hXDiJkUpn8LOAZOTU0iD4Ze4CrdsaMznPCmAy6KTMDDQmtfphiuSbjYgi+Mur
9oyWRiFIkjZSJumpIjSCT4pCbpqzzzek7gXplhc70Sp0hwmiqSqGa1HdpGh8WmFz
f2W5eKnRd26Tztj/aeHcFtS7kcxOacNi75U2e78drzo=
`protect END_PROTECTED
