`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wsPCzXgVpwteQUGFJ+z3cOo3AyYUX8Fgq5OKm71mU6PxUyuOCqFjBk2PJ+psdcxl
CIo0QXjXyGaFU3OVK8uMnvbr6K0eJ4eA0PW/qTJ8cLrpgznTiLQlCcBafBkgMvii
eJNa9FFHt2QAobu4gzmw2FbnqSE0REprXAfL4168MlhK6YlN/u5SKHyorkLH0p8z
hcH1EFLR1wHC9pS8tboNbNzUkiFrh0Asmc0hkZpKyfmmCoQL41P7XwpbBw30zd9/
a7kNFQJfrChcddp+NcNTTk+myGEpIDraGF0BPFmMWZCVmvCas5sKsh778anbWd0P
bQ8DKnp/hjhZdILTah5BD4G2gHXVWCEsUmco8Qsq3cyS0+pVsWx8Wo7Ivar2ahY2
`protect END_PROTECTED
