`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nO0uNI7PMQLIdLUR4f+iWaz86r/ts4bWUjy8g9X9PcXiQEI1n6/IgJy7C53DqdWj
sY2AbP31Hi7QdDc12uPjhRSJB6CeyWRRQt/VuUuQijLeLeJB9D9wzGCc91FgK0p5
mi1kQOF3/r/isyKFt/mZqPT3BJ6pWmwX7HKuwCBBkdKEER9K+oOxwk9WygqUSdS6
Dnwn4JGwuY57BpzfzV2ztrz9SzDAVS3s0L1iNLEZvGLLe62L+trkF5edIdxapnEC
2HNkfWzb+1lYeQWngJ2vK209Lf89+KEloxnbuhWu0z+0o3Ugd0iSJqdzvOPyOWB+
/TNluyZbXZa7sXXsZyamfEsBbrinrExfWCJy/4GBkCfsoLsI62RmQXSPGE+ePhHV
8G2Lxk456YyCfD3tcrpvdGcJ42/WY5DJI0DSx5FiKyQ=
`protect END_PROTECTED
