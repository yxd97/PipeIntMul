`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Upfe9fM5Z1NOVDLNFwHwH8qIbM0s3FtI4tdIBp3Uf3N4BG8ohDLU2CBbLjOmthOl
kDJy7IN+p2PeArxieKNk0ivFly+d5wSV04IiEQwktMJ1KGdEdm2UZ9U/0Yo8e3sS
cqrfqnobw3y+DXjg+w/KVOhpj+vtA0+ikOgMZTZcve532Q8G5OXstfREO2ytdvie
AGw0QvUnolbbEbLqcVpbx9J29Ted+pvy+z0LOEYHyVrr8aac9F+y0LWWpqeldfOw
MCMcos2PLq2qQm8Bs93XoJgE008PfIEzWvbWmPVu/2MQNvGHyyql1s5OO7Y6igVC
zJJ0IwGrPN4HfgaDbkOWQpuLZvgHl/eJOEhlsSIzBrlSUy0OljKkyApRvtCTIW5F
bJI73is3Uj/gDVlmdU9MkNNmokz46dE7N5C2xsu8aZKFSy/0DbMXxpItR2+P5FT+
kwnRa72GsLoz4bODhMg+XMvgfPxwfxKPf8hGKGu7Q1Ns1YXjz13rBpcs62FoOX3h
Ot6JDJuXK//o+bcUD3fQts6+ggDFeeQ9zoilSwVOaQuouXS62znQ6cZzabFpoaMB
H4cJS8hxoMMfz/a7OrFPmQ+eWkqjBK4bvms3OGnp8YcK6DQ1A19gCDNXueg0T9Yl
ObRhIxxZ9t5DPjgFDFfdKLJfeTAkODJqk+JyKSjLgh7J9txBxvKUC+dRRARIkWKM
zQ+QcQYaRYnk5XTkeyKl+NRoqh3gRg5sXpz2Ag8fJf1FKw3/lYLVJLLolRC0/jlr
iRadYNPTLlY/iT3arr9PEXfr9TAYnWeZpTPdQVuV1s9SjCzBBC8cEHYo5lGlvb12
Mot91HW6WCBVzELLYtIpDv1EY0A9wrjVOoXIZ4WACWcSkic0B1ZjUvbqxaNwizTc
pOQl9GDEZ6//78L3GNGkPyHefFYwkBQ+eGAE6+Cl6lZynmzLyPoypmsmX/F7KBwb
DwF0U7noZDJAGnDsEpv9Fbp9GzJ958v5tRRbS8LhRLlq86eCQCC7Jz0g5TBARuLQ
`protect END_PROTECTED
