`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdMF8z2KCASUCigbfm5VtQbE7wQbmeDCQ7JMsxgn+QNUGOSRxYd4wCaVqqcKpvwQ
t6vW35doXydQC/vWLQaoJ959qjovcXZF6X60iFL/x+eZOFeREmSPE3HSPthBwfmO
Uq7g/CadRULJmyDI8LnMFB03KXcSjE0bbo4e8cjooiDGHzJiamRuXlAdz3FsRXC8
SeXnUsCbygZBpEJLcJc2ds8507JMrQS02cRE11mSiFFLKCoSY90bzHw4vpDwl8QF
aY1ojROUHpRvaFeb8ig4hraYMi7iWQVPIMgi4t/u0eNOLMil7Qbv2waY2+t0LcR4
pmefts+QfNqyhv1b42t0DvGEmfP6o5TLknKxDynhVoEVVmjkDZYztiuWSHjT2+Kz
eM13k1+g8PihCO+clC7xMA==
`protect END_PROTECTED
