`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRd2Iu28RCapKzF8AUxVT4gHblnGVewrFCP6Bh5Tk2MXuIlDWgaim+QZc6ds5vJE
yVJuRBSAGQy5qHURX+LSCs1ifRDlGWUm46WJzYKFRzHX4EZ0uEGf4Hn0Z3nTQ4Jf
NMIkbuinw5zgWSYFTzKA/C4ybwu2KIc7g5mcMS2aKOK2BHqRve7bhSUVrZg0mwwl
v2TxZkgthOos0Jz4XgryvU36vytXBRAwb3xtwgCYO6LGE3rYm/SblcRoFc0IQdRX
cP4FBgMgzzDF/6tH7Zxrr8P8RDLqqIdb7/jgse+Io9+lpKS+MeAiIFpH5KTZHw6+
6OM8qFN67n76WpfuE/vPeBpk86KVGGEOD/1zlEDuwZC1/WvIa9zKr6PaPX4KK/2r
MOIfpvx9fuOrSZQHfw+F+32a0zNpYNxfoL4q4178QOo=
`protect END_PROTECTED
