`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sE5e05P9aXhI9tkBf2YFxMzisCXNDR9KHRIMbEFFg+sgbv8g2oj5Twpwwk38YD08
k2Z0vpGl8Jw8yz1l9g+OvNUqstmvYWv0cUompIbWnhtCnIh6bfdk0NWKROZPT0eO
5ehQp6Y+JncC2scQ8vbIkjT021zG/BDp6A9ygjs9M02s97VGHavj1vPfpwP4gGGq
amBB3f1hO0H82IHHfRsLtzD6xyJILZ6X2EwqQBPH6rC+g61CpqxZ9z0b2r4GVWTh
UcueF4f+qHDQPPlNjKG1Bp/EwwswgUo6yZAtfLGQuQJsA8EjHGke4cV3pF6KNW10
1Ppede/5MrX6nWiW3MXNkvHAXzm8ZOJkQda+zJmiSDw8Rsgstg/iGQhxsYOxuhPR
dTFsBGeUY6Vt56Sah/J/p2j2mwvGaQXyJF3Jc9gfUTnXEDYW5LEQ6AN4Nb3XVaN1
IqbzM28QSv65TS2WPkRsSmCh1sfd4c3wxAosDo98D1BKJVr8gniVSz/AhvM5LHKb
k+8YjNSvzJJziaNps+HTZDbd4+NAGvXjSkQl23HnbBDdtJhb49mrf66fXjHpXCcp
QHBTmPIrfp5dc8TPPwKAgDw15v+hE/V7rMDu4Gjl5rsJsAOECft6ven12NoXIZpM
VmBHoXhPbQfRq7A6CPjZhA==
`protect END_PROTECTED
