`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhA+1vJi7wbFG1yMnQQgYTzpVCoKMMO4W0wKWihcZHHQPW/WTatNGdeSDJu4rPgb
KY4OVga9ByXbeM72lvk1SH9xgHADNoQlk8s50jElbwB505ZTxWs2qEXG3M3cFAAb
4yarc2zO8QUYpkmVyey4VeWMnQ+1Qt/lH9vrpeBMaKg6PQAP3fAav/CnhpmwiqQF
CRITPTqYspSdlqoH1T4FFnksIu3H84an/xQIRnD2UwXlveJWPER10WnHkbjbDV5B
BLgNQZk/JiDhIvVtqd1F8oVMMk/AdbMEtnoTcl7k9lKif+eLGUViiijPQq9wvSf/
JiePr0F9CMonqCEW8rTxIBHw62bEWOJJT7a8gQ9SihbvXPY4X2LMfjiTeHiWJqPe
4kqYiNGyxSGGTAA/ry6n00xsAGc0hvQT27vU6hiWB9KCKnDDwH/rbbASp64uWbtA
ddT53YN1y7iE//hR5K+0RHnV2+KpHyu96opzENLvm1QbKNMEWc+quBvzPYdW9wdj
5TMNIu/pkDfkwExOM7ZdLQ==
`protect END_PROTECTED
