`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWTjdUNOJiTN/L/6DHhf+2MvWsFew6fm4UotPfb6FK9a2H9LIlDaIOz3JNh0xXbS
nxbF5BUtztJ9dlBOgFvfO83O2qW1uWQ3YqUcviy3MipFBrl4MaEzHsmv427MBKwH
ALWmxyP4nneqRkcu95clOxcFiYmnPLAZZ/ZK6b/RqVvrF44wFEoCndmmRXXY3Yhu
8I52whA+7YbKzUM0x4bNFw6P0oI8KszK+CM3HfF6Omv2tj9JO61uLyojLvoGPWOn
yqZROkMimNP/c6ErrhRN8WLHwlHoAi9XwI49Vf6KsAQxR+yv/pApxlXeniynO3W0
w+R+FXxiPoDSeSPHPRgpqJRVMbYOxEezDrrra7Ro+QzIBKKvLBwBeUcrUrP6OE5+
`protect END_PROTECTED
