`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaPG5DaEEa/e/6SmV3TdOjBADJtpRKtD2hB947xi6KBUzWqM1NxK/Y3rfeHd1Gto
ATo9XYPyLEBvfQglTOcDrXzp+Zj9UapUdxyWKcSNopVtO8xgW38mN/AqvlNcdqUh
ukE5bDxtzh9XdoPz5lAL7ndhgt7SPp2pW9chwGF32HWdDHErNGPxDWWxxG480zZP
EcMlPTM1/1OGgBYGDQeTn3mF5AkU/WbcSrgL1Wzm9ujkbSa2jqWAqQp2qdAHinme
/x/LZ8uT+bL7errORL3OVRk3ruCvHBW82pFXF7CCkhxGE606d2WSH3nORZJ3pJW4
hdQ9j+OFBcZdbOUaURiZILwWYNmy3gR+hso8OUOCTwvkyfJnPdgHqWj7hbFnudJY
OwV96ygd8MlE0TecTo4dwuwAA+XPO7VbJX1ayodTyJ1LSjrADjUrPhkiJyowbZEV
ZsJ1yZe6itLEvSR7p+UrjgLOiO4yTYsUDabkV2E40CxzoLZk4bDCpDh2tyry+Qxa
hTERg64flL1++PSNdkmd/IvLyiyidaVEf0gGaQXysk+12mSQQAU+Rdnrf3GmWRMQ
yDkeCynOMV+24gT54zqPP/HiBj6k59h5G2tolVOHVNLM7lqHjZa9wD3p013b+dIz
kUUFkCIBfAAmttuBVpufZw==
`protect END_PROTECTED
