`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THWRabXHZfyYGvOHew/0xL4q8PzUVRrPanutgBtIBR5XxV8RIDtwYZv7gynB1eW1
RbOxcZyIChQSFW50FaPHaINuh7FkHI8olN1WmF8JRwqbH73miZaUlJtqIWqdWniy
BD2t+2BsUa9uEGPBfLSaTg/JO7ECjnuzHbuAsSMFBM7fhBOnt1lZrOz6hw36LudN
1pxJX3RUcaYAI9PEXgXXpaMFbSuRy/uwkyjNJpoK3pIJAbe8D5jb3xtmOOW/P21I
G9xg04D7/FEDoKCKYKHE8LnqB4RiWkO9b8XRXwFndRMN3BDWy8FSQhCSB7p2z1Nd
7Wnt7vPyJFCBEpsyDPdaW66mSHqqsiIw94CjaWGvnS2fa07iZhWkMcnDW2+hHBce
tGgMTcWyg+RSRrz6pU1hDJ/dscU3m9EEyoDG3ZkK+w9a4Q0TdE4ksNS14X1xiirG
dNEDs6tvE3B8nCnIJs11DzTlIGIGnGAePS0Vr0f23QHQgPoIFJc7i/2z8uzePCgP
rFY+fxX2drAAv6+uCFNsp/kCf4MD3dviHkuq1yoar7r+DXiV0XJEhtTEyhvh6lkV
QXfsFHV25iB+4/Byk7X/Hutsb3ZIq8HqicbedJSjrURoumWgT4Dxuq7V6dAOAMa4
GlNmDmRJMlzx7HKkezKQ51GLMKQCXNzJ67cuwJElrYXlkgTA05cEa1bLJQODXZYj
gVk/RgICRPemYCvu6cpd3KQrNONXJhor5eO6k38P6+PQt8P9kJ/EYMrT9MCy3E4L
yQQx9+fChljktSbBUH4A4IL6T4GLtjnDxFsX9IUogFRs5/GZUS5r+ODVCjxnDG+f
P4u3Tb8fsD+yS3uEU+Sa0A==
`protect END_PROTECTED
