`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sn6KgROsZLIUhm/QIuepLX6vHGWozM2K17Px1YeMa7hqsmR3P1PcQ9Ha/Hsxbskj
OziCh2fJOxUIMZ19FQ/BH9LJdoJa3ZSKmPRxSPk2gSUcT7OEboYws8xFw9LSNdGZ
6ckNEgC5d7S9IgJBu5M2b1QLUJI2qH1xpZ/19IO32upYG/oktmEcPN0oGC1t8b28
4lfhTYzZ70dZT2qC1lRFhgw4xVUjxZGy8s4ovu85abetuVZ05JjPdpTh6iIIwECp
IWs4d5OXkwbSjuHvBL31xLLWcgEpb4iDGjFO1Rvl4TSCBgtobuuhp0I9lWP30Hp0
alyd555bDyYo+22iPIR3WXc8K67tMDxJqaLJ3W/KLZBCdHYRTfdy69HmsCkf7fRe
nb8Z/pBjORe2Gj88h89s3clSweuANjj3Qnk6pISQI9UCYUCuCO1GciT40HBUW4Nt
`protect END_PROTECTED
