`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
03mvcax6WO2PK3TdFGC+/ZsBROsdncGOITmhzQQ/F5b1C7n1bYsBUCQgY+gMQ87P
k0/adYQ+B3fFwDoGEi0h6mVyR1ZFClHDvo/gTBKuVEM4Ze/nY1LhAIO60XjObXEv
OHC1OBVsErcvQYbFNJEB80aEgBTZFpzDuLHwsIR7kkN64QWff6pPuBV17zaFFCiQ
y+eKrlUe2FYk99Wzrig3IjOQVXJoWfT91eKZb45947AQ9ygqzitG19N3vHEoC9xk
KwhRgJBSWhhYEVqRqDUtmuEwNmMZVN7ynwK0xKXWWVe39XoswcYyKNTIoRbxDEia
GoiKZHyCCmaBYO1SVE92GFsK/ijZla0F6WHa7MXXHhs=
`protect END_PROTECTED
