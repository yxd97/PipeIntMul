`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbV8VlWM/MLPXiSRI8tFVoQETbNm6y8+PDiU6dHmJKi42KbfaaaaWySAmQISIMG3
hseOmf6Iumo2NqY1tPjg/Rl5Q9qnZPHrrMQjz4hIPvo4jwwu5tE26z24qyRYcEZm
PiMCFVu844rgTEvKDQJDdIzk2fYemAHO+KdV1nhjUkejcIk2+Wg5b030wsAv2kYQ
4S47LazNaDncZGvongzXboZ4DXpcubcq1KfhvRiW0BsC61ZtaRD6DaOXHdVXgJiB
SNyIdorzt2HoilTzqE0XYP+PaH6WXJKWHGDSoD0OmZjoXSzQS5qNT6UJOclqjN/K
FqbZZjrfoJLmo2U1BvcArkhcF2xl/HLqhMZO/8mZ3J69VNd9jM39JLYwZXm7iL8v
ff2LuHTfYgEdkAGn8RzzRpw45EcVYW2PkNQAVULZJiZx8anpYV6ewPG+CyKMqKkE
WBqPsh2RRRp3eKnGeQ9Vzg==
`protect END_PROTECTED
