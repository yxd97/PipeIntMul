`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zRyD60W+2Asz0Wij27bRtZfm0stqL78XN7Sed3hNGWRwVMiBcDRoFXDLHnmtYHwu
n7V+unHSeNAumyTmo2m+fCMxkaFdcD0bTA/HR8+eTzbl3kmdPVXnzBFIB5zK66Q+
OQKntx5A9g0XPsG2f5dKMilM/sNhIlqJ15XpNOpYzAaqqel/1MpPLsm9o9xDfXHK
8BkBHGCIGEJ7CIJLGuXqMOVHe35cv2yIoM03BYgqcU/VAlypyV/rv+nsHP+OEfwm
LAiEfF6QfrN3GEOk0qGz8CZwdk+WJvVaaeXBN02/1L/+MDtDD5WdcIW3x4i9ALXi
YbJnymKzdFa9BPKx0+rP3QMfFqpQo2kqGtSQOH3FEsT9PpAk27t3w3Ola7/ebD0V
Q04IrCORe/piVUZ0dbd+0nHJ43OMjLKb1nEFUdsRv629YQPP+Zkn9NN9VIFgkMHo
`protect END_PROTECTED
