`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u52OH29N9kyzqSLiFDu0gnRDeIQdsmys0yWGmrxqTlqS/yZ5bkkVSFeSmtyE5V+T
eHHku0DF5JahPbQzDN1BlkpSwfd0u5WHFd7srhCqTjJJMLtcM00T4XXMYlWbP1jb
yMZ6drhA1fZRrQ54JtbCwQ==
`protect END_PROTECTED
