`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dm55opX+fySrFccZQc9djGghwyB+2pSXF5QkrE6a0634MGu+jBCvCxWSwTndoR2O
83PlBxbwcMfh+swmNPtf9yrvmYuHABI1e0Uu0nQlhi2/Uwa5XZbPJ6vfGoJNc8OY
KsYPTBaOGjiE1ItBVhPhsbC7T2eJeCo+WJUPM+vYWZy3XQdF0vIN+F02ecU9ZQPv
6PDnMpH29OaNBglJCck9O5mJv+hbamsWWVe0xusEqibNnyQBZffcLZKZbk7mRi3m
MQ+ikl21H8ZHUa+r/TuxnF6KSNX/OIYK+EursFfpRgZxQYnabzgG4HNJJOjWTzol
TboF4vx2btQAZ6bo7aQQpdp04dofy8pYAPFNzXolYNmPDDb0jkPUTnpp3BC5nwLZ
vPekgYLOhApNzChof9xvPU76zU0svvMrlhLL1hIC+iQ=
`protect END_PROTECTED
