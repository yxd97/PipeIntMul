`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GjBWT9sbGK27T5LjcSNhsB4FcScY5G20/0hbD7CG53cpZ3KeSiAJjH0q5NIbGIIM
/5vXsU513d3oyJj2a0cp3qOAfg4ICK/BKkDf4pR7mjbpepaXlAr5oycw3wLmGkFg
ZFPbkZ0eop8rPgdEzHf3/qsmM+8W9TpMoSyx2SRoWzw7uCXvUbUfg1hlHjJbdRrZ
kjnRJLjtM+CwG5y8N64s+maomG2jF/ogFC8LffzbGmXc42x6wDvwV/U1ATO6VIc1
rMLEsg0SkUthg/tam7wn4FSq+xfrUqIkBczPsQPH84SIwOm8lSsZr1FE4p3eZJNT
d4+yi3ETUYdWEvy3pvOfJuwq+rW/pJ37QNBbiQutl8Fq6Bj1pq+7X02lbtOcNZ7E
aFvR8l3XZe7fbOMhzcQgfpCYq6uUYg9urvnQe92J9jrlMp0yhIc3/caEu72b5nZZ
A2X5Po1edguHDiAHbMEah2ZpX5/a84zP60bZ1MidWq8z275XjXxZYfDAH78ze7Yi
`protect END_PROTECTED
