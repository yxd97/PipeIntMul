`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uaw4SPR2KaR90Tmprdojro3ygZO6nLcBM53XfudhZSaMGb00Esj2ibeQfsMKLCRt
X2xHUfKeyaLQJMVLhgsBkd+1k/m1dVbCHz5YJqLERAbFYSUtE7tF+DwbaL9SFpG1
M54zA20XED57eFtmBUbm9Z29JyQebOVhFXtDpY6pf3/FjBKPs1v/W3DU66lHego6
9emMiY92nP0BZ9qriXoJMQJ4IYwtzQSEcHw1dy0d9stjDFO3kIykNn8L5t9RmUQj
/d9fD5tGe71tdbq2cHZ/L0Ifh/IUXCt5421dKQxckL274xFCtOBSBstFd6BBuQok
Uytxd9hpH50kSnIuKIMqVd8cvUrqXNtJ7+qi1SFeCwdDk1pqGyaRvarRfTH6lM8n
pEz4j2qhFncrBwIrPhg21SFgyFb0gVHAxFSVNWLK5wg=
`protect END_PROTECTED
