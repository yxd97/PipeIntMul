`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0iN/SVxOtp2ueoMHcMbqjPi+Cx8lB+1rkUGDp+GQgN6waE8WVYjXWXhr/kHXjY0c
ZFLMYG9B6c4aHMycgvDxezHp/4nomjWnZyDoHsxm9HMQPj06SKddUMFhy0U4L9rJ
cVE9L8tjAKDD8siBacjZM47rZ6azl95KjpnLSEakbBar4UhIXM4p7xzP8ZX1unuQ
g9PD8iM1w24ToOSVDafKV3AMpHvKBHPZtweV84HxqjQcEwqWgRN3E7BuHD0vvtC4
D1ltF74UivnIM1UKP2YWckrLZ2Js7tBi8GNWX9HhuQR6SYBTv6UTL4yGmwJwa7t0
L6etdpueVwW4ddr/gco0nj915yHGcV4VT6wXb+baEzDy8qitv0oEbq/Vcu6JE/h2
cyVaf/zYGqkMcN+w3WWahWWbfl1XPmFP11iwx2YtJ31jvJcuUIWRD/XqN4nsRkEc
JptBOGcps+lU55RNoKFtlJBXFd5TuhS6+TTVVNHufcomHH05icL0+vhMQ8AM1bsF
6WyABpwhKJ09W/iqCjNB0W35YhzVwtUgraEPpWmlAclFPnYXRYFaD2NcSBTqV5ym
TomSfCMjk3DS7G8MTDI/oAEuXQhSWvt9leo27iARMypjxVMOLSkiHbfIjLeNyAJK
gmPsnZrEQGWUA0Je+4xhXILEbGb94sHJYUJ3ReYJPICyceGpVus3Q5S0v/KHjLwU
VZzc6K9MElZb2wOTE+8H/Lb9vGYe0DQLbfP5ImLMBDu1IrH1Jw3RExlMfejdhIes
RynTAh2tsqKOZqoBaQSuU2OPgob10CgbNjK2TpdexoshfHZTDc306X73qz664mEq
XYS02p2hyURZQyqwyrCcL0hDhJLMp8Y+qwtud9WVQ1+zYQU6jRau8CM4aPGg3Nhp
`protect END_PROTECTED
