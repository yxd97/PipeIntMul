`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pUgr+qKVm+9/FGnKgpkAzORW2Ygh+BqbEHIx24ImP/iwfhMCTBvwPiPKaqCGWA5N
ZTUueENqW6xyZR2bVtcmXlu0QDWGLPPOILavfGX90Mvhh5o9DPsUOFTJN2EQYW7R
XYAljnML5jKdB/RqqDSorHAql3d3WOKP75VNooRiutFllYXNIFacJCIzhlBdhxa9
WHCSL+x8O26ASZEtn1o7g82nia5CDlsml7pVD5NhI/CD14kWp/pJkwCcteC0+70A
Il/jOqKmBjwVcgC+iUWMfgWGqUjif1+pI+Kj3SVGVo9pCkmHtUIj/zHLZ+PY+fI8
`protect END_PROTECTED
