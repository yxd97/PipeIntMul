`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVuAXKlA0DsE6Ralx2uOvYlt41ohN0uGsTdKovMNlQ8T2SltXz4rxJoRMtBZC5iw
+3VfrD959lY81d8jf27BROD27TVqEbFE/7JIlnn0ClaTLx1ae5IHkgRlumEQF2tc
Md4LTp1H1ufpcy3foAvD6AkEiW5j6cU2e50I5wSOUvLsGimivBL37JEvIYhG+Ryv
0ma7S75jLLddXemVBGw92QDiDVjj+AfAwKhtrqEfjBo7ZJ/9nwrGoOw1tZilbIDn
7fx0hLhAlIy35vsj4Td1eKZ7IRKWLWRWbAJ7rQajGyPevVRUvEy07HEVURKXJLFE
Y7rV+sqPgHidKx7fNI+r7QteTgNSwsWFognABDkGlHjWnq6gFJd6a/TxgUhSnk9A
c/dN5uyxaFDA+WbU92jkvKokQg9MahMJYhZwYYDPecWlpjar1ETf6Bc9McKsEqBM
braUyDpt7sqLVcjQuRp6m4Bf/NBenjWNBarQlhuKP8K64yKdwJ4SfXFXbVREGIS7
6cybv181YC6XJ80Q8k5dpa/GJcG4M5Mn3t2RrI72POz42urtnCs96JDQWFKc+Rbt
YBYqURKsJFdLEEsZ9a/UUGwNWu1YO5N8LKPWCYWiy2r60QnKmQZS6xl6q7cW5qd1
lTcIMCqMc2CdDXiKm8YWq/wDezG9EZJ3n/aeEWVVD820H2jZYwPuKMFehMG2887t
AnK63tOsam0KCY3akDyWTMkg1kbS+JvRUMeB7FFlFRnavaUt+sjPE5faAOFwn0qK
KJjxAhrkmL1ggMBrWCRY2txiyfXgUdIjUDm8xkuVwe03+12M7/YfXMs8RHdNYuqX
Wrrz2anJFYO+yExE4zmdCSLFaZ2UUS7C52WvM4uNC70RDtv5ZW0JfMW2eMR4Mwf6
4QxKyh6uR01p6tDMteb+yQBrTGjMa8W0Wb0Meu2X6/HlogZujmBbwzxrpjCrrHX2
u263pwzKC0kRSVQNKa+591heoLDSM1xFV1iscsOFN4wFXQDAZEGoLk74moG6TbN3
EJntHH7UIyNzkyEmw/nE542+sjOR9+mhdgbnreF59rzShx6tZ6J0oeYMjRKrk3Lb
ofZNxzAJMU8G/PQagCpbEsSt8ZMv+Oir1DhbnWaz/Mdn+3X+4JVTPVEIkTyA2ZKM
6jEN+dE7/wrigvuBWFPTuIZ3pmQkaJtm/GjQbA7bHYIu0YULG0GL5CLvjZHOxZg8
tlDu6Hhs6Y75bJzOkeXvDapD9q5YjTWrD1lCk4hs60/YF/D1Zpk+KwJTZ6S9EIFC
bAXWQp1YYKqz5RmeFyNXB1gh9WilL6lwE1tCtA3bnvc70lXnBdbBnp1M5VVQRMeU
CjrRG2HRAmFqGQmYLgOn86/PaS+bwFU3Ph5iHG7Ol6P3MVW4VV097apcG3YV/wfF
AoNyfhx4dKKJotjFFiIveLqHPHvyVlO4uXnUBEINIS0Zttvdd7RuTlZqzeLIQHKN
L+/v6FqcufrFtHiRyawRlxBmSP+s5dwGfkh2JWSqNy+Y/9EobYCa+CbFyshdqUd0
0gJqAF9tXFe9pflINsI2xTDc2f44/SWCwQbUp/wf/k4MWd3URBi0v1bzlDkSU0MP
5VYB4LuniHaOEaBzrGGaU8Cq+XrH+74tdXrP3XTGxwdk2JXjo8SRfGMZFs/jL06Q
JAAWHcAanowpsKHC9ff4uWTYltUo2q6UYGnilBO8JK9BJEsO2cpbBCRpDBwuG5+j
kH5ZQwUCOH+wEcGIKpfC0+sMBKZG7/GIh/zERrm+Ega1taQr+ZRnQIWOaioXdpHl
t4nC8DbU8To4WAu6HHU3S5bkpFSmyP1cTBnG0Clbqdyo206XRQOwUDgU1yXzI8hx
vg+Kap4JTIwh71xp6qtIrxNlPrggR5GOM0y0QGHT43JqZTxrJwDkUU+aee4ofguW
CEG67EUssNH00f3ylljrJj8/uJQPIwZODcueCUAEHtxvdyCZlQFEgcPpqXhay8Lc
zIL3u9YwvcXBDGxAXrK6XKKuiMzfom2czbtT3ONoykXXMkWg9dGH+GLE0YZDq+Z3
gTdSd4I9+zBWyCN9oR0BqUQVcHkJEA4jsa7ed2zjS8k=
`protect END_PROTECTED
