`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mx/RvMSPm0rzzdM3bjUDBYFJjxBCrUjnxBeAZQviwMUWelKei/v4C5ue8xLoSmqs
oLPDs14rLEprnwZJw71ZMKtq7VuxCLCRzHHQYEJtd7D3Y/V2zUIbYm+PJUbOq5GL
7ocgYv1qjZkmrGPW6E0v3pRko/e+Uhtr7eh1RkFs9xPAr91Zdq3iEXB1zsH0o02V
zYqyvyyhzaQLAY7WN5yrWUgElhJNhZ00GEBMRadPSE55Jc2hoHItbsU5202tthAz
QwqIEt1Q+OpdzWLQMgDLO1fZC6kq0ksZd4t6kZRnuo7pOuIVf9Lue96vkyhp4dce
2qV23gLMu3asJjuzwuj4vSa0nqE0dfGtOKmpcDwG76+k/S84Fr4SNCaIcFbT8opH
czWCTFkaSnSFFlj1AnEpfGhzxcd1tjxZHNto/jIWKAbvyBOBe5AveoYCqhREcjy9
`protect END_PROTECTED
