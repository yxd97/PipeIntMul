`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6KC0p+Nwbmg0zTzSNDSWyJ3EogeAOT/ReJvtd8Q5HI46inMVkVBFShaaEnx/4or
JPPs4poy6Of3yTNyvEmxVvIp8kGrkc2YrjGlYAyh1QuHyWXwRsbc8BJEehzjo/fO
Be++rdZ3iFDsNwxyeF1ggdNZKWm7mqEQNk040m0pOuAZuBd0JLDfyFgBV2Nnel3e
Gwwb/F+9guvtj1KkgvwAlKK/msZbJRZW1trSW/wGaOaT+/kLn7nADqCcJZ4hrwps
3HGa4K6Qkecao6/5QRa2Tc0HkUSOOQhQeLJhkKIwsOznCLOR46ahLhX7QUNOv5OU
TeIquNEneIPP47+2x6e7dPI6wLyavCcEpMzAeJ2V4FA6jEXJWVcUUaiITO40fs8e
pxXKrbBKsNogx8n5vv+lu9EUbzsZREsor+DEH49tQgs=
`protect END_PROTECTED
