`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46DrKrTbMFHq06wHcyGnzmxz5+esTufIRoB2L8cerpUvm//UsNt+KEn3n1ZfJ3dK
1YJVGfc/8k4bbFJ1XaJ/An66ceSZGloMz5+GD08ROStQe8O3gMNiawIFxQJm9SQu
VWrmMzDWLRflS6G6panD/KxCgrajLLwabHYHoWoMeW46xsapStiihtDGAWLNlcXa
u/sN+TE/83JZnuIaqcX/7nuewSyRMWhoE2EX3hzj2Gjoj7Q2KwSdiniR+qD6Vmd/
uB45wdkYbkz1F8RiWCewJnJrogSzBQhMYbigkuUYMw/86CUCrwg0i4XxerXYPlVL
p8PKVn/KBZOJL8eOGZbvCrOKGkCHr8Y2bzecRuHMk1hZS7ao537geuoBE1FiiOZK
NqP95R2F1jVnlgozXYBFRZMrdWincbqZgBCHj/a4iqaUHZP0XZRhjiuE81wA7qN1
Y5uYn1jm3HIulzHQW3hwVzzYM0pBHh4OxJ06y6NEVWjsfJQ1oulED31i6eRhwi6K
ZU8GDerJTRo2/8LHqLhTPgXUvToF7jt7/Hjcbncp+xcsuIoaKuXuYwyUHC9dX4WG
`protect END_PROTECTED
