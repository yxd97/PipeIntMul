`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tOBvynvc3OztdqBZqccceBAoBt5lzvTTU5FUV46BbEEp9caG5IAw2lJ9VTwtEZPC
h4UdYxotEmA0lVuiO9XD4ErnXVYPCag8kIkJjqByz1Z9KkLaaQmyJcQrIpTPvd9N
Ib6lnMr3LzI+Gf9dGAuhoAmMzqXPhKnGz6GGrZMctH1REoPBZDeCmQzEpxzJj/5v
RtilhkIQ7XP602iAwDpnHP0s5VQOufP0VXcfchoES4OxnQu5/WgLsJS7lyoKpqax
t4bZ7QnE6oqhXg/3pjSFml93qZYvToEj1HH4b8oeHe3heJ58LH6h2r/pfNYu492F
T1l7URsgTtDUMbj+J/kGMcC6poQNFf1um+G8oSWXnAussW3BfEzQD/T4a14csyFg
vcOZ3TFmKd7yrtbW9Wz67cR8unE8XQvDM7kfL3xeuUU=
`protect END_PROTECTED
