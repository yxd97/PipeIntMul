`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n73lpWXXOXyYC0k9I4PS2Y7QZrMIhxhZ28q+SQVCowg2j6s8FrDazp5sZ+FOt5Io
Pp/umf4rELCXWdisZCgQsW9oEI33HrU9zAtrXsmxfUt/ty9QY471C4x6AM9eReOv
n7fkzbAx6eyy1Iz7i5D6PE59bAIQYHA+Pu8suhJyS9y6w2Vbt5wR9j3lzUrDebwP
crvvTPL2pEMAFHAKokGzBhYufi6HZ9TmR3RjWMLEi2X8jkmcGBNlZtB23+GbMtqr
M5yF5l0FTRqepmBhPrx9TdZuPB+0oIFNOSgNi90serqpkHXWLlNJ3fQtxQ/mA7sI
SXHiIbM6dfIUQ0Pqyy5Rozn7ywiIXHuLhZFwMYsz1dVeSjMFPnCBPIMtVYfYUATH
U8Z2VHbMs64DH7oS83+oMwyUgp4t/KMcb/7UaNgEg3245iuX+HyzXYkvjnq7X0qL
J8DW7PwSq8MzGO8QWpjoWnK/YlL3AI/ucDAJjFx1zS5WOnNUpvdxCm6A6ADtPtrv
2myCyTv844ZyET+oFxvejtLHfSroQRFmxXIsXiQDNDP6IsW4u+3nd0/DGDWtGJGl
+YTghxlrfJJ37sxYZiHS9cEv9RlYX1IgJyjwReQesqvCmLSENSUyIQ1CvGhR962b
+uLIaY3dqhacApuT5BWi8O+olmy2YCfqhR68WpRyaovSCH2xB4hZ84vJMTXBTZKC
z5ES9bOHukE97DCHMEpmBzsRfJNBzcp9lMK1q9PAG41WhHlgD8Ukv4k6q8BTI2XD
3n2souZLhpxXlq7idO1U9EOpQ+HVhEs63ATbcgLZoCXFeq9K4yk05rdJmZGN288d
zjflLuzATVhsd5Zf6r1zcQ==
`protect END_PROTECTED
