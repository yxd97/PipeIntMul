`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d881qrTTPJepwKr6fcHqZ35NyJ2kGAXmTBZ71KuXxzBjqelLJKu34Fm78Y4Sxbt9
R267G6pj8r6c48nCnP8sd2rwdetQaA62l+CLt2cQDkiWoAXVKRQW7O4sPnyhL3AK
6aiFbuVZBYtQiJ+le0RjGNZfLbmaqX4PpQwkVVaW5sJPFfLUYKvOx3UGaTv1fhhJ
qpBdmD033vYr5PbommSUqq/BqptihcfnsAIP05+9O95H0xL50B5JmUYhM8ojxMkK
iA2uk14wB2Anbl98gpR+Tb1r4CIqEnqzVeOvllzlQduXu0wM5spw/9n8YVXKjdDG
Gsj+12aBLF7tU3tRbxNABx1UC+tKReggdNwme9wxilVm+MHehy23jqDMEuzulD3y
nGMQc8PZ7mVDpzW2xM16cupxkIQ1CO1UQ/1CVdrP7Eb1av0A3cYHpGB+MmxVGIT6
mRvTAQwV4ES2NnIdd9KWxJ9tRuv/LlUmqt0KOc5tNZc=
`protect END_PROTECTED
