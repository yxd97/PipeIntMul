`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYZt5jxOEmDAz4OX/rY3QFgAtS1eQYnJRxXNBSlFcOh5ulEJjxBXpghZp4vXCFdH
5MPRR6nRDjTqiCD18MXG5gOPZ80Hqi1f3PJLjc5PJMO1UOXDoSro8WRMDVCfAHCC
PVfxh4YOWR7RQ0F/o9vZJD5rsqcFYerVCvvaTwx6GqnTU6632ZfrCLidA5gVUF4P
JCfceoIQujYse0nkHw4cdVILiLMquOJW/gcuC6sHr1buxv7rYcfIRdME1Y24EFXy
8YnDJ9I/NACqpetGLzDwzKWzd75Ibor+RilUEIC21sDSNAiZPVKGe8xtbNXmKVUI
q95F0Z5c89xvrl+onLeilX/KH+irUYevSfxBX4YrH0gA3xdU5+9eztwpPMao1US4
5oULcyPNvI1KGIUP+I9VCD0iuRRxq9Fk8WuuxvxkOhwv7xlzBBxXaHxZAkQ5F+2e
Q5Tg8TTC1YQd2O5glFzkf/pjp1rB5h1GypPGENMcA6x8U3Sd5bfw1LS5QOWcONK7
NLB8bnJ/RBj4346S+6Sajee8FUvA8snJbeQVKLlTYWWwAOZHzwYqda+TGSfPo6zz
Mkp9nXa+mhQ98nkgyw0NWJzu+YLsWTtWXLv5nNSCxz6XvmQdZlBrAYazw8ayJZMA
tzZ70FjPgkEbHgY2UD7s4Sylw0eu6BpG9XyK40pTkPBYQCSkzLPnwirbb9pVyXtQ
AEi0ZlXyJA0FEg5QJPJb99qr75NAq4XwlJBef88Asq+sDNCwm7serBChrMIWAdDd
5lSzakkdXACeeaqlm9oOaTb8/OZdKrzCY3vr3wxdK1DKa2P2pEH9Y/3QFAy/tvXx
Vr8zU4mkCQ2JQAyK+w4ctyjFqCw5afVS+DWyUDgW4W34dzXxadlGhuIb2ht1Pfvq
s+6vbsq8QaiUK+xJeiQ1hufNkPTJmQNpm90Q69N4vqCFJbVsRzhXURsH9QB5lCVM
zMietuOoRpUldp9sd+UOv2cuEltbXmuJr7qE2C5Prfs57Q5uiVNDxVcKbGk4doWl
/ax5UWWkDvvNRigvSRanpEswuXY9ISRXyciPY7hmQppSt99znm9F5v95Tba3KuDc
iOwWLkrXvGy25b4bwJzo4EKdcjXlqpEGh1hRef/QMK72PLvree67sOf4D3AuOij2
vSR25VQCeHfy5lLX0iLry1BaZQlDWBArLsY2mCKxKLMPjsunSBuLA77h4CWQSUzb
6kRjCwybUh9FjAaizK8z4dT/CvG6WzRE607fi3i+w5jOR/oqFI/+581WxrhFbr6B
+gatspbExJdP/70ao/lHGulBdwp6db7NJd2YxEQlyn3W3ZKILz1gcX6UkKHMGGh5
f3VyPVSq+OCa76KlnIzBgAU4rJTVzRQGdKuGHVxV5Rf6xVcvXZpHunEC1jrrBm2P
6O/ewU1l0ZAq94P45/VXsshSsRIyxSJFHvVFdGLmvrpA6uvkGa8USXZc40V2+6S5
G8gAsHb9ZSXyWRj2jlNpMbYT6Vcb14v8NF+/zOK7q0aKoIYozdR/YPBnZzTwHuX4
dzLqcFysnsyF4hhpeIwkEdiwo60nZCGyLzjfbQaYTo6eRdGAqPL3Z0PhBxBGVXk4
S+y6PvlDUZGRrc7fXv3IvurIW0+W+TfJDiOU/RXJZH0eJ0Xwh+PiJUVMD3YVH9ok
6kl/U7bn1ipNbMcd9ZVz8udLRELK1rEXm6rtkQtBkIZ0vgBy7rRxTyBSrRsPexzb
IjyWFpKDeuUgfJY1H81/D7LIrMi7EmJRO5q4QcMohwHkaLykJTLWdHvifZQLfTQL
Mo7tUX5/0Z28hgh5tguFdp9ReWhzVi3Br6qc80B3y8YdZQAZgvkXLIkAJkIfiD7w
JW6w/MCYipvNqnqH3qwwZSfewsiDFx4HAY5imU8notMAUNRBW+lGJsStSQ/Gi+Pn
1TxPI31NIUDX/MtTnDuxoA==
`protect END_PROTECTED
