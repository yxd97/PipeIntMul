`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEc9P35iN8jp0NSIMTVJSTvasHFTYWdcJ1Fs9yuB7tdboGAIEVVmde4qzHI5eOrc
muNIvLNe1i+ujxqCVCLH7kn3iuel6sJkyw9RPPC/bZ5PHFPtsR/EYDMhwMXph8rK
lBYSIxBaAR80D2ODDrSfU07kJ2RHrKOzmQddXV+3blqGbpXXU6m0AtcwKyt5ghXQ
KgxG/d23LGh1HfaJx/Z81uG9WqrUAjdXEBtQGT7gJjRPs7pjKSepfK2eQRvd4IS+
0P/EFzOE10Ia9lwD/U4hnEnsS9dnkSs0J5U+sAMODaFeQiknRkDIsB63fomtRJje
ws1brgrdfGdAts+HA4peiDww6QBG8CBEB3UhLpdMLbCF+QFXOiq2L6MM9ZzdeQXj
vqDSICxI+Eonp+2qH8V3NpR0BToxkAGkBu1xg9wKDZr56+bGohVZuTSY9pEZQD/a
KDzd1C3D0thJbbTfeQmdjfIkZ0Qednqwi3xVBOomUltnpY87lYZG0ZDpuzoikSYp
eygRfpBfLCoP6L3QhOrN3ebZYMoYEhrTKMlIzKXRH/LmmMwXo1siqJYVaF6HXPko
1c/QdSm2AMEM+96X8nKo5/WYBuJJZFKTyNrkLKDBbRZcTmAGXj0gSHH2Ol0dn2Sf
CBJIEeu3/7u3pWJdhVILnRNY0izMkbX6FHZ8kFFWzisVjV/Yelaci4WNKiJ5yjEr
JE8MB6WfCjNDJuQlhCIKKs2pG9dQWH/EmEmd0Fub4EEtDaeWxAkAOEwnhyL87Sah
vUH4grX26evwJIlhz7aZOe4r2ezu0OVxb3vlLOsAzaEUgs0pAF/BEyJYsW2z3suA
AnFJXk1yodiqqQcMqW3qD3hU972md2I7wwBtcxqnaDDiT2n+53QTATY89bmWB53a
PSx3wZyKUbivlh9a2ImUNAeaI6rvHbV/pu5B9cHYkPT8OlIfb6x0SwBmHw/vZS4n
pWbcn7ElmfoWeX5uKR+zBi9Iu34vY6Me+WJKCWNZgfRC17eaI6YdCH66lkupYBQW
wDcVVH25FhiO1Erj36pRpbRh4NxxDrGxIGshYxLx62idocpO6sK6gULzmqrrVrrx
`protect END_PROTECTED
