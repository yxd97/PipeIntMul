`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1iCTF3oFtojp3jVwAgaVMfp/UI37Mq4yFADQ6PeAPe1R8QTfab6LRrxFotenZC/A
vSbI0mVBiAL/33BSVcnWyTT4TuArhMG9aeqZuog5zYFpsFSH6FQ7Vsp+E9VVbqML
WuNrB19Vt9hAHJgrWDYS/bChvLoVC5dUPaxU2Q+6/YgdicnPlatH/E4HndiPWGxc
7j38TioL+CFivc867gEmJDgNmsu/0KfqOxvp83FtK8AfzStbvra7eqk/xuCpxtL+
8m5/zxqEEutwIi4wk4L4jjyatdC7AkR+4jx4yrdxUXca1gdn7YbccZjBHGVHbFxK
NxWZiRqPr3vjY1gs8Cdq8Q==
`protect END_PROTECTED
