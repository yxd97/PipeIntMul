`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dRPjL/Ss8ODLQFGTI41SCyOa3VXq59ArrSHYsKIpT2zRNvc8NkPWH4jPtWfMEFJb
lrMJDdKxAxeWrUcHx/z4MllpC/usg10+lHEGynKA/5SJ2haQl8298IIPECvxz3zq
h5DAe7in7xaFFsLSYaKPVej8/6fvSlrgxlFYhPp0wuX0g28Rs7R/SLMukStpDIZG
D25Fa7ApckvKZvOCEN6qkclgfK0ez7R0vx64MbVeZFXGX93GrIbXc1FWlq8QiAuU
hr8tDWYurSqP4l0QdpIhnfKCv8/DhXPrsmqpkqe7QxxPhcfSTW6fOS91Lc4ywAwp
YkM/+OdmlMq9geNW8+xED5gUM/lyTdfiDS1ltkWg9a3PlyriV0rEHFVdd0cJ/M3N
4xnGisjz71Idc1v0yvo6w4Wrg2YDq70IhfCY0rq1l1DLTzzDKDkFRhTSthH49y+W
HLQbYgX8FSc+VmDCgab/LbkAT8jbDIb6uC2kdS89EkggGpVt6WynpxJM/nG5rvma
89IArVYTeMLCTECcB5464jkcs8dAyQofhO/tAvd3am26XeFJO1mhqNhJ/tJsKphc
FU07CoRI7r5YnC3sJ0RuWJ1t6FSlOvqwR6gAjJ3vyQPnJ31czqpHT73p4+Vc4sgB
u1CYZA9k8t7mhjur+j5/GhbAPdICtuyEl4pNpGELapLvBuyPHYL3QB0xqZ5c/ACt
TV400pAi31AiakiUau3qf42itdC480Gqi2FyoDXX1EPSQYOIBQkujEILlgZyx92J
5hZPLAo3py9E0eChnEGSxXtl3XhPLkSjs8+spAiNV4/BIlRBcbwf43dUAT0FQKD0
mFBerNw3mTLM9SfOhI9FnmMkEQUrCVBJuBemW8zC61s22cbhw+TynEzZDjPLSbNl
Q16/jUSJeaql4cToXEsql5vvAx95QqoRJ/AAySdInwxP7KHAvYzcL4dK7gXGSXQJ
vKd4UwyDbmvwHSBjRriaypSgBeozo/N6kmcwWT2zDrDGt8EPxJ8GN3d0CfwR4Aq5
Cy3UhO+oTLtw8l2yh83LBl/V5ish7mgbgtg7JpJrJzIwuK/a7OWiDMCR7d3tamEz
3magAy5WSZwgkx24C27ymzHBiA+DfTCTQmcFVhwZXHlUG9CjakX2A/ZUULRHoQ9G
PjrFgxdlVKs3SLPvvtYA8vz84c6zZuLUI/NH2WCgdda8QYucOi4orZhma9R8kVLQ
DXFdRS+NDsf0ErJPRKVb3F0hXTXiwgBTUnZkXvd1jkBVDYYEU/P2mRS6Xl8dgn08
IV/PygHoFEiQk3dTyFpoWITikyF4S35xqZf3BtKL+9Peq4yCl+pu4sQpaHrouK0s
YTzLKCDJEzjfR6zDZ0BVVdyb/MRg/6NQcP10EVMijY1gQAZmPmch+FUmd3gfb3PE
iewUbfvxnYqENk7EA/UCiKKT5BRFcLtA2YBq9bOMToZjAIRuXZ4aH/3xGY0sA0cL
0pWsFz/JbkhBnwWsSwq1eeXfY2NhKMVSQBZFryUxaDSgcJb0AZz1MS/yLkB5kVfX
Vvwa5JJuhnTTUUJjsQUXydIEd6Vh4czn4ZvXGDsEtSt2UKR+KHTUVDrDc943Oc9J
l7X4qm6sD3VdKj3PBDyxCMdNBrF19ZWwVIQnKfO9269NNajwOTiBw/ynNAlhqT2C
oYiMHwAFvPrQpSYwg48IzpxFctwd+U7iyvpVkjPkAMiybr11h9kEsureEIcCZ53k
LXiul4Jp5T4c2R4AK/ova7PMU0elkP1A6tnYiOOcPC67GWnTzN2ABbSVliwfItpj
25tsX930/UK41sYMtQDWNkAlC2NEftfbvOZYLwdWg2O2EOzZsvmFvZT8/LLuvSaJ
MsGRgLbjA90keHlgEI8tmtT4ZO0bkgsf40sgBcoFaZLEcvYt7lxjhbzoo2XOJBLf
9Ji83D+yib/SucLMKyJ03quDZnfXgiao/6iIMnE7CGcTmelzIrfcg1fB32Uk4XEj
mK7TpqQAXywV1g7DTAkICB4jy4+WfBSU4RnHYHrBwVtg4gWAr367ky4X166P2r/f
ctjZWWkK50S4rnQJU64D/xOMhio5G28JVFO2gCnAJq9sTyefehqoQjWh86MBLFRJ
GtnSQtNMRdle9dkC0/osraURwkphoVu0mVDQSgX0GE9GXP0RFA9Ad5e/cVq/NFWE
d0VM8f5JyLajkE8gdH/ywKFwucmcAmIpn4jkVr5uE07Br6SBNSqsT7DgXmWWgjwp
6mqZkt8z6NIk1ulSQ36dlx+DmviFAjuVhmNevphITR5wLnuIOLX+jQMdT9dAjZCz
uR5A1sr30tqJXfOCHzA9dU2kx8j2UNcJKQK9BiYCpeuQYk7Jjaano+GJ7UVonoUK
Da6OH4Lo818dlhBp0teLK+4YxkYlrHEHQ8hRoAPRAYfGM0qdpTmVIzkKaNI4mEMZ
VGMDXCCLrrCNPcn+KeKOC/hruLqQSx+kXQTB/KW9Pax4keSxvklQItQ+IhjmZIYB
1D3GNugZQX3e51CqWAuFrTj1cKuajf0kL4wg7NmZLnAXmvVGIva1Oc0ynwgkzXxm
3rC65YcwO6m7dqvudd9L1kD34DNLHeoxCG+GU88nckDXuwNwuiWUqsbqOi6lr6j+
BG+1vfVGPi9Z4PrElQaF93/UxvoNqz4ORkMtw6IwtliQ10sulCazr+BTGLT2jMl1
N8WKYqeEs8C8nU0Gt8J9H/n6Gon8yqj6sEjZBhsPrhuAQr2tboQqsrqEyJUZDfhI
OGJWC0t3G5UEgOR0YxZwbAnsYcJ0x1jjLo3pOicsvwKkeymPvIM1FunDo3KADsRH
XPAAOITElNZjC1AyMkLerraSEZxOAtha/9GZfkXPiK+tVanzgmMcfLzK9nyXhiHo
TsKwdTe9Qxrhpl+1WxmmlOnTTXJf+WACPJBIJV+fhzrCx6cG6LbGPTpMAYDX3NMp
gvW2Mkf2n/2HnR0kXMsGwDrmbxt/90Ci15C0o4fMmxl87VSV4vDM9ejS9/o8lAVD
X2ZsMTTSPnpYSlvzF7N/w6GNjNSCeDTcY1UoZZT49PeGf9OR8KFWWLixCByCvH9V
QDlczSUUvdrurQvxScPnSZj8topxa6nQlQr+1zKKq6mkbmhjOMtmW9m6dhu9uTAT
PFU3jPz3VNRW1rdhTwwUWG19Yp1yqyGlfKAcz+IAyVjaC0ABASMobYHYnj87Rh6s
JqGZh2PCbFU+XawUj0WwA9+LIKwbl0UI4V86U2KIqbF6mBE9TiKn0hGL7LYvcjh9
qSdmL/vx0+9PezJEiLTenUGe7GzubRcWxxhv/Spi3vbONshmodRTTu4qpY/vC/bl
mHkF45WKgQ5TdWHjCmxNwekSxEkdPn7aQR2sIXNdUhtPsuHUzRUEpu9pkXgpz7Xq
R+LpuAarSpP3BSOhLVuaU65xQ91pBS9xH3JNcXDnfaEkAINC3r/POYCckoS0Eh7/
y5ZUGGqM3RPRjyQ5Iz0eZBvvYKp/jziGEmDkzlFVTIka+INHObemW0n8WrmjAMki
01Ab9ld3yEvGDWVX2NwX8kN9jNVRdqng/mhyfuXb94oA617XmayRLeGDI99Ykd2u
t0tsHRWwxK4IOOYs27xuOmrDRmpuUZLcyNznt30dNsGHxB8UW5rYKMNblLfi2sNX
s5LzxBY0Ig6B13elyoiuDuhGMC6ASvUOqWRkezAFjBakVkXstVAHK1boT1rWBowJ
aI68AzOoU7/DE39J8aUOYfbID0gIi6ovvqMOcUYVkDXW0DDDpAhWVDqIpMk/ZO4j
N2ZT2Hnc8mzrmminCVczR7Fu0A7v9Xzim2jS1gGYXKs6iwQzkGpTdPbvyo3JeQRo
VOS1nha68W7EHZysO5++lje1bGjuveUrvPD7NY4pGToKX4GuXehXZjvFLxB2L0sC
JnTe0vnh4zBtWHDNbwZ93bic7oj4T/dqKVH5oyu5U+ojjPCdnmFBgD1pBGSmvyr5
p4XqGSk0cYsjYSAAmC/g4xLiyYQleroeWXx23SDXCxIbHcV1r+4cAEH7rmddnN84
O8NRFLcCRM0YGQeTkzoSlb+GrMcSLCbVgO8Gukrmq9p/fwxX08+wQWbrKmXTYxpr
iYI7ZDYMsfUoNZtQpAcLJclY8dByhH3jVyq8SNo62cm7v/4sANqZ+XJF57DkMihX
TD296Khi9Fv0ssT2NXgMkOCjSOSxNYsHOa7wsQHXkl5USVFoGSYczZ634iaiCBM8
U7sxv/obbNQVmisJrqcIwcHEjEmWQqaXJGJmbQP8+oyr31xxOWPgcWM2DBicJ6Lv
7o0XXDixiRCwe1rGScbThXYDJRE3k1Mlkq4fW5o8sRZbgQFGFIW8TBS4Vnunm004
24ZnAJfEg1jHpDetli5QmckgSsuGhNXDvNm8Tt1i9TNyxZLqLIZvilxMawUdJCis
o2GHEtsPZWxGoHHfwzsP3C6bW5U350NG3b1Y2mLx8IEK5qWtWHuNqNvPMbEgeJjB
uvtqxTS0epD9F87a8qzfJiR4tF8N47Djj6cCiwSpUifxScN/ZnRp1fYl01rvUq58
JUvKKKJibyEvZggY42yEw4k3vAUYa1hCwDMvVrwo39U6vGziGnTs8fL9xryhY1RC
2Qm93C657xSBX/Z8IBh+THsy2/pF4KjH1WJBWXPNX3f68/qM9/XPpSbDw42b688M
HnACetHiBhW1WDfWGnQxAd5esErt1S8/EZVgpefmYjzvNaR68W5bUlic4i0xUX65
JPsHb12tn/3J96TGM+Kd33h/ZVQzqAZBC7nXh0dZ3zevjT07bLSJO7S/AytDAxIl
ox6QAV6XEXN8zjL/3KV423HRrWh66B/tWfNuF4NADr/JG3Geo7izVENLm5SuI4iw
X0hgWxDug81ZQARcKxNKJj4Xn4YGJ6zipPafQ8QIYaCBJqVUbagx/vZF1RyL+fQ8
Aa81olUQAStleobzaHooq6QMqaZJ6oyfSLhi+gyzXDA7SO/mJdFrCgVDtU0mQOFz
RSHdt3ZL9x9mV2Vf8nsn8UxBoUNjrD530EP4CC9/KpIjP0z3ubcY+k5UeYnFFkWD
ll0j5oi1dhU91VBVXBOG/sTif7Pp6ww6HcY8ZLSMrBWVXcsGzxbEwa4fQyYIHpwp
7Ox3fJGz/T5j8ws0ZnEPWkB13OPxECSjS5KUAQi8T16j/wLyHyU4XIW1JYMv9Jjy
v4KUL6DCwc28eMqWrorqxAiFMenvIOBPJJ5IJdIK3sLVjlKBi4GcWr7NDhLaSJ7x
FSWfpb12XynrnIwqpDEbR0BuiJ47k9z5KjHdIEQpwGvjseIJLOmzPhWUlblig0NA
brke0c8H7w8b+etE0p5xVd12nQ039R/zAKfON0JEScT1H0Vm+qhmdE9sgYDsMWwn
N2YSG48cXpj0E8DU/mq9gkh7ybhoQXmVLFymKJcuL2acNub2nZPyBF0pmk/qEnC8
GswN4iYjDhNQoN3zikmRo3J8SDLO3CWxVPeU2FWN/mj1TXvQykbJtdCsHBa1VH0X
bH8q1O+8CVDhY6lSQvMGTc3TJgXnCdLTRXzSJLWebZqz+pAXa+5FClVRAYYOAMD8
+tz9Y7baAc5XBlzJx9ajTZ5PVO8cc6xxzE0FeexLvrrAqt9KGncEIrbljg2pAygL
JxCEfPjTzAQsApcsuYsPpqy0K1GH7GmFItojsiQyRtc1SH8rKXdOO65bOJR+iaf5
qVXOjW1ANi7zs+Ur5Ss8pVOWuwOD963QjCnZXiQM3DWg0vFlJoUvJ5hh977kE9za
skfgIuBtDMd2nxt9EzwpAV9AcAr69HX74Rrp6AddinkDWNgk4qDmkjDddWuJ9cD3
j+qrYBOPLTtdCZBTCV1WPyCR7PwKYDLO/IIbJzq+FLFfYyIzVUmDpYerh2AmU3Uk
nSB7rBi/xGBVOMltYGFlXmNLGk9Skgcva3Os6G6BGcN0+G8qcOFvPe4Kbnc1vF6S
rXPoVoQkgj6Qp9Z85rDaUhjUHn2AKeZQGsPVVTEKUn5MJzCFyamCFm9hN7ADcNWI
QmIJIAv0bZi8uYNKQargdSllFskKnengvxZOIjpU6qEJ9dWI57yOcuj1JPYRI1Ht
EB8fgtrEUgtr9jrILkmW4M2zfQCScqEL/FPaH30vedqgKLkA41O6YyVGU2FS+EU8
dtI5KVOMGWuiw2jdFXjSyyD4XQRTFCmhaY/jKJEzCORsTmgUVU1KmcO57ijFSVUY
SwsjQBgwc1G5aN6QtBgL8vlTpHXnd0KMT/bGzfZ3JIsGnBrVixffdyzv0PjdGKex
wO7o3cQrJEKAmgBFrJbA8yAbBVKeZ3wy5FygHEzgHvSaF4e7/o/y8g8Sf0t+lYaK
uLfhbS1MCLL0mXtYURc6mGs405AhJ6WOr2xrXP6fajgEsqGtldK1jII8+cGYD8TY
L08MRv9RTd/qzl2k/v+Q6lyvlfjBv16vkhSXzJWD5hnERsW+bh24dzdWGiWDAv2S
S45+4/LNuvo9m3Z+j1z7q90384+hTWVhhNSRhB9Zmm1HSPwS4EVnB2E8u6Lix2YW
/HTYmsncbuluJGglOSud9ceaDyMzU9szwO/mM8biC/dZ6XJvK6PeSOzjxV7MpRcP
nuZSqjWPpf77dsEKbfQxqbfhlonTIE5dGdrJk4bEQy6jFZPLNSW6movqLuPcUjx3
SCkZ9cbJq3hWAFMuwXsOtHxgUV8aCYKM3KWWpFiEZSjgW56wd0tV+mxzS6tGtY+B
9avmCoWXsdB7I/xRBG5XAGAEeevB+1v87ysWY9W3d/gZnfMgWf1rnkUh1fS4x8VJ
GeVjuet881XEA88qKGDWR/YXYRR6NhlPmGLD8dCVMJPmMEL2AdC6YE8bDgYmWP9b
rjBuMpGVUOn5JTPHOn46zvdE263gDbp261q9NfIsYJwM6HHMRlWsq8x0LT3Lx/q5
3FYMTlyPxGfzAE+EOT2fKg1hurC9zZ+KB6IWoyPzrDFCxVCMNWqsMAXYaJyz6rQi
LMwWauqZX4qmykDKyz0rhWdXY1FpsmTCl5dC/NYx43o47k2eWDxbSamIO3kd83dK
T3mWrhHt3x7Bcbu5bQV8SK+1Zwpvz7O3OLdyDVXNzofqdXQ9pC/JWE4aEdm8N6gb
UHt6g/GUlTAaqmH9f7EAytsu3CM26afTjCRhrt0NPw03z3Is7dVlCcdV6UjzFvxj
DEdzKWdfbJGaJUYPsHuCM1ZJJlbeY1SZZDCFieAXBe6DGRyKrurUmqU6wPTeVR3L
4pBVfS4+GgdhrrDAsWxQ3PKSfTzwzDOa33yr5BueDCA03/QM1uguvc42Ik+RUJnK
gnSM+jPkpfmBA7mLLt/pVSiAHi59CRBLYhlHjpJHtEdJEDXtIYk6+isJkNrfSSnC
9GiR4G46k+fmBE+OaJ8wKOQ4sta2B17YoAKrqRruP/ZRBX042dfpYEOx5DnaR3FP
MRjtRkHHxnAN6iL+ZWWTDiofpGbgsIHdMnTywe1RQYXW5B6AFXEQaGBWOCE0gDru
Eqvxkl0BxSq+gGGsX15YbMspdaOVAmeAVgPtMh0lfHz8YbsTmEWPesiu2pICeuaX
FeiIRN4KUpvIK5/h7rW2GwoV/6YDb2pKn0MT6I9eP42z2e2phKDpJXMqpy5Krl3L
3NNsJcPFUEXv14ECCpfePHoIGaI6XcdRpDPIBBg7OqKu+DSBrZf0K+VctZVNqB6C
g9BAYpFhe/FcoOqHIWS3I48W3YPj/t7ZFHCCWbIyC6j8mBB27BbwN6u5/xhnK/Zt
8WUOwV9vyXB3/3+H7y16K4cyZLaJw3VPDCClJObvJtpPjQDhbINRq3QMYfrzn34p
qFPQf0lY/G9Gut+NrM6lgmL9vXLz7IysWDrDJlLyceEiXufkWzcxVsAAgxdgD4bf
SD6ZT0q0OFlS3n6GcwX8bdzd1gGP+CudXTmINmYH0wLgwdnNRsq5g90D2n6J6w7X
YTarVwUXVXzTyCNaKB+w1Xv3uR1h9MVPbMnnERA/r5FBXZ2xS9YULTcsv9UNsZqo
MDt3Hd03BWWy8bAn0eru8ACQbyUmMBlt38kFRYe2OzabdkDvCubegx/3MMr9gURR
2wS3CMvNPfLTomstS77KsvGvPbdhHqhJBGsAaQ3LgwSVFDMtLk6xpAGxhah1c5gJ
lfyUwmqIokAlkwk/k7f4d/LbnImwvnBlATtsCInTpM2OAys28Dqd1lWxRKYG+0Lt
q9dfNUkK4mjT+vgoEF2MH2t06/CE/vBJljx/bwKTAuJnVUXd5TeiyMn6heCepwad
hFj1mSfyvOdRbPRKavClfS5/LKc1tumsn+Bhd2fqk3IsUyGnecBatbmkTX7qV9rT
Is9HToox/mOS/1so2l1utMs3qT8T+/BmPOnrR0y9UEXLIgYRj7Ds+/IUqaGNL5PC
eAO1HFrD3ddPEY9Sob/gfmIgkK/+v33qtYhkXZuh2MwhQXMtcRgT2I44Mi9khxRP
5iIySsskswTTV257CYinZZUhp9YAbXzN0ClpguIUdmvgkBiClPAjRbFW2HE9kSUi
AHhXGs68RazkzWWFUsZz0fhekjY9kLh2DquDMuwRlenuMvIV74Qqwpy4JZBFP6+w
hk/Wq3OBbxWbV6lggNfzMpltkYPh1GHNS+G7UE2iWJBbg+69QYljLf60bhAJbqQs
Xr7msPOlBj9KsotwjIx8RFPwjZij3jUPQJVh5hCeQMlkNldpRvfNwVp2hJ/LP6qX
Zzz5bI0ek1BTxoXHwm5qrIwW8LrCKoUary615NMmWBnD8Hbuh+mJtLkUb4ChGL74
ZdpM8RJT4ewnCSOasZ7EdkBtAyW8z6qX4icpbooH+c8NikTMwZFqQXf3JYpJCq6K
wWLXf4UegpASQgxRl7txRPPt6MI+8+uUBA78EhkZK2KunEfKT8dAg8MnqQDHI/o/
XrwhCpHh4AenX4pDdKduSI4eCnSQZ2lgbMme5l8u/XQflIr/zPAsfC+x7a6RRgO6
f1dVe9KpCcsyLKG9ACxt1vymVI0ABZY1PkIrWIyDjwCzDHJqNR1KVqsMp6r7drYV
M25q0z+fZsEB8yjlseovNqO3biODAa0jEKRkZoOiMo1yFKLR3OhupL3T6XHIVn7+
Bzn4OwSE1xMDPr7/uHIPhxC/MfUwC8xZ7Fyc5J+jisqnnahSFYNpgjrtGE8GDiJH
9kDsYNKktHc6v0y+JgG/Iy9tH56yEuTgpFQXj0tqrUqPMUasrZZaJW3+vMycZ/AO
db4jo0EWsZ5i5gWENjwmYd5l/Kq5kjqCONWR806GlmePWmk297AbXRgKt/bkxSDH
Z2PFQJtk8QkBx1n61fbA7jgEatUrU3v+hA/i4z8i6NEe9Tfq+3uNSzs7/Xagdsov
BdJoTukFKWVoQ6T0XCsAQrh8QuG2EKeAvHjC4cJfvXyNNUdJpqzzGEG5FGfYc3MN
mZ5ZWscy22WTglP0BdVnp6jy2wjfK/dG2hXmyQ8+PU+ZnPmQMOhGay0k6x46OiPv
2JIZQPP+Kv+xmqNYdeOIqk8yBpjTxkHIBcf+54VSKvxrNdJWTriz2VuNzp4KJyBC
aY9GrWx/bOxV1RvkyPn8oCGWJPvq8pEC9mljNJpCFDrv1uMTVwTWiTxBz8XXlAGa
nIKN8vptzKDFFeST0NSJSjO54+P8AMZNM/qKYAzh0CptKPboqMS6xnSrpMD40zGh
jhB2uXQSjUdw72wtBm5ohr2HU4txp5vXe81bCt4pAqR+sHIXYO7znMHkI2yMePQY
GCL/KCNXut0xjA1Q+XJOT3lpTPdDXkJ/yKrK7KhBqYYq9Dsp3yjO9CZY01qoWjTO
S1tESd3M/yCQlIHRUrCPdKWolHG0nANnclY1tRcpBLU1ZAiY/2N5f7f57B7FQr4r
2EP8VPjR0uq3O7xaqP+Fhp8fL2dssjiTUDdxU3Qr9L5rCA7v/Uk1xyGUb2CK1vRQ
s5maWjPO3xsBR4RfyTgQXhgtk93rius6LHqtGDFYiGIqdUtstY72TBds7n1XL4Fz
l6NzW03GW4KLajXdxFMJGbch9E2IAtE3ghGbf40QpIwlXciECyiWhEIS8p7k85LN
TswRwMxH9UMjpKe9JX3JOHktxUUuKKp+1Ut2oA4N5Qc5nwAAjIOcNeQJNPFXo1V6
j18yxn0vxu4HITCrkT6td6CDitYNUpQJEDth+FUrHmYhbZ6MNp4Q8xx8X2thHkwi
wL/rwCPPHkOpxmanPFr/i6oYSy8rR3i7aU5a3j5dLQSGusiRh/B/Bi2vHR8PQ/Kk
Q5DmwYymBUUcNZFb1Uh9uRx00DGux+S7ohEZG5MHu0kWRMg2cMArlL8/rNsjDxpn
TiFnCEABr7paarUfzWBk2oU9Im3Jsd/U9o3v+7tbUm8kCXDeZkgqV8GGjZbQn+cV
Ddp8Q3G8TmwdaOiHqb0qx1sPy+zTEcLhgaZcRAaRuEfh0ea4NVtDAVdv6mqfxdiG
nlBdOFHaHFv/IJDTArZG9+0QMk/A0z1CYO/4gbOJiOxbTEa2vZbu0JmkAqWRmerZ
NXGDCco8eoccoNpfKyOVf6nWXyxXd+/RCjKhuL1C8UxxOA3/I9iS9rZXejPK6BL/
Kr78FKNhSCRnjdou2enzMryOkaycLbBdHJlY5JtMBxkgi9ULxn0CiZD4Z72ubDk8
eGyOlyrXJyD7hIUmEl9ZHbU8g4iTRLJEsCYDx+5Mw+DSvOb2V37WemAzw+h9xENc
Q90VT9tQrls2pOCSc1qwk83ieS7FIBWceHZhYQLQoNAcUQrX774sdHTIr2XmDmxN
3E3c2l44x6qmlq04XT151CdtkBDdi9M09qa6oMAggTU78tEhwrUIKp3Gg9aktgIK
abne6N1ohCYMe7x1bcV3R+fzTT/OSPIvlx5fFNO1/HLfJM5EpvmynDh5QDFpdQmz
Acu0WSYGUQHw3xzKIakNelYjCznpUuTaRSCqAw496GQ+7qyGlPPsElj+CMyXpNTA
yosBj2bGZX25vB38IpPc6mSD94T8v2v/h6NQwwnNFFRzw5NOoEBVl1Dbgvr7Pua4
VppswQA0Z81Z1JEzUoWIkU4chvqgMqOlLI+x0csDR0f7eBvXG1kqUFyIx6daA1AK
tsSFm765CQwJc5WBMyOoXbjXVya+mhq+/5kwyKXKUN6tDuQLLiQp6tjR9QB84sdm
hLnvObA2LG4j1l+4wF/GmnGlCvSXiFH+dZNZoY5Kgyx8fV74/dLDjD16vuqYkb7o
cPZsY4V1/NwT3+7+s829w4zpJ0ruZ6TSvWDcMU/3b+4Zxdg9VgQynWZqIlIZtloo
hlyl5092oboW55VOCOS018zYU5o2jsTshRhHSpMbO4trh4CMHLyn9q6HALwiGAWU
5kE9ySxyLOBRtXZm5GRAdTdk5buYnhFQ/QRYOM5ODZcMObKC/ui4VZ38jDhO4QP5
MH8igDsWe+4rbpSU/5X4n4TvORT1CD+aJY1UN8A5fO+zgbwNQM2HjZGZlz/mTFVp
5/0ldKKeV40tzaBrPa9kdvRzjnC8OHu2cWcvDZx1gHoiUY/HHPnJYaJwSHb6Ottd
kF5KfIwdckdjbU2dUQ/S9R+MRD4VGXubjjnfSmH41uF45iuKXLcsHsHgNgkYIsUf
VveFh1WY2AVtO7TcDVvdhUWh6lXb2AMklWW48UOjlz/lmWh5Nmv+TPbs43saSfEr
LYGm507bjOt+B6+iy+sSMLSN5yV5kgHCWdRchloZiwnF1uTt9hDuuZ1Qe5izELWT
rrWUhwcqEG3ovGz5Lw+N0xXZKtYqACCyZgmO/b3ypLHyYAx2PHxhdsvPD7uOZ3s1
bTfO7VV2XKpzqAsbecXNxjobVlv8drvKYKOM4kQ6OuZyJ0uePdJhXJhLliPCZMHJ
w7j7vQVc67SIXz3Hq8K7vHGWd0/OFUcqnrTEbnF8q+dPRQ9Y8Kd+nt+t/lWup0ak
xlNFNMVhUMpuDVhypdLcrQSpwpq2Ms1hs9rJTOFxTNiqxa2iujmvBCFgwWF/IC7P
RG//iBKQden8DyftZu3h/EswcpXxod921jL2poxBWBCI+/II8ub9hGQnW74l2Gga
MGGw6MABNWUlXx1J1zfNYOLa4aRgUdrXZ5L3b6P5seMkT7/g2JwiAXfgTEYJFIKR
8xDhV6BI1kpdBcnh4X42AQcSSPjh09IrFE71Tt9hqo7L5OWyUfZod+nvXKLFuBK1
R0QZhnc7cMpAL2WSCO1feETdtaAB+a09XCWXnRqd/HukJjageuvL7UrsMj7E3SYB
K4Np7/6wnH6CjiSUDKHwZya+WMIBJGlNzJO8DeMGLxjwMlw3BDaJchPQ1SMbfb2s
yUZsmfV9pqxrBmRVJ4BaBzQoVdh3VO9Vhw3hS6ZkLvTHqUQiqB8GN0ATInATIHms
QRNovGitjI3KryOtsU2quH1ysXJ+bgl88XcVT6SRsWiYJF4w946f5z2VAqugvXdl
yZI8xHH0Oj0iCA6RdStpM4KBBFbe3jhvvigt8eY+qeh++/3peWFCI2zhTCTIgGsU
Fxu8s2Zoiz2HPhxzoRe3O2LGmnVVnmyD33HWEXis+EJcmnQxfvJL/nHDSx0aao9P
yvxaE7G0RFIsns3xaNI1/Cm9OrlQi0REie4X4XpdFrkiClJMWCYKMRdRwzg/vIvb
ywfzhhmAI/SM7Xk/PwDl+NMhpu/lfrXdsIbwD4MjJQWD1yN/49cn9hxulOFUTnww
W3WPIQk9xOGWemZ7vo1XaaOJabZlc++HJXdUh1/kECRS1Hk5FsLtoz886XIvtgnk
SmiUADj9bxl5fO7SqGXkkHh1EerKdkCGiu6ctq+FquOCaJAlr9wH2RqK5i3qxMTw
b9lYRX0olvA5i7czoU8uP4HfO9mcc7UR5vXqxytUkhKL2wJyeLPFO2j0C6PrzTBw
cLQRPP5J5WMwXZygLb69PtQn+39jaQc8GwTWlDMvs9f0moZWKJXjkiQEYNQM3UHm
VHS6ihAO8YR0Cuoc6CDVFx1x4aa5yrOWeDkwHBOCry/yulwlBbWXQZkDz9W2+MEw
19GZIy9TOXII6CNPcUWvc48A1Nt1+oeX387MEVguUAITpn8UjI7ey4M2NH7PQryX
tTYlQB5dzi79fMQPtOoa1F7F/lrsf/vW1c5AdIZJmgyN28pdy1fCCNGOC5gXKENm
i6SYsIksHCsVkV6+jEP/gZXrQFwy2f2YhqR5D9WSb/JhJg4l/sIjnuUZ6covkpXt
y4zlcgfn8XwaCiB62kaCTDNdiUDdpK3cq53LjB9uLWXWjQ91UVKZCkBeRirT+H9T
9UfoCE2uUHIR0oEmbhyppd1ky2JgsUWZpE8eCUVo9Nv7g9QadE0sSgusJwjbBYnh
b810tSIMBKTfI0hQd4UCdaEJGY5CyH+I2+EX03Ujcp7+SNHwavJaz1UO6DvcN+rD
e76D9ziCUvAM0bfqF090NnY5Pg7Aefis88WTv0mtHycYGvqwLM2vLA7sdOw3oCcD
V2bm+yEfiTHCoTYl0NP6ms0NefTY0FLPO1uzwgljwOnNaP0bIQkpugcEy7LDAwqn
QhQLinner+JjSFZIYHlUuzExNtFggmmvKYsCjk0z4sQWkTYqmP2Wq5MidgJSFgTs
Ma066N3oPj4fXYqzQHZtPAv8pTg36ifAFLMiHTY+CLeKdnkwrCa5kopgp/xl/f5w
BQmDmtRAC+1fye0a+Xge5IvKJD7z9kpLZ2IQ9rgbUI08GwhMihU4m2cUqOfVaT1y
NBj66Gjj+09u/e3imkRfwLPw3dVcVRqWhBtSt0K8ZeAQcnXdjioHdNnqDlcRTJdA
jDboNnb1/k0ahxozw3H9GtmXtRQ/3hWOLH9GujwJKgJnHqhDxOQuSTgCAEOij+9E
CGcydQXdFNcrSZ6Tuu6WryFoZ6aXnmVG3hFd6Yq0FfqFjQYvNpjMBaTiWoSN9dsS
po7u//XLuUSWREQTfOxq+Kw+0Kfd4mzWwJGjWQ4+glwAxYNPthq6VAkwBeYvzNIC
9e81xKbY9gqPz4uVE0DOcjHlbhzrG/+IEUvC0kHJmnrYQeBwHRhMeuH7tq+gGSAP
n8NwuUVMkT+Og5RmYD5qB7aIORurlMvssFDrfgH2N+xCiW6ap8cATdktWSJGoVCB
fCXrqrzd2Zfq59PCLdQKbYLPWTmtUwUL8ODI/r7oiQnZ+4ZmFrxdrkit3IXjo+ES
SWaK77Ckvp3NEFTqIVvXdsU88M6G+hIhLuET1JKzl98t3qZSoQvbilunn65IyfTx
+JfATAK6CBGV6VHGPRO3KymlwYMqegul04cNKqSLOs+CHgp2q5hpXG6IydyTCjLR
oWjuar0016EiLMo2+m5+0hNOpQ3vJcfp5iAF9544oDxveT7G+vaMNk1VegQlWGQQ
gnOWxdgxMWB/eircqCnHRWWdtpSvLqkzJ+bdX+sy94tkw3JMF1LwsDGq16RKYswz
WvgxpLXCdkYZqZl/+FV3ZqET2bNagEes5vkrmOdwEEWcp3eU1plQJNa5Og7x7E1H
kpugpOrDWhQoBoqVT6ck9quPjaLDHh/IvHrKk4VKGdrQaKj0D4Ye9FK5bW41oRmQ
XCTeqz0MkyrbKEDbXZTu/70xkEUfY6jGTfa29FK0pKfKTBYc/huL+dlvUWNfjTpd
wOA5hKX+i9gEBDn0Pk5INd4fcJCrTDjgttKeWbA0QXCMGlZHSB9EqzP1DTJIT85M
CAB5tat1/RFhlfH9TkEvYMS7S2uVvgG7sV6F5vbmWvtf2LtszQf6aeIR9y0pW91o
pvzoaySZRk1Qoblc99IVXGSftBOcVPKK/DnP+YCietbZt4E6RT8mxOZIYhN0Cw0h
1GUF/DF2LQGuF6V6BT/I+LbMNWJWBuh4sgTP9lJS7Gx0R1au2AKhEqVfPj3uk/Yx
qn+xkiBCKkHmzn+jyZXQRqX6qSeFdXG2RLqkUoFEHBGof2nNqrzK6vDyx5pE31jn
WgSqfWjAyBnHAwVJ3FjEEYDvziOB3CV4V3aD/cA+udWrvYNfcL8wMPsljt/vceMI
n/kVj4LKsHPWuWyQfnWSpWBznNhJG6qy78VIsth7/czk7wL+wIGwu1zeNPYrwGps
C2tJrHSn2HSN7zRPFVPBJFfNIHFEP5OGPsK5v2Gc0UjIv5kKQEpo45TjHAS6navo
jzzEZNHbFezzWTETd9xE32L+L6wN5XCmOvYL19Z2RYL3dzaSlngge9CFULyyXF3A
hJTJraHBJXO21yjQFNZB8rT8qYPsc2fy49JX5iy0TjVl5ApNZfA7J4qjGxS24ifz
uJ/QXbSILTiWhlNhFPAo/kzZj1IJLCK/LFXf1d+aNDrobrV1/u9zARTSxwXcQ5A2
J7JCwDZvXxi3PtSnyBn/3bnxk1SSff0wGURd6/kmn3ykvOiVhR4G8lj+NmJ7b9t4
zDehCd477WGYfn8UxnlNw9xz3jcAEWN4V9KqAncEs+RXF+kfcqRIiy3oUDTD2EF7
IujuyidNzaZXgXZq2OuaI+JhZoCK97AC2g+R2pRfPIVG8gfCtaoZijVXR5IIwQ5t
Vcxi0Rek0chfqfrcBwLWBb9fKw/gAME6RfFxfWDOyhxkF58c9psyn+sYUn39cg0N
AUYzMh020lVK2JEdVfUtRClv+6AKPMugdUQiEs8UpnjYYCbOsiRrKDEzQaF++IRU
FjaEz4nIiWlziPdX7J6GyLSKabr3AHI/9HEdN5HuNZBABT4wd0TVY5CQ+jsxcayK
daIcwJZuXHSXqPTytQno3c8rvyIlYsUWBZIxkdV8ZMIuK0nOwNFCrwjedei3uKqb
9bXQRi6I54wYVIwB2INcPWr7kLaKcQa0GsA6lW3Fzfa0yPNe/kkswIkFtYoeYF9j
DVNHxpOrdkjAsKuRbydrU5CRmqgPd5wBHOg5lUAASfgjXCHZSOlT/9mzXse078a2
cl8Rk3zg50WAQtNEEtfv6pDnFADdjE0sDzoOXC+Qp3f1TednTO5+KzfBNvbQzAxb
tvan2z03gIOoTJEdOWVmXPUBBJfMQ+mfuDZCbMEgiz/KkcOrDWxSymY89u4kI3RJ
yVtPDKjpNhGdd0sLfcmRnOLV/h3rcK/su2GbgXpQgpjr15rKg7p9HKj/QaJNBzBj
YyTpmy8Sn7CsyC9yoOWOmHpQ5ykcOOEJ6US2/kXrl5m+1BTcrEDZWKOWJgCSK+Cg
Mz8C0IxGH6Q8O/KPRSZV7bk0wvBU3J8Guh/QIAL7U2dgHaNataUFBry8TfdlO1M1
qe0wzNOKOEUACQV4AyWHbeH9xOJTiyZe7xR/DQonh/GRWUO3HkDr5sH7H1rhsvmS
DOcjTOh0nxkT0SnSKLfArSZgWtiw8il0BuRELuasDe5Wm6Zy3t9mAIVC8lBCBUd7
+1T1aKPhX7UW8RDPlOJpEY900NG/69wpA8JAGRXt7sWJRpiOJZ2/k9jSPI+3K1kc
3qS/hKXprFifKZ/rVSanyNrmB9d9e0zAldzAPfnq4ZYFxrMI3fzgew4PSs3HrKWk
YBRPm/ihSJyCaljMiDH536XPshYEoO2UDCBfjz+aQMRdrS85enfKW+jlWQl+VShu
nDbE4cpQqeuzRBINa+RP9XwLA4fgDUtb8j0A1LFj+xVU/wiXdmTdalm0/mpU+EbT
V9j0N4scJkZWVPYR4yN8vi5fAzXziVDN6RmQJNNaOSZeOxh9QB9vclaF+J+SNm0h
TjGPb0dRy5S8cIxe8TGPYMVxSUaQHi6hPuKVr8KStqAxBfziWmYdXg3k9hPSNAXI
2wjvkyvCEU1nwGh65Dl9y7z4qTGMoW0IBcKUT2jwllg7R3aifsg3OoCRFAburZ01
546uF0aCEZtdTHArB5niW/GhNbyg23UEvcHLhM4fWU8d/kq09CQnGRE7SFtX3b3c
VCb/lc2nz9Q8IMfcaAaPP/tAk/K3CZjs5S5RAktfLIuTUbCRWzQzP81zhQtAlT3N
9Vcaz8cuGo+qUTTcH/pQ6aay5BzB0LVl1YVhaxnm94qoO17xuohOtNqHhQ8UatLg
YcjQeq6+JdcMKL6mCaqh2v4W5FgKWsLmjmQjpj1JYbTLXJF1rXDXoHtcUhFFN4fe
uxCAGs/LqXily9eNcQwleSf4m8MAHx09RBO8O+9ARk1P47Bp75JqMaUP6wBAyxvz
WG9XdV2O+MnKb26+MxofXZvoA6T6uk/nRfT0AStqY5eIqZag3T0x2rgyn76FjzLy
/mEThgyu1btvSPWzGI3dyiA8L4hTkOFt2EAf33WHjLclclJl/JMt8pEXpjdSk8N1
q0S7Hs4kczDKT5sMHKjOeBtGMGYMAccSz+dNgHiU0GIhclfEptI6j0jv6UBP1LfQ
XVQLDi6Ky0rNWGvc00V4FCFyq5qRcRMmJypv2SAUqKP/ThyQp91FsVMK3HuAwTIF
sZvBAjzDZziKvyEvup5eckI00kbmUC7UyuKxAGxMp7HA0IAXrdt3coiuPpj6HVni
aMOu7tIq031yEvwdJwyR5TeDYXrep2auRXCdSwhTR28qZz5o1kTcrD4etIxu+8ZK
4KeqvcyY0dN4T3f1q4RwoF5JbyqK+tDcjymQUB6QHyOWL8x3QIWlbQ0vaJkxyvTm
KEb9m+wLsnISPKFlqK/fqqowFd1/sczGMvTvmVUQ5haJeCwcTfiLJF3n7HvmUxXF
hR2GZb6HG2UBQZMOtK6vNzQF+xmTvOXucnW9OByMCTVaL1kfk+MUtlhsFzvOXuEK
NjABw/y9BIvmwYKFZEWS3O/cP414uUrFMy3RIezV2UQZlGlVFrqq+k3xQhXWQcX4
tzp6uMbhW2PXtEAX4WxbDCKxzKjtbp7XvGd+6AOyZ426BXHR35DYgXCkxMhrqdWI
knfyv3vofydHJSENVizSgfTVyQOYnlnUYa92ECUs+QTVyEkS56jqbM42mR0Ng4C3
OxFRxuwQJ/iKSJfAPg0jP9HbWOkz9lU6S6B1+3daCFwxrYgZFJQ0y9ph8LLZ5Zwt
g6kdZ9DsKDM8lbu7DitRYYs9IrAimyAOqOHpleZZuzwy2QbxgGtHxFmzRWTU6n0U
OYTGplJXFyxUVEdgUOXDm2+jBVEXv6b+45uq+NWZ2X9XlbWWgVAg1n/7/1sTr8Qf
6QtYGCwjIYi64+Dfcgn/NSK+QLeEluYmKMQIRrHNjJLdzd03hGSQIa9y+8YZfpHF
avd8CJWK+eIdx8TG445nZnFXjmFYOQV4AMLbrE9ad6kwxPc1vB6RXIkekDqTzUd7
HtNAUOTIlMF3m7w1Q3GSNNLsY2FTTr1zwt3jrNl+SIz4p81e7iBTQTGlX3y0cXZk
irw7S5UrTHbdeL8WQoNTvHiOMZpgDzIzFG3Cp/dzNqYxOWKc3v4fipe11guEjYVn
JJt+RHUXCsGDGlDIA2MIZeLj0xT1j4XFYmBKrcFkzquciSjt88zblDUw/kEhd2W3
hBdWz0V7cX74+9Hl7TcOIe4SgYHh+JGIh9Q9jxER2NLCnxVd1h7MV6ZitTh6X+wA
RHatQC9V73f5Zn3TZ0NcIHBLE9k5D3fjYBotKh4uNoermQmbI4twG1tU+hFOYA8Q
tJgKsGwtokDJDJLfubQqIeI/8wm8LjaOA9mjHJxGNAcZKEgvig8lFvKS2QSKxvIQ
cIx9/TgTdsMi4HpUetKTh3PAUhpa51ZdpKRBZa/FAMKxPqLfljt5qIutfPiNm1HU
06oKC6YjcZVL7mEHrJ9Dg8Cty+SBFzA1+TXh2ARmNbjKjJk1b+iw6EBwj7guJ9Yi
1R/ABXAUx/JHomBZNFChhkYD5z+3T/vfhb537/ML7nvJFO+Fc3nG/rpI7hbNuosc
wlo4o9wyHEWDyz0PfcpNrMmreaP9Q1lbMUWOPKX1srjK3/tQSox56J3AeYSqmdbM
ZWfo/8PIX1eWAW70MbBA0E40fU4DWkgx17B1WDve4jjd53wTEnfH0QiabzuFQMWw
dL9Iv2YKJzG6Vj3+mt2nYVkGX6+zAKakxHnFNyc6dgfuxqMecNCv6rKFTUnC0sqx
fmD0bXy7mbTzJhEUksZc+IjiYGXsVXkFo+JyhX1ucT7EKyU17Nq/7yBR7D+z5kHH
CE1txFM/cp3utD2QRxpXWqv3Alz2/PXN+hzje3kOSO3sMMlQBJCWhWTaS4xG3t02
wK61xdhQTwtoKQfiFp5kHkqbmPm56YEcAEJ4CHsbKEh0IqdVaOwwCARydSqdClE3
LP/LQIp+rkUrdE9ii4q/oXBfCV+Ma4MZt0wEYsA/lZ4MwiCCExLjEVRr0tDqqvXK
7cDWxTMFOI0ePCJZlKnUsfbR5EpTXeqYwPCng5m6ULPr7JYMBDdHy0f7cmlZ7z6F
1UnduDZbtlGsF6avdLXQrbu64zxlEMTkyVKU7ek3Ofxm0PyRWR5BGhF77b6fzpL3
Ini8ySHP2KzSJAarXbLynOJVZiI03fXUmpkCYA2PdTo0k2CfQas2Xq/wj5+Ek4ue
TuaNf/B7Eer7VK1D6DoAXpD6AYpWIOHpxnDWhg0ECuXvVu8Igj+dvBMJyKdyPQPX
T2v9WBvM4dhVbxL4zV+zOArjFGdz78Tclk6mY6qtlauLSQIGlHzjAAUFTZEEqO46
atAi0YiS9stH1J5z5ImKD2ofHMQxob0VMNR2CIGw9HosT7g6fS4PI+TlJZ9NL52s
20qNBjd2V5Nny37xxkla4jo2d04QFa/odCGbtXmHrDG+xG/GPGq3oBgEtpFUB67n
zByqnXAGk4t9l8e34BLDW1B0rbDGfWXS8Z2z8fgP/ijNr5w235TQYGqUTJCY1e+c
0bywKS8+hMwUiE99HZY5fjgF459Xfh1cLhJ2U/cwLqr5L0P2MwnZptERVpfstD4s
jpA4esXgos38FVFOuflgJ5Ubd94Vt8Q33TTJV+X8nCYIA4WyMGP86KyRpm0nBacZ
RwXeA8bXr2Xw7pLeXlT1Xlkj8RHWr2fkkJAyLDneofTJpvRUDV6lgc/+dLkVGNSt
y0XuD+iWhaWrq4tO7+tiWyHZe1iskL/P7ziPAU6aIpU2xFduk+jaoshT70IwKcsm
TCsiHDp0FFxlVe26MeZnv4qcHjMl6x6dyM2J6vjtiMItMpVi7Tg9l/Ew7KlwyYbV
OZOnq+6RHkd+V2inPMUXTgzPagoZdYWBc33/i4GQhK0OnfdahR7VDF5BC+UciFAP
J3ulHYVGnR53rvzeLXTLioctGMUjO4FwAE/OaQRrkg0GGK3vOd8Ydied7D4AzFAo
PEAgQChTfQQ92G+g21JQZhY9bT3ItXwMaz95GC0ytrdYT7YNZ9gqOe/DpOKF0YGU
l5Rr53lWLl/0uc2MZOVGvIOUc+Iv33gTKkrqh6HXX/jct+xXv0ikyO9AuzKW79wh
0SlVVr4HcYfWZGBPbMTRY6dpyqueSmOcSuLvOop+wUtFGxCp9g3zl9iGrQnGEPYt
grFQdilqikrYjf9sAIEM2aluZC20Q4G97s46WfSSZBYT2bX0OZ8xCz6YJLERE+9j
2FxoQztpMX6Rr2KgQgFdGTuMIM6cn61ZP3C4dwtPro+QbPZMSyB+XDurEgJbB86I
dHBddXoX9saJCtQSB+i+/+6659gr1GZMQYZLmAPbEe3cPrjScbuda7+iyJrtjDwS
FC2bsMQnEJv4D4QWwwUieNVx0cehyHCYiKAY5ECbeTUx7en3gGE6w35Hu3jVK7x7
TxBdndxSz3FnhL4MhuYUA/AyLX++YkKMPClaOqUI3Kx8xMaPYnuRbX1EfxjerZED
TOoWY17Mc6DTrB74OYFeRkUNLlBn9NA2Eu0EYa2S2WNdki8/qyzGhSvJkdtSCLcR
UK5OKFYO3iAYW2kl4JPE8Xr/WslUNU1LG5fXTI/TK10MePE07OBlziM/kzLijixC
JuYN9ZbP5Wh4apMFWx8jNlswB5JXB4VPYH3jQ7FVw8eFw1MMB18zAo+8LGDBdqqv
rynlF4egr6ukVg+5Us5/B10E4lKja1yiYOR759MR0eDHJv7HIXkJFkyNGqXPQZxp
FAea49+7oy1eXceihSkzTg2cr8McOLwTCWHYiqcLA3R9cSqb3oldJK2e3XuOx+6/
iEb+FPI5g2XsolnC/vFBvW2+V74Fjciy91WXIbh7QHPPnfSt9t84fRiA93ykEha7
nnV8XqvcCrSfVXSTlO/OKpBV7uFDxVzbKQncyn0wBO+0pX3538CMh83CzwYCGSsC
el7IMXzlAb4fkajGoHg1nETsgyv/HOOd+eu1YJaoXNGO+4TRbihJVtAhvsqnLFI7
lW7W9G41zrRwrM4wZRj8ESeqzFufnrisiEcV9SMfjmP9++CAcnkGR5aI0uunK+wm
nHZl8Z+V4CDkMqneUMQLhpbarfFYcAS7SKnj8XTi6P0lrXGj52DDy205z6t/HbGf
49T3HgAElpwbS0s5GMEQ5UFvcZ1iICC8EOghuNMjW6FdktN/xXOAME8bsjNgQciB
OOsxRxqvENxPvHTUCEC0K+MO5cbNpeH2VUGNmYCUFk0mNhjUDSr/1dcMMuoJoPv/
ZwgKGWGDnO7S6DJQ3gyFsJVdJI4mhb5C1piRKJhTTj645WbtxNUIapIR/ilqFaZ4
LYw38eYV7A5GPEiwALsFd/fWWL93Ozli6/Er7MA3SSDOhR2PaDlOdK5/15V0kQkS
xn2mFAbT5Vwnxv5mJpkaRCS+55gnYzas4nqS1FRwPUxlIFLG0N4PFUbB/Ud6x9Gb
fac/K/NgaeMLLAuKkkcJet+rWh0x5y9EAPd9dqC4hKOpY8Wmx+8HMIBWNyw//oUc
TGOUB9zwK8m9qlFwsLLvGpo9iNUo+zrU4W8pkylo4eH+S3RbFuqhwTA4LS7920nY
89JwY/LHdX6ZtjdaLqux1jK/Yw2HzQvXEBPDkabyqd6YmgA4nt+SGZ2RPpsFCGPa
JqyaLEwI/hPau74jSvVIrVbJHPxpgUbRf5CW5kqThPrBsBTpK1FBQHtWp5X55DRV
AvM5sFkFvVv0kjDpcagIeFodD5ZpRVWU04X4NxNCtrQBtDkQJ9+kzrXRfjZADbuB
SBGsI0xHKYwTdlQtN5cg2yjsfZL1qsKksML5HcG+Xdw3wHJgKdMBRKQThXoLZfRP
wVGpngxw/iYuIGNdlCTt0gMWqsAye8M8S2srWM61AaxJva2vmaM4oiUixSym2Lt0
O4GuEoGvmB3Nlap+blwBl62kZwfULp8TobDc6goFMva4AIOqZR78K1gtbQ9DRQSs
iPp5327Pjw14KB3T02la5f4ZLdYUjtnGAHIVS8rO75Bp9YlBgzXqaWRoX8QLQCPe
I/aiJ1A5ZrbG6f7XQm3oIKBTT2VQZSaIyymN4zjM4yoy5jrKcIsrPNI49GvrluSk
VBlXhzi8SN5OhRl9bSIbcF0FgpBO1tbfwu7rO6hXxwKTbZhEi8GQ5CddfcheK/kP
+LFY1v16hL4W45KJzwNOPhf47O1z0/rokFMk78ZqXYlQT98Mbw1rlodxuBO0CNBV
tatSYgpBgmfCr5j5xSupEPpRJd2I+cz09M3n/7RUbP9Rmmn11VWCLuHIeqJy8lX1
aRIXNijOk1mma0q9MtWUv4S1lx6s07sHK/Tuu7/ppAVVPjmaF8nQZutx6MTmbsfK
lHwjuRrqS6c0k5DNK8kN6ouNG4ddZURpr9R6CM1feuupOuT47Pyyb3NcH5xL7GaY
P6uKFNGY+VegPDn7McZYyZBTXMe80VpViQm1zxaqA6VeWbXZ6D1IibQQISlpcg7L
FGzZQcJ559Jor6oOG9ytSxPIvBruSISOi07pinMprO0h5CnPeIeew3a9dfmb/fPB
wjOLKAz++UHq21JcESY8RjydvdwfSPmXNwAwWg0jLfvKhzSb2giGpKy/3a/q7eYn
R6pMzindZXgP/yiQ4PJYz+zFb/MzvBl+v7+SXVngsWGzm88PzXUJ0s3u/f0AvrxZ
zMx0Uh4Fecljwh0FrZdi60OdoiQKByL0VUboPWaCMp5+d+SKZwa8YA/LvcmiGi6g
/hY2ObTK3YL6JnVU97pNOubWBmQAgtGqEMuFUoa9n3qbE4PcTjhFQHsx6PNk5vCH
KgISL0HuXjJqhWGsYtw2fXRe1Mq6ZznQGZ66L/5qEdGiH6kI3ixaIu7q3Wof+lCT
JryIjn7lHcICpDVZk+LJKQGpN1plEv/ntEZlRFmG5gd8Rw3g1mYCtrtuSc0NlnwC
UIJk+DB/ldTpQxO1nxfYYK4zTzJIyq+LINXwdWWib0ObdiMUZkRjhG1289G7xP/q
YsQxFqitWgZujT4gbpb1zHI8ViBpA2YrJyqR70lTjJcKCh9aI5V5gxrP+XZElaR1
Ed0HQijwr0+EApeh1vGcxBZpOD4Cxre7FAF5Qmjpal8mh451wfOoIRpQ2n2WdSFT
71WV6T9qgIREWxvn5vwLBHEDBs6lVagKwXaGFIMdyEgwIryxETBwr43Mo5gAjtzd
JKAwR3gdhcAFyfNpZeO44G0FymHInMUgnTsFD4gfgqmnh+7qRzTb0AQFC/GCsoT0
pmbnYRBTjgG17KOmilQ3ntpmx5EJKi//BA0+/fCJCQP13mx/76Ak1GC7lrInzjOJ
MzwPAw0nZ5Gx60uqAYdxqSevMuPVJBvmWdGCt3AAx11qzd8vxMeXaSAhcVwHN9XU
0H4V4mSWd6Bb4g1gQeTgCvPM3lbz9Op7TvahbUt8oClMCSVSOUPLmWVUN/vj3oEX
TjzB1buV1iFG+qgtQIJ9uOQbSz/tw6L2WOcJNo8XJJvhQ1+R+5ZGCsk5oojZMMoA
Pp/i1yLs+imzKPldNyIoFp6JVyUGyYO5Z60QiguNgnUe6L9gEnM79HL+uitoiMrS
Ap3nq3CqMFke2PTM6w9dqqLDj9n5M1ZWeYFNwB6+pprEWs4l44x+HgKN47ek5lGW
BtiSR0LXqxIBztGxVO9kGnexlwsaJ8Nv+6EdT5Is3ybT5s5/i2aCH5TsVwzmRnfm
uMLG/YVsfNeEw/72M1oi9Emr82NWZT20skBleH1cu/Y58Jy6f4thS3CATO3q1+XF
H9Ot/FVdyTRRiD2DD/CjQ2bFi09NilJv2HcTw8Pe6Pj3M/uhlM/sVe6XrYbhF0u6
Sed0X3yqm/rwIfT5xlDABtgNU68PluyddPvti7j1XX7tuWmKy7IJgv1jiw67vV5O
F9YH+E5dDo71/JhEhWGbh1irTLk6XEJKqzIjTaEbeQH5qbkSXr0Gtfqn/GmBwN26
UcopJLA+AXkeMZuR609+ZDUiqG2XC4xIrDFI2No7Dc55jZ3fj5Jel9rYuDi+y/PQ
DYoKMG8Et+5SokO+bpsL2DcCESlTW+wECr5AsYwyllhZLXJwjW15Li/We01Y/pKz
ykyKJyEENyzLd0EoF2455JPNFUDCo+S9qH64DGLOyANgUA8ZAj9A6yw+jdui0Egr
BBRaSxXK028PBrXelnQvag0YS1VSkL4QUmkRyXR9MnP1te3FA7GJRg31Udyaka1W
DCBPWP45qt8xl3036NH/GCjvCrsTX49TMfDOij3EAskSbgIpg7FdbwTXcrssLFpm
FD0hx2Upz2VTo59xA0zmHNAflw+VRhK70TaS4AnI8msKEuNMWqWMedmdqvVndC77
r1HrnfOvK+SIYUQWh6wDxH2B9+KKxDCYUshQaSZTuW4Wur3pmSJ2piPfGLpNB/jS
vNsvl7yY1r6PPioXFB3odJLs3pUonMlEVfQoD+6oRVv7o/ipJUxpJGfbi553bTju
Z79GLfc9gS4hrAQzzMffAi1R88JsuJNsjoDzHL4eFVXgI0JMpuSD4KKV+Te0JRzT
EeU3Zs+JOIQoQG7P8BJWPEBWp8i7w2A+0SFM/HGWL2hnEvSg853Gu6SaZ4g7Nj2T
Z6rvjUmnQXGds9lJnb2zNw8RctPENkEJJCbb4tPcrzfhbP02HZ5wIJvmLdhe9Gmh
5UlvfQkYyofc81EFEurO2GFwBNCccL5rhdCAjbMQCOfIwyCqqsJDpZqlG0gN3MwL
JBgu4uoYmjwj4omzQ8brCWvCjuAew4Blv3dbWQy2ZyM1JZBDz5tkZPjcQYTgMkkT
dAph2y9xNakRVNvJk+jh4/X9mkS1rJ197yn2qcCQ3m6OaeZUEnNGfpB+lEP4UX+q
+jbeiOkA73MY9sL2guxSbHD8gqjwIeZeu+LbtifuWRLlzbjD2Bi0rRTrFxrOhrjS
DTPU84auDE6FKHxJjxDwvKDIyP3kW9BhIysnCGWCWAYNG6Lb5C8sNoH1jBaqzsVC
3p51NfKbAKeggqUf1Zx5MQs73sPMzu5Bos+8Kgr9TQ5EFPSPDI20bMLUOFUjqyz6
/DQnj/Jby6GL4oeAWnVfjDpO+bIZsluRlfZDvlyNi1kusDRrz0Dv0gJJAquJpk0v
atTbRC1/AVimzQI8KZdwv8Tq/TgAf+g6zqRehkvjiT12loIjKv7n7OKxmg0E1+rs
++GDyBPmIZEaSiGWvfbU3bmWt7hOTWel5VhY686iKsgZuSmk9o3yQPRo80ljigAL
/9cUDxsV2yEMSzqylgEPo1Mg65OLRf5tG7rtGikoOUw/22hvpSR/ctI/GYmBpJmj
YB7zBX1zMPS15UaHSy5ZLnho/bVq7u4F0e96LGYtvsvcUWGQn0oOyfmz4yfVudOB
qk54oVLj2LBmutFSNlnif5nq7KXkYpnNwDRbPAYixjAsno4P+IqPzgeW9Ti3gSDf
9ufM3KcBfp7RegsscxNL49aZvj+MTHVhRJHyAOXP19MeEevMeyQSy+W0AYd1ch//
eKaaMO5Wx/2CBNQpL9IHpZ+XaGnje8n+46xYKjDJI9GpCQi4JZnlq30pIrO2QDFo
WXQ3mn5ZEhE/bOWeRiTarBCagsuIexOd5AJmXUgh7jvFPAQVYH3VnhpjqE2SSLAN
P9bErMHP8tM7nwKKV0rIuqf2ZrV/E/rUOd3m7KA4LkZAde766XUewmIit8VNzMIW
hLP6yOG5xDFEphE7Ds4dMyz01zQrC0p5jb192o9sbKBF+C/xlo+GYscEWVSPOSS1
w5VApbnEbC/xT1d73PHB4l+Gs91TNts63eEakwxS+J4gCg4uTvhb5PlrKXpOEvzC
eFtMzQn0g9uNsEawvPrkW//6HkTmNsKfW4XiIhVqDK4tjdnCbSSawITEo71DxtGV
nto7DbuowhX4fgOat1oLkcsFLD8kPuJgg/oL12AWLvsT1pPkrlxbtyQBjfsS4MNX
rWFJ/XaYNl4wpYwvdq+T+mjWDZktLV84Ota9lov3v3m3yX1ALc5RP6mNdJIzwFGl
I0jDx3w/2io85YyDR1bQiTfdCOqbj/ct06JZnqP8B+uYdHth6tikbVJx3pfxmyGt
e1P1esDA8ZxqxmTbGCbya64dIqya503lxpOrQwduTh1iQ/2J8CDGddukpwtZWWme
SXKW35hFic2g6ZqDkxd8GXoPKrAv0q7F2hzhsiYPRFc1EbPWVOMrRu1lU4fLyiOw
9vO2dgS2Qj/4U0RTdC0NXv9RFzIQKzB4PbHkqa/R8VKkFwQx1TXTD4OyLxAGKvXD
UjhmsF4TcfWWrNkrqeONu9HFKmhBarCy2mcsF5dcsqF37e11+aFLpIMNgmTglHro
/1HSTiRF4DHUSOuRLBds3MBkur98/cf/wr56RBYapUYE8fNePXrz41o7ossQ12JN
hLCDVlezy8kR9w/wpUaxSe5yHTixd4iS26q7+Dxq+jQYTvioxAVdtXq+YoMAOkLz
pY+gF5xwj2mIXHjkmqlFRBtbPhUaV8leLwTPe4sqj2tWk6bVRKwyXhweojUCZdKS
ZGtcTk3rDdAemR2AQnFP9HoPaWDBePCdPcbRSYIdcYCJm12AWQaJ1f9khHglk48j
TambTvgvdbffXr+dAcyLStqkJXHVQ8r3fW3axcKxhyD147P2NuTJskJ/OjyUvc6e
zxhJ50GJGkWL3zN6VhlQ5/B84hs2lid1w56Epl1nbCIIwJurvDyaZCo1mLa0rQl9
qZOsQE6hx1KyjtBafID2W3qw7aBwCjDaE5wRkH4u1BkSLTKbRN8FfEVLDf1tWtIv
B+e7zBha1GD/gMc6RLG9qcpFYQduRFciibDkSOsqVNU+VN1g93iwWf+Dp69NlBFd
Tn2gm+MnowMAclrml7MUqKg1FU90bRNTsfirLAKB3wMRSTqMCZg0EXkPulGA2oq0
1wRkCk4cVJzQefGis6Wa4QD7n17INDtYG5YEXyagwAFuyAsxFSVhlyA0ZOmFIW8o
uyanQ57o0/nGrt6g2q3judjnjljcBFLpukb3SfOn9ZMJNrNRXkIRIu29q5T3PJxt
e2FD21VV5/1eigWCs+eGFk4oWBcRSTvkJhK7KgnU54JsqGKyYNQSvb7jeybydrO6
7fSXzBLdu8X24TQtatrSW/sNWnTKIGd9xEsyO0JC85vALJ3h3IM6LcIw/rJdQSO1
9SJ8ftU80zlkBSPntnQoG+0oaRhrXgD6/4Qp3HmRz1nE15sE0vzQd9HqZEdw45D6
fzkB7M1dXvIhPEz1BY7v59edBaCsGJhV8lOSZn7NxCg9+WhpXOuO2JWgMxnqrqgd
D72Pr/nSeFH8JqUVeG7Nl6YZ7zL1CtykWxly1hTyD5A9vJEN0qjOHz0JPF2cNaZO
7ZrJIUxZggkWKs8g9YP/R54BYFsi8aqK0ijeBk3hvYmI2M2EB9l3CytqPpBPwNW+
mTDWKb1ZDxiQJvEA5wyXAjhT4Z7Bl4JUvhA06wSBPR/7hk3sEGlkaiBVq5wtjlC1
vJufMAcKS37wRWAF0w1fPMp44MA7L7A677riwBIdQsXm3tv7YfYwqRlgFNX1/0fP
KIlj61Foo+1//Fw8YRAQIVBciBDJW0zyHmnziGgultTzK4DU7uhCBy9V6tHJTXAn
/FEH2KgJyzCo4BvDXrnJ7gAmcecgYGJkZiWT4fwuUG60vz/VpMk8+ybim9Wy0cKr
AbLZ/WiQuTAOH/ZOIZmU+hsqFASbhvwlzbr0S39TiMcppelSFexRUTO4fGFhrw16
ASku20mfA8HTtB2gtgGJAkdKWJ9r+3vGXb5ftgS071HGOZF2/b27ZTGyctnw7QOM
yrzAA6i6vAWMy9levD0bzgvMFw14AYQtqk3dO8EXjLcyKhCcZ2lmaNnLtX7rdQuS
hlHrceVVU/g5Q13y/y9tGPck9Ryy8Ze3Y+1h4dfEPDn2wftDMKiiUaRR88ZHcx/M
JjdakECFJizfgKjujXqoVJQdSxlSYWegbY61e4eQgTkUi6f1RLkDZ/iPyyBGCnOp
i8SqGmze1Lq/rcKRRjS9dd2GZLGytGK8LhOmM1Nz1vart63XljEyEiYiPnA16ZA8
liYSKIeVd0fh0SNzF+3IIoV59Y4MJA8ULnObaQU0dOqOLvGwjhFdzjGKcInUTtpA
TEoVA9l2PhWapV+fi/KZd6iyKv+4x6qGuSF0nNfaKFVPEhAhXChySxIm3exEGp2V
F5THKAlsIVkSQBTCBdTCimzXDsEqt7ThOBNWDVunRTu7CtlSomxo0sG0FdudGFMd
swR24Vfw/MwUkx/3uh1OF0uesyMzWkLh82ne6Dx2W3akDBIeIMNnlKGCnGqcHXqw
dmTthv7Jiuj/v2SvIL3rkR25R8zkXmaH7Am1vITo+9G1iXmVGOklPP2U8L9c/mop
MtT7EFFATWHhLqWQ/6UmwN+l1VEpgeTtOAgN9fX2fKSI5bmWz4sgxAOtADkckk/Z
u9v/4mUdoXVQ47jPVRP1+IZx82fbk+rX/Eru7xFJOfxaAMCoxk9XuLpyCIOxAbOq
JtqM1EcW5CBN8Yf90KwgBJOsfJcVDe6sQO2I16M6tQCVVjU320KerFzosZICsJUS
w1s02bMaO1PsOPDth4+pcbawlt6zYzz6y2Pm2aK9SDNR8PL6AA2XBX00QNYnvRW4
1RM6brnSmoI9IMl6+j6I+/egpOuKpqw8nYgPrl3URG5Xi8onb22xVXekL5A15L/h
9nMsU7Kpbd2dTxLDNhM1tae1rwmvflViE7gGoXV7tiEY4cmmiPQIyauv8rFN+Q4c
bLxSbhyQAnBsOyjrQxN20ozMJAQP5zFsLoWeTVdhUqMOOpggHL+RBKB6HMnNPmLN
lWnmPWTM2P63ZFGUBrBFx6FhWCTLW58Az5zJYVsmeIWzYfCCktpKWZ5NqCrincEB
p2M+MLJLxJ6V25qi9lJzkPiUGUwBe9wV1ZQgRhvp+IIA1nV1vxdRziUbPmaRfewB
8jIosd9cQasL7mqDz4XwgpOvHOEzlT+YsehZyi1cwcW1tAQ/cnHX25+dkq4qHxrw
S9JpyklXNqOvxxtK/amnobTHfAqS/LRbZ1TuWwGcGllGBUerOvF2KX5gGepXlth/
BoXwpMrWeCof6CACExkyGfnYRHTnvjhPjssY6OtcLPQ47vpo6ISAPpdLQx5yV0ay
Apoad6MHW58dwO3dS2mug4eqQMRgyh4wBT1g7RddZnf75aIhamw4zffRg/QcNytJ
BKP8LA0bPe7ijclThsrLXKdfmTgfxLHzKoMyF8BI0yAxoEijl8aaHRvDnf9Blk+a
ig0XvYkq5E4VXWqYJykEEtcxhyIM27n1XbSutsKfekufTuIlebgzz8NdZswhyNPf
a8Z5s8ROP/NxrYBviddlzCJakZfsxFh8jJSHemp84+Ci06bb6XeB2BnZ2D4NsA6q
S0z8ccmH/Hb4lbrn4asDnGbcl//AWIOW/YE+whtMHnY899G8lUlB+2/Riu2oPPSN
bxdMq2+uyguJMZfAbBQCcCZYxEsZ9/sK9wmOjbGHt1MvEX3Aj55GlOEWstkUd65Q
sBoSxIiuiPxjrCArd+fzGivKGVfUuTFASscqqjdzlwpGxk086wG275giBOfMltwg
l3CDJ/XHBdFCm6YMzUJM+OydAcXXQMdOQREF2bgU6YoU0xeIfIL0rpSi6QNoWRVF
BuZJLugikFPrQY12naEl8WwpgUSOK3sdjjszG6EtrZo4pUx7KR4cEUEI+PsM3yLX
JD/Ykzn53jbrxY76FRWVKBEw79BJo2q4q4sQSV9MJ5PCK0JJ3re2JBy/z+Vy2XuT
016b2g2oHQPW0MqpxdS7MyFCRHzAnrQZKUOahiS1xiWmaMZu2E4bm2/6o2tzucXJ
piSFDQlj7gGyO9wVlzp9AleJ1kLXgusx5IBzjIHSFMfFFkmNMBZ8M7Di7FhjCdri
NawbJwG/CzQ9B1Vm5QbJ4lpk85V0Cw29XLnc7PVU1ehp6KQmZKxT0k9o10ZsC65O
KgzCoKn7i68nq5tl8djEd+ibWWOc+/3JwzUyX9lv3N6aB85c33/1oAg6Miwpp9qF
2YQGNNCMZrbvLgJPASnfTSiH/34OeMxr+wcBLMIrCYWobE674l/WUyH06D/PsGPN
rjZytiap1ZZNtjt51gIWBFCSbeUrBk8FKIgcfF16wG99mNot2YZzH0DyMNOA7bvg
Mzoz1kxb59facYyiFTuT4ifXaCxaEjgDGR/1suc4MmFx8z/ZG85yd5nfe6ZYXvNL
6gOy+CSAieeNe1zIwVUlEAoVT9+d/bEHS5Uqv4sJ1pP7inH8pHCEXOCakQsscdF2
oaKqHuguZt74IGhsiVcx7qRdVDSVEVXmoDXsI1zw5pi7yQPbzzbCbsvUpxleqIZ5
DXwI+vqnZROkesB/fwtrLe7hPqAXSNjtXMNy63/f9yAAF/h1nx8DwFVgca3zhp6V
dGzoqxLLi1yb1MmAERYEd8oD/GWzbzOjno/FIndpRSWLXeYq/xv+0vMHrOFqXhT5
/uhUK/S0cFHSBPCLi7MkCLwd8R6LIqaEUuX8xHm7DZUidLfs9Dm4FDfKhNaSHZvs
xh2MqYkPWrcqKlpSIk7iMjptaaK7XrXeyz44l8PZSl69yeLnnoo+GLuzp8ZIuhmS
UhKMwCxvPwwyDJL/xasMRyXBLuNq3l6YFNGHdtynofG9fdZp+OU3tTvr1/T9i2I9
R6/ne0mDMBgQ5IzJ5FJlFtXKHcFC9RfIOo2FGvf/yR88/vU33TUDOjqi4/IZZL48
jvEGVMs8W0cGDsEk9LnSnpRRxcMN3JoIP6Bq5JNM1p6bfkeA+E2avhKpyWDW8pPq
7btTp0+qD10fx+v3W5fvyfPPxDcLFL7RHm9rPxje5HELemlV5w5jMPlZk/a6ImvZ
yid2WxmGQc6frtqTdg0wH0nFwMLkwYPayeHq+7inqa0xGKewAM8Wqg4K06fktyyA
IL7hmjU4P/cFa4FW68bnT1GorqRrwWCgON8B4XgJ0vsalyJNMQuiRlMJo4HZ8oCq
qVLeJlxo9schgcWEk6WB5hwrFUd32FWP9El35a7OrznmBa27FRPmJQ+26QaTTsGN
on2trQ3uRcBvI7PCOIekWM4b3ky+15LJJARwkLe8Em+Qn5l7S7bVW8t2T+woNuq5
ZXkHQ4i5OC4DIPoHGhURwwtPK0UCiSTKinTIvGCVqC0BaUWkwrtG+ZlxuLY9QhV0
SDQyNfNPkk7GowGlMx2vMvkkZpbXR3PktfblBDYhJfRF2F/DInMWdYdvdGwaiTVs
/6UjKcwkGSiq/MSsa3IYx9/4V20F+LBD5UHFZqnVqjhoF937yXN5OwK3HMYnNqdI
KDvrjgN3exdQrMD0fgNwAtF3RJF9GorEC/xu2RERGcxF28B78NwzLTcci3mJqSDg
2AW061UHR2uw0Ewo2T5FR/41Fie6HvhseimGmdrl1t1AOVHik6616It0CXti1w9M
qva4kyLl0xkuJ4ClycnMko8nUlUNmMCo+vyqm9jW3JSu2Bmb8U8gjKH1BBkpWia2
CLzU0dacUmWxFFJdEJ5WMsiYVzpXxyvrhfBIJbQTMe6uyjwtUAO0Z/wgwOC8aEg4
QvgJjyXYTWWympB0h2phGqjYfZrI3vh4koneMplc3Nxf44Qs5zCwNVIvz/7Bgi+f
gMXi3E4fVs/EB9tVw8/iTnEu3sR4a4Ja//1lzyi3Kjo/Yr8vIMqfkZcv667KfOAA
1bMy28h/UoUosU1JHM9rr6pPVOvBy3bUvFS0g9zdhowmmQzgTICWUHlzX0g2SvUp
r3pvmSYG9xtPdLKdfB2/qxlEcCBE62MDMqt917st1AZu6us/rAv7Oq120TUC1Ssn
1wYIcyZ2f5WZQ3ETPsEzBSCmD2GEPP0PHjqdfgRurnG8Ge6cWRwklGNkPTGsSZIn
6k+ngy9cY5JPQczLuo3pFj6kvRlyaUis0+SA+WrH70OkBaeJ+JvJSh+M8IoV88gg
3IpYFE++tW8B5WID7PZpzzDYReAPWrzDzzhs8iTKjtsCPstzvhsuGBlSurfulht0
lj7LNQU4lOwIBMbAbP5hK2rGjLGIeGK4OiSdHSKPQP9WC2WohMYdLU6IueOoEfne
YOj51GT7iGMDMZd4kg8YPOibdO55G9rLbzhkPPVVdbEQ9jZJSqvjVDhsu557++2d
PP1ylSieYdNO716Dc3QeXisiGUKkHksbFBh03mFCqe6zIrJYTJvz7yE+AvT1XMEx
kap/124hj125DBFybyqeNjvD4UPtiY3zmrdAanB3bNZBGpKaaV1MADc14rjx5aoY
SLWdJ3G6w/ISTJaVpymkewZA6oSC0uITLK4BNPDoeSm8rcB9Ut5TJrgvpRzLLpbc
sgdDG3qMpw8AUKxVtTIGuzAAT6ExgqIPFpMgpr++evOLdvEafHAkZzkrfrYE0/UM
48CqnB/ndWNqejq4ooj4FmDFpPUMlZNNa+y0B2pMiDuY+WrXaA2+c5TctnzUU/S6
8L2FxAHuws/7HVU1olg3F7bfCEb30R/r5otHMzs0/R7idr7CEkwZ+usfrob7TSpg
mQWbEahwVFJqsi3Q4hsb7gtLOHOL8EPnzx0hP3EmvEZNywhL9E8DKnHWo981MEKI
QvyNwcmJ6x+nY8WmtDyXjiMR4F+cmv9K1kCNcT7SJ8MmFQLb6e1HrX5qLvZ6Ykqc
YUXqEBWfODNTDVdCawOoGCVwhtHJtWszoVkL+IWfK/yBk86MYMfcnp4T+9gd9VSW
vi0jg8xIeB3pBMUMXnCCWmJmu+fiE+JuSdCkKQpiZCFuoBQDtwP362hfJ0+j3yR6
5MzyRbaURm66GxL1pOnV/W29sH07F9jmYmNWJQeNm9/v8TMBDQFsIONH0FR7T20f
MntxsKsRYQdvszK28GqSuay4tItjUO8w2XyWztu9nXTaUavee0pt9o0aBhcX990h
o4p921Sd4y+oCtpedSsjabkC8uD25C9u3b7fKMo1KeKPXXL5jMy79zcCZ/6dCs29
kpdkvhuYnPfEucjR7FNcU4spwak1YJ0fPrkukk0FlZEwn+i4yLVpg71DSlx0sMrD
hvhadeGWGttJJtaIgwjf1uf08KIKQ9PhnvGQVU+myoYKOdWhcNMTNpTDRtZaTPe1
r0GEawn6xTxZdyJFtTpkZQfaMIo3lYF3vC2F/ZL2+De62GYVkDjXPbJHcIu8ECKU
qYZtnc+eEVpk8Vju0cR8hqMk6amBLenDBPMGutKStW0XqvFs9i007apf+P3MZ+sA
T42vWOm/OUHcYsLkEkGS5YRScBg8gY0mZ/EbphPVBRw8PqdOQVp/h8TW6GAGMnvu
dHZ2cH9Orbo42ZCjfYwfP8BqYgBZvfx0ndfyIFrdpBYQOTWI38oRyvlC8spJcfen
/3/W4mbCz5P7sgxhZPvUlolV7i9noAjzIKcI6YE0CtQo8cE73F028rswIr0y6pDg
ZfzNfqcaTkcKZ3pjzwraA7RZmsO+sFfhzZNxLSKEja3MG9E+9xztIKZP9bLTq3ut
ZMwYP4XqDdlAS0MZFXdS+DGSoDDh6a7qzRtxwZGUxVnFnCXZuIlwT16HJ5fVw9vu
85wb3ZstUjE9tNp2tknWJ296p6vZ/u2j4xtIHjd4mo8pO4KqvN1b3F2Bz/rxk7A/
3gn23K5n2vGKQyC1mq3QDNyVUYHoS9Cn07Dl/MVxZLru0k1LQTzjcMbTXWG947YG
SFVqnbKUKfrNqlbdFyzxtLh9fQ9KdbwDmhaAoATVxWrmsf5fFyJOWkd13MJNlq4c
11sqMknysEGpJsSGMFKzYzpif+Lq7YgjwV7cafjNKvz5aXKn77YFCwPiWGMgIpe2
1sOWftA7t1u8EQslFVXWDmqj1Hz33aNkS+tjKAsdV6RH/rC342sJiO6nZS/AhYmN
WF8YvDrwr+vCY9bCYuAv3LMfsLA8RgfUQan4FbN6n6TUKy3wBH8fvYC+g+0PXKLt
AyTVM01+goXjPC5sjXjNpVH6u5QKtzRB9X39d846Mp+0Kc1ZX/O6jgnZDqfl/HWh
c8kEAJTsEt7ltJift+wv306I8sflm7dxTQtdZC7LlaYOyRuuLSfy5T5coDPVlka7
hkBV0PjsHAEX6z30dbXJF+4NdRg3HuBnlyiJRIQgQ1kOUV6Gv9zO650fPCR6NkBE
zR9aWgpWKiHaYsUjkCAJqmWj8/qC56IlBhnQCq/Utx52zxKNgtlhZExDs1Rda7T0
nptnMX3E9uoMcczmm5VvcpXNGq0ZDQDl1OPhbi3dczEscrccd7sLkxATYRmpdQqb
h8prrvaRTg5DJpsx4zNV292PoksOld3vHEM/BAroYH10vjg3CLok2f9YmnXolxI2
Os6Q2Hmv2b6C7IX9hrDRGtQsT92tJX+bu5tj6NX8komsFvawEzSTYehgT88lfrUG
JtsHWwkSB/6ocxWMOuOBvRoJ7UoT8FCV8W0uH8X/d110j7fg8o+qhfahDkAbO/PX
HlEVml7j3qexPLyof9uoTncg401NWZ9N9oZeHmmZ67ul3NZr65b1E31u1DyGyIWS
OrNvhp9aGdl5GbFF+tbec9qcvhZPdWoWU8DVKtuX57s6oiDCSZrPz+Ae/afB/Dmo
uANlZ625xNkVudT7jQoyiw2McPMXkunj7a6FLdYNAtbbZVFO1pV2lG+LGqEmFegY
X3fbrMjpIo09Pawj6TYIGtug9On1ACkaE1N42jQvosIYdX6ZvlHvfRKSamw1lEmt
ZlT10CaO8JPlqEArIEVgtSv1Dp464odOb5jN5ZaEfFzBcuEEHYJ6vdXzUb8OL+Et
GTc9h/EEp84jdxLyzvprYBkyUie5ez1rkMyLaUM7ROzZsTxmEOyJq82fUtDWFDCy
kAjeBHACk7G1dzTpM+qYrBet6LsrPcm5iZOSp/dFVNKH3hxiaQJ0UpzmwAylGOZU
wSU2WqlvgbkmumjlngCbAuczKU6YsBlRzxjfpTqk08G5ySIcyaUy8kz658mlthn9
CqGJjEpL395SBY++yQcDv1fDZt0PhVCmVsNCBKgpnO2m1NrGh6myHeQRBf+a2Ayt
E1TfvH2nAO0l/fxiRDVF7/Zrkfuaj+qRzoFfm/sKAf8ZGXruGCWrOXoZE6KE35LN
V44zPXLTRKrPECTprp42xCxa6E9hDKLgbv115v1u5EMjcA6uovajYJY8kRNG98pu
2IS30ymnF8pjpfpQV3+EN6QgHVGt3da62OJOWdiZl2ya/nnjdLIDYxyhatyF1ET2
a2YKCe4IdEFyQKh4rAIUY9Sl7Z/kmjeqKJ6XqIq2drPsui7S3tMwvRF1mkyFgTav
b7MzhaRAm0Ty74nOLV2rNHCj381ySYNh8H4UfanIPjnY1e2OAulZWXs8RG2EkPqJ
Bb0eO+4f/SKU2chkh2u3ATZwlTTrM2SVPN+y9c2EEunBRuFyvl13P0orI3vHQqSq
oI/rT6W3vOGX16Lw6av3FbrEbGEfi8h7+ZhlmsmdIdwxzgM/Ua5diJBB73tvtsc+
Rdfc36rzCmAipT1rZ3Yc5ya9RsabavLjMyCs6+RSsMJDJ0zhOEpiIWmZcz+HOpnv
VZrxlTPn2jHZGd5dPsljmYOL2oUOt+HwlBiQAnqTtF+/ADSKO9aL/CHNwTAsLbaW
34eVslbRsghP0mUbqNEEN66qjMhrYf75kxtrFuzdVau2OWX840jDYP2ak6/ZxmCU
nGgymCG/69AhzcTH4tumTgoAoV342fxQ1vHsYebxYb4ZmfcpOZArtc6VsJP8Np1U
Q8WaP8eAPAiIiid6m3WYsWLn6Ncxf8+CFPrWFx90teI6Lr4Xg0i3IZRyi6HQ9BH3
p0d3y+KVYaxAwt3cp6msdZbdPGhk/5+2Zz2c0DnvnOnfjl1wHoy0WGyqcNr7g181
lieoHVOgi7R75M8kqLt3I00sqmFS0hnCimgqdJm3pG/8lxHX5wvOhNknbZurPfWC
kYaMjtAitByO6peFIfiWBiYs8Wy8RapRMeg2scYA+5alhERTisS13ci2nKwlYKwW
bgYIAF8fU04ERLpKYsTKq3bU6buNYCdUB5DdcUsui4ka72XRbDMdlxZzK34vx6Nm
Jkim2XrCKJ/wDxhvqrVjF9rEzRswGXj6OJQVZRPcKdF+nthUKg7a8M9U3ntdcepb
8Qz4EO3Sp5mN4TCAyIf+OVMpuCgMExY5Y4BeQbIlLA41xXaOwwyjzPCUw1lW7+Wf
/FzRkOChdd7OsUhaLGO+tPSchtr18iXrET5IoBKvFH8CVDo9JAYSLpcZpYfMnnSh
Uq9rMQKmlPuwiTxQOeRXB8k/zVoZiS7wQy2YeIXK1q39/mctAum7DY+/1KN93dmg
x5aIDaPd74gh1tCHJ7w1GnWdpoeEk3Qzjd32CQN7Quo9jaCJtTdR+FSoLMBJu8GD
Vq5fu8T7gUWZdfbFJJxyQ4Vax8Phg0nLyYv1rKthvrIKnvBrvQQqCNBSD7vWB19/
DMYrmMhVWK2hj0uMZl3L0B9kCywO+JVhL7640sy/LoTQmYaA/yhq2O3rggdzKlF5
ZOMCL+ZpCbryWuXhpzPxYt5u8ud169mWVcZXyv2vTdo/okwMTVq1Pe7Gd1JSIz3X
sacVqTYDd6iqLfl8Ve297d7ZmtE0yYMwk7vVBd8U054L/G3EXlCwcjFWV3IlDrcj
OsZpe9Zss4SofjrLtK2yg4xIc+YhHmU7q6Plz3Mv5JaQzdgTbUmuqZso4wr1lDUQ
CYj4+6z+fk9Zx66UFHngy9w2phM9OKnaxnxkYY65f87R7hGKeviBWpqMW7X8iex+
fPlq0tMNByydRjseFVWxDLJj3ZUkrDE6q3h/pMm671GG7eFhK3qkzFQ3soDQD2eF
5EHojOIdPD+DHy6w1bRyeLgONz8Jj/D75SKjIlEVqjlYGWBVtdg8XMV/sVY+s1MK
C6sey8vMCAIWdY58yoOODdPw/GPEIy+bHTq6Cm9s3s1OQVSF9bFpi1LINZsRMbzo
kC7GUfjS0UbklNgVJsrsb4pHxuO58jljLJYMm2Ttu2KloWgY8vjSyFBMmRbxjf8M
H2gqBCJtR5Lxk8Gak53mgriHx5thRs7CGFu7CLE9emixAy/pnOskC/hp+AC57PFY
ht2HSSeWI/So08xFi3uBRr/8FFDtFGCuzii93Wj1xFls3xt56RDxKnd1DVWznqut
FwQ0i2zG1eeHqUy1/2pA5KwKNE2jaVV78r2S0tEEwi350YaG+x4BWGtfdmdK7fZC
gwPykhb+K15Ki4eLGk/Bts+cIORiokFonwdc7JJBISHAZFOeE5gQGXorynILSz92
rUwn7nT+cuoQs+8kYmtmRTal8RQPNumuFhFuR3v6+Vwdkg+cl3keAljKQW4My10D
0w5JT8z/xPTd0dAZ6OUNFbF9l/suFPl6kGscl6jLTU6P6ihYWNzDdR9A+ohQ8aJf
bOvlhGBSVhR8Hk2oIur9xDtzYsFAmf6efgK/ClWIaKQApXLZ5D5MLEXf0+uNjoBN
shxIz0rbvOAQuRYPqOKjJeED0vQ3mTjQvOGc21xWCwD1DzGsm0XBChrltqEw2bmA
MiLj5X8x3lB++bq2MaC53MJ2loQsjsWmtDQ/4JIopwGkeNXf2XmcWlwpg49eh41q
O+C2brjvgbASyWNgYZQAm9oF+7KkQCSjkMBaCZ14OGARmpBy3jfuZ86MsfrG8yf9
DAyw24ZOlh1FJNzIQ8cjgHTFTJlmb/Lio3ZjfeJ5aVXCNRhkiyrlnKFWKK5P7HrS
yj294usES5RdQGf/j+or8KmHZkV0eq2/bPr6uhefOME5CTga0cATInS4hYgYr/JI
kmVzc1Hxh05h351CbirsgCUSW4jgiEedYRCW8jo4Zd7sK3tGySF7jOJfYx4HTU5X
8AGCwf4wSnB3uRhAiJws9OI+tZsf5ErY3VvDIOLwz3dbrgOJ0AparC7wLNp8pf04
lqqTnH7JvXEKumEweZ7D12vMFHrE+fKM14u3BVzoTv9z1sIPb9Ax0PxdE9/c7j4w
X24ttbql+T9ZAcGA1o0cD4QKEnoiJETYjqqeYrGJVpkNYPQQJtipn07y+lfeT9Dl
bH5xLA6+Qf4lNxQ8YueUorCS3IPAU14Mil6bxAJc5vQcjS+5/5TV84aKmVyh6M5F
Ky0QeC6et1Si05sBgOZjBuRwvJc6Qn40IkfD8XmcMFw9tvqPiG0C0Rw0+r8p94uI
uA590DxorY7rDB31AFp6eahSdNv1CHO05nLOqvhjzW3ppuAkE9Tvrk1hJWOp3qhF
qn5ZDj7NYO6kr01haC6LJXv0wgdRbBdXguOC20tF9e7xb5fa44eqrlSGCkdNNvrE
QPgsxp/k4yTfJN8K9Y+jGbMBxL2clyNjG8LGBVkAMDfGotLgWocM8vg0B3uVQ0XP
cLKGfmPqaYkYhyNKV9AMsHOCoiFq8seyaEgX7Ck4QaXC+UNLn2H8eCbCKWWad07d
zfe1X0NUqFu2DO2doFtt8GMOpixJKlB2AiNsXral8kvmjPMGQidtDbIrSUWv1vLM
vImQJMUweM52eI3t91J/ZekQKh4TlPKeBg28bJlAhfq+4IcnfGIwta6jk/EHXcip
kFjlsahADg3bnAhTFZaKzD2W2LQonAJb8zRZBtP6ZLY9lph1GoWaGAtyq/v7CitC
tpvtI9CO5ZIsaI5F3mXrTMgF9kycWm3wRUQLeIlTaeNNr0RnCex5Hy9JkvhVlq9D
YUbdPddclEd4wvy4LISzVblEnyrgqmEALfRDh43Uxnz8dn5d/j0qqMkS/EmSAijE
KqtVP7tgIBizfk9woR4VM2wWTD1nwsyZg5lrkL8+ogB5BHL4Zths50AKFrD4qUPI
w1n9QSEdIT79fGmTZDmpRA2ZVF/gxV4qPEi/L9rtLywU67dWomyuPAQzR9bWg8Vv
OqjkxgAsTpTXVsqjvdrfrFJJtsYyfwCOnFqM35P2PVZ7H6KsV4HQN9I9Sh0GyUzz
A9VmN1lohw2zf4+lWyc6vAnq3j9c8amsXu/4kyo5XoBPIgRSZZGiBb+09yvlDDwZ
rT3VlfjWFu+bPWRKUGZpxDkYTVnobbx98CzwzL1sKbGPLJnxNqvRKjzDR/E+ldVE
ai+0CQZqRzekbWQ05F6qKPGL43do4eRMcZFx47CdRYp+miKYe7xKKTejdBDj4pz4
60cp1Sofh7+c36OcP4JY70MpXxupUTyJLUyB7k1UbzPLZNQ5tHeJ3OPCiXz+L5sl
RQgBRJnEUHZk8I9QftW7Iz0Suxmxro5SjhMJGvuSDFFo6NPdShiNWzYJjAKM12Eo
iTI7QtqAa/Gt50OE8MBz50TuW42xF/clpcKwiYrC+qaVnzD+hAhvCqhQKx5vZ3DA
Grk0GkaYMz6sozsTbxfC3ccFPIS1jgEfMgDBk8Pl5qClfg7Li/04MZ45N6S54MqI
acRJD6X6Tcw6/kCNOQXiClAqjF/MVqk+ggDwHu87zYO0qZd3mVtUpZpvlQg+aklg
FmpeeaGI3pYUViuyoo+vfyzTPFW9TvJ82xW9z+GZ1RH2e8k+EAgDkDjMrRJadFdD
V33dUoZFpK4JlWtsC50Yog6C3HRD0ZTspcIhtnvNAvSdNUKKq+VCIx9ipYUjNTlU
pEAHa6bekZ5CHHTqzgm9d8vF0djsV3H2A+VocJlfh3ACatFblRFE7ULSSAtO0Z7U
u7WbMg8x8meSfOK51a0xrSNewsvJ0fMtrFwZRxzVeHfpiWrIaqZjsH4vEZCz5Uma
eLufZlomDncaIV5YXv3y2YlN3Uj3xniNLr4T8hG5LZMruQ5oeImB35/FpJoOs1O0
zcSov383B05KBDMzK9xlFwvoHvY5dUDUkGnk+cghic0Hu66A6La/4g/aU7/WJtdR
TDx1RJXVYqvqAVEdubtysTByR6KgtYw0eKBsjGm0HhXNeU4+inUBG9lwZLreCARD
wAUWUVTryL3M9uXqzbn9pOQkANQyLwg1ucPlPsTFGWQlIXmGom+397pD5xSxEKW4
Tuh5PXhh9w0TXfamQQiLFeCgnvuGF6gBPWfhvN8157uQAx8wUz5paJvcCKrIrdsl
auTaO+8kCEs1EEkzex3EETmlTo0CgBRLBkYMz5/W3I1Owl7Hx0tYj3IMa6GQ4eRa
0g9RDB8OCGkJ4fZE80Wr5bAmq96z3ThhOjQrRenk3rCjW04AHpYiHKX6I4e1rFHq
WxuWGcpuMjPOAceWQ7nk9NQMG2C7t5X0XYgaz4YQcMF4EntkWAlGBe74WqEdghlf
ycl9yguNDc2YgVHsyzxBIbfKxr7EzNfgzSgKryxYThElS8W3Zbj7MehabF092xky
Hh0lvWlQbzQb6HleGhv+V5RGY/Gp5WSOnVTQtMM3Ji8Cy1NrShoVrBZ84XTapBFu
cjtkMugOHOG4xqAno4XIKej24lzmyUf74eL8ZsJ0shfyiZ8dLBrRVONTOOqES+ov
Lv0TfWpATFumpppIFdvnxBJTyY6zxLNHYsu/wHnJg4HKM9UMuQgJp4A32I9pC7XW
5mFQu46tWwq3HCgqeJsGMnuK2zb7u6OaNNCllxB0wMhkquTeHeuz/PJC3xEJWIXI
wv1Y41P3igE5UHyopxyawr0zCkNjt2NBAZVe2KIkx3aiSXgEJZcyMryKjfhnj0vz
rs4SbmWFDgvrFFwf0PfCJShmsrLGUtJL3f5M0iq+ibUceRxu2ofG/W/zmWjoKNRq
kemXDB5LAmPwR3x060WibqXnzjfaRcZ+rtq9t+dyYZUKJu2EVQ0AdCT6DA3f+ddD
ycL6fnuT63d8L6TFHlrFGKl6M8oF4POpDVLghvgcd1dGwbc/WcmjoLqC4F5S8+NR
FYsH0JvW5Ayg7kr+hLm+syrmF/peZPV9OngLNLig/HdXfH3y1Em8Sv/5Za+rGxdt
rhbU0MULlxkyy951jpI1CoVNKX62QT7rdITxfH4Eg0YrRzYxKqL8w0CGbOYmObma
bXQ0ETeHEG1ujeOlsyEcXXAs4pmAogkE/H8O1FIVZpQR+7X4qiqF1tfFBTovCHdh
XcDjQtXqq/G0e7rNgZ4BfDzvoGpKyQ7fDiXtNqUa7xHbbPJW2vhFLiN8YyJq77Qd
oT7G0qaUGNVaB1TWpP4YckhFyepdvdLW5I5GwPPLW4BxqTz13wzMw0nK2qtEI4Cq
8T5nCtbdy2yzDqg48CWwlLYIFvIJpR9X63LETFvtn7414G/CUcdHBbhr760tXqUD
GrXSvQqe62G+03qsZxgtQatiTPHxz5FDtMp7n/POmz0sAH7Ne+I/e+GuyhVLOZB9
uBS7JNP4BwjznzDUCsTrMhrimAnOCwrzPWYQwwH8gHgOt7qkjVjUrS1YWLUNwD0h
SINwCzTyV6ogucYdVFq/RIQ/4q4FEctEdg0aujhehvFVieRepimIz8dmCCONmKIv
Ca21rE+RWy/DtjfY0buCZOpKqqXWfKCzr5BAXfXaimJt5/3SHeA5tUUB+SwiRiRk
9bTo9yY9XIXjfIM220yowFx7bpkD/8h1F84SP8xL7rYFcUxusbTXGCUODUC3vAT8
J9GgezxEeaOX58ndKaR3mFhw6HSe6JatPcWb+lH4qzot53YZ7peu8QK9V5cxkZ1b
1JqROFnKp9FjZRL+0qWFe2suKDVdJ4PtjU2Gfm50iTfZgyV/QIKrWEx1r+LAV5sC
olgzOlG2MYf4kXiQK+RHcedZUc2qS8Pp1RU2v5bf7qBkNAGSPL3VIn7UrMMmMptJ
Qjo4iDTuPehdAMMoNjegvgGNDd+zsDsJcHUULWjIbiCLZf9GKchhV2ojyT2PY/cB
oxDcdz5XLQoZhske7fbGvYJihrKjG6c8sbUFfOFKUCw+zvLILEUtmLta65uCtH6a
cXSDOvmSrd1Ww8lHixmG9Eil27DeI3xjOIj/mPX3MFqC5h1U/Lsm2RJ7iuB/xzRc
Lzle5QN8z2dV6FSmfLY/SZnFFvYbDCxtX00kQenAy9/++LtYz81IC9HyTwf+kilt
EQosu8RR85lHuxmprmiAFhNxpDqGUsIOkP4CnAgsy0EmgvWT6xXJHdPT7tDhZn8J
aUjQI7YI//AvfoXT4xgyFtfF2w1n1ktUw1phDNanMt+z+CwQcOiCpkTysmfNMCiL
zVMYIM6cwMDSSny8lMhJxzWaluF7DBnpiM570dIPPwPyDoe5OuG0rx/5zxF0Emo8
jmQZK4btiLxHQeLBjKRtzhJSbEu4UAc49DO3X/50Ilu2iWLx13rspC8JOQ6/gBdR
15VhNpcbZbIoQWxw0Hf+36bBcvaVdw+NXBWFawzxY2/k1+juiKH9sHBUBMcV+NzV
1EZaJuQBYRgeA5379e2XXJ4RNC1GsZ7erkq4Lr29+iMZnyvEPXQB6sdiLnveqQyu
wAZqsUc2Qw8v40MpziNyeaqMwMOvX3tNZxn7hjeXEliJF8Il9hVCUeiTJdiKhbY5
jJxW6Hpg0FedShSzO7bI34D09LoEgxBDgXTaVvTqT10TqNxnzd5ZeQpuAETPquEL
HnCqxQfXfUSiK4SYs/7qmSC1zVW5I5zZuQ88oGHa9oH8Db8DHWquLNVwFJ6nVhpc
IXvfBD9HulTXa9I64xOfF0elE5rvT98fpgqxwW4RMmwlikfE21x8i73a8llZhhLq
NZNZd7zJPxQ8D1CI9/UPatdfZPOVMLdCka62cIH5uC/J4CRDVLrDen4SXsdaXEJY
2l8B5u9SqxkDcPxmTvS7oIlJH47Wy04Upw18ZB0q9JFh+6ULSGf32UhvnoSEwScw
lSyDhgfh4nCvCQkJ3DemG3y7+4MBah011rbAXXKVoxnsRY44DuKDVUxa5zEZ4GXu
f972+SFmbu8KBbUizB/zjW81+gycOsmfujBGqbgJa9Tc9hCQhWlxjnT9lVHXz3pm
RPAdlLE5xfvPQIrclibl6RYFfmG+GnFScclCuTMwcha4BKYxzFueNpqb9w57MgfN
rWKk+mBuw9g3QdS91JwP1LowOL4EkS/uLoCscgmEjl7xc5TnHwW7P6D4R0Kf4Qka
fUXGkGkrSdg0E3Xo9AnDVWwiAcmMTjFoNQajUsD0FTEWk2VTKrvWEMqYse5TSPEG
Gu3RvQ8z5yj4IGXWP52Tj8c0xC6+DvI+4MtaBKxUoxd1ObB9iqLL3cjSARcZfHVt
VDGHSIbJsR2DJv4U8KGWVMtvBK04wWJ8NDwJL9TzmAH00wILdlhuPTW5UFCJyzaA
`protect END_PROTECTED
