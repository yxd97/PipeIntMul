`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vYdu8puB7LAzpuVwmjknXlFN4phO7yt7LY8q2hgzpAuSid77PYwq+gVUygz8RxBo
atwa0ln1XQ99agLpSdFiC2/RMZ688FmQVeUUAEGKeNX7Sers8kTDQNHftLk3R068
rwpC6xkswiZ0AoOFqP+8z+KG8svKE7LqLnVCporUxrDyxotPG/1dEYgZJZbAIR9H
o4gty++waKUpHKrtoLP7nSwmaEP8eB/3BPbwCU4IEjg6ocZAZSOYOpues6qbg5xV
KLTlGL3fEUs2SkR2Y4JzRHyNb8DKt/C74YaHIggeh+m3yxgyfdSHYCfH5sF+9nBZ
S3/LMNhOBrJx8vajNaJVA/Gtzy0S0hhty61CL9SZnQsnqVaYgEoyDT3nZJGQhc4A
8XZpQ8dgnJiN+rRrokGFLg==
`protect END_PROTECTED
