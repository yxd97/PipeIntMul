`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ocbKk1m+hHEjEKK+oX8dQtBg97zQdHsp72PG2QukekxgERppEoaq7crlZnpdLlC
zq38EcxyZqxZ74PRPAZdw0BtkLiTQ5FjjnZtebCOPLotlm2fo3i3BOzPwOyziICr
pbHKB6F75Dp6veOGK9WwakgW2hEZW5HF9e3svCQokarVwA1LRvpVliPAc3XGz6nQ
o4WqEJ+fIPMHJ0OHL53sq41Bfw8Q35Rx27DOwGEfZ/ZW7wgSYwlisZ2Y2gt34i6M
rKiiVCkKp6x8h1m1bZl7oNmvL4kpOAknN6dpD6K85RWe8JF3d+ooQKlIWC3iCHre
m06vMukhrIVbn2fSk1Rcuq3I1x0D8lnscKT6ydp1ZxAX03oYH+gmgCdL3Nu2MVHY
UMKutjqG0HKVGp+1NvjKdQ==
`protect END_PROTECTED
