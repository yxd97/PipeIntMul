`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRpEW5izrMqzOJHukUuU14BrA1ZJxqA2dVX+7UYgEvCEupLLl2LksdE6t+9tH6pB
cDBe1cL5dkMfkKb9LhgH2oYVdeRDMG5CmyH236waURxsw4IsoJrE8PXp98ZE0k0y
/WM350744MjYQnzZaeab4xSIzfbRDyVN0D5cc+1xPfYkZ5G7+FMx2O36Fc+ZR2Nm
eW7FMTPSBAgG3lEvwYD8Q21VI6ZiZaLtQwu4BBpxsavPkrGvXo1tcFO4oiwxnuX0
YTZtTXcwe4HhXBAX2rUaf4X6LccQ1KTih55PpTbRdd1LuDy3tXAsT4NAndduknk+
qeiZF51MyrM/Rx5XOyaH/Q==
`protect END_PROTECTED
