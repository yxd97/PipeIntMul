`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yEK08JkyK7dNWLvWPEWMGVH09zRdv2YBp7MmjRcK2xm4/vDuQV18pNKwrt0vkab4
+elXcR1HR4eSBfss8TWBf1/BOdiiDTqsQ0HA5O6aAt1oe+6nrfPPjsLxB8IsKzDF
N8aEcIv+QBbAbbxVYzRi8KPRvU6KzbCkISxYhTFaIyb8BenhJBxRYcONMbEWJEoS
JUlByPX6aB+dNqck30QMk6+gUbnHamZgNdN3dEqZk/hw4zBBU5CBR7MZGm3s8KCB
DcU8cJkNQKuqY41HpCRQIGndNx49o7ZyOvxItYS/zuUmFA5f2ypQ56RnorYB4vHi
6Qy1Tz3MODJ4CPApb5+oPJ2RGhxI2SlE+9ppiaHhJVGed4nIdLxokSbMNUBoIzSN
IuJzAPw3Bdf/wsuEEwK9caNTYVPODX1O0ShCzmbUnSbm8l7fHkl4oRGI6wVnbHZA
E5bwJpkMKcaa37eFHZxryijoLe3YvTHX418QPc+GLKuXcUuK+5Nu1vau9FDmlOdH
UmKpj/3y/QBIkttFjt3KYWSYQC0l77fb3XZ7Ug5qtjCPNkiW3OWTLAxoVQ/RHmZM
G1XfI4fnCkvqa1ZEeL9JGcXbSLm8n6KGuEQ8YbbTD4OUt2Ww/Ga67+suR2cG8HXJ
9zOzRqNsc7q0osMJCNOSqnWxk/4a41JD30YybdqFQ2b0VUcRS+Ag8QLV+yL2xwqt
qME9Feif5EdWzntjHKPyF2sNKesIdvlAxF4/JOIKzEGOCIv5AJ2gRyH9U2PslRA8
x7shbKcZXzRjsJ6FIBvWfT79K4svrCq6Po5v2jpLDfaJdGFWRJoGrbmiMWx74Ade
nuWrN9ZkJZqOT36MSzUWZLwN0mSNWY3hdLWzxiGUGl69Ld8h+dXqu8XHPN7CdqC0
vnNBzMYIOsJEWyJiyh2XIL46CCw+nXGCtdX9TY68WHumomxkbKKAIXcu4xLhdEfi
n3ssvH/ezAp5+IMjrtKza2/Kn4RoJMmP0hE2wkgkEj+EgCNqwfUoX0IhiABJsMOS
ELABK55xcygWzlh07d0dgw1vlxARX2mZhfmTYO3PKDy7n7GFTukqS4Hq8zN2Lh5z
tUWHXaXKV4rDPyOTiQeb7TKUjegTZAcf0Fnr2XeOkC/1ZdvDmeyo1VH0TDtWZJ7E
jzgcd4TXy3FpUGThgdazlcPxqUlwLxIBUJxNPdKmEXtMGk7NKm3tg3oWgkqG0vgE
hWLOAKI1YR7Jq4OfhxPpsbI7IzR2ShixGh1ZPPqzQmHlwB+F2tk+BdVFYG+XH+96
DrCDdGDqPEAY64qdfOtUwUALNk0/63X3TdnbKt755rztVZRAWDgGkSsNNw6LLYqz
NYPgm8pRMjGdvTXAYNs8hDCfWnGQ4HBZImoX7jjQBbM7Urxs0EwlKdqqD//egGmU
DiGbSwfiQ34jQybwGvLN06cPOG0LFg8bb5EaF9zun/o=
`protect END_PROTECTED
