`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cRiR0QZFI9qtDpgupzdeuIOk7TFMjGuiTzhFV0xuaBgZg0Ecu+nAr9LfSgFc6IaX
upLR1fdy63XICT7JfQjPYKceUsT4lq6zZJc75hdZEVkOd/Kki7cLdXOXeiZ/Gdc4
a3U/Urgq4q+3X1FghMWyEuuhX5+uCCYcHhvo2DiK70KIL5e5dvt8w2Ataeqn1Aad
J80JPV6xRew4vCvc5LxaHusyzY4gIiEoOVxzVirgeH1ViY9DEbqrZJN1rzWaIYU6
4ORu1OreSP284VsU3wcEYCmXeT+TuMHry02qja7PBZn22O0y0ozBodUMfFGHf4xF
Usw7fbQiDtV5UL3e2OKYVHPMV7uNPKjD1+0LEBcnh1them3dwBZcH7GxfLQDQZz/
`protect END_PROTECTED
