`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fn/D0p6uGj5Omr2T9MUXyfoO/rP2amMd0ZhjxExNoyVuJenIeWfC8ZvYrj1w22cG
v02JYzDsMjj7HWP9/8ZbYiNSHTCNZi4XqvZP59SgIG9SphpKnSY81et6tFeTndNn
vYCTDn7TlPVYSA63SFzspIeMLac2C6JQp/CWkBPa7GQQfWLvmVDe/UR6Xc95Nhm9
T04vtfjHKKUVBCwtOT0LunwzOcdVPOAd3QjfT6K9nXMswsDWnQHPiI08ESM4V4qD
VrSiZpP7oKHIkdcXtuew3XKtNJDGgWfxh/+XNmzOJ6a0DUXrgl8ySDOIarlKv1Tz
x/6n/N9LCo/oTCfrzjc8v7Lr8I8VsBU/pFbEPqPBSmctSpLHwG+Bkiev0711gJpV
fz0l5TntkrbmzDKcOOkLucYySLws3l87zbL7jRu/MYBUpBay5IOGxoc7xRHAvi8D
XcapBtp4WyteTfRqXvWjMChGnqPCvsxjYzGeAkcDsB3pV42RJk8cRqv/QwVfZCiD
s1Z3+5svq9yo4J58Vt0A6s7RGiiGSUqHuUSC2RCf50gc+kpzwuUYNmbPRj1/PdK4
8MPv1ypidLMGrgFYsGnVYW2EgOsC5EllBJZBcXoFtwJRRUnMrGgV6IK7C3oHU6F+
gn2/eIS3Un00eM91kkJFGxV000P8inBkittcVHsdMoX1UrkUau0py4hVNp7U/Heq
lcoGU63lqLfdzbYeyObJP+bSZ1q0MQiYy4pT4Sv6C6j7ao2bsmCB2+A1R0w7/9BO
shFETeGaxCz2fmT/zAD6XA==
`protect END_PROTECTED
