`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uzZfwtY3Jia9SwkwCDnnegz8n9KjYYQVSKF/LFAjthSs4so5oOXaG9m//M0jNxJs
2zusVOsKQZMFY7hfjIgaHIu5U1CN0Vu79bU/Gp+fJ8YeBGc6psejYDnf2Mveovg2
bpaRLdu4E+ygl6urYN4ByIRqo1Jx5Dm84JhfcWsddeJjFApebnEoKzqAFt3bRY6l
g/CsSdu2mKKpxZ30pLfv+4ES+5nbZYJ8sE8ZTK4vqHdd2dLt3QuA9BbIaXkVQltM
M1x5OU8pN483BgarCI7y2mPqGcwipQ33RxjQsDaALuDtSv/4bKbdw9hPzwquD17Q
cj5Ql3HQGro4kQR3q+XCk4L2VpFO1M0NLFYO94DWvstP/Kvx0zd8gk8HdFLhTEby
BL8Jvdte4MBs+iAvH37/tnIdqVdAZ3JSiFC8HzNsnwoVU1D37DfxeBb5lnpssl7l
XQ2IuxZQlGV+P1Pgo1jfis0sWgqE70EXaBcyYl//y18hbH1279oaWXvxKxwxDND8
2X6eEd11qEygMDTIktLz3R+N5/Z1P2Pr7+Cpw3k+ATeSTRIoZGaHiHP1pgL9spk0
hXg6iIUGZT+vrswcf6l2tTerQxuBhs8fkMgt8GLP4kEG7ddAw04/3G6V1+3GfH+I
Vc8WypD01O/P0x1C/oJxnT1R1tXg5zQVNPFiDeGFL3xI3UMqzl8Yn/Rjl8Xh/vHW
8cyRj4x+6TcUm3v8al5PMxkz+9+rju4cII5N+Gm1SlBRRKWjpAX3VvNcsbc19brn
/1U7Ovx140waB2NBFjzGpe5j2Ocpk0yb70sv9wa/4BcFQSQ3y8Zo4IHZWc3NcziA
WGb6xnJiO0dIUDHUJ5h8UIO+YhwSFry0j+DEeL+7lG3h7o26r2Lvzf99JS8DbmBn
m6I+Dp9lTO1qmA1GYFd8uhygEKaNoopWWjh8TRHUSrga/A0YjMnUBsDutuoeOxk9
BTUQzpnMxAzAlGpmGHgobrzmaP58F4Ifw+DJ8DXXE509IDktnPtucVoX9xwmkJv4
1eWPqP/lpjcMGexcKbvj9sOrIkdGDnpjeNVqOOMZOltJ5MnWvxJc6b8mGtCX0A7I
iQSeDne23gYLO76iPWgUgwfziixmNJqVtAHzgZDzpJT4otHmKh/NrhMEN6TMxZo6
Q5fj2hWNHaxEH/p5cGP0sxYZbPZuHkvgVrxRqYjUYETPXQbAAOdD4FapNvC3rCpZ
J7wSwOLppPIvG98w9MOicFKx/S4oD+OAyfENaD6/qfQGJBpy4qSfxsicIzZ5kxvS
xjyi1Q+d30YHLtwc+gaEF59qi3h7h8WHgF7ivKgK8uk+QntSsFs//RGjzuM69Qju
u/TG09PMRotKolTqwqb8CYNXrHusCDbqGjPfXr/MA5kAaupW7BIhyvdHaj3XJDsT
lCr6RBrUIbYjzZUp3vrMwsOoli3l5G5CEmBPrq4ryWEc06Ey1tPXDt0rHn7Ibvow
2mqxlsQH5duKpZArAHC2ev1VgGwwYz20zPrmgdxHmPMFiE/Kj4wUUKJlVHXLWSif
oNu3Aj5ydfEOdITQsJg9ic5YuNM+FWHAR58FyGLBuveMvZZD3twO9H2jX/iuKBMi
ZzUMsKRUmqkY4N6bnItlxalx8XbilmRIe2xyv30LKtCqBnPqMQlpATCA0g30CY3f
6F1dszQFnvvNThcxm7Pt1ls+FYh3bN23lz7vQhK+52zI65IQG6bW4un8HZ9uvRgh
2zwMxB5nFcr9hZW1cErifGpmgg3XGjdCFHGC9kyaERQSBhmi1Q178UMlxcnzSKiD
Ep8lcSJKlcsjIQgB5h9Y5pyr+Gx6LvbEoCGNjrWCw1z1k75K/pvkk+JTcMtApGze
sPE1EARz7/AdM4qxFykn1A4N8mNSqfZ3DgISmVVhgVRUu22lN53YDji9HHOEMsfD
ezoLLekemjGDreYLxmFKCFh6d15oeVMefC8fT7Xov+aiIwylxim9XZ6tE9Y9aXIS
TBjkaCfk4XEj0UMcpEhuxmYeM5+vbOVqwk82CUns8xT69MEIPP98OpkYk0RXqAWX
jE2mHSYNOnRrDN75D+qzSIMenv+KQxZRhWpVAvsDHoSAKqokyO5tggsZwHO5Q0k8
FLZz0j3+6z9WG6mJZFQqQ1oFIHSf/PdeDqYeUr4QDeFzj7Aw+5J+FfK7rNwWLQPl
LBWxm6q24/8GGoj1QA+co1a/ix6mtTqXgPVLoMnkq2Hp7iDaXj3WCunqr4rsP30w
LmF2TaS8n29+kavHCsfgSIQpJo/bpLdxDxQdVFteHARtWNgBt5KxXq8qasv1XITT
7PRq7qQi6PnwK/Q1sHZP8EbF2o4GsaFBd72NPcd1tSl+dlLagWJgsNBP7/8bGucd
jLcZwFxI8oGKBveVEeo0pJKmx3OCG8KYgz3NxxSEkjKKYwIf7CGHjQs+pwGycZK1
izcoYsTNN/OoyQgG+DGJJA0IV/oki6PwmN772n6Hp0wVJc6QcqfEhGqypMZ8uXAW
aaRBWjTnPbxMfkdw9aN0oki4xplmUuakvU+lmOH3Xm94R7h2sl1Ldxueg7xBWTey
CHqu2P2xN66c7v8Fkli8xRUQx4vmDaNHa/j31JIBZckpfx4WF3O6iXeU82iPEU9B
jaAez0TxTRQxdySxrz38Us7YzvC+jBEo7oPShWwJE7FJDPi8Nc5c666Jnbwcd00V
hLn6U5qo1TZQJyCO2GyQztsQbjCTYRVqcbBk2+Pay9y3ZAWRMeprNstT6w+8ibXA
xnIdlH5dYqv4wl/lWpeIaguTOZMW2saYjLlQd9ex3wPJ86oQVFtktchRtqSA2dQQ
0AC2am30rGwU46vEqSRuk91pRN6UJKI7ZKNfxladPT4GqNitO4ZQK/eRQujAGDNt
ZFq9P4/em27QGQvlJe/vqz8gQ3hQDFd8QEln617Ah7069dC/AFdrK7uL+PSXVTah
u28A5sMhdqJ05/GEIXH7tAZRzestoWvHX2Smp4xn3mB4zYw0z3pxGhIGNchwTgjS
lncFVbZv4cEVUmHFypzQ0wdGl5DE5nBbg4f5Mn6/sSKeTqP8WLAKlMP9u+gWWe53
qcZF+Apm60Xlu4SEupZ8XikDj1BVe4ji5IbWpt/idojX6QbPNBCBXQot77OaCHUX
nh0b+Rt85MUKxNVd+0y9eExHZwqqnZNnPtodaydxt21Qtd0yxamvMXpDRMsVSmhT
WKT4S17AJGLckB4rsYUexRPOois+jLJzHUzCNWifpG+Px+VipMo0IZCdxl+uze8d
t4OfTgfeT22t5bIdhqp9VeemEAjt0MSS5Ou5nB3FJ2Rh/HC1EHyqnPjQ2y8bjewV
KZ3CW4mp0AxvVocQBhZNeEtn8ljau0MoREe7vICoPVmm1xXuqMn8meQMgMuS2UFl
BwJFwiZS7A88OpYTwXiPJtI1JIqBuo+Uh0Y6NYUBrjl/RfrhwhGgqaJArBqeCcFH
1ZESwt6mQK3a7dgiGSOo8RSsIc3mHF6roQUbsKJ0xTSkBop97eEGpx98jEntdtVI
be9NA7Bdrj+ZnwF3lw5uJcqCn44fJAveirlYnqBpoFIDrc2k+3mEKb9yd9N8MY3+
xW4pATVbpkpQoPFgmJ8vQSVf5kl+dWnA60eUsHOnKn8EmTx5U9GpT55H0tfRu1DD
k1oTIg6Uqj6jE2X0IGGNPYfnoDuoBHWwi+aShoZXDiu2mdJfhZ6XIcCBR+8O62+c
`protect END_PROTECTED
