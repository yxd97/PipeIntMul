`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdpt3OwUim0965ac5TaoidCdqqMXUQ8SKOjNbIjoz/j47AwxCcR4FMWBmM1ll+zl
m/G+v5SIdo6pD8H9oPAmY0RTJm5dbxoTxuRsffP8R6wmlssvNB2lGWcrIeNX4cos
ZXTPC7w/LkFDZtLK73/4kO5kWqT2Rmj1/Cyr9gpfnR7cnpOQs3iyE/DpBywFUWqK
DiHnjv8FnMv8rRuPpzt8M4YF8KWdkxmz4x10WKMNBqzvHVOYXVDaEvrSjhrjU0zb
4TTCP5qbQ2/6JMOfvLpC+MkdgQdFv1vrjYjpTU4hNpnwYeVYjHIChBBNfhgmY3+T
X2uaibZRXAhnw6CatoUTQQhnAjLEZjiDOZh5y3ElJn7BAMXFccfHdT8sZZAdciU7
RrKXmz2WJs7gMjW2oyMHKnQTDdOVGhK8wIylijTJfUr0WHNDJBAkoUpKe53HZw50
hSGyuFcW4aqNQteeANWZuc8QhSn/PC9xMv1lSbViKkx0szXOQ4QwRi41HBMjp613
ndctDULxj4zdqZtODiFYtLERNu20rbSjeMpFtDc1rLyahrGzy/3InYkQX2PXDsXT
+hZ+Y8uFRGYwmPIt1k8XlRUPf3yuSX1wq9yIGlhb9HvZyHCxvGz36DRTNZ91VmUf
d30vpzRv1HaU0TETLE/8QvgZZ8xxzFXySTiuoku4rs6dMTl343n61Lpcss6oIBB1
uVbii3uY7kDpo81snE339cZBmia5zOG+qf6A7QeIsbbW6SLpbQa+uC/XoYlqBv2S
pKnIEz+yaBpQzqwjHLqmKtNaqVBkoKZIDSW54u/JwbJkvUfGGIGLCYvoSpINun43
wsRz4BrftHYfAmwgOHv/RDtLzBw27Obi5HnJxsClf5vsQzGBb4BFgals0FAMmwPA
asgRMzDKPAG1iqUVSri7YO0gHaKvwuoV+HN36NCwX1Au+8jeQS63PYj9JHYVANVz
OqbZLrYBivVOmsobJ2H3vxjULQ9QpAIcdMdDAUkUviBS5gymo5Fcg45makvFZptv
5y9j6RSq3e+1LAM/2jv+pLdoXS8RuceVHHJmS/7SGN42EdT2JcCmq02vgscUrW8S
zMoo0fwFOCwm4tf0sq2ECTOM672RddBhlMhDJGapPj84wCLcLvlh7+YLJMUpGlcK
QYUZVvumnyzjUqarkOBm2chjoWhp2buPYvKvWUZ5TQjZKNR/lFMhnIY55J3TTz2b
/6esO2nl8E/aE0Tni8ojsjCjQ3PMFnZ/xCPNZIjv2jIxaull+0kuUm2R4BIaT2dv
`protect END_PROTECTED
