`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5c6dk6XConHrvvx8J2xq08LIrstAx+WZhh7srjvbGCIMKSQyGAJYf87vLLCc+Yw1
epXDE9uqtEAGCD9akXELBku3yzeJX+AZEs/l7vPtj+uM4ATWkydcHujnw34g784Y
Y2burvzT+3ch0hHhYYVYt2WpGXpHLMqZjDWu3fMOVVhUnl3TbbtYMbqQfQFPXdns
l9B1QGBWrrG17QLBhUR+mpi/qRkbXS9F80rcsvHKz8aCZkJc+B08QNLSu4o0k7sc
FlL1tkl+zCrLl5Mbus+aZp1te5jK8pyLbToAHfKQ6AFIoE3DjF/fpznL1noDkpNR
BXa9HJ2GVRSjCnWrW8umHM3g7upyWkl4LtXWIfSf6xcv9QlVDmocASAXvC7j4Cs2
UQy7Dok72yppBMuOqY5XX9oAcfQM8t5DTqWiu9ikstrOYp/ZsQpB2fy6WmdyLOs8
d88iuepsk4br4txbI57eSOwDC2Yit9p/0uOrvLjBA9Q2qF/05o04aIalbEL3sSiz
envXRtX0CsFEm00q/R+RKK3FnNlc8MY4k1KToxTIYZFs85P29ebI0VG4AJIMuUoN
att3YoANtpfTLysUP25szpQ/BzXKsXFtD8cVlegUpHlMfLSxHN6JGyJIvVi4SQ6b
fzyHglIWaB/XUb5LYYP5KIqIDvRZxEt0aiICU2+wXN4xDjUcIj7eruG1Vbo177by
AaWXY6iwhx/DPtCsNEqOtchpn/I8b9XbRV1EbenRSQAnTaGMqyMhEP/fX2a8/qFU
dP3ltJz48ESRaoHpi8hV80Z9Ia7XGQx7lHodD8wTUvtN9U1YE7mDH4kjpXMr6Zg1
ZerSzcKW9tAcNdAV/F7u1mIzvSU0uD6Ak//AeSr2LWzFEGhFTvFIG08AmgrSc1nL
DOsUoneWFVyA/RB7vner2RcLk7cJUerCPYi360yE9oB7/DMQSlLdd5aKquf3qeQR
4PCnvGuRi+pBNHednI5MlPdWO3wpYU2rXXDiMK7Z5CVocILjVDdtt3CaxqlE+G3C
w2omA72nJ8Ed6MPfMq7I6HlpvCk7dFMX5QY55U1+sKNTpytdk5pTGpOzbyfi03Tx
DtYq4QwdbJdxsKN22QvMQyE3v8naMrsUISBdFI1Pl3PiXE2aDmjBKcW25LEzuO8f
IGpM1Zl1jFkO8R0Ae9NZdtbmscZWsjH59mf5bKru2pzcNjQrweGl601EIr+t+3j7
SQPrnN9Anre0BBdc5em2cnzFPmmA/6UUB4KcYJZslqasOkA6me6VdKSrRdjd/0wL
pIQ2xba/A28b1Uq8M7/aoDRWWTgK9D+XEjt7BxmbzkoWlzdTZvKj4EGUq3exjXnf
k78h6oSRSH6pJyUfO6dx9VEAkWFgK/tO5xOxm3IZrZjH90A+1asFCs4kWcPOIEBs
eW26VmR5cmVzyYCgowr0HeYHKkJQYvl6FB8Mo2ZfDYRlUtf7qt4kuQzDy0KD48iw
vQgiY+VEaVVHqA/xjAhvkILCxnFHbhH+CDC1k8iQWkk6cpeJAKFTyemS4i4dslfw
iYBa3Mb9uxjNjciEzqrq33hmF/Mtvm8MVn5dmXNzD7cJyZxRnf2fLV7iwUN3iDOE
cNUCI5nnr5jMgMi8apwH4jqTyW+ggnG8S7ZhA1vg1g8fu1qixu4asYcH1jNUSFuy
pstCTlGPQxpyGUkm9YwfFlcGs97DRlCim/74ySy0cK9Ktrdm1mcIwuLZWLQ1uWI2
5ZJjnpa+2K4A/sak53vVPtTrZCH3z0syMErp/0N0RvjXnfhyHpD0ZDkWV9hJjwl9
HrPAkmcWwa7CJGRQ3F5ALLmcdzAO2dr6V2+zVgGCQDkANLQtTiLgUZOT1Jnraobz
dQTCh713AvrrY1QRH1Gub/ZlrJsr5OAivB49jFQvq8On1RXXQXPU2z+SLPI4TOLH
tgb+iL4MzFnhe594WnbCzy4FzSh0e0asFXwgSaoRgljzb8ZTkMlI3avuCwxna+nz
IcomPZAS+GS25gNWjgW1FBCFIm9mnz4nro4vESW8eLk=
`protect END_PROTECTED
