`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TpvD0I4NzGHsovhE+9AoXaB0QbMkNM/a9uVtJKtU7qYmHbYo5mSlHyE5fghXBKxE
Ja11WAXiZ+HkhnZ+A/3IdORGrRNJoGG2afmprBEw1RqNXDRWU21ouoI3E4DiLdZW
Zuyeh5h8Tg0hZqIQisOQtUpBPH59mcP+Mok1vFIWw74aVDg3UTKjucw53AgowmV/
Nu9aGgimDpLHTHrAk1dX7wHA4j8gALe+/OMQBWMcsjimm7shwyYiws8FT1U8teS1
xtqpj1+PvgksaZm+38c25BCtk4WBM7brYCQII5Kt63h4VsJ61GeGihvfp5tp7Pfy
vhnjw5y5sQp6h3i4vPTFPGJ72xt9Wy8vF41b4OVj4BiHgNEJexom6tiGC+K5Du1r
rAjEW9mG+2g7ed8loKBKXyGjEhNv4DIYA+DjSebn2L5frrGXmHO9IZKobxqOTmWD
A8+73Io60HDub8KeW7O2+lm3zhbXXwj40i/9uHxFkEfQMg2dJhapPK8t9yzlhgjr
`protect END_PROTECTED
