`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4j0wiClLWJ//8CB0xBP1lWYIRR/dzt58g8G41etFPhHFSiDIpq96zNEmsZjgxmJU
7kc8XeNYCTsPNBVVxnxJqTOTRX392co0kQqgmwnoeCESdCR4EEDvAIAvohYbJCuH
n62GbRL8cl4aC5MdK8nHrXgpKZB/AQAoeh4IsS+Cd+ik0G3NX6pq3GpEP9e+nQzt
eR6AlP/4kSi0MdpLbun39sV7g6nIiVRocqVHzitT3Brx4xGTr8law8Dd2bLQ5VYo
80PJSkha2WLqR4aw+S4DM5e4mor9zgi8T+35hKXQ4eU4TPY16YPiB3U3n0+KsOTE
Oil5oIwmIW9N4jLqq4AEIfeVe0epD1poNhYOtz5MwtdWVf4/pqYDgQOdgChtXnQ3
yprtsbmq1kHfCrrx3vfXmJsxLJmeC6Jf420J+w4SoSWz7P1jEFaydxLywHPnYmUp
XFR8SpjEVrO4jz/bX48gIy3tIkzudjiM3PldXrXfpjAReIGptrCBIdYrp4TsIvFg
CHmp7QW7A9u+axGRLqARc5TaMjEfuS/sYyYiLRpMSRdTCTGlsclvyT6Xk2K5tF7I
8xcMgEY+c/2opQbA7xO6+g==
`protect END_PROTECTED
