`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z3IGENmLyt37n05EKk4AkPd+dzlIIGCbP4V0upiHQZLfGLUaSKP7tupZ6h7afOI7
2k6XK9R3mka5vBLCaI1+eBL25A0zUjbp0zIDDxJwxLabv72cRAYAbfb/xiTfuNci
GmzpJRA9oe+IKMa5VAbDxbSH3uSzkbHFIyBOGnJyFxpDQU7eZCJ2NLswtNEWK1iE
4C6vcq78d0ievdOx1Q1yLKXqoB5TwF2ttgshUMFe77WnWpf3RdrkCvIPelcX32lx
dhn/dbZGsJOIacaPuhXKg1o2GtH/OD0/4HtX8nxksEBC+HuayhRBBFcqeVpwhXGT
9yVLWQCabYY9X5MYhGhhdbjS7outFDP6LQqQMtlxCLq5PK0PyHMFF71KhwirNn2H
tEqTh6dj6ZOWKNsuUfPlc4gmjasc0hqhbS9rSdAYQMJ3nfGJuPdnLDUiEUWmCGeT
cOoBwvDh2AWLDOImPOOhhjf8lViWvREVDKqy+pgBi61Rf77D1sDgxyiJ6OLjqbcV
WEeRumAyYefV/THfXT82ZaY3OMmQ19CrZiVv2QYh7kQRudgGg8VILbYoaRUz3G6/
ZCJta9cUO7NSnEq/8oqer77ZBnhwUq2H31UBstMUv0OvTKF9LsSFDjFraiiDmSrR
mJCpBuIK0yXlyT1PESDTgMsEVNstOC7bB9dKso0MjeCo5SxNSDx34mOHAF3ypA7+
llBdYMbDjDtLxxg/9lMji5E//yVnOg1BZk40lXu64CVr+k6DIMEEtOF1K+GSjGPA
QfOxern1k2X9Bw2Mn5pXu02w8+xPYDeetyA2uFS56VOrL+YPFdzKv899tGFO9P1g
l4iv+m58C2dh7bcLRNjQRBqCh+Q12WzYcwO1bqhbxbPRuIl78CiUqI413ccKLoOu
QdDpeEhzvdjA/Pcj534tizhPEK2ebKFq1WVyuVESPTXalTI8JxBZFxn1EIuJUayb
mffiFopsBlLp342sEyFvfMuayzUsc3wdHnHKyAvFVhZQYULbkZA18sj5alzsBBQH
VYRzCk/whqJGcHcB5QsUE/bWck3w9clk+hH06Mu5UrXg6MppEsrwlXOyEGhako3w
VMGXktkg3WXA3qRpZkgzVM1Duwp0JSfU5bMenPODTILqYiohBPv1RZodj92QaeeQ
pTR1qUmFM3GrfleF22VFxbpwSvNrm0usQQ0U+Ni6kdczYVckS5iPg/9ZygEb+Tiy
ZwveY679qaZqr4Cx8L40OCdJ8p87IiyDVkqvkxQ5uWuILvzFhsRXt8gh7p5LGj5z
SOUBixnR9LDJIDdaCBAGj0YpPDztmemebW7VJKm/yS7WyPykGMrDSQlQGKJGIj+k
p+MHuD9h7nicIbAPABmFw7K1T40+aCt0bSg402nqNzSPkeUYeL8f01SvH8r3QcDj
9JYX4d4vWe18b0SPLOJGGYixp5RojcmR7CLjiJ2sT4kA47KHrauL3VzzUwvKimL/
fIfFUubHtKfmPughiUWLgK6V/mGil1r5Ra/36yprj7zHxoGGicf8V9yPxFs8cx8s
bKyONL5USUyPr9OgUmKpmGRRia39r4nABH3ZrA7oVRJlr2IyK7sDj+oQtluIwHQz
3ukNLQVSp58fjY4QaLpTrE7Q5DKOB8DnonJRKE82DY1gD090foFxh5C7cpBoP7oc
`protect END_PROTECTED
