`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fiA5GJaSt4bfylfUUZjefS+M5SdxovsFx3pyAkhmbtDLsWdSCTaSwrkHK6koYAsr
jQTgK44r31sOWbIwv3Ad+sOC+JpZvx2Dxszkup7WyLjOjmZ0BK+3rtKK4UgBMqHy
/nJeROH+BAotZH8fhZFUhEX3YuMZu6pGz1qDIPQ3ynoQSpIaBNEgs6qGlCHlWrJn
otBc3FAzI13bnPQ/dZWkMsF7BkmKA10/VGcb86ecnqRstx5o6Vo/PRljGuXC75u5
xjZ7XIDxHEB0GscI4Jj3ta8QvYoJqbAttf7F40iPoUdY1ij/YbD6UH3ByFGC10v/
0mMppsvYIKUpnq4Mfg/YWRzW6Mx2CT5WZr7EqX5/FyxlXSd5aKk4nfl17CvHU5/0
bWViddUJ6hkpYiZ/UVeykkU6EcYEFtXo0JM84NegpfzKLx1mQ1yz450O2BQj4JBV
mKVi/0UDaKG1Ku8zWI0kdgnUpo6sUhua+uRwMQIZQyHhqUUfUQ5ptUR0rxxPyQ12
zg/2BML+d0zNvsgZdY+7UJ5sIgNQyEHOwvvyrLC+P1XoZRKeAasH551KvTdtBqgc
mKGagq7w7vi4cpoQppA0t6M9sEAG8UcxjDdnh+PEihjhj6ejH+R2jhpbzFYSFUkh
Ereg5U2sgDh1i+kucBWA68m4jPo1oALm7+6Qz+F1cYMDLpXJDuQwXiyh5znau9jg
r1vtM0VYR07FS1m66PREjGNaRvJm3sCqePXhPrZ9eMZnrNVJUz1tQty+4vAzhNyz
`protect END_PROTECTED
