`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9jjphbne5xHV00tUYyEC0ruOiHaUB91s8Bg0p0cg7p5GjwD+y5xfQKplzV6fXvZh
YQdCoLcYT0KvPpwKc+nK+tysJmunAvEyoaj3vp8EZ6a+V3nsxKA3huoAe2+tGSJ7
wSiMxE8ejhTD03LhC4md7rbLGtmd2yMF2rDBy5oPyhraJtICZOzCXqc6WDGcTIyh
sVKFx1lhvIVD4X4ibPnLZzJH68foMez6GelRm1FT9rgCA+Z2a/9RMz3eBCN+EK1q
Dl+/cFYakIHVC4GzTsLyxthuYwgHFbzDLEmCynx6KrY/EuB5nFDH6oxBSyv6j/c+
F5fLEJcdW2XVitTmfHjp1fyZXKmXDPvkKlq+byk597uQbG3/37kagBNdey2PuUuK
E1JSiv9iEuktibl9+mJfjaFEN3aNZdSZXC+aoQbvmol7dlkM9gL2zISHePZGznPC
yhM3gDyWpqWfKLNMVPyAFifXox9dYimAA5oj/xNobdSWuqSIkpiaZ42kR+g1y3dB
l45yizcjtwgLSaRZnUcD/oqtjoxLSdEENjaCKAXosiLwHMNdNzRZRzfjGfH3j5pV
xBWFTh7FV/UKcNTOZCgYn1PVTHwoaNFxLtFDP0015oVXlLxgFlPFmWbjJvCuz83E
+Ict2X/kNPkOxqonsSeesVDxea+V/wiTmD7dq4/wJpJD2nrpH+PiK9pf3SDsH1xs
3fBSaTCG3Il6gMlVGSxpj37QCX9W8wwcTE/eSLseZkqAYTaEgovTrij91YVwauo9
O8nynln1jFcHHH4tesMTETrdC8zZnZkbXGhXrDZlg4Ysp0WjPRxbl/ch1jGIhmUZ
1KfBCP+wQPVvT5yq+W+RGnymsEl4YjBObyvs0JtN92oPq2sxZ6S3X1vmOWsCjWAW
KFZP3PYXgftk3WUMm05YHKN9F76aH/OVAy7PgcbKCpMmHkTOiXUj4Da2yvfCtZfM
5tmQFimsUACbWUwRfGKKptewIqWFx9B80ETfkheExBUgZn1MsHzNvwdNN0pEzduX
WDCRZSptuL+CVO534x1NwA==
`protect END_PROTECTED
