`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OD6I9mmpDcJYlO/pN8L7dH9CfoHZWaWzNwQA8UE0aVPfdR7l09GCEBegbU2DcBlC
QT6zgedWtLC9EH6/3RaihsGyM9XXtK+77CiEuf0fs/zHOFkXVE4OT2lilQZ3fDr7
Llt342KiEZr/AdOKarrYaTgOQ/8lL+5HqgqxQUUnGI27YfoqVV55Te2kSBhGA6u6
aYt8fCz0N56nZlDQ/SMudX08ZugdD8DceXqy94Q6u8t5uiB4SI0q42Is54eYfW7j
ALxe4b6Dvi2hycWtSTf+Xgv/renybL0aH5rzKAFCRC7Ett2bEX6fkeCgbdGoIWxg
bp5p9Y+VR5As6hv2yA7sgchfXFQWBo9CZERDiT85YcGK3BFboCnjWkmOklXHh0ip
GHhFXcN4sHXDuSFhqdvdFzWh8qF/oU0yjCwWZt6FqQg5WxA2M+kUQZ/nlt90Di14
ipuT7CtSh+fQnQ4d0xw9HinOJnJB4/jCXzUvmDM0ST/hNorh2pDEk3Dd8/zAV+7I
REqRHkEWipimw4IIcbSfOZ85nvRq1ooehqLPKAp9gJPLzbIr7nSnfWZ5o53Nbyra
r5OSDbQKBzdVRU0ha8GjSjZKVd3Ffn4F6FZ+mESjICC5018CN0+iMPCTY2LZs30h
+i9dIU58wWAE80TnG/eQY6BQk3rb1SJN3yq74Xa3rb8c7JhstKsDlQFBOEOHbsLa
2lYL655E+RqNXHi0ImRayQjbjpyJhDF7x5oYJRmEUB4SL3c0gZSRi8YPKMAMN67K
JUol14j+x46DEwRAjFIQfDfxPtKy6V6l92wogV+Vfc+9lz9yOKa0cJwW0dZCdUxp
6hpbArJHy/F9fcijaC12NoYdVw3YbzT5/w1uttgNyn+dBAY4sPhQHESVlfbRUuz3
2NP5bOCeafMSgXR7kbSvSo5jOmG31W7lyEZUZPAHy4t3+7K0pJpHOblcZf/1BPb3
ZqvAJ7i8Mb77rX3n4Uh5uh2K+BWb3dcZicNuNDJAF1htigvUxJMmM9YIeVDLb1+m
qAhz42qyC5hpDoBI9g90/JGMLPKYzejyGABbTMa+F/kyCMcH529rp+iW3ReO4b2E
k8oo0DIyC1cMUSxwy5uubIg1eDRos+pursDXP3tf+1/oIO9uKZTwXRfErO484NaO
he0GiVxRbv4W4HpYz5hekZUmxn0EAP3CgKBM9WOJQjHml7tE9iODjgMkvaK0lbzn
NsXvJk3MDCKVf+jHNqs+vALuPzxOOLUIDddZjwlaKrT0YDYFtEGhYPHvoNjJEQUH
F8w9Vpin40f7uDQlDieuqrMDeYOkJ1vbs+DjC84q9JUO4S+GogzqCHB/JJ02UcFH
eOCYzaERAY6NJAt/xJVYQ04TkkiZjju4JNptvB/C/293zE1NeDXZZd/3gyix2L2S
z5YHl+KGQP7aIl/ao8OC5w==
`protect END_PROTECTED
