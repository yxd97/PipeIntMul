`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdE0l88sHoBFQgM7jiSMhhSZlDPzgA5YtEVwoLlnw9zXACQYnJGODfcoE3LIRxWj
EluL4TEuoDJVo9Mk6TmLOnVAnUeBkq/0P//zUxcSaVg3s886a/FXitWi/dK9H3NA
kyg5M7uv9R1JJYOTFWodQB2ZslWA+IxLZBP07GEGG9p5rhlG9ED/goid3FOxUvhx
cnGI5JG6kjicjL5Lva9CoTFPOQ61XW2pX2wNO1VOl3V4TldeDCol2ebi7QV5BvIG
yA5aLTeL2FZnUGm1mDsCtOZMLstDVVYUlst4MeHQxPgR8ae7b3HbqSFnQCEoTb3D
zAhmm5Sc3+zXifu7t1jit0BRIsvzOn418QBrGdH1ru1qXotFcE2yM22bKb1ZDUpQ
`protect END_PROTECTED
