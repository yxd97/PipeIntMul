`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ygusQoW8sbdCeK87nSp9rK9keo4HSLzfXQDBP1xSpdRbh1SF3QBExMAAHvCiHeGc
OoTJ2KWf5umvVUZm9j6WjNuXTNUWv4KFVj3PGzTxNnbMrC5AspeYs9sz4xwwimjI
Bxmp6uiCmq8TbY/BkFXCTtpP6jL9GowYJ0ETsuIl5Y/xll3eyXl/wm3d/Dlkq0BC
YtQ905C1HCqP4d7JczOZrA54DkXTF2QEftv2vMdJAdVezxfcrk8MXKz8TWSarGd0
EUPEhZAFuk4ecY4Mx4zPKRSZQJ8II5eRZ99c69608nd1lrd+phWL8+RMRMeabv/e
1y220S0/HNtCEXbIFxxE1HHuXBHNDvBnuo0nfTnnXUiTL7th2OTVxnBjgGDb58YK
p73zbJdRTx12/dlBCUkdxGiBKzNRT3j60kEB4KL9i1LkO5mnB5w1dMXD8UUksNcE
UasX+Ef00wvWlEOQ8aUilxS+6KBKJXI//4DW0jKjvdqsowiy2N/O5tEjd3bRfTbC
UXHKD6xxRRGJcWe3iHANIgdnQF1jkxO0c61rNqPS7+B+hK4/CLVReJlFqosz0QVO
sQJbrbXquCk7PKt28hYZiAxTM47+lGSu3iHRfe/rSnhHS/ILrdwYXvlRUFM2br8+
LT5ZM0YKTXet9JUKh2CAXg2fDWPO+VL6POE9thhTpWM6q2KV7nJnY9OBOnbrQgAJ
ymTbjQTtxJYZuWTRiPdR49bnpnXDniCdQMJyTMfxd40sJkTKgYSk0EgO8Qj8OEsn
HX9V2ZLGqu+yXR9O1Lg8lnIV8VRIcX3+CRX3A3EoL3c=
`protect END_PROTECTED
