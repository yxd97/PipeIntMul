`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q04ty6iaOnMcqcBFIs7GHjUa21XloqEYocoyYcYAGipfQHDPP61ZUhwM7qEYh3/T
2XpycEUEHxS7WCdxjAWt9O9OoawgIAuUA9nFPzMP8/9lxYb8kV6lmvFHoeSlSf6s
/1ieU1WbPtEO2UgQAWZqGyEdKsnVsy7RZErOPz3Bf8QfmpY5Ld6roFKCwMRvRd7I
CV7IZtdjr+S0FhlBMNHbtus4GkOrRA5xpfEnBlQgF/JcgJf1OcdQF3QWhJiFwF2c
AqeIAU+dujSnUFQwe4O3RlyjT1Id5CiIiIwWJQZkgtX3xRB7AOwKBE10l4f4yozz
4jiVaNmPYH7rIDLEX8ZyXvM9FCEEKQ1x8RFw49o11oTcM8MftoDl9D625ADw/0pz
3jZuMgPDp9tN9W4ndsePdk7yLLSmr0TJvFsetAbIKN9hpG+gkyRA4646ioAhwf4Z
5qE0Mb/hoeV2eYxbgHWp7zUEjSN1Q0L1vhQ+T051xrHik4xdlSAapp7ZjAG4utjP
AA6LxD0eMSJMiIhGkH+rltiwk2Fqc/h35LIu9YRI6Q735WRKeNGIsP4JDXD0gl3r
EY4KWiCJFR8A1kJRU7ILcRjiqly2SMCOws7XxuDBMI3mRkyub9MbQNtmFpY+Cm6T
lIAz8FcrUs9wLfnJt9fbWF/wSwks/Cq9cpeQ+D3seLN/Fz60lKPuG/Ljq2oz9iZJ
9ohyNn1JJYe87hespJUkA5HHQrGZP8FPsId7LzBp6C68axHtGqlpmx0FbBXbUR0s
VjOv922nti6KBv9GDeBlNeQucV7zASXj6SJRcME0jQYzgrB7nw05t0eYMhfLCZoF
tLmeVSHy/iGyITDn5oO6XWZkIQv+JKnNyE/OYd/NuOwJfKGy+Q88WdNkzpGRayG4
L+fgFBYPuaYvunGwQ/A8hcmMy98EWmcOfOeHI6eS7PSpoJuHwwO+/OoyGq/E2zbs
qxESgKAQeWsGy8tMzLgaGIqxOf1x4GGyZjtKohVZlgg=
`protect END_PROTECTED
