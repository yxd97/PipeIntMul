`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qfbArxRody0KXeBifPpW6lK2Z4GYg76O7mJ3Xxaj4gtR/5NeLSCXdry4OiklwIh/
XuH40WWI4NVVhoHG55tXt46iDT8wgyoP6EPEF0xx5/paZmjmCN8WUDgSO06wsaZo
H2tLQBA7ZSvhZNlpafnyhGyA1IcQqxMPt7WGGhWBZTB6W5AT/CkEjRYoihHDrQI8
PfARQZWFrgM2fI4pS0XhPliyhJeLeDEFD8fDgBY2FlBMh03CCJfkYKDyQYd5W3SU
/7HPpaNX6oXV8ouq9jAHrsO2BGm79V/lB2pG0HHda3ZeTSP/xr66dgLNgsvU9BeL
783QYs9wwQe2PLAHdixRBmyfnT9pK5ag1rYlUHqHZknriY9FBPnmJDnZVPZAhaaA
ynKz4c54oIQb1Rf6jucPCQ==
`protect END_PROTECTED
