`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
igT6pRY/w9hqNEKFzxOLXgi8YHasWot0CV6zZRfpyz5NHui9mntCBYV0sdLq+13D
gVLzm2ZzAR0CXT03U62ZmGvzsiSBBgTAN7BucdbwWYFjSTwb9POEZ5blXiXiEAfA
PGH32ggs9SkiPe9VqImhE7eee1FN2SMecOWyHP2uZCUlzvB7CkmRxwtI8PgZWPDB
SgkzpXbjz9YWmNLQuU3nzxTC07Vvu+1Zq5iIT/TUvDMK4r276ENbIlCtU2LeY9om
UAiPg3+x2UHcqH+qHb/FAYnEw2fER/cNxr+k6N7J7PPYJ+OEXfe5zmrUCF16eOKh
4JDuKHt4trfJ85dVzin2IYjGW2r/EviAHiOxdDawqKEarzH1dzBlKWHTkQP9kzZt
yaDfimLPwCJu21vQ+aiidu4B8B77B5Hwd7cmEFvrR903DxNljaqtimYUtW58ql/X
oaTzkZZKTcwTRNVfb50nmsJdmMPO7tjZk6uz1vK59DbFFKZ/MJHkw8eBdA1Tc1AL
Pji4Fw9Ec8YthWjyRhqzGV2kjz77cEMQvTWJIa6rKBA0oVv1G43G3BrScalUchqG
TDtRWg2jXdvCh2as9sWqLgJAy+8HYkQWI8hoi7lnOd0tgcbsYm15jZy2gPBYKQcD
H2+QYuPVD5VFko7Vfc4Uy5xtURL5WrwbgIxkuStHC59fmuozNoq2kwDPLKuSvaw1
kqIewndHbbTKb2EA38cikYVUBza3AvOO0VBnoFhBrShyk3kNB5ASXenluMOfKfIt
nDhDS+1KCI7PRu6Kkv2LEW6rwNhjOrxE7hvAEaiMpVKvaAtv58NmSFOSf9IxO6jw
mwx80UNt3K0LgAJXD31vYg==
`protect END_PROTECTED
