`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYxDolnvGv5rAAB92rBX9ghoAiYnFGbdXdNaZnC681CQTnYmrYu8CgM6PECOpis0
OgL+1754dXHphzoDX6Ibx/KmOvFk+Ct+nisk6zQdoCNIMgchN+7LLYCqSY2W/V9P
G0YVQjjE0/cYZ1uFyCpmVPxqZtfwwmjr6esDBKmbX6V6EUt3FXglbKYQDEuQnPgR
HabYg3riVKuGMpqwTj8yH17V/R2Q6R2Yn8dpiYfLv7ha2rb7tc0zpDV2xg7xNRQP
mzkw8m91mU+lqimX7CZe165o926lhLwYSCDvP4+OAzwktbajQ2Ngz3iQ+mEjiPA0
t2P+g1uJDgr7PO5rvr4ENCxCa4Imx+0Y+23mlpWeWGx0xJxtqbHFAykKBXbNoB4J
M5hCAu8V8sMaJiTLrKR+vg1wVPyWjg7YjW7wCl8KEtC0yjbGcLq4sPjq7U/nkob1
9uNAUKEUFWRE9OzPaBgBmTjryGO56A7sqgflnOhpyP9jtZT8Du6HgfE0Ru0qTrS2
KhuXLpsPP4Gvu5EpbE6yKw6HV59iiYpw6ohKJ5IuyYM=
`protect END_PROTECTED
