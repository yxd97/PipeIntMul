`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DeMCsY45OjyPmL3xVedXVc/qRSvJOP+Xsv9RvfVWDOshJmPfUeFdApr+g5gslkRD
6+k8PTXWr5hg5crdhwN+apGM8sdE7mLCRv4uZqrSFwmacPnk3sGa8ctfryOm5Deu
ifVwqb5ZDiSEgvx4PrfRzS1S08Q0/G/O2Ls58tIWplW3JN8QG7X9FFdHUZrOT3PK
ssY2LkqFc7S28P0BQueElU3a+estoxtDuHN52REKgn7xcNqlVOy1wVExkvkRiax6
AtECtzXck9bs1zcRuXZngwAOU/MksLQ8Fpk6879wm2Q=
`protect END_PROTECTED
