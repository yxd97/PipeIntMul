`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VvGIC0QNtcbaeeCYc6yJUaHNLInXNh8Tw/e+zi4ZIjRyoPhS4/cxG+aslAgFafw
kC8SQuBW53LShtt/5p8baSGpKEVdQQW23aWxHvbJmohEMMtY5XFqj8D2VMs5gNe0
9+KZrGhHmtDypRAk8VfomVjzpk/yaBQakS5ncV5rO8MvIXAo3bkEu65EVABhJq5R
b/4MEr0nfaU9Y/hx906TqvaDVjAt36q6a0z+gqQgSH9dgmV1OKD6lFp3zfdDCi5O
zif6xOViBfeT6lMRv2X6Y2k6TVQGFX/Ls0vBdau+A6DodeOLMdzjTKyiIysr+ZCi
TaewNgGSqNXTvyNNyw9GtVsMBJ2Xq7ydA3kwuTwWJoJGqKuZru6B6V6b8gc+16+s
9mPehClo5zAuCd83pz234hnYA0B99RsNcjMq5AofD3OgAXPXXfey1EHwkCJLSHDe
BD8mg9eVVIsCSKCnBP27oA==
`protect END_PROTECTED
