`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/UrDOsIaXl4aZyBbCZESkJZ9csfvUpmznHDgl29xicPwvnbxvFcz8smFgOFFYTz
0YDNYP+5CatpeP4ggRx8Vw7aL4EQa/FxBmwMBs2aUBH60/w9zayLVePtRoPiZQt6
cTydVvDtoN5U+PPr8/YVaA6jKi0eXNoxFFWt2cZCQAjFlPyYpr0hSYoI0z6oJb2e
5C/qAAO51/erKpMVaPIupY33X6Qb2QIZ3Q9+wwqm/Qm+d96B3a7PwLe2ttrXzMkT
LsPiIcNYKaTWvkC8bfKPG3KyJMN7d3tsa1GD50uAqSVyoaVnBhNkZrKZEiMB4BnX
ZCJp+83CeqiKHCUkDXLhEOQZO+7S5nr1JJS+3A3tx3s=
`protect END_PROTECTED
