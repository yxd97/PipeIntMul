`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6cS8wj4/YDazV7bLE85iAC0gR98oEi/3fIiQWk6ydC6JN1LHfZvcXqrMHHNICZj
TphyCdhvB9BjniQIi/fjkOZqMjJWjvYX7GoU7IUrVuLnywCYeI2k3Wu7wJVSRwCL
PSiHbDkDhVZ0ikoMc6IBeVF4guL+FGHnaD9I6svrxK6BVQQx6S+kwDnhkMu97Hkt
Dsz+XsYzmOL9v8vFT4KL77oP5MLiAeRHfzazsJUzkLh+U5FZ7MjAvdXBPInxq5GS
i5OnRLuWezi0973y/kzAlsbK82nEUaOTYaPHI5DHCtwnzNltFmBMhYslubXDZpVP
kb9o5NX1TGVZDRzbEajKxBNHt7MHnQHIU6qvLLRSDGPtB3CcVpNvOFjyhT3k51D4
0XPgxWT0xQwyBarws8gsQtf4Eu+41lfqGy1q3NUtl+4MCbjHEE+SDI8DDDUtehhu
O41fHkXomF3rchs2MNyt+3NPQtT5Yw+smcMD5rJ1FuYVfPUkA6wmWkS9NVdyTwR1
JOAlkri/6ICsqeLHvG1N11my2bFW3EvcliEyify16ae9BOa/Dx7tLXAnhlaJZOPG
qmOU+/gQydy8u8e//qi1lYNqzTgeZWxGPl2FJfMfCrZzVXZMJ5A+bMS8917+fWW0
MLXye+ttZRAyA+pz9/33mJfvhae9XZgoMzKzJzcUQe5DndGsmUH4xNf4DUL2Y35t
ozTL79l1oHcpeYnCta1dPYvjWut0KpikME7NRvWTM79rVj3vaYLVqEBCabc4TRSl
h99GbYt/S1jgCyQ1tdDNCWee2bZvXcjdoJia3aJd3orWqf+WE+rnd81ID7DjOLyj
38ajphSkx3RSNwRrO00GMIRLiZKIAyGWP18kDVsS2YwrpiXvB3KSlhMFpo+PS8gw
t8++zwzfPLCOMEgrHg8E3YaNktLvDtBSH3D6BIBLNqJDK45oLDa/7ZbJSZuCqQ3x
XH0CUWlblJ9fxaCopaa4lWlKK7LuppjixoWOntN7hFtQ4HtU+yr0ENrmwHQD7+LH
ixjUwv5f7noQXIYQbf28Id1T2jtUAhHnMgCuo+VUoBG3xUGvmhK8XyO7maW23jR8
VQQC/gFxlZ5CxWh28M+4+9lU08IL+dRzB8ZlcU8BTWFKVX6SLLQv7D6c0OllXoPp
PnzKhtdcm9IQN/if93A6gc0M36u9Sbf0276IbC+B/UOFKlN3R3liTFKf85dcBQc9
OsCUFrrWYLI4kqawpL61NyDU/i6RRNnfYAui+I/hYKyVkaUjeE2z/tKg92d6PwuW
rfN0xX31NJMcl82AeRWoYHYTHro9CCzHIyyfwtTHpg1makaOJntS9QhCcMUxljXp
8JFDw2xUJkIbYq8+h9vQ73vBOPcCL+1NDojBivgEPz0SJtkfgM4sj9uV6y0m8ETR
PUZhatAvivRgCrRhVXFsQH34vrfMQEHoAQIwO/Py6rIpxI4zu/HLDcK3fuVv1Ky0
srW2wudKLjlra7XgvmPHu6gYA1j2uwZezDHS/E0hMsTutgGlg43tG3lfFsGVmG3/
sHBCgUgCYP3BaMvgMl3xubzeDcQEUbHZ4PujKLYk9KIRXKjfgPragri3dbcAyS4I
S/kYfYs2zLmw3oDPRmCYy1SHzk02ZrcR8YAi3jITynlrltKpvs56y1K/l3bwwI1J
rFOMT9Pe5E+LGoUXp8ELSp22B9ETx6DwKZ7no9jAj6dBbXqP4LtVZxE4DKEASkn0
aQ3K/RdrDD+4ex8SXJyO4pgo6k8re4f8cxf6MT0XQ9kiT2WKR+fGTjgfwthm7Hhx
W0L4+02DO96Fs7xtp+C9rA+a59/lESoZIssSXazL/NV1M7kUSmWRBzkT1aQnBM1N
FjfbHR1LFjeIue4O9U6e8x1iQ2OQ1HKn4XNbWICauD7eBb1RsVOWQ0UQg6ffs8jv
COfIdAHN2E0D1d+IHy36SqORT+bIYkX1fk3cTq2iUlpnUKKx1nX6b/6cf4bFRSwf
t3PGV5fgSwswFDtLEdRn+/DpEdutGAiMga4PPgCJG6O0nQ3HW/eiNKZb6Z6fEdKB
`protect END_PROTECTED
