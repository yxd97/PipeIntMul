`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzNThZxsGPCQvSxQJj+d78DzvxoYSoduM1tLWUuenIokPUVC1t4Jy6DYFksCZfyA
dj50GEl83PbfU3ff8rh+tyWHiPxozMBZYqOm/g7DbPyAViOmiNfRMAqxFf6l0UzE
gdSsavJBjUSAXvW5LC5QXKv61tBt1ieehF6D1kRn/+p2obDpev29xckllm7puPXO
S/fPYPNmHp/q09UTLoZ1Is3ixPZA9nkd94JaFRluDNGDVjOfXG9dhChDsRn9SHpd
TkRUe+sVqw3u9LxLQWvFGnNpqjCzfrYG3L1KBuWdMBMZJnCFIWTaWyTOerbP2C1y
kkiTNR0XJ6fouF8deyb0jxHPpSH8TDWilp5hiCfu/cIgRNjzheLhHiwibFwA/7lb
+tPta4xJUJ5888+CBzCq7BUWJJaGv+/mm3cDZyUGtMpJpDpi6G5VCFNL/M32FuIb
1Ivj3qXxcMYEm2sWOrsxqDe+6FmsAB1rwXfgaW1OUu97DJof9+bjKe5Cdh+Mhw2x
J0gUlfeYTArS4BSijgFpd9sBFu0Qq+SgKQx4Gl9h+YYnZp+RM1RFfLPfk3uMEn2R
ZolKf12kArZpjYspOdUIDY/CORJHojyWPH77GfgYYMeXcFZaxhanu3fPzC7Ue1Ka
5a7gvwSUphdocQAcJUxriq9ByeVpn/9LEXINy4A3rWM+/ytvQqMr1te+iIqWBET9
+IiSAi2415kraYw4xkZVNFQi0Q2wFbSwRQcly9KSkj3RHhCXoivMEi3+Oj8NJ6s/
BUkJW6SaPTn13d6QK7TDG9NggYSg7JQyfChlWG77CABX9m1Oa3pG+C7MFm731I84
KtFMlcoMiv49Dwk2pygdY2WMmoG0gjctkfUJp213JTHRgzQevTQKqdmS/Y+ap3+S
I5VWDAeJrQiXsrgOHA8uI4Kjll3xX75Qz9OgEXXNRYd1g4X/drCW8Xm7TWCF0ytB
MhcOJdge+Cj3QWEF+t9rW235bB2kbeZKn6VsAvc0dA8h8bUAN1X6kJvnJfj655Pn
MT7v2FibmZJId2G3BvO/+UKmragUeS+WTes21E5wmf9bxS+5NlaCn1ANeJz2QKx+
NjHBi2MF6qjL4wZZGIWi31elOcGzzFyDJssME4eG2e9itYg01fyk3Vqd8Gv7z1kD
acOM/a/NcAt8yQnJ6pvLq61p/rTIMy6Ns0omojC+Gnfli7e2ktYvGInvM25uXRyK
LtW2qAjfsy5BIeP2ERYQoD7tN2IDLRbFZTLmzWLyXgrteh6SbVQZli01ytvPm9kl
z7+/kb7SDCzENHwGAH4scuMjQfYfOnmYk3bELphe3llrEAS04Z2vHw5DAzB43M1L
ht4ajr7bf+27pWUZcQ+nBvL8U1jytP8uPjKYT5J6AK+itQO7uMbsZRRPJQZLRS6R
qfXBasSeD3ahFMEcNvCX0GbIBZUdhu8OG9MX8K3cya1F16CFYXo9BkQoQt3vu7L3
5DTrjt/S7t7TUgJus9pxUFZoMS1HPASYryHATec47WbC6Bpl+YG4XCGmwT+HHu0n
VF1wkgVSpAwkt9KIujg1xwkzdXG2uGOY06igfm+nB6pKHoLeQdJiRMGU7CwgdyXu
`protect END_PROTECTED
