`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovYwsKC/g7H6OanjB1PKtcK+1Xodhei4ELsNYkfK5U5NaiE7IKfyBaklN/WxC4CO
5+viQO4MHtaWh0DRMKD0USn0wYdsg+7OWYvAXFoi+ZcYaMDcU9pGRztc7n2khi+O
itTZyvI0gF4vpyv8SUIQS3lPmRjh8nbkgYzNGWFtWGhmq8NhEVzu2GeoSljFNvC0
G4ykDMbjcuVqTeBUI+b2FolV/c1NmyRGu27x85I+2NlQ6oXTpieydSZcFn51KWn2
7ClrJbczBWvUpjsPO0nd8bbXO6LV/hLCUbBHPbbKcVk4NUt0HAdNsq2SOXcV0ywS
4FFmWd5twM2D8FGrVanoc0gEJ6WQSEOILL7MAACdrPKmYOaNM2Z0mJ5nrDE1wX91
laLNFkUDA5cV95HNTeWJTiyr+cPXInn9O3DDavnyEme9zCZsOjtceotRoSIYjA91
00B47v/4K8LEN3ltDsXIFjUoVAS8iMBRMohMhzTWgBdIYsgm7RD63zO4GpWqe2E9
499Kzn4DWzLArGxDZDKztd/BpyBj8GIM5/xjjpeWJTW0wr6R1Hgt/d8DmJVMSN5Z
Rmb9n1Z1YZkmaxWnaFUy+T0wMi9Ajgw9XP3X6JN8oqYQNnaSZPCTc000d42JgJnj
Q3e1uYGVwo4pILHtDHgntvaG2dXq1n5JDCwjoR0Nbic/j2sGuKujooLeScP5OgEv
MgV0HIZKnI9FE5LwBE8mr84HtYiCC63agGO8Daq1FNnJnyTwQ+dWJL7YvvIFK9MS
F6yg/J4DxX2SlPazQRh18bXNr6Aob2ebmdbLCbDCAScSV3B0rW1gf4m/CjQmGdaI
B9cVUc1crfmn4uZV633ClhlXEUp5uu27Zomu4HcrkUE6dAV1XSG+g3+MAE+QypGV
+24jf5jkFIuFp/0W1K7Fyg==
`protect END_PROTECTED
