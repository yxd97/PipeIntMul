`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDdi8L0MGxHrrpPjC080nP4iOAK9XkE4ILslbejjmAdocLvR51Q5f4c7whVIZJId
4IW6OzsWACDsG28osj6KsRL1RbDhyVDZpj5z0plBpsY1w4DCMsR76YDHnH+CDjR4
Oj1oL4eT08TvyXWh42HYo0kuwkuZUV3M7UrjezE2EdPOXxpWUGXwKF1p3ld6usY0
ha3czWb4Z4SUedmJ8W0cMhOL7jd6vo7Tk3ya7VgITBqeFHcRNKB5zpcNXaRaiLgE
OdFi5HycJ2WP4OifvKvNtcPGiR+1AyvZ7wgEhLvO+caIVgxwLbPTerPXo8BLF5mJ
rAuqi2OFFSHud6tL8Zhf4wn0uWxoaVNd7j5ZgKm+P6aUnMR7NMo40T7sH3HS0D0v
exwdmwSFHHpE0lwteyS+s21SsjfFnnDe6R8yBgf+MBB5jrGt3QE1Sjl1YFt/I7eB
/IyEaOYRCQZ16iWQAjCcqymAVl/1iiDeA2syfVDVEEt0RXywA1iPqz6HlK2iMEok
B0QsJGYTszMcjbFF4GRG7ky6zZGN6ivvtwwA4LdYwaflZS1n3zrpxBDY312IWLzQ
LLcGlRWQdsJNiocD8xnmzBo3w6HmlyNUl3WtG64n02PL7TpxVrYlJuGxXCTNOxzU
QPN6ftEazpLtYWw1GhwkLPeQ19GdeWc0TpJJIlQKPQrs/dXBAZMqjLsVAX5BRGih
eTCIi0VLRiAt3ti2ClKxBmdE2y9hRWeXLIdfVw8zLgg1d15+ER6Wz98ZKnWHTgX0
oURuwNnDHfzjqk7Qgk8qw1qMUgCPCOfwOCndMK02D4PLiRPGl1zhe+p3ZEZ3fgeV
mZDGXyvV++EiEbcQOjMPaTaVF78YyUdVHRODCy4kfz/145mRdunf2Z/CaXfXt/Z/
9EqM3K3VrqqGaDrxH9xmFeHlyg9+7OtMM2imys8mA6yZGXLouE3+8ZceEQhWiolQ
xf88/MePiQq9kFpge1WoQTUKx5gmLLzMIJM9bo9SpfdKHxGViFGkswkulbNOUz6V
W19CJrFsnzBcLsDFMdC+AMNMcmTvovrr9kpYgwwyxj8KDDpal9L1kNycO5vmvGZ0
DpCxIMejybvUSitmgV4QQZVIgw89BdReHvp3yvBzL9QCSNUAVhwCU0bJHs0bJvk8
ybu39VJS+rtx58n3PwMWEdC5ZDRvgdIUi3hFxZ/5DO2rabqdpblixVZXOzkgCyBO
q/XTKL+8rB9MuJhi35wS/iWQqzNXOm6MRPBB30oQBYy6uPrjondfihByLcQns+X9
I7/mQI+Gw0y1D2h+zw9ZMGcIV1TKUmkQ7rmEXYRskhk5B1d27IYKKDfKc3MuUPxh
l531N+qYES1+MVG8auaHcfCh7T6u1Is43bKVB5T1bhIQb7d3KJGeG+XGG/5BEWMj
3yxu4vNMMMvK9D1iPt+U7ZQ/NJehQIMM1Eymqc65wXHU0p3FliRTjI44q7oGok/p
HVjU2AMOl6Y2b2eLD1ecpAmwzUOwuFM/xROJDFgY/fnmNWdE0iETdGpHF1XHxRMR
ZNYjsP13ot1zeJMLjRdEjA5T8LxJejf69gmZ3MSLJu1xH1Q7vqn6NYCFohsqH5Nk
SCj0RmKfK5Z43rCClXrbT9MYeguveWoEysYy8nob3+c2SIMBGKzkfMHly4dD0DuM
sRodJc6eU1l9TrWTSn/EfFpFeCoDytk5GiEYUrN6ty+zW0z/VbazlFddAFv800TZ
VRy3UTQpbE1NRbn5MaaJkw532CRt0iZt11UaBFo1qy+gK/ZWoz5wbh+9saAs7CSr
ODP/a4rzmdkDBa3Vq+Au9vvJbe8mx99otklet1ipHURtwvlqvwLgYC3Wlnva6rOH
yNyf2dm/dxqFzztUYM/mJqqOPd0FgIjAZk2MU8aoBOTOxDn5tNzP76IyDKvG56Uc
Mn1M/X6EcCWP/gzpyT03ftgVb/PpgtLIZPh95M3tH9zS4CkWGY/2fLSBsxKhan7d
sGtwnWSqhlVa/Zl7ljrfpOon4Zn82vr9Ui9NKFj0ZQ3ok4wOUz9gLf+0zPld8JIj
zsiJ3kGNq+8Q71P2tJtSoRuCPbYqIZqehmeBHRCO1XtlxxIDXWWdUAd1kWUWK10z
Ce9ZS9kANh9Hhu1ulCcLjKR5E4St7NDF/O74p4pFDPBo1wF1ssNOMMaC1inRrifg
8/5Y4fY9YU0o07Ew73PEKxNtVpyN1LzN8QtWj8MUSckU6Rb/dS/ZDC/thUvZBNIz
`protect END_PROTECTED
