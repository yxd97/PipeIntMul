`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2oYJqe6/jmhJHU8lzG0PS4IZePgG0cRZoWJ6c1C/FzKnTeBXigEkoK4133vHi6j
o00hjDjkAoqanEx38+6QhwhPfgv7Mn0477ZZLJPq8epLfzIq3WYV2GsBQIlKw7V+
c8gBTxZ5BUjDD2nLXI7r2kjSh8KAWDm2e73LDs08hU5rEXNCIlFFXUZ+D/c8rvl6
3JnnzCoZZRyr6ap4GkfUiWXjeEQvwYGWYBozZ/tqxo/5SthDUYj6Gd921/JRhfgQ
Wxm3hziRbGAEETX1VzaNzi8c3SjyFSORQovjXNwQn9nF1Eb18cuqH9LYgyT7CNyV
`protect END_PROTECTED
