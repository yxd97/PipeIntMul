`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vh4dusYUJyS7ouyT60j4W0bJ3K779OM12+oQ4cwEIbW6GbO3cmwokT6VA54TxNi2
zwq/2YfMVpwhqXqh+5MsZ6IDvMKLtkiavcyzcqgjfQe6QqCbdniuYLafAStVnnSV
LARe04kpq6da5i6PRsimrAXk5KLzkq5xWXTci8YZepcMpiPw9+K4Jq/bOJvmjhim
VuaMiBdCiKWDw7KUUW0tl7uR1Az026E81nKJSKVOKdPNGZCOQqYNCLnPCrYpoz3d
ny8wkGXo41SUYYK+TveEuFm3FNI2ERL+NbIDGFm0m2xVPLu+tPfTDxmpjqQEa0X2
CtKlegJsCtRzVp2a71rI+GuIKeHko8Q8nhjEmA5jvvzSJe8tY+gxE8geWKESt/81
UBTduuGF2P3U0ygcP5sXqpSqmma1ae4IUKJApST8FvU=
`protect END_PROTECTED
