`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3EDM17Bma1KaypXEUni4KQAowFt1To7pBsAP5jXkLhFX5kBCWJvxntgz6ZGtREz4
+APK9oOru1J20Ks9ulEzpzWPzHYUEbg7UXPqMXSzViCeKe26wQWmfRe7GWcuADso
DYCJGjaVzSnmxY1a/kYpi9DXvwlD5L7HUvEWw/mgc5Lf2QRdNGkfC9wNsFUQK5/m
4t+RLag3dxq0zxv0Kb1Yodo/S0WXkKU0REOUVnu+3KFuytCkAZAe0PclD2JiNnlg
bFPygO1B+n/DHmeTXduqwmqKCUUbWvDeT3pH8fYExZ7A5d2GRQMaoiYz6dh6Zu2X
5pd2II6pwqoN9kJePBYTHFW4R/tPhn4VYppt7TuXo8Re/zak04hu5K+kqicIj0dF
CmQ4lJHCiXGRzHF6ABkiTw==
`protect END_PROTECTED
