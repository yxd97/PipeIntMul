`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bB5aIYroc0uDHQ0+0sS2abWWZ7/98irr78Gjsk5OKuZbneuzXWnNv1/WkaDooZjm
gL/Sa0t11JQ4VhFcIacfiwqb5oD4tqfquVhH2WvVJRSjiUHmSdptdm2e9qUw2+N4
owII9l3DJE8nIe5GncyhX6dtEkx0A4lOlQ8+9uwz8+sXf7mRUyQajnQgCeAsPuYY
1b9uddboLpa7CRLtTsVycSKpkqE5SYpSqJpKFXrJ3eDMXGOzkbUkjWOnq2YYpxj2
JT+vBHJ/n26Cm65opmiENnaEIvILJ7Gg8kLWIPD3pvLdjvK4T/UnyqvB8FK075Hn
Ziyu8snFNdge2LF74Etmi49dHL1+ryJ6du2E/Zy2L6xn1kJKZSRiOoQEfES2O9SQ
dmKOtuWWYDL6mDrKjCFTrhUol53RSc6O8j44I8GW4dGzhtC3fpTaDn5YpM6ehyN/
BLjahUtt8ZfELCc+lYiEMJaZ+4L+wlzEwMCrdczkbVS8Cj2ICyXUhnKqxcszG1Pi
gzO6clMJKBCKOvsvzTY8ejYXzLkkseeIwsuKUT7nhtDOS95nMvJc4fbotEawvcT+
3N6GNHcBAb+xgtFoin43H0SPiJZF0Wi4pE0i+YOMSpuzeyBHJx+A8Aiw0+QCtCgu
rhjis3RIT7Nf8yHAkqTzqTyGlbk1wG1fh6u2RfD7kzc1N24K4LIeZoC3JmcMQp2f
uGANOBeynj/4EcVNJGtUjJC+njD/blYYNKAGW7QtFiyfL1gnt38mWFU6p4ZRnwPE
Zay/M1DTnUMceOH15tjtmTLzX+Km1XCfHZ8NZhmPefUADFm6g++TYMpeHJ27nbd7
oOZ01YyOKk3NY5Jm/k0uan4GJeAJqLX56WtnsnEPeJXDPGj4Hx3PaY7X6UD4A31y
QPTDAE/hSheXC2VqHdSVo4wYNL31KLEw19n8Mw1Mwg1ydrlDKaUOE8BbBTqf6r2Z
B1fMVuKBI1i818KhcHJh2a9+2M8O7Wn6s/425OIM5kg4erveSBNf7vCfhyVPEu1r
uClZCfpclDdObJcLbYdcGTUpDMLDxii+p0D6tH1GU972nI3cB8C2cgW8x5sHKHWJ
zP8y4fN/Aq3sDV507f26QOfnd0df2G3+C/L+SIQxOPtQcyygEaP6y1tlYQjXTi3D
pydc2x48/sYlTMj1c3qUAv1MMhgSFUFpG6VNgIjlfrmiuOdQgK+D83khG/NEvqfC
t4MpA7iZ77oHGTLdPgMsw7WhFyw/TU6oZyEwCAYtORIty//hn5sohvUggrcGbNji
GHVRGQDiRXqg+BJCycOlyxH4fDhg5KlbCCHfpL63GRZZie5e4zLF4oq3VuVy5HDH
UGfo0LHK3Ev+VYraKPMzZianhsqToR1c98815JzyCu1NwkLf/NBF6JzeOQi6GX9B
c68LWQphDCJDqsC4r267ScsdZMOsCa43tbDTrnC6oAfb1jJOIyiwRWzHizSL6qCY
bwz28zek3fhNTQCd0Bw51xaCJLLmryJih5fhjc/3cFkKRln5oyMyDXBJNZI30pPN
kGxmZl2JizjBASY8eaDS6appAaXZ+gwHi3gTZEIzuAApLj0ZsNEaSolPo/ZPpGNh
OjsOKEPvjszx2v0vK94EeEIgpF7ELDGDI98bAz0wAb4ZF+MZXlBmqd4R8tyy0dCd
g2l7wKg6mo4H4nW62xtBjeUCLkSzxkZqCXeB/qxVNgn0qDv+GcOX2r/9GqxJkXIO
2rxT3mt4eU9HOSUDwQ3DLzJ6wlpx4FyO5EIuNCITABSCaNoNSJuVurjmDnNzHBfY
OAdl9qwKcyXJZ0QaTPXgwEnoc9SrU+LRAxdYhYk04IG0lcOXiOqDk172Lj0y3Ih9
yJBLaHrvkuzxoXCbjtM+RWJ7QtlL+yJPYZOC9FVG86gQ/8S/lJ2LfDv2muYqNrjg
uK9mb5IFqe6UkTLsc/ofgQ5jvxWjkqN5IarSf5tNaYXTj0q5lU58yxDMIRBOfKgD
hbP12ghOmCKOsAZ0Ni0dETDna9bhVWMrHcX11AHo/A1G99Y6okjMovWy2ztVzqWn
CI9heRzaQWVlyF8CIOHvglNQm1EGjzF5Hk5Ujuka0j+sjtkAuzJqSxWvpvatdNeA
r2sdauqnTvEm7toSmfRtMVE8lEYsB965i+mLj7ifWgfDkG+WyBGGj8swcYmMozfi
7gDDuufD1zatMj8F41UZrzqYixjICSTTcy+fip0+ejIOlUJOShsgTHkfGmgQyRFY
i3CJyPdq5anmqDQjbzk0fP7SosaMEV5KkrYn5n1+lOaH89GFKHLgQbOC05HOPtQ3
PPWMq3A9vBNqcNa1y9GMboI5yXr1eEP0XuZobNk0zmuvZaw8JCJM3XwqC2pjmiLs
Ozzg1ZKR0eJFY0bfdD5vSRXqU+o5MskywtVoDqWzWVVLlcteyLHrSWIszkC/He43
qMufxQ/CvX4iAGtj1DNzdP1X2IXTzF1wGZTH1oO+fuLZQdwIKhlkFfWHj2u96mK7
+LLDn7V9XjM+9752PQhrBA010zLfKqz7IWwBghPTtc6xzvXFU97/Pp/t3VIAxnkx
QOsEhNbvm7kRT5tmpy0Vv5a38OO7y77/mRXgUk6ARJHFHv8/vorJRgg+zAIyK79m
2J5y3M023B12ZHe5CuOKgLbU6hEBp4V0+GsBW68ljGpVoRBEG3rvlGH/uZPQMjqc
6F2RHpUDcUj4FkJp0BpWXgauI4xaElCZnLHKv03UA6K93bxwFsze79V1kj14DPcj
9xHIHCIyvudTX9wXSVZ7RMfFXrIyoVTxxRsHXxexZWI7PjKoaQ1hgaeDQizdQkgb
HFRMVgxfqsexMxtSrjStlvsDiI6d/m5b33G+fol14r+Jhibi0EsFQGTyReFlOqkj
p2ys2IVVxXlyNhf8PprOqYi/1jOD8Lvnyq8YFsYWuBT5mj3Br6qsL+8UJ8aZg+jc
hum87wmHTKpqzy3wDGH/vvxQORqIqeZ/5w+f2YMfMzTsU/oxgK6JyARFsl2Cg6+q
LPlcyhw3Kafl0aI+C5mPFt6FimGun8KfaKSOE/WWazj2W4gL9XDEhrkO3DCj0vUT
M5lzxwqTBek+DU91LWm1dZ5pXF/V+exwsWT1x6CzJu4P+PtK1FJyVEdicwDKCyQV
QqiTWvkeM4KV0KMdUvUYsmhCMz4lFMNm6Xz1sks/AqonqU5veqzLb/colC0wR9P2
qUkGn2GqUSJAA2GZvmZ4kEp43/Sth/QkU65YQ3WXnKObLKepHWn9uYGO5NJagNI/
RNHjWan2VuYANJiZneuptnFaWYND/G8GwSCITzCJoR2MSnxSpjFiikFdyg8YKMsz
papmclhVyrzgBRf829id1CsoNvolDqYQlFkdUtOOLDSxaoeXStUJDcVgdpYGZ1oC
WTUjCsZq1RozI86MbtbNwh6NjlH2TFYUj3ZMwMyIPFkVMohss86N1eau43/TWLHp
OpxeyQHEt0dM0CbkHBeMJJs3LGu9uEy6/OmILZK90dvZYQHxesCYPjBzz7/ppNOe
4lAZT++iIpQzLKSN6Kf6MFK/2IK/1xg1Ta0H+PG+VL26dhoXTQUmR+iKlgIX2r/B
Xajxiho4JnYxGtJaAbLiVO5bT30I0vvYs6M36FIpuJXNmkIbtK8lcgiciSF6yxpN
y/2hCaULUpBX8o3aUwoVvRQtfGEBjr7GEuLTx2b67vj6MHN0jUZ16aloIcWhCZLN
jBSWzQhc/KdZ/UqzT3htXeNCBbs7ufF9abnhDEbpZO3r155wNJ3V3jQkhulCLzFA
uwiJUWazGFKZyZDXIKSYWZje049W7MUAhsFdnJZwRBZdsDu0spvF4WbPvQgcptuR
RVw9Oq54bWkcavEubQx+G0FPlNxY4EiyZ3h9HFAu0FcKSYvE+moc+etP6wbxXD6L
mZuo+eOcebgP8UxpR4TI8993X0b/VHtdktt1yLhqArlyEsz4A1Io1VECzsvn8eJL
YP+Y5EOb6uManvliY1RZ8cxjQTmWvwO8zjGA8VSGqxOqKY296Q1El3DMEed5Fbbs
tnfjfnt2schVwiln3uoFEMj7+S9wpS+++1M2RGsVo61SNtYK+Lp0JWxvSfaj5RCN
5ctTROs0btMDVaqBw6CK2OTsd+s4DZwvpXPisIQ4yFnuupKmfyV3UrJ11sd1EK2l
zPRyV934DQbevclhK6plN7wvc4QQPFZcR6plFsBccAErXi8f/i4l64ySJD46iWb8
FZIwGondBADxl++c6fJxahUFBSmSW9Xt+86k8OolPP+ocMpooEiqih9SRpYPlDqX
+y0OYUSGow8z6DUEFXZ8U3UEhj0auOiomsaYrzVJYV5p7hfWoeLTHYuv3Y35fBw9
0/+Umo+akFN9Zw2L522/Bqg18K2aRvFTPaSSJz9ICAsm/404QXUgkCbrMtB/FRTS
DDJfF+zLIoZ2G9Dhm8LbtNEhZjqtw385+TzaWGdKw6WfB6+Ppr7mXD09ZmuSi/lI
l84iEbV3uHMXNk82zBOpDlj7nQfDh/NxUO33hWx4pFPOnZmqZ29Is3kXXpwY6Kfs
wdXoMtWORqcqi1vYjuMzUTFwHyA9VC1jsvnNVX6nCUFjtRVKz9nUfvuaFr245Fk9
sirrbaETMpzrJwU9ua3cTOU3nb10NA3UxfnUOkvu/PU6/akFbcz0tXKUE6oEBbHz
CF6Z0JnGNY59U8V7norhYnL61BsDyePhQYWto2fzjJ74dn3+vqGSJwvTZAyb0ZzG
oUtjivXic/e0UeYplhi/MB6r5WJNBAa1HWMehy3FYhYCbic/7s7SlnwvWMLwqExM
fXz5O5k1B0mwbWteGuM/aMoLa1fwPddeXKj0+MQrcCRLzQKI+WyqAjujUKiUD4XO
m1Hx+pYP4jzwe3EIiXz1dZtAsjVSN+/VYNONeobVbZha19q/JZm9IxRCJjxPOnJ6
ftp1qohno7WdrVQHhee7YW7RXJG0f/7sVF7hnirA1FumgY2MLHVal6wdfhvp4Ulm
sEbthqopic+XvQ47JDqewbCC+Ab4bBut/NsEoI25h4lvdm6peGe+397RoSpMlXBn
XbEpjOz8vWAYCVh80+9jLqKhYCaNcC29ILJd8ULeXDaeGn0Y9eamxT+8llXYQPP7
lobnUwNWQYmhvPeSe7c1uGT9hHeu9jHjX54piQDj6pu1tC/s26xWeqUm3D0vyZFZ
lFnJbGw3n6IKqpjp58Lr/smpTROVYHwoRhZSTV/CmVm/ZIP5+zIPsSDa0FEci6iY
ObhgMRrOxUZfr0jqhSb49uSmE9LvJlMX3QoDFfzBePbAuuVTxEO0qgmTEPo4YYEH
CqVoI+UQR4vLGb4vKPFDcdxG6Qsh7FK/GYU09WqEI/HQudpCDn2fDvjKfUDgnu4g
UCAEOWANI4c7zfoEfQccFB207xxbr+KzLJWS4w34cAHvv+YfH6rRaRJBrsloPFab
2jMj///VFo+sE53ggEs8osh+H1AOszwqcHwXeEFxuoc3WmmY8zfeTdscTnvozq7J
uF6n8sCqusxolqynp330nUuhfjgPTvQTlNwK3LY5RSTid9cVP2wly2YLxjS0ExFb
rL+5poQbfh52W+oRw2PUF65OIHh/duToNsdz4obsyo2yjcJGbmYwRB+1tgcfjLM7
55prKyEkjuLeyL1CH5oJ0PY1BadPf5UaHih4eIpArbGrL0g8XVxvPU73ffU2mxXq
SFqugAXr5fDs8yGTLlpZBDWw50Ya76nXr87z3y3Odvr02IDvMY2Lb9dJJDkoiHyv
LB+jEMR8VBDkI/bYjxHmgZ8W06rWzWk4g/KDSQAXV46+ll0WoKh+45RurX2+n+6m
xz/hFyvUjY0GC1ZrPJUjdCQNc2jDR8dlLByV+pLySTCGQLFVt1+uohluv0TO0PVC
Pz/0NE2R3YKQcDVipUKamMg0UgUMuHNVTDq01GMuBS9CLYtLdLmN0HKgIzU5PJLT
Vy4sihe/Ryxa2AY815Yg9kLXssxPkZhbcCNLetUX1DXFLIv8S8dUozGOMi8OPWkn
WnI9Bzu97/Kqu/zXD52jP2NRb3NpKJFN9smQlEL3VnP/VTMDFfxg/7XtIZFKBFcn
OMIzNNUU/K48Es8FrJBdqc52Dn5YImEJ1e4pyNArPY/hR2BX/tr9F+6CMVduE9cM
keDFNb2Pc0ccZcK5oHrVKq9f++bmlVsNNPhx9c7DO1DQ1gB2swNXKX2K4KvT4FBW
PIGvT1NPVA6qjv7Thwj11J4GVtme4vjGA6NUThcXg8Cq2sXWZ11+BCmJBmzabBfw
SPK/XJQ4F+/fXr+ecxu6HJ/F3p14ESG1yxV3EmyTQ+Vl0+bx/2dkLYRP0ZUoHbB4
HJ6mCoWtEj7HNOaEAoSKadcyR/95bzajT9TkzaIdQnZ1UkIlrQE0wAoRpsyI0tQT
m0mmihZjuqrHsUXzeqfX7Vww5K8MJ+Nkd52zTuTJxQrF/AraJyyRoT0rykKtFtC5
YZrunmAcOH4LIXe1tmi3NQKCn29wfsjiApY/UhF/w2+xHc3XtOgZcjISwnopVsEQ
m2+287Yw+QQC0k5xgejD7Y9E0/SUIy6N0Edzx9YduM7XEncb4BT8orcL1qTIcbDE
Btn9D4KiI5VcgqDlkWnhbwPmr9/Xsu9TRXr68MRfzTWRfS9bvpD35qZIW8+VmOi3
uikZFDdQOO8i+qyv05ofbRwCE2W2lmpsGmvJIGbUEwF+0s866vj2lEzl3DFwRIs0
Qq0+KJiWwyw3LRsg8wqhxPoryM1GY73PW1adi7oX64ACNcNI1HFoj9ph59CPZoYD
WMr7t4w592QU73oJqVrCZD6Km1/kbRV304poRLNc1BEP+nAkVkop0CkAb9ID3g7L
b1ngdYhrxj9/EiZdwh5uyNy4wDdnr2uZpXC8p1KZ/ZIU4SuSCoOpjqOZc2QYwkSS
WMIbuJfKSziNpHKEQRdCjuAPaa3ln3Iv9QE80tVny34cWU1dHt1Z0Tfa9lhafofQ
nt/sxPYFPzcLQl/L0QBwfZu0jo7//afUTfFT49Nni5JU/wJaKHPn8PxyEshvNatx
Vg1+0iWfL6mhfNAmAJ6fma7eILshNQXUL9qt2zSQ2ybCHpuJRNoQlpNIyByk2TKL
xec2E0hCBzv5/2nQkRywQBaq4olmkeicE1j08bms6fgakqJqidtuOfPqQAmtFByl
Y7zaoAwf7p99VX+sa10rtQdLTe3xgXgXFSg17ppEiYBxBL1zLqVpuROUZ7qDvF04
xpLbgh/USyoBbQzuGFX3FloZktvr9z4w/usk2vq8rKc0sH5jtqkutojDplQRdut8
7uNvyt2LjvMQDWAIdcigKiEJ6ILTLr7eqUS2EKnsh2ScWc/e+c+qj8gn7+EqJJXN
3wqj1f7YaTndtboxq0bCAr0skJgLvixmp4sxRWQJTmCusOEpek1UIBwEQPAYz0gX
kRoQbzSM88aJSGsXNIe6XdfBnGmPZXCw97Iu0v6UoFKysaijlbhOwpfkM/FpWKJo
Uk8qKZHj6K3fAYnIq+QDurSLPKVZHfOBjUllb1hgGip9q5z/OPSKZFhQR+LfpVJz
tC5b/WeW0XnZU4/FFoDNsPCQdEuD+U8FddNBBu8ap7+1O9Euiv/e24495N14lRlJ
pCtypWPxvHzR+B72/h/ghGM9FA3QGIsbL/ZYywmvpe9lUvF57Mdw7zTRSeYCTFj6
hpqUuxVdRxL2DAPXH2HXZBFMkqPp/xUK0OdJ2CrEOMrfVYzw9NqJk1rwzS5hlTZ1
ww5E1qyqQBOAVfOUBXWtD6b/Mr4+yV0X7KpyplqVsZuItYoB2aIIoGQ/MPgKtf64
mjjCRF3X2/XA2bWA9YadibuVPJzSjMMB2ZouPtnpaIltse0VGA1fxG42pTDYvwD/
dgl7/ycH0ydNXcWBWOcCdZI6YSLd512YnmMWWpV6zajrMSgymtZYYl49UBkzb1HS
Ejss+sqejysFikkT7YT9iy3jKQroczXd0oVSl2w7kamxNtQ6Rv8a/S/2UtY+f+Ng
ag8FcIYppH2JWHrjFfN1nifywm/XL8hAVT/Y87YJGdda+BCh2ozt9f+2s277MWzf
CuM20Z717mmAOIJ4lPlrjCt7TPWoDQ8r1qYOVCVVckcOSyALhegrcNrbLXs1zw0P
SVGQsuxEkoQ3NSMl/MBafw3tZ3wurkOHhQCVm6DRmsYFz4mY4LdQq+q69q5Xfzqq
unQ02MEotatx4nj1V2WJ/xYSkLp6F9YqgtNFbVO3QeDoWpHfDFDxxxhS0pXypkWe
SGz/DMrZijns5HanIq16QIngxSUb9u6N/w73dewqgpuaygcgUFE5db99X4f42NcT
W/W0PF//hVubwbFRfPcezlrvsb/UBq1wgYnh/4eMWi9PEPOiP1rjhbnGlPu9tPwZ
npBRY2Vpu6j32TtrUrs/QGc45aqrKscJdo79C2MPjfOuKDFrgeiOn5Z9JtWFXEpV
lC4alzH5WMtVibFd1T02vszyfFnhK+U5utKiYmgoAGUcdbZHu43RB9V1eMtlNVfn
FtplqzxggP6jtkJYZlrHTrBjP55fFaKAPDqYo2R2O2zl3qJla6cJIABuOAmOQWQI
gEStmxB9X59E7RcRHWlYppvOEJPs8o9ftOHEM3ZcIjNHva80cO5kSQSSue2O5X4Y
nC7D6RCJ8gdBPz5x8xdkoxHYRQ3BK9BIDam5xQflXZSqb6P90O/9ZWtcpmqKXZgg
wGnk6G0tX+sBG9aJrQXZKsHLoNleq05ANkJ7CN0Tzbv7ymUceYLdhqbfS5jhWB6U
TrGNaUZYe4Jz4DrpTsaLaNpRPykDqDeuf+6S8mmJbbmAuiAPs1F90USUugkXdMmF
7H0K9XqlZUeVx69ptsnofDlGETQBv9FPAnpcqhbgArvWbgduhTESXt79W1BG2rOL
VE1nhIEBQeH/isPPQfBkkj1DT4LAhrYOA6S/1h2woYwvu/B5R69lJshSvrjK+H6T
0XwdJgKUu4cb+gHkXPC1LOe0oaaiqGHUYM8FAJQzZDJrfdHAppw2hvGEqXgZHsWx
jlaLaT/zJ9sFwkgXlPMsst7B0+WZk7tdc56gVFnO691k7wkEuiIfjDzXZdvzw9pb
Pm9CogtR+/INjJ0uS2MgQRr6ZESqr3mTSzwrwmHI4D9tcPSFAKMORX+gJVZuAT6N
DLAThzz77d+Fzpa98hcBLJwFBtmVZfPYhjEQLZ4UJJrh02Ei2a4ad2RW4uUxXyEE
pguGggivT9/X4nDSaAflizTUd7QVIvDGxGuVCwPl5HOVuUoEGBNAavA80uwgbCL1
OKs1ApfNO8wpqQoCUCsk+EzRHuDhFPPiwDeOrYMr62n16e2HDG2MlBDJvB1OIYiy
B75Bp3I6ZUweVXNk9ILuFYSZhP2JfF7yGBgbCm7qZfkdSZQz3HGeqKvPD599HSz7
lFWKXuHz0pm/Iy+bJDpmhYQIEVO+btsrgfVMZ4u9Gnh39Nt1KC2N8KXtPzQvWbTo
u4qJ6FVIGT2Hf+/phMSSKj12alQ6RdvtShyJ/KtLNNCBWUPvCrGDt6fVMHvbULAY
J80gru3NNIDyw4aaVt1T3PpTsv9J6cyWie0jjg25nKDX+YDW0YP7Srm5d5OPTrDb
IXqBXhE5E3iLMmVT5t0wt4qp7Zj1j6hHR85LJ7DEOooadPQcYZ1YOChimsIC6E1z
ILqdSWMY3BnjWCQOKLEGsUb0MIWYMMuHzmhkjnJTCm1LjYmFoBNmTS9LOtqvmgLQ
57Ib6FrCOpXxN+nt8HC7YMqIXBAQdIHCvjCBPm8YqJgsOoKn6ywsKlHkfyMlFwxE
aes0yjQHx+07w5rVXBAUeLahIW9a9GXO7HnFk0GX901hwU3jhIWCejl8M5lb+/LS
QFwF8MK7VaS2k1pxT2Qrv8IalgbX3Ncm1G8Rhih9l8gfkUmBF5Nqd1rS8oJyuHAT
imbYZ95UWaOiLnzmAPWaT69FKfZ6jxDVFDTrxcWjsWYH4NYP3pcq7wAs/1VNijJ5
cX31MZ/XezIyyhcUGHf5NVlXGiWapbcwWF1A53GajwVLhzKdzzWVNPVZFF7kOe9N
1FnW2wCW9wYmjVzjK3+F8kuIocQWXHQLhbHEawM7lbyB9FcH4x5l2fad02xaM5oU
3oNU1OMPX4Vawi0VOowvMrn1GlC+HcFzQreF/GmrBb1EX5IAwaQ8FDjev0y8V6qU
aB7ylKXunUXumvoa1/DgfwRZvmfW40xQLhx9NfbQIu4sNViV5g0ZcQUDuLimQtpI
TThvgkS5Z3B/slBVLa0x+RRVWzGwi51tfaSjicqwzUPnoR/4DVINWxDAd00rW/bL
6wpDPCGXbL0gK5Ky9etARm5UyhZl8Xn1g3WTANPAoiQSTxVid8KULaMxFDv6fgje
hZ8hBqzUlQr07fftwOyiuagdRscLbYMzDkzVZkEj22YAOYwfZ5gyuU4O62G60UJm
/5zI8KSYMOBmy/4mhotH99dDl271YrRSlvqumI+hXLX9I8Bii9zS3GFmwRaHDKso
naykWLIAUG7a+12yrOm4NNGkuK1BypjM62I7NxkOEPthEEOk9xdHr74VK8WnvYN2
lYetOrpj7v/aS2ZmXZ6Ck1E+nBAlDasRAhPykgmbpgwaiTl1JnQuKpZABwXKA3dl
VpM6mY9kunPwbrSYiLE+ElfVAatGVY2kd3gGx2s5u4+S/7vHe3kVWZMCpQwN2l+6
jfoVbnz6gpn8uAvDSHlWZ8oZJavbrpLGNv5+hZTPMGxqHNqm3EpL1GqVXhL3rq4r
Fe6nCYFCdskzRA+xLHql4LiMvNHvit6POdg57/MCH1Sa2rspjKDntSH2+WWdzXQO
EZnWKTjFam2ayrQiNrFd0rIJfumoazMqObzLFCso3YAXPiE0EABPBWyhqYEuEafP
yfVIHgUeVeIpOUkGDgahmhzs+R7V33d1gGFe5RWxZ7y97Y+vkznD6jXqotXZAOI+
s3+ipItiH65k1ehLpgXFsEyePSS1rAz3/ysu+gl2kWjwafmA59hKRVw4FqCJewV6
V41iQtEbHsLf7/lkUDfH9pk23n2mqi47faNAtfUthLOWD8AUznBljmkBtHunyDql
b/Xs7LgeTvdCBnJ6IyiqHDLmb67WVgGIGIpiAgKF+POc0b++Zt0CNvI7MM0RkGts
C6XkimJiEm+vEANcz7o7vbSBLwFDx2bCqjOLFQDMV/h7OIxRHuq10Pj2MuqOwnsB
K+GVTjfiMqDduha7YQPQXWnCrj/gaYrQBoHPm6DNZES66db56VAR1ZHiCSs0/ajy
43JAqVJqzGQjOwD3tircnlOooElRfKsrbKKfyM3i7A9ZcBJ9cQ7ob+AGDZVJZoOg
hJKiDs2qBYqw/hba7jhdLkxJt2yviEO5TsgIik5P2Uz1Q7Az5kj2xZ16PlqJ8z2z
hrYpU1gIhygXF1F/pzuuEHNvGOOpHIolu+j/PsGjlWGMCwPimnhdOy2s2WwAOLjo
Jk0M53WwJNyu70XDeFK856GXoWMMXwcthZPSh6qCP3ZVT2ZLdu5pZkfpSlH/GsAi
+UntnI/czcyAoHNFONhgNbEH8ZRcFp7AJT4fWUjHkbNoOyqErXhDOlW80MhxPbBs
nXwU/McQUJH9nAkLtK/0aAhWnN/YU1SjWGkmblU+l5nx/aYIhVfHOf/LHhkmmSkh
SUPlDuh5kRZg3t9iys6fP8qX8klAPPAceRHGg5jL+2PgLp30g9axOl7j/2pw+0e8
HBNERLoK4CBEfcevKP04+tF/g4LvxM2N6Eiu0uv/HE47GxFJFJF/i4J89WvVPJTq
Mrj4KADy+q4S+rvLpEGodUAkAfM+3oCKjX7FyF3fAUuGuyPUnY5hImQP0AoCHXy7
6rfb/dyQolS+yMNcgSKP/OvOuzoaqI0Srus1+l7CvCqlJw7JBJm37n44kgbGTZyT
h+vTI1BMAKr9kzAhFQsRDSuW+FaDlxWq2jiLkB6rL/4HekTMR5KSoIlQ34Ru3ClS
NIo0zhhCuo47X22fSC4LBzQ9PASgN131d7sDDst6uB4wR8x/f+19DD20VirQVJaS
V6WW9q2gaXMAW4u3If1xFjGehko6HpFoHamjFNGI+3sqpyobh7FXtfzL/xeYTbx6
yN8KU3IZlAa8pCCY3QzjFboQkpmGVJirgaoW8auqDJApfI6insRt2PhK5ERDdgFl
Dhs/pEkVAAvY1m03/R7dYseCs1lPHF61tigxVdrfYnYgHPNSir9KueRQrpJ53wS+
PnrsuvzrXDwL4H82/Gi5b/Mh5kdnpS4JMsFLet4kdrB0IKvaX1PzTYNf+d8CuhNc
vQQo9DeXfwkICejjgu+f+8kYpx8Cot31xIMEAH+qbprgFUce4XJDenv1IUyQCeXq
EUy48JfsAYshHT1gifZG8rRYCY+emz9EBW3r/pLEp+cN0twNZb/BYZ9ThTTGm/Ll
WjupHcAQO5mTDMxqoWyYgEvTyCC3xSUkuUQbhA0jSMKCzE5WLjVEXS1AQrRhbfLp
c28v3X72ZmHNJNo6pPdTKiYY/QRQNWNi5gyaE0I9TcJrF/omTTASFU2JmZLy6wHr
4JjDWlSOdZQlJUx9gLx3AZnwXDn745bRNcwdCqObUDiUd91ocN3gFNyh3HJsmMin
1CQJbW13xjC7EUGM9G0xz4pS6fwbeAv2DU66i2vG0arThcixSTGkLCCUTAT7jJcL
9LjIHQH0kHEpFHqXrn4SAZlI8r+xSrk6z6W+ta0hIidXszNlaFKXBv8/O0T9NNK9
wWxMR7Suqb1rKg04VZHhnIJNGLjvGHKK0J72RzJrEKoMy1JNFumGU2KvCam6BwN4
4sPYNdagj44vdzpR4zdTChdGOdDi2xARaEMtl8JjCChOu99i8aTbsJ/N59XBJYYh
stR6AiSklzskl7qUgh8lDTZnZmT4T1CBjobVNfEwGVHBLrQSWqqS9RZWKRIgYOh2
FinUD7EU90OlMHutleKouWKwx7DvDGq7afqID+zrjIqVTI4KNeffiz3DDE2r99XQ
dWl8oCJnGq9T84YH5/p0AzgRAUTzWk0by+vqMKRY23JO+82ZCYsymdFJBdtpJrxi
84omgUXnXH0fWAU4ArYNTqDTjkoHfXiRPtBuvbEXHU6eylHtgHu3KhN7hjtIQl8y
eR2IJGkFXRS2sWddwWYbHLCyJc4UYtyQXvqaeL7s0FRJft640hIiP85d4w1kgqyQ
LwGyE96etG8qfvCY922tAX3Qeh8SjFwd4Tob6Ewlbq9WCoSnXwUGJRM0Wm6JbVfR
IUZm4pfoVmgsXqv7qCJif8iuwvPzi9qbf9MOtnziISpWTnpq19W4QGX9Q6ZrO41d
cKyksKbQJagzPSvR1fojRTIFXDULwOMfyElIwucpFdh3+p330Q+upf5EOcq3RXG0
tcQXvFDpLsuV5v/rzXB4bQsVaWoWLrh12rau+EPcUYMigmRVpeAB/FZaOkcyQTE9
pgHPrDlS/T69x+5jTHNHQKf57/4+WYOcI5dnwqFT1DzA2gbEyu5GgwyIPsKhFBcO
l0PTBO9pPMBaVl3FoRI562VyXyfYL0TqIO39dBuHL9/urheId6R2AeFcWNhHQ0Bz
ILKOpn8fam9RrOjhQbkgSh8lfL/UpkV4XxjdSE6a9zZImalMYbqiEE+rTge1SN3Q
JPeycMlAWfU9qnBVbDmuOQZJHaBsM70nTK0SZrm09ZSLYBI09wd1yNh+cgyig3TF
UNtaW2nuce0r260hzi6Xx7HwCX3Dt0GlAO+x0sLnZoD13JoDTIjOSvbDH/d4C5Fi
qCUzj+k44JUtRsMhJqQ56ooJWU0NTfUZRCedbnMB3fqnH344m3RAxZzyBmcuFcmG
yjkUa1r4OANCW6PaA1EEpUGJAn263Q5CDNQrXb93T/6nQW1+LUejyteyvDwgodde
7SoufDlb1L7bN6kpmQ9UXE0AS05NNAo0cSndzp3BO7FCFLiYelnfm9nP+Ew01fx/
l0vqu7oQYhsssgZhl23sSom4+sYpfP9zapA+TWWO7oHAjcICPRQHuFyeVnwmdEM+
wMLVaTfPD6AV1esbbDVcZHju5BiGPcng77vYvUBaMTz6a+jd8hvYevveB922ay9r
4DeB9tUHzCEYQ03P7304Fim2SRntv5hye4glVsbRO/cLa4vr0nsqgaaU2nlOUz3W
KIMu7MqVd+hktAJIYF2VTDZTkVZLaGFKYO967EoVp4ZX7QMH+QSzv+ooYSFAQ9Rm
tm3qfgXBl4SwBCQN/QDEtP7WSZyRfs+jzHFMUchjAc7hLaDkGL4S+9jVt833pUE1
BhO2SNiqn31ALVvU5JeTTIMM3H98ee8S1QAONEpQveb2o62MZI6v+pUZusU6g4FE
THHXPHTMtZXxePoLcmbl5/gRDsJqDSqN0gzYSN+1WShFXgZ2P+4fiX4chIQrSYEg
YB2gHlogBtEljrVJQBJwLdWtDb6wksol4fw8y+ZP1PMH/jExh2jvDSghihwF5MP6
eJUR0gWWejF2w4CUbnrm5eWvlYLFTDixrnK4rLcY6jIxLCz60Vd2KkiyGzS3q98W
e3gHI1i5dfmfbQnoPaBvRkejIPAdVFJMuuCl8w/InRmGg2MWDyYtw2/7LNgwT63D
H3Q04vAlelZhYcw3PWxu8qwWAsPeEqIo3C9t9X8lJhiYx0uXBS2hl6b12RocM/vp
z1XIPhtNsSm8gArcKB08iOBKmkAu4zXGAfWeigXB2zvNLG79EtTZwLuTFUrYHam/
V/P02SjTtLnwOrFCs31tCd1jJaXuNMEcCRODX5thLBsxXRZuQuNXzIcQ9+vM+tTC
+QdNetbIBcvTKshXh+RKB8+RYM0gEAFSmDgik4jb4kbZstpDpeK8jKCNjQIMP3UY
jfmCKDIF+2mcpcNGhBtjyI7G4aCiUo/us8rpVeRXFa/wKT6AqYqoLJjzpIW5jyLI
kWS/6KicAbjT+JDvPXzkOBb+rauRMX6nEhNjqr+gdwxlbWPIRXOTUgiXHqQHzQ99
D1vybR/Vp/LiK0G3ex82kP09JV5XiGZ18594YxFG2fMnxqEtL0CfAKeL1GRtB/5p
fVhzu4cDmqw9AjplTVVPMsyncqxRiWFmlaRo1rU16A0P08CuT6RZoOByoP9hISsa
vqZBskEpNwQf3jCXG+Wdf3awJK+/DhCUUUv5nGZfuLT/GRGZHn7zprL+AGRPU7ru
vdYgptHOS43fwpQACdVVjr/l3wDtbJxivgussK6Eh1Nkl/MPfvAJRMEPRLhDRgqz
3E35eE7G6otSb77YUlf4Z01RngfaWLhxQ8vunDLsn0tkUnN0XAU4tZur/WXtIBkJ
9cj9jvQrDpWjaUX7NTtyZYcu3LC6mBskO5Sl9GhWK706uepm8YXUVBIOc0zeDU1J
Mt8fD9iBqFkt/AgwrnrK2DxZzb79BWOMQrrg2taBCRsiYh78XN7zgGXw87te/QMk
7E3fmhotqoCCZCYtaUCuwaqb+VI34dY2X4VdIz/PjJ8TssWEWxC+vNbyMQWIc7Am
aoY0R1Yp2U/oZ8No0Y4Q43F/zjKyzz+MykM98quqql7sYZu7azUWrecwaGzwu/GV
CWRIp//VnEkQa3dgXFG5PkCC53nMm50aVHAGG90alakQXQ0hv9fqQBWv+l4z+oZt
tbDmSEvnAr9YbqTc0q6Vtg9K20OmKXgmGuPcS+7qljyKsixYuAgDCSl5U2PuBD8A
EkdJPpXrNG7KtJkp1na3xGVaGlFZ4Weze1PtQ0vm/2ljvAM60ilpoLoaVMDNa+Jv
zEOcyjDhF7QAjza48e6m3W8lc5lDOB8d5AyV2r6eRsaSxDnmthph51cgczffjcqG
2HR2Dl+1lwpbCbgq+wckOpPJPaRkerzAXu/1mSVcQIB+U/lfJd//t30HnFdZPNxQ
wYp32/1wbFG/McsZYaYf3BxOxZDYdukMxvkh5O/pzMp8NYL9wHpjiiIbA4qOjUGx
KiWjA7BTTRPLdxDiRJRBvsq3Smw3ZmPcGVIzSXDGlVqbPAh1YMfb0X+K0P/ULkHx
WlFOG5Cian2W2w+v4XCTszEgfV3iZ5z5H5mRlUPJGVwbLSJzURdpHBpp9bA1YDSE
Ftqi8jzMKrSNLvW8jmkgRZuz9/OZ1z3Yylv45BTtDLDkWiCAoCb0P3rk+ygT/z5S
4L1ClRzwJCKxRywv7WG8eFryLLbt2PAqR7U2t0CedTim2hFvyJAsaY3spJ4t4zJM
pSXmk/s+uAde1uUkZMtAiTf8dSfSqAugpKHHuSGtNuV9TlaDsqW4dne0eE1pungq
sMnpELkZ3gl3TLFpR34usNB0U1buqHDKLoCF9Ez/gqG7ahVhvxXk0BQDzDKTzwzQ
05eZei+sEosDg/SU1xlez3aGGg8jSAsirTJLfIL6Zgc71blidPVL5dpp1GXMHt20
60BAwVxGKtSk1jDweoMMP7tOzzkv50Cpr10wovo5bHnRE1ho0qeKHd+BmX5ixBHn
2cwoRZaQQXgowdh7+p4ZkWlmEsNvnhGe6eylwUq35nbvBIW7MTe/bXLC/BNVCfYJ
ssnKhoT/aA+AMWmgn2V90uJHk9NutCzzOw5oyzkUsQy+uOKo45+7RFsj62A3LI6n
UEkqVhwMpJJLtYE0xaCFhR7oVHINrnWqy334mIzDRRV/9DQs4TJszUlveKujhgY8
60r5jtnSXWlfpKmBgdhLv6nis9CtL3k+TBqEYnSiaCHEM9GtyhvXPPDtUHXknwVy
9f+Ot6Pot+wBqfwbxbQ5aKwSkb+49HLA7HvkW+jztcWWInf8BEoqi77FCjZluuDv
V60gTLX0T/nH1V2I4HQP7ubJ+xG3U0iLXwPbVmQslYSFQyO6TW6uEOESfWOg7x67
eq7VdAQNqRVgn+LM/1LrULtJD04WZkgne0lDPBX5ZgvqCSmt8pCvtE8q+xGAYYv8
4/xggPI7BpbjuTIv70MkrkZn5sCYVPCLN+fAwfVRJA7352kY0ag4lrtNDWYiOe2u
9dQXlJcJvWQQFr8TXOkMdT0pH0wMNOdi4iZb7crNtMuzFGwUu/aoyo/EZSXfVHr0
tPJrOZV6O5P7NoXbhEdL6Uem4PdN3M+8O+PokiL19oUolL9TJfoMO2rCD272Nzg9
74/btqR9jnCfIxZVGxb5NnrObZmfYm+dHH1k7sArkl0Qcf5mJ1k+krscBkYp72rk
eJUQSKAvlSYprJTJqneyY+OAluPWdFEFkTki9SqBHWuCEyfrOItkWalO7ctRbs4P
5kVTsNDnxp3MQUX1hzMkWaH4usfZMS6+xhVTNh1JrsPEHOfRMWYxhpF3Fhk6fiiP
jyaJrz806e8F1N+B6iqjTod4QT1s1FF/MGNjjtMXv9r40+GcN0folthU2S2ZnlHk
HIlCj2fXjQVldm7UmhLBkRad4cbGcQwjtKTwS0inpnVgFtBwtGEOkTAgOteWLuMe
x+TtgxLqVJZ+bt/MUV7MaWVlriyq/m92ynEQL/jiy3RZFFXqNJ52vaBJQH9CK9ME
HLSbP25nRrkWIw18yHl6B53mcZEzH/RmxIMekEyEvfoz1CcwdFov255tA8JSLaRE
iB5nsH0PcSAWmnpXR2NScHb9mxMFdEWG7dhXkJ0KgHD0VF21Uj85IitVFa1bPgOH
Nh9CqITsngGS2jENdr+osbNgtKBei38pef9yFpCxIFSkKuSRfy81i7rapqnkrGJB
mkhsdzk5ivB1JOX0JX02T9Z1tJeD2r1b8WsHd1XnbtAKgbMSWWezKbw/am66mXwS
zkcK6pRPmeIGOqTtane9OEnTaC/VFesj4Z9/zdVsmMUiDaqz5DFlcffQ9EGfsDMW
reyLJmr6xFB48vPYBUxNgo7qoelfuPpCwynnTLEwzKO+FaEJ2CspZkxr+khmXmSR
aTe9Z4cv8zl3D2PKMDsF7IvZ4C+kCgvgcbxSgSAKbED6nsTeigw7GA+EsQGBn0m5
d/8PQzcnatM4ASiz51ew8ghpmgqa85kaqMvT8s1tJb/K5lu3wiavswkazup4SpgP
R2SgEE/IgOImRIlrdIYNDS8QWFAEx1gZTxDI3LPVrj0l1OWRbroaSMlSxSY7u8E3
pMCrzs/Pk80UpP/b9qnevw9JXcRYRvbfAXaZyl4O3LkG/SSBweGHclCmjsN1c97I
IIe90C0KqravGYF22a7fKDAFWCTMuCtcXvviGE97nKKujDx7cxzs8CQj3jF7t/4P
V95Fy4I6B/ZmN3VsM+aohWobXmurrW7R9qmoT0NfglBbhuXPTivaaZyPU87vIhUu
qSL+K08KjrkVls1WmDvh+uCuU6xSJBucZXcoeYJV6TptOb4+2kow5y04OK63KhAi
40DD0U86/jBLsAXWUmhNjIqxbuRlLTt5ifnIlcwp+QPq++8nDlvMfS7sgHvXmxOt
lni6XfeVdqtj5hLtP+G6P0JtVGKVM6wIjYcpKQfT6CcUPUKTjW7HOcZrcrM02Kpj
jYhF5+tETPnVcUksARadQkyNqf0Biwe1fm1LcilnAlEjBGlATbkXCa0iBiUMuLmo
N0RaqSrtTye1cocWwUc+xfmxHKcuTzVjJKKtblSpSsomnmRXK/CWPKjZe9+/Nhgm
5bH7LA2EMrGAVFWFkNkxDc/VRwOtjXUEfiybn9u7CE/KOdsBnLkVok/f6rQrNtBL
PrOG8HMikqkdZy8OqLKKnZWyS4UCk1kDciDzTzmYJ/SWEbcL2G5+ZJmvk0A33Svi
pXLYQC9LoJlrBJVj8ZaiVQTvwmTc7zz180F2BBsG17S00fAPb+qjXhCbDQk+4+BY
XNbBOmwOly2WjOO12S/ff5fjnSfLYC70wy8Pl2cdvApF+rKFw+GGpt/fp4MSsNjD
tClavNgylntVZOKM+d3ZM4Nqq5W3j408tuHPUAft0c+UdRC4pArn3k97lKKrIbEt
MEmT8ouiQwnAaHOaTqUQw5VVTnnyXw7pLisi3q99CwnMDbTd23Q/Z9Ntsd2BIWws
129WQPz5H3kZ71VAKElqyHQn3/uK6CD7uBRD/klDypt73fQG54MG0kEbvulYywKS
vSWYDsOivOU5j30wjS2Q0cqQ2BcYyWsSPNgiQ6otRQeb2RgSFJ5cX4fAVzNdTnWc
cDYK8pI9E3mtHyw/qcPrGr+buQ0mg9QGKIO+QCpzc4JXfI6uZoXtNn7g442S1kkL
38M4QihP6/L/EZbxyOYsXYbnMeriM2b8uzk2z+VbvXClKohQ0dqSb+xmqBnE7NjP
1H5SXuCRteMe5MSWPGOWpItetcZOcNSfZlhV6YRH+mZhX405PQZlYdprswvYAW2x
JYqNBcs1zRJ88TXqZsnp1Z+Joz+ZjlwK2JgJHmU3Ucgq8mHRlzIPGFYrMDIDhIKQ
MuCOVXZazX7M5FAE6pVpIfllQbM34L/ircXASSSjl5KCEnzUkvaL9lto5CEpxDZD
Tb0DTalqBans06NyHKXX1mclRUIC73O/2JydYqmmQxb/9EzT+fVn/D6VsDTeborz
xNODU67vWmu71fXtSEkW8H4Lx7XiWzzThTU28seRsd65O9hBe/hxcJMWjcnuHI6r
bi7i8n+3Gi1hGgdnZFkuy1MNbZJFPjgiI8U/akmsLHgtlPhUViGhthRgDF+6qhr2
YCfbEx0TxDYI8pdhtg9wHn3VFxfnL8Wm27FWmfHytolM63H1IdujJY3L5F1ERh/5
a7f0ksRFoAX41nSGJ9VMWM7ssZkkApaFyzgjykT/oZA+Dtxl2jnAtIO9Tr9V78zJ
qDQAP38VBoz+oKJzzRKlnfoE/R5h+oXBB9fYnxVn6hCDff7KIiUFGngcI9LXUkcM
E0hPz1D6roJqkmgNz+HSS0hYeZchoEV/GyOL4GoQTcuZA8fl5VvDCYeZVamSwVfR
wpRK3+XXJqaFz+CZm3t0X/mxdkizAu7q5J2cYxM2En1+cXc6mtZICSQrH2p/S5ef
70a8KYxDKKR+q6u1mdIqKupL15ZpPvwiI82uAjVGCGZd6rkbSLl+r4Cft1GotdtU
pXFGqAMfTUwfWDDUHc/cp3aQRZu3v9gQ9FO908Sm2bvlXgS/QtLrppJzw8MF5K3V
BNjKoOyjJznw4QvGwSWvPxm5D4oOcYRmWYQpPGJMSSDnYa9KBOyryrz1MWqB3rn1
/53CVqjbtUC2YotnAPSq7i6tz48QiD0kA7BQwgTlRUvvB9HD7BLi8qX6QyZvwUu7
TyoaJlbdOJxF0s8TGuqyTlvTNAWJL3RWN7n87T5wIKGBTSDkReuFXKs2oOaQxx9g
yYK8XEL7+mdayzPDb8RszQUjHpkRXqSz1bD6ueVOqzs5Yx555fF3e5dGXqQ3HWW/
K+qucru0iR9tBTH5EeolHGhKI0VU7r0uoEb8eIuXG6FBY9yfEi7qobUqZ0wFmSie
0fHuDzBSnfE7VYVlSpdIwPMFDCJqh9eqEZW6Q77jJ8mYtN4RWwgfzmsHws093jRT
rH8aeuVmrHp3xwWMjAzvNpMNMyWyy7Q8XMnhyNcUet7Oaq1ub11/psKCqyj+9/qE
/FwQzwADXFV3fTu0ORlureD8f2n2l/YkJToFILmC1iECseifRXPf6vbASeQz4fPm
JvXMZuW7uAUKJ4tVYh9cENRURzkzxBMFdpNw8HcmmLGP+xLt80fPP/Xe99liF76z
KY4j381kaAC1ItA/MC2TGfgIBN1MmvPH9tm6Vr5ZA35gP2+3DzTo7jg59g5p+mDh
qmEG87i4vnHBDWLe0PIDoYQvnxb/1Y3rTYdRZTTx7ffieowPTXinB8WmIWNJb821
5TR89Uw4DpMTjJOeIGpPGPEQo6wVnTZrkBaVMnv4YmDVgPyambGLMF5nbXn6FrRt
3uDnMW1gFhb05Y9YUpsl68CdxhkYjWyKdWLqVPUVZynkPDA4wfwQe8uscqLmBPaf
GeI923eNmVkuzsempnKdlSvTiRknIr4VjnnsZ/lH1wtfJzPl1URT4t0VlMDS2T8g
u6XprVM7ivc2g3XRodi3vSA6NhAQstsg256qzEmXGgrpxo+/HkvKGYFVjJjwzndr
fg3RYbQrBI1xJ8ywEpaZgImpXvkDWpTTwrp0JKq97e01V9RnFz+dlIONVjCstNKT
1w9RmF7cA1nH1gK7tHC7qCNJ9oMkXbE3cYnTXQOetD8b0Q36eJARyRRflmE/As2p
8uYRyFfjEr/fZWOOrU/i/BfMJ7GKLA4L8f8Wa0acC3O4mrZkNe0zK9Amvhk6FQrZ
HuV+6ce0g38b3Egv39A38uRzAYWVWXxaHIMJvOjtZGYe+wfeobywxnEQlakvozbl
LIFlOzFoGSI2hsJbp4OtkZHPzEt7UlL/BoU1B+XxGj6N64EAcMQBwYcLqoLbhC/Y
9XdTwJPaLEbEin7mZ4laggNptty7eeB5Qc8JxYmLBNII8bwsh9Aufvf0+sJJoBog
tR0PCRbSSSDGLnjRuj9NdPxowV+QRlKPnNalaENPdxI01BXJQN4bNTm5cN7In+Hq
2ApXR0dcQ/7/4jvvvVsp0DgHJ+Z3YKpVV4KU+lAMB8mzU9gPTOhf6LTQ4pgCzNZ7
1AVC0gMHjS6Sz8Y7SjDU0GFAq7v9vrgffY9+BSAxioizqJgYQnk8KcqX6LOQ8gR6
W/Do/L+Lqdw6liBpni2k2b5v46Mu/cUwJLnuYnLn3V9g7UAdjKgYyQfebV2xzdT6
EZRPDZqGGDg+dRVxdaAM1xITWA/7H2MC0gRap9n/IU2GzmRfyQGYbIJKrWLVDszf
iF/bAsczRhr4NBGAMLrCiaFQ6gGIbwKFCrL/YW2Z9CXm04xQaYzMCB/+1v6D2RID
VBlZyZrJDoepRICSELzWkszZICeuG8Dr6ONBjHUBt26XQo37JPbcU42aF0agGqBe
eBD8oEgPPpsilq0DtrLJ6fqxvqoE44YkjgyCykBWCMk40wb5ZAdpKj9nf76SBYb2
3TP7ZcCf8UVtIym89Yy7M03MwUHvU45rn5EVud5R+dR9Pf/Fz2bVxyUuNL9qwaGo
6d8VwYAyyrj9uoeR+XcdCL8WcXG31eqacddEMs90hxzajURisguF49z7Bj6WV+GZ
swa82C4fMy/PqBFifROg5IA0Dc4jTz0hngFKy8h6AwKR5bGJZXKGaHthiWj3zznE
nZ99qQX0Rsw+zv7Iolr4tmt7wM4qYph0ImLNYUU/R4Hc1Ihjb8JTUWiq24mraqY1
PBe5VCLDuRhoU/KtwCBQa65vAsMKQ83z10+FRNsrpVQfG9DXMwGQp1H01WRHZ87l
Pmm0o3Wu56uwX36q39L/h6RvaUUh7IkYPiYSkNSLlDK1fw9Y3U7+ubMUueULzEpb
xMWU6PrEdL8Z3qOS+sUHA0h36D25JDGWryEHRxcHD5t7ovGJZvwm7/zwZDZ0SEWi
5R29JO5+eVqYlmXHpQQtDua3Wap6D8xmyOXyAegMyvoU4cfTsdo6p/7/9Gt/kuEy
sUOA3qsecl6iYdXDPj/k3HYqhDa/raAHc2KJQJN1OMcVNisZPOZSPR4f1eNDLWK7
GMLkZZZ4Vq2BpKWGoQln45ez0NZmUiK2LrVl9ieUTq8HT9ujeEINVRQ559iOnk2Z
3/Pfw+qeBHe8mPcelUZbyQaK0GUl0VHGgwd8Qhi3N9lxz+0RvjEPTtIdT2x/UIdc
dcXVqDIh6Vd3Mne1hoyiTVKiCK6Diq9jQMPM4ggTMbX3Os9qbhQlagwMXRm6JE5p
v/o0l2XIVEoedzqcMsGQzj/Z+47JlRWPDMt0tOfJiePrDSIsACxmY8FCovoIiTZx
1+r+PKKgn1Q//igLKRx6lbrqScAUGB0Ol+R/JtzFYCgBq+Z3eUDb0HnEYglHYBmy
42BSXz6DuDOxf1tPSqeauaF3QF9oi2G/6JKQp/wxxRHoqgsuYgIRRyBLwpSl6avu
Ml7N/vW3Xr9fRFdFCNgw/ql5VGMrZOKqxgIEvM6j2p43r8DzukkvijRjMmyuFuI9
+CF9zGqdcXvFsZlYGbT+5U41DGFJQ41HaJL8xXgkktte/MpdWYF0RVlpwzYn/9Pb
n37xZCWC8jygbZmppoOvfq78p8j3YaUo/h4N5b/SU9LbW8PZ3AZZ7JBSfov9Bh7I
/WpY4v2wNcV0p6y4BSFUDLUKAnPIoQhYeRc4P30iJzYrTAmVOw/dBUPX+J5CS6C4
BeiNgnSgSu/LU8uRTIBORvDYVndAtiuI3L4zFXodI7W1n+6QKI5aYyOQZnzSgkIw
l75fnc9XhkxkxhOGhwoBhEq7p5ull6s/HTv5n1dgJ6nfe8aywNAPUha27/S69vF1
JYZeEz67N9jpFQEs5cMhrEHEvD3jpmoaJtjTUsjXf2bEjzaZCj05R1WsASXW5/ed
VRG6YagsD/Ba1UBnc+8O4pTsE+gVZ77WHGGB/LOz0u01k4qEKwJ+mFrLyLZCj4Ez
RWYff5kOD8aoiWS6wpCq8mefeeD4VUIWmdMzG3dfz3HIW88wNNNmY+ZQpouxfnuW
6FywYfMi/cnf0SupbOICMXfsmGHElXbb86p19g1AICVz4wUReS/ZHTlqlfyZgyn+
GGmU7oQRueE4ZXuJaEpZouZJCi6mjEnjW5YmKIB7w2RtPVn5cUBJjIDFK0WE0PqD
HWwcFyeDMtz8JpPmwhr27dJeLXdZnm82II0Z+jc9eg/MfiFeXKPWaZQGDVx6RcJw
D6I1H1Cv4uVFAQMkG9fm+d5mybjRC16qkTA1UW53a3rXD2ZZrSHiPDuzAMkRO/K/
cB1IZy7b7qhoad/IU5RCZ/RYfI4WhHgrOqUKO+rS3mFqOQ5PHJaE9KU+uoT9UcT4
NF1cNwFwc5U2JcFYCL53Za+UKy/g77K0PekUtVpeHS8otJiGtZstUcDnlv3HSddL
nIxyydD/PqyY5L7fi6s+ttg/VtMNM7p8HNNiUyI+Z43S/uwjWRI0dZUnDJlXoILf
dEhyiOhNUAQwCZKmPheA9vUu01YkODdbsyju7fBNMFAj1DfNxwyPkopT6onwVRAE
woRx5dbqwhQeKSoTgstmeoyG/nmmTYyL9wLbY7BennVzR3a0qw2x+8KIzeyMx86l
YADTSGFv1McMC1lK7mvhNUPiB5kz5s2hE2rgVqcibqZa4T2IUkwzEk4OQkRqK5uw
X+dxQlQQh7LhdT6Zn4RH9UDM5KXDa+oU4wlW8pFqtvaoU47rQ3LtKIeOsUccYCmo
ht9tQQfuf06wSD+pfw0uHLHxJGjdyLKyo9Cus53ufZmRPrK+LLnDeyJtoKDsMST7
JsyZRjX2iHwRZmwRCyYFwc0peTjXYiyXYABaCkUMscafW53U58higICPwjQWOfZY
lHN16I03OIi2SnHLRgJuEXyKkKZUM1KVqpEEnaS8vgY+WibiO6bAK3dpkH4CHBye
MruvaUBiQA6atDmxQfGzjKsXqrTBFC8gPspfdIh4vEcgwRJSLUlKJuf19kxR+BaB
4FF09FlMONg4SpgIPjOr9V7lS1E6/86Qx5MGm8aikC2psx73+5k5ntURV77BaGqr
39HIEVCaxdpUs7w1eSEwDurPGw5n5O0vb+gLTtGf93E115C8/edK3UZRkSGIYr4f
Cga+TC02HtgvsPcQfLCGoE7cSH40ETzE4AUomvDhcWGfXi8kXnC29lcuT7RGxizu
CuRQfzALEih/SAmfpjopGeM4pN/1AQKbkVfnhYnzuZQbs9JVwo1FyBNb8tfylAnz
J2JjPSBqrhhS2g4jBDp8RUtxTkG3+7iSuEr/SBMHAEZSorB+ylXagGoKSKQEIegK
RKn70NWTpI66WaUJWJ81fBhHyR0ANK7JS60ljGKj6AW+q3TVc4GYL59Z7jXv4PHK
Q3ZV3vXaSLNjn+AtQ0/skuNCQWcUkJtd7fGL3ULZSLCiwb8JLEMwXD/bgEiZCR0d
RIxCj9lBEyc4fCeuHjg4mODF7Dkwx5mreiZFLGgJp+96p9KMENGvUN6iqZOxBpVI
OCTTgyJ22hrGq1qF/jHdQGUmXsZRB9y7qBBVnxzAX9vUXCyKOo9B8zlCNzMNYJHa
9xOC+aZTQ2LxGoZkjlcDnPBJh/PYc/jCzPifAi79okSoGSHYyhW5puvObdVjh1yo
G5GCCkjkNFB914u3arawfZEkTWLGOu2KgXz7kfdTzHklhYDudxFQQa/q6JqVtoVU
jlvfiiCXYBdOwPdXJo0RKgA+OjSQ1y+KzpZInOi9J846/eaWBtrYX9fkJXbhpgXu
kYQlIgIO0Axr1rmV3MslEjlMDoF/em2q2kA4rItJsXwH/s4sqBzSyWSq7Me11KFg
jbOij5B79IL8KlAKkmUpiNOLLOL3fuh+mHKBroriObrYucaz1Y1W5bYLvmOdrrNT
EpuqtgWSzLJRcUXpoTjNcU+6FctRKxTqibKoumai7p6v94MV9pADjwGdegI1diID
CYixipKZdnzp0Bzwp1UCqZ1YMH0uEqBr4rdIlX6ht4+Q+JVIBSG+T+3saqEdYrUo
3qq3Q6rtripqr3NCBrFXwVa46bhr8AT44zUFonBMya72ZIsSZTd+ZqLLM6GhXj5p
NNII0FAY+6Nfio8oT8Nj3QIOtx68bn06prCjcInOlC7eGDO2n2ZZE6zEGKqhCnP4
ZwswepBFwefr/rd2EPgWkBo8I6FoLTn9CAtRZc10u8GL/sSHn7gPILQs8asItbuJ
jtTQ/QX/cDyB3eoROyowseiEmn8jsNNkPhQwxSSJIOnPbMHQhXHNtH3ed10nuP2m
gr4D2vN9ircDXpMm5/9IwgZGI7Wlf30lMVGiM1+2qdokaFqOZdoZVZm3Z5U2ZHDB
G9Rolxi7cg75SWhP2E4pPPIG94yfdD5DnaVgauy+z851KQYfdUen1lXA0Lo1blVl
E2lsYj9KWtCLRkJGWSgKxgw8lK/iNf8KD+iC1BMESAtJMHHOBbTiR4hlOQO551yP
mbGBf5PN15/4GuLQxiNj0p6DkNwt119/2ajQBs8ebz4b3yNUMRHGdKNw4/w6HFnS
WWrYsqFxYcM4FC8dNlLbiw/6kLO2sWQwpe2VRlgOUDpXURte/CSUZ7XFcTB/bkCA
UUv5HLzVRtSeaXx4rtBZTRDxuuKSYLSrDCXSXscj/mDPvEnZs/ucJe8zLB3ij4iq
zsLl2QCbOai2rIXtmq2ODUJx41jm58kuDRjk188CSMd5RSDo4aJzoq3JKN8BmqtI
NNI8Ouqpe/+A9JFIWCccQsWJztlCHBKAg796cxe8IyofTXRNR93TvzzlmVgEeqXC
d5ayVtRmYpKcx1txBXbErEgeSiJZZYGvTf8lPTdQtje3azJ64VvqntD5KyQp5P45
oc2DEi0FAS4mjifTr5hnIe46LQzwudDC+M2sJbhVBxdSBS9fSgFCzPSjdbDPx9Cj
ac3+vuGW7KEkFsjZFfZ098YQDzgcnj6fkaqvmcvNiFTyI8SVNsTThD/DkqHpf1cw
BE3f5JlAc54n6VNqtJHXGbx7F5+r9u1sE9OA59K2zFMg/eT18Tv9GG6ZTh6gp2i3
m3LH7Sq+MvajLA6eqUz6X4Oa7jXqgCIZraTM+ItaZTGtqcGmHEwbQGeaqUlsTwgt
v+m0+qjeSAVy3U01aD08yjZH4tyj9zwNGD8GiL1PU1WZmYypDMcRtrgGc8RulWmg
JQ/SVy5zc5pe/oUnDV1xTgLG7cjgnToDc+mNILZ8K8UY3iHdXtuRPUdRrpZrmajI
mPrhEQt16yfz3nmj8vfd3mPjKVtsuovkARghIkOKcBKvJfjODIJt8bjz/S+B0u1d
0+VXszr39pTTpR3bQnFFXWIPpg1CYiG2nXLKkG8D1ldPrXL3/YFbx0IJl0Rfu5xg
ezp+cbDQ3Mx044IYuXxJGhXzNcf7ruuGZZ2TDxVtLT7UxWMQXHkNxlOnRlxgQFxh
XzKNPa+d5ZyH4TmkPl77wLe8XuLPMvf8Rf/9sn9Jf/6aAildCwM9nTqBE+MXZudp
sZIQTvANcM35DACEK8sqB16ksDASY1LdSd2UVnwW7OJ5x33zvWR9HuTm4Isb0O4L
Xwe44R7CIC+UHF0B9EurZLhHRs/M4a8R8gLtshcFakvdV24FgNCAz7RzCarCeA9H
TC9DqxoIuzqGBj6jbHAMOhcVd9YnrUuwlZ7w33+cyj/uQkRpHHF/Ns+jiPtHXhrc
GoSFEniq3YRTzT/0c9+lFKOMtRCy8YSrlrJH0JOLxFbjnQzeV+ez1/035aIFLgV3
i/B/f+Kmirk4CUt7YL9SjgaCnaBQeuFe5KpNNiCu+XGtI/aRXwabS4hrvUER9KLh
bGQmRbtAMnZePPm4fRpCrrUt/9VwzyC1tVqrcxptRy31kW+dCv8ceKsS+L3CXsss
bD2syXpu0zsDNt65ufQcIqOsdFB5C9NOBKhP+sZ0AxPrw6+gNKAKfVJywP0cfuMq
+h7SsE6j3qbWTZ1oBXcTswJyr6+Hte77K3n35tyDGUBWFNCilkb0pZHA+QrI6kUz
sJ21T5n4W4a1INvLGxeqVZMrf3k52pdQzqnDD8jWtR4WOCE4wEF1W6x/JRsYBLb5
nuVNJwkonnoL74bERLpnfbVSDgGvhBK75Gb6gqw0wMI12t0M/KaM1fT1HP7bq7OZ
utmZXzgf8JmAENW2h/KWJVeU5IQeTi0wxLHsTxNOOpZu/SJKj3KSyqqxfD91TFJd
KnikOyGo/6bzxwuJcd+w/0v7f+xCTmRCY01a0oX4Xjhh7xNAg6h5NhFPeNB6N80d
O87YGsR7yI3suVF+rlzjpvix1eCrxM3LPPbgBazyudQHQJH8/bR+aXmjvlvnFer4
oSf5V+MmOzD9+TdA34gMqykRGBO0Nsk9atfADoTU+bLBk7QDbr69hu1YMnIyGl4u
ei4ahYpuPwRGR98XJJnCZTKhS5jguoRI6+HgLHHxPdtrnajKdD8l7dKq2V2ulCO+
W6ZC+CP6TAftxP3Fl4+J3cjeRspYxbsNSfWFMjFlJ699g6laINLoQefGthK4iL4z
kI6ILdPodXZbHZcc3DCBMpFYZjcyzG675glCu6kC4jIu+J6xYAeCK7i9EXHBEsbz
ZzSddtcgHN0UCi/7KbqUNgcqiBdDi3/HyIHbUla48RIJsTheps3ARHdec6n51S+l
evWFSC8mRwPZvezWg7EapEHRzGso5NkcT4Kc6QGr1f/wPzS2Wn4c3EgA6JEidl0/
0woDM6DLPj22maOddoYoN+2f5m7IzODGzccR97wsyYUj9x4rWrBrkWt5NTdJSbzp
sAVLufij7ndam7EFG9F97m6IWp4Rfj/6fqvpPFLYjGTFkmdosaEHiQW+HVzIW126
o/piz3sM+J8pOm+D1jf4vayf6f8KQOojOwSr3kfJFmRGnAErjfoO5AKSkKWFXPc2
JmuzCyz9kt1ETWko+F13Z/uiykX/TdkoOw/6gmTNZLTQzQtup6yGdr6eBnfXvklJ
iB9p1lGR0sKQYzdM1oK1Jzi9sIzYkNerBD5mUXLPsxpXi1WTlOPOB1zhvEuK2MyU
/GFRJI/nHzjfAWjT/ZvksPCsoJJGziaDqQp2Ds0x11xTIrpUNt0675AN5MCUUR55
RsmvWF018Y1ityNCvUdZ6DaBfPTGdY6Iw/Q3vJH1ik8ACHYw/QD/Pw4JwKUBw6TA
5KtMyc+RhXrX/5W/+hZb2i+SeZXC98FHCUYHD6jr1S2VnLZ45N5BEKK3tBUp16vF
TmZQPL7BTXEkSQHE3q+1CyAI4sTkxWveHekrZwNr3sXcv9Ntr6d/fRw3RSmkyPJL
iRLLKXn30XekmO3TByhiDixrQkROyQax+hDzFANtQ+N+/dRvQsJIQeMmtYqFjJbc
IZrdhlZpHprElUYcotE4WOcx+UI9cxsUqbhQHbyuDBZZKuEmcw4KT0ZgotL5UZN0
2Uf6qmcGHwTzst1q/Jzf6KS2qBS3wtTX/KmbhgygOn17wYz6SLqriON7Ty2ezGnM
ooPdshRRpTlFk4fbWH/j8/rShZNOM5XM3niPvd8BmOr/tx/dLQDc88SwFscc5wyc
3ir3a6efZMwF878mLOSGroXJghAVv0MTNobERpgxvXSth6ymeGccEahJa9xYmV0B
KyUY/Tu33VTfTR39AWXPvzYc3UCFT08UK3IX24nQMJo/xz3c2RGs1z81rX4x1It3
WC2XJsc0NNCSOTlBkh53elDpebyXC/K4dXAK739vloKsOLuHI2I9g9B+/ZjPuLvj
zSw6n2wbOYrg9ZFPt6FVlGYyg2hYj4AvVuZOQlRYhsFrgQp9er5yOEDuDQkaSjgF
JgVVxLPmTdiwwsbssvP5zlbgk9nLQcHP/Q6SKJ5Nbc7TT2yD3F+saMhcgycWQp97
vp9W3acf/wm8xiRjo/4L1aUjvnRScbPbXw+vptymOi5jeCNNNCflnWX8ZQycnl6f
V6K03nJ+OtEWTisdMRCP5Jlj9+V6BcmTIspww6tJePzO/Zz3FJYNO8QqAXkCSLeX
3cnWp3KXUcKFbECfARsQ8K3C6lSVLbq4CVTvuxlvUbtB9OzBe7m9s3UNIRUcXYwh
IUaWqhgp1mMwvcW1Ms1Px+bt9qSW36qkn2zG2wz1IgYNS5vymY12F9Y8XCRYhALj
38c+T27ETjVzVBca19AvFBlBSgTHdx8zyIkO+lmqt+DNDEM4huQUHI8CPws3MKFZ
zLGQRSDj2uW8hGtGbVDQtcTWHQI8m9jEjRlGmXfUFzpLaOILy0pEHXysTgbKru6Q
m3wuqXX/bvf0yOfucaZG5UG3mYEzalfmxAnnwBMHcBANrC2V+hU0ykOIvwgzGRrS
mLR/4BTnSJzYmN1Kk43blUeStpVZ7V0vDVQ1QGvCWmccl2pA2YM+6VlnpLOgEG7E
Zm2F+UoYVxgO5XwJQME/omzaFX8y5kQ1jmJUesuMRY+qxEHDYvRsPsrH7iqx3NnD
DHCcRE/1Cqg1bqQDHhSqKKkteYW42LRMtMHagz2GtxUq2+usKCNfx4Icr3vn8Xv1
xG37+J0YdKbUh6XfWujkB4h6VuNtMaHzwBn5IciACBPMr0mZnLRJ58N+MpxeL5eB
r9mA1NscDPosz8MRCDHp5kFw4r21FxLVDEvsidK0BYvGekXjSe4jCMBIrHzU2Mju
3eCCrchHWDtitZCtJmXe7Q0P5YnLiMp3i+Bk3UX3bt1x/q7kaCisx/NR551eynQL
+0nc1kf/K8Jq+kqqANmxAspvOXUtTexE3AtmgTZ2YtVLpkkdT1xkPZ/AjZ0qfdj6
wo76enWdqQl3JRf60H9A2K4XC8vgcXMxJOfAR+4GLEfdwoR/IjW08dqHBWArOF/i
snjAiR4kymNTVO4/rP3U7MqHsrjFYKftu5qdXH4rYu5w/bFOl8ayMLmUO4rBLePM
ohaQvBYesWeNblo7T6t7K171IoTQcQaYXzJmZErrUavjDxlj+hpUWrIpCquf5C3L
JP4pKoU+XSjBQ+iNMOrPvi1p+h3v6Yt9kQVQZ3qdCU677JdjzNo0aLpchreLS+8b
QStrFgDv7YoAjk1pN5IPvMBKi4QFzM2wBFmAVVCe4zUv2EeAFzKH0SXD4baI4X0S
DAK9Ih1smFzRc2xDvMAyASUgAb8DPLrOiTXHLZ3bYzKNQdRNepWn1lCDYneiEmGK
xss5jnVmkQ3BvKbkvPepBPJUIxbiAOCzH2qoGxu0BOGBajO+fggL0ttNZ3TphHOB
dO4RlgoIsrDAHQ0n1WQsWjkMkPgENZpxBP5+cnbxOlzZuP1IL0Yb0v/2aZ0kGzBL
ljhLi4JWHduW4zef9hTC5Kw3u/nXIRtwo1+WlxyyGzNLhyyI1IXHWSm0hvjc4cyX
HlR5g/025SzbTpjZFg+LkdYNvwbkZE2lxxNUz+ru6Pm8BBapoiEHaXEad0LZyYW+
l933qTJt32kUIEN4IGZVb5UqYX2sauvTL3oP3LpaQMx1js3ploFg+2jYxK5C9paA
/eTEuEuywnPZSSplmKaWSJRyPnz0e2dXnWHHz+2c5ukNNCsEJjSb2BnnFiJyFAp2
Uq9PhqDB6aclMAqgHQV8MbaVgmufhehPIeAQSc52uepdjzEC56LtqpJUpPDrkY1I
jjs3GN0kIjIOCVpaiH696ctF98PWjp3ACo9I8IsnS5fHwCUUXiThjR46oMcP9O1M
qovnyKNrnm5pBvb5bsTyJKiQbloYuUFQ9+Kp006TESNKw2A8QYjJUqTaNmMg8hUl
UqNPMDrcRpnCI2MkC9m7xz2dw5eMOkx8u0JhFmARbWdVNByYXOxPp+VSBvJ3EKgH
ryWI+EFqqo/Y1Iroxu8KtQUXez/vufwnbn/qohv5jmGbTgr3skRwZBM3u5840CUh
rsvgBf9VqYc0PZBQHW2+glfJqM2wkrPgXylNIbZS95oooTYXnIpn4YKtqHeMO2Um
JSkAAMuMOZwI1v6m5A7PCp05byzDt8nFQyzcNIe/heYsfSmQuGwIP+9aOf0Vs3l2
fUra7iHx2czm6W/9wvg6o775F5Wqu245VQqe3N21IWQtYOwhd+2cr1DLx1ckTaPL
FxVv9Qw3lFVRysVT37VGUT+noiUwpU2vuFgou5rXCdqrXEa0MFetXULlcCITRdbT
kbcW2KqmEX/BOCu2EjB89I70DOr2rD2zFTeeqopKqr70dcdVhdfwRTIuOJgraB/N
YVG3sgi8PeHNyVCfAN1krmDY4SzxeJOzxcxQT0Lcx9pG3kXZLKxfM+vsmzAUE8fw
wR/+Pdf4d8hEm+Yri5gRMOHCJDjz7qGhxWrCu9N7KtzFdgfYLzaj1YiDxIgtGkjU
XW+ZL4w4Vvdu5YlLb8vZdizTLzQ/WjPKRZbcEYHrhbRzi7tMYlVhlj9UDGoYocKw
6xB2j3csgCgo+vu37ar877LLdcHcPbQ4kzUqLWI/ssnPA619sTjapHIGkTFEgLLy
38/KRJkMJGGDqffJir7YUOcLmrZh9fQ/f+EPxmARHQBRoOU0T6kL+0yR9Rq5S/K4
hin4ADiTVAuJ8Bj5vV11XCj6VAyrUaYy3S0B3DxY/oB6xuowvoZqFrub1G0g43Tb
gkHRzt/ZzwMjOWvq40buwJAu5UHX0MnxLLE39Z6TU1FGdBrbc8n0EuNMjSHmzR4P
cXXYPOqMjAMjDogOfM7C6bdEAi2288pzk7MBtByQ3YLAwiLnuHMAhohZnldvVnlc
SJBzFIB8cW+jGcQWG72hb/zYjNkqxnvHs4fz7cW/yrKjD8nDJNxygmJvQ0o8buSH
tja1RP+SPU/Rsf1bYu2Pg7nM9bJWzGo7wD2LyM9KfXjkdmqmeeGxsFoSJhab4Qym
DVqDdF2EgMnE/eGl9G/JRXfSdJCKs9BA9aPE8Rs4uFWaCFaL1LM318d1sInbApMD
DgIcmI+C++LxrdSMtaqn2Bg8p5nva5Zmg9BqHwOI1yRevOOkSmKe42z4FqdUaxXl
GRizGhlsMz03veMT4ajO0XMEvU3bSqSt1RANYb5gWx4xhpjhLmuQHqJ4/h72r9eY
1QiD/FkVqcQsjrW1DoVQklHOzkkMH6hugizTwzMrfsftG6tMFJKBfPZ9FQID+5n4
mzV14+uZyfnyka+0dL2C41/S0eAuCMugkCg6yj3RYBzLtw7Jjy11bY/tKyegth0x
1Gq9WKD2SqK4hygF5/uKDLSe8zKCTvwoo/OSXQ5DURfFjFxdPU6tQ6rRkq7mR39W
dH7AgY3YJMMjztf+bCusEpNYhoNq9n88veEeVfS5A9pTEK20IahzJB0SVxShTpKr
JUR4MF2qWdnbSqu7i0W4JLxrJkbKYLRQxdfIr/eLyUv2BzyxH5adrk8b4qai0zCo
5Y1OlJPVJXogD0YAh8A7Ga4yUHiduI3NyejWD3NGfCCdc2oybafk9G/XLCwXcVQz
RvI3cD/dj88fdPCUnkyezNPAfn2o80i3Xjpg1XnkADquq34dEG7QXWWryROoX4Co
MDIkV6l9gsNQwQYP32VMrmvPKsYZf52sZeB89b1jaxFmWFbUpDUY6TMaW0PO8yMd
t0xpH7igRRkXZzeRJucY82WutCny5N/rlzKVtc2YnuNLg5hEY79aRHC3WIKEgza5
8rqyHkFd+u14AAksc2CCNHvsH8OcFK/OoEbFmMzYFAkotVNaFIEtvytYW8P6thpk
aW6rGd0shpNWTb2DseKPwhZoDAmYUY5UzIp6JREFVCcmAwBB5pNQM7fMl0toPLKD
7Al4POVVv+EjXklX2t/KtHoPPDExpjoM0hDPoWsyP1ciZasQPnUWHMS95LCZYN9t
22rGvi3fEGAyTYA2vclCSb5xOtUbH1W7nfmj7WOvAk5xzbWARaoPQP8/CTdIaJQD
lrRGQCzWEoPgDYeM0NNTzqDSXhZfMxXdTcPN/cFfZH5C1fw8yvG+zFZj3QUYyVgO
NZoJqUsbLVKE91W3cmfd9/lj8Lsjn5opbq37ROxv7i7oo8+cJurquzQ0arTYmfyY
33TT/FJRMiuXeOeDxG6W/7cfVATnRs9Q7vsBsquoHQVGd7i06x/W+hsouXTY5qnX
5ROE7HHXCJsGo+60G+HnVbjK+97nDPfwkOg/Plv0XRYuA+e02sqVee0F/KFdLtpY
Hc0/rGw2tc2wkqYF7bpdsva/cdWgp8P+nq+6RuNfR0lSi3sG+U18Sny1QmK3uKPJ
8vrgIzIl0fGRMt+DpT3p08zmcSsb6v21CTSm/M/xqDIzgGsnPxbVrGaPLDquzHTI
Mk53hz1HYAJLBb0v/uuOWDIkgt12tkNkMfZoBV6scCrZyqVj0isQNkWf3xvnc2Az
kn5vABlq6yzkEA/cjCjbJQF43edWf4S+rNdy/rS0hA0COm/OWPl9b1GBO2fbQzv9
G1YV/o+xtZ/unXVyUXM9vHDA7vVInIqcBEDZexRc3uUXd9AotDFlr0zaRhihTIeT
XGRrxEyT9B6CFdXeOy8J826nu7eedFox3ntQvxSQIffRWBlWAToDAZkpgAX7WqtZ
l2QCRfHxBRsT+Wzd5pwPgSjS6GNgN7+UVa3IuQdI90OevKg/IEVXui/SJYD6yQeD
Xmzn0jJ5YBYFwUICzqxTS1eI3BhsgED0b/RriRfBZ28gW6nh9JdOA3wSBD44FyxS
Qtypatl93CuMthc9WcJS4rSxEIQeQg5CJzExJNt7Ib8vSVhMTenfV5SBlKulx3hX
QkBT4kUIoYyL1aslinSt1ngy2llJZM4FCgHipuXVubGFtnJlg4sKg3lq63ewTsX/
BaNbaq1uA+61Zn3KMR3FL4s+7qIscMAQR0i4VFT2XIDEk8Brj2YpXeRCsZa77Fmg
4I+8MaoGMVJ1tXxo/JKS1b4TPQoPz/4SCQy801mGuCD74KdBQJdW0n0TE93eiL1b
c37NXf1+f+iQ5rc1tnMZ2it9O5jPwTs9xfS5ld2jxSG2m6roGada8n+ERzSpbrjn
ehCjg696dZlgCTTyWpnxJN0nTTvFpva1MuAg1qrJbRd4i2v7gr61i2UHw0fgw4+s
/NO5AiF0i8/Mq4UrPPFaeNzFC2v7Z4+hs9pvfOe3PHWTkS9pgZ+XvchlAET4ifqo
dpdVtfOFuu0yZo6TXG0B9a/fwPImfXPznm/2pPCnzMOyv3+4eFD7J5tgo6z2EH+Q
HOEpqieoEynh3oqBNqJ9DvcrwbBJUdRwQLniSJIxiaCcb0aCEj3PB7kX7l+ZyBhb
PYhHxi0Q7TXN5ccEdXTZZHAPCB/ftvfBIr2R7vYcyo5HaRgoNHNLAPtzbUupr/zP
1/LxLDI/DWCbOSWxw9e4uvO7uyfE2oIIw4sPQM78OOqxw+uOR+mJGD/t6/W1J7Fu
PQJYsF8ipakYckOVLEj8myKnwqFwEs6715MGTII8oQxO0RcA5ybThHi/SJKIVXBW
3RKcgwKxkp2Ynd0R76pF6d8BIU+ngmrtVQHiP1aSfz7WRS8ADuKNZIfXf+bhpWTk
RLzpbrt8H8yAcDnV3+AYe8yAc1FjTxvmYcW8yicTZ8h5cZRj5ZcLznca0TPVL+hJ
b+RoyKZ9NRag/VncbnESuaXon0hTV7yZRvFYHwqwcuenkTy5EwgmC0FC6yMYUxb8
i7+oNJQ6fG8s/3BN/7RjNWe3PmfRGGAgc6pNj2635//hlibBj1wRyzEB7I00PlRr
s5SUwg5JxyWh2Heou/CsxAK2TJTdfIY5MkXuCVTgrBNXR5D8o0fJWvoiFPcp3rg0
yVFGimwI3pjd8dNCVmEkQyU5GUhL6CoFphgP62Kh1Nh6sL9qnkIgfhYyPoxSRazS
uSbqM997HzAbwD8RsRgqC0Ewafe/OuQL+w7JV1amuvoCJzuiWb275MNAyy+pSaea
h4oF2jZ5w8Rg16DfvDzWJyDpHERa2/MbNyFjWJfWNqW7Q2hJD4Ck40uY1n8HALIn
9sYsDNHDlWBE00EnQXn8uyIQ52u3+gWwfxEazGT5rSNalIzDZeRjI5tCin6OUidx
kvlvZGLPxnCOBMGPNN72PK3NSfjohLdbPwaaJdfaca6u2f0eKhegIGjGRY+tlwkq
BUbRE446llqxlMWXFaGunbjOPmvQEvIIJATzon2Jo/TKA8LwaSSc6z8kUUDZcfOQ
NBcpbEJQenA0/bKLF7yJYbyDwyT9TnReTf5hG/WVJby56F8p9x/A2z1NYjQKqhEQ
7dBwSuiyGhQ6AKapQcp6K8PiV7r1GKd/FHO20diqGb/8OYRLdXydsP4bWM6FQB/e
LB9iVg33N5GSTYZZVsGCJRITttC3XlbAnI9ygNJiKzVjJS6ih0vrCkxcJMhWC+WK
fWyivao3yzQN1Fs80gn2jR7T+4j5zEOoHBaZFsjApzmBadRsCbtOEmlNz2K0juT2
I96aLXX1MdN4HsFam+xF+Y4JG1N2UfBMjCceskQWSBuBa5dD+PF4nhIEyYB9kmjQ
g0rrTb92yz870R8fIwUjWnab0Ule/BDSqTPAeL26gJ7Y1KFq/8szPkoRIzPotPzh
9Xmk2qRktXdfxb1u/YNNQWD2gar4Rl4aFtCR02+XhWm388n8HJyOprwRgL4v9fX7
0XCNeaz2ry19ERrRACf7n9OGu/EwIm98JwuE8Nd+h4gQeIkCHXe8vAPM48u1of1t
tR93Kqe0H0P3ENORAf8o9qUlX0kWkZJq73fRblrhGFdYrmTk9BGcy8VzloCnTTfJ
5lRMYQmi2+9ndNL56fq8qeaxb44VsfCKBNnnzLrJFVzk1tlYedi03oWZ2I4WvgwS
eh5vEapI3b/1oK6Wa43JY95dtsq/M1CEzPL2aKmk+q6V6qykvaSFe1rB64nG096S
viBAIdCPoZsCsUl9dHIBxL9oZzIzyQnFMrH7kUJFkvt1DfPbjTQtKZYW7B4w/uT7
I3hO2xoFzNz9JbWYwnGQ9b3CgSLmeuFCgKzRwHzRC9OLNm95Q76nFKEDCHlwCIJ7
RR41wL7tfWWweqyp4djKx174pFXcpQquY8FqCteIIAOQSyea6nkHmkM83MJve0jJ
m1C7CVvYvlXUgoHbaPamhARJlCdvxADCARJ5AVHV+rDiCTsFOl29Yrwo1z9QvLG9
/cqGJ638JJLUrb14snyJIhM5TOMQyJDR/jMonA9RSBZfidFzH0ejpquZdJVCOpOJ
9T01ksp9zakvTA/wrMlShCLzcgHXzix1oZ5uG3Ryml+mvB9BK+tH3RMLMFmQBTQf
YeR8juPlyt2MW/dwu1NFPGizMyeyfZt5QSX4GJe3SY4L0tqgblvZ5KuZpC9QvYZt
2GSqe+VL8IV4wev/B5mBFmXAprmwrkBtWeHIPhrQe5E3Pe5/HuAIEbiIFcmpasi0
ORVlkecZewotvjJShjPnlkBKXu3DdlHr/HEAkTJAqeBYDuMeMqTjgey4NdU+OJei
gbzdchEa/XgfQvXhIW/fxpqJFZheZoaMZv9YbxVnHhshZCqWivaLKJ2ysEiIdOoX
Q8cGWlxo4F583Mvwtro+xvsV/wQSprQ78WvxZG6o5aBNgnwQw8HjTvNeMUKBl0JJ
zCP0F0MU/8Bft1qdvN4+vj2ndwcUfeN07zMMs59H3fcvgbWPGWbiFa4R9DKvqCnq
hIN7+n/UD7taGBXvdVT2lqOdeq72yPAqwfYYjrK8roG8Jdl+zHqfHxrbWUzXe5vD
uNoAFXaUu+ydZRIhpA/mB8oGyMqyq0T9vIT0gSgTBeSxS4NYiqQLKWiuMMeiBkd/
jp235BwoD8yX9gecegAuMAG5//U0FNT1OncEuWTJFMZ1kInRoL3ss0hJ0UXHeESp
JFgHIJaNZ+H15+myLUXN/I2GBKFye92s8KGw2+LLGFBmHrXh0SKyHeai+cCNJw38
u2dknU6EUau20neZbyt9o05J3t/NBTnYu4xIkk9PR1JIBr9AlgPU314+DZAjcTOq
evZrU1bE0/f+IcoSwY8Ijm3oLceyacfGpVdcPLU2dzY06fj+PnSXwIMa/v8OlGL5
2bxSdl9WJBapIkt1UW5keupnsosyq0LDMjEjXFYk20VWmyfhippL/7abgIi+0g3n
Zr852fa9Pu3g7H+f+sYLicLXXHnfugsGQiYn6upnI1sZe8BjfhslcjPVVygK7U9G
/XGsaidakbqc2OsBySEMZcJ0SD9Kz9h6GMkmzJK3KS1gaOJEV1uoRp5m/7gBh9BA
ePOWMeJnUwtCW9Waxi6wCttkAy8isXRg+a3wpzTszdH2VFR8zcgH6OuRn1ZIvV4C
SEzrQu6snHy5XRNLR+TalUOiDKAFWPnilf6PXA1FlLPmotUUQqziyJqYzY0sHzAL
zqJfOxEGIJtUi3M5pIRDMa980UgnNgVR0uM/qLkrfSHUJO09tE2k8fYRz5JNuObw
5GMF0qAaEt0bIe9hi+gsavy8rtM1JeLWJyMtqMmySJ5JkKTSCk8ZSWUgPNL4LpiT
yArTHUSTv+etVdP0ox+QeP7l/Of9m3SnChZTikx/kgCaFEI9mb+IYFEoRx7LX9zT
8b4HR84jBVKCO/6hU5OnlP4XoXkFkUmd2Oo8RNMmQpfwsxA0XO1zQJyWcAU1J3+S
ukGTKcWT3kfk/VhbFyN+1vEAaCVw5wYUQ8tNo5hSX/U1EWaNbIt0ZkSWhER7PXb7
Iuwc7PzfadLOcVNGGYYLCzqAyrzildhOyqQsQMBFYXZOjJfeaw89x8n4Q1KvPi8M
xZuAexYUmd8jN7IgzzwMsVmcgDN88K74SdgQ0+K0aOap8l/gfT/1fK4giaOM6Xrr
+vrp3s9X8k020s4DjBPNSPcjSlJr2RBojKaLJ2ufyXLNkk8yjuTxA2OtpxP4pBzq
SgbnJFQXl7kouHRzUTIkbDdWbCVubNno00k03PHytV3cgD1liF8TpFrOsawo/IXI
3Llw3IW2xyHYHZOHlrUB75Cl3hjXNUKq/Pf9jteHXEeRgmcri2NOuGgw7pTRtmA9
AQ8vJFdk6qYBPMsXrqhK9kSYAWPKQAMbYPjJ2/2KcijWcjkqmKXf24jJExjJU5dC
Dshm1NvOuLsJXP0bRrN7GtGZA3/bwr0Qnpgs8U2aCW0OyDZwmXb8HtQ5CsNmcKHl
67JUqjjimh+38RtEVh/kI4uIz+VjcCcV/x/Tn0wGhiSM0efwJAxYM4cwh8rdUhxD
6HlL9uv1VrzTWSQ+kacTf0L5JNKbLD0TOlOZDggvQsKdMYpf4NtBR+nMgPUtby5A
PJsxcrK/9D2/ky80BaE/NXfvH3YDK4CE6bBLR9750b4Q9B0axJpfujHlO5vVvHRq
sT3UFixVarz8mtW7nTjd7Xzp/v8/zLm1kGcBHD1LtapRHhJBOqYyOp3QUCRsj5v1
CT98xEJtjbjD4WPU2RXvmRxZZG1JAwY903XdhFYdf/Auxm5tedxsDi+X2OMWXnD4
m4Snn96Z1o/lXTPvvHM1xsL9/7TGa8JXfHA+IKnZL3bqYu9VCgNEqU6TfLnsJbvd
GWSUKS4Z/xJOs8jfiagKejMzWrF4W5mUPbWzPYnhZNIKTE53RVFOG5YtmSHi10BE
KdFbCpI/4lF5gWc1gO3UZYNd+grhrQufC45I7u9WFJguDcHvpkVfbapkkFbU0bpE
XdAbJ91m5XU48qGblm/tKndXhGopGu3T8Jw5yjPUjDMoB4LywDCX1gksKu3J20el
XOF3SrYh3oUY6d06aC3ogi+QdhgZ1KZ4D/AHRjeMP0ybe3GGvBWPd7Rc056HEgMd
KT0o8l2vUuUjUVBbFU7lIPMFiyZp/GR0kdnMEGGZXKA6016BMPg0VjpC6fh+cP0M
P6SUbxygWOvaSmbTt0uJjK9+4Qm1zCEX7gUvTbHg4Zukp1X4+fXhYHqAspEVgYm9
KImRQpLjWSHdWcamDMNRlBqw1uOjF8UtXhYm7ujicTTJHWZEx6WMvZV4Js7tl+75
bRxTArQUk4ddEEO2zLaF6Ov5qVRV+vO3SLZ6MO6+FVQkbUrFlqBHiarPKKEFEZoo
Oyx7hf7qJGqqHXuEawsIHvpQmjGJAJ27LVC6Paawge87iZt1NUTmiQXX4URH6vcr
eoYsdlJsMQ6B7/0wYoWyHVvLRBm9degfrxr9WBbIOtjQcFUQFlja+5r75UGN8WGA
78T8FWWR7bvdHtW3I6lWLYSQMc6VgF6m38WJUhr9FIkVpU2HZ+gvnSuHq6qESrTs
U1KRIfACmjcGhsz1j4BYDo0KvsHAWTvmpCmQuzCbHJtxpCQz7hSf2gi2oSqOMECI
jDJdAbclufSQoA1L9oUEJycS2yrnmbvIkBmjhSbGpz4cjHgV6YEmJLhyip2Iuzk1
yX8EuQySRrgP7QFmBbckpjtATy+EaQkHRcK62Yl7rh+WfGITwl22SQhlcT7tI6J3
NvkEZLvKyVwOhG3tg41aPMBo6R+hDYbwT+qAsglNzIh6SJxdB5ATwNEglhlzrNaz
4MelwfFhFzxfZbVavN6/AEWivf1wCe60/wz2xFQYwSoMR66RsMoy+57IJLGQ+8FN
/IYRUktfn9IodCmR4Batif6rZO8wdNcdGxCTVSJTCyPgi2hB5vW3nwWeA8gNPYty
g8ZttUKhp5fAIwKcqAIYbd3jVlb3+nY9aRI9edVk4ougq7ScSDReiHYvG8dw0J9Q
EKf+5fEKb9vsaqCGPMUOmOeyRiU7dYE+lx8TVSM+A7KxPZgTu3Wx0xmYmzsp9X+I
tfCijZuXClB3NJ4HATmcTGoNI6X5gQeU6IrtIWtpq+LO4ojU/NX1S4nvuxq/dn+y
rBCEvq+a3+KFc2rifSIpI708/8+1G1+iGN/9gNO1eVW7/Dm6Ga8TRpHBSa9ooDRG
VMXsx/QH/fGUoPz9yZPA0ewe6yCfzdzXG9LJNGJZsvAKPcc4MgL6MljDFvBmzrUB
MqCFhJMnnzhQduxpagzLzrMBOvjbs9ToFfR7PbcJHiovz6Jhe4SDqezYM/eVa1hG
CuJpY6QRdG6efhdnp/h0IBtZ8tdE4BSdX81UUacNBTubbPzjhOAZ7qkdwyf3LqxD
/9dFhihjR2hWc9NpoJCVLgEvSCPxWxtJjaDJDM50csBekrEdvWyaQX6c82/VOcPn
Rz7Tg8d8I4ZR2nHQfnDcgL1/XryjBV4FZ4BQ4L+NYLhAWs6DjclhdqueZMzuGBzv
+yHFwBFef0QaiDFhBX7GHmgRBZywF9/FwrbDzbX/bDQdIKTTTuLcRPyDS+3wZl7L
GC7P0zzp45AFRToy/iSeEvZvLc2ITC00wazX3YexeyArjtJ7Jc4DqlHofQDyBOpx
ASvQCdOozxwQ8D4BGaOz8i4RQOrcI/6IYOu3XTPpW5VLoe+PqMJyPpfNqMC80DFc
g3r74vNS//Q9L3owUsoJeSNN6Nb+Ul6RNFYj5r2O+NhbF1nuvA2D+D7JK/jnwtsQ
EHYLezKkvBmYmpgjMezU8jJkuV9HNjieqMR6gHu4TgVRXb4wRMtiJrd52dbpYvHe
uEglEGtP0Z3OyKZJe4oqz6Ds2Js62S6h04zVG3aQFtsASvFPtFVZ+6bnF6m2nMKL
36skrKlxKdu5R5rOeA1vHtGWlHMr86p4aI3QnR3sYTY9faS/w1EhXcOXuEWGmbhI
HZDiM7jN/iPN70xR65XUAFj3Il/Thy0aP0a4UrC71VIuNdfiXzZK2H4Y1KY88tEB
vF8zTHl6pltNrOQn2mUAPnpHepktQl0LgkbeNokjirHZJStWUBHWSkUUIZW8oPUB
cKlwuUQp5GMNbVZI0TTOZCGjmiIcW0MA/AStpkpzT5BzJm5MFESDb8fbocTPQ//Z
qCqfiWXMqB9PYiQsgjoT4oTFZdRVigpKZXkjsqjntDugq5JBe/Mrzed0zjKx1gOz
wAcpgQ4Hw1ljgoRbE9NYZv2fKRJOQDew4kY/JmdWJzfhb5H2G0BKzne90jt+Tt+D
nAbjaAgu6gyx9LQhY1cMfqq2Oel/IMX/N3+5JUxxz1MbXZPvUG+asGhmOZmgZG6o
q5aTuCPqsJ6AQgjxT6BmdnMz3Pnyl+xYuT5rkysq5uCYIN7AjsXx4gI0Is4hNaBD
mZZh42iEApDRwk0rAC+t6MqnlWCKAjQ+5dFskqDHowupk3khdMu2DcrzD8BlwL0q
yEGG48aTWQ3E6FnMlGgqAZ0KEYpAxUNWznNNuYE7vA+j8JZVaAuB0O+PzWU/DC9n
W3tpn8jKUO0RV8HVWoi1+GP0K8mCGzA6Xs1ebnIz7HqlsVmDp/DufSkLw7nbpZpL
AGwNM5VN1P4BOql6c2pMfWL5nD/nDOQb3sldCX8gFdUqIGPi4iwyfV+02vhWbddo
f/RxXTRVNgGjC02AWQRiFl597IMtIAksh0xceigTa2/kIOX/gipSDQBQADJLo/dP
BvZ0lVpXdr2kc4eJ7ELek4w3rVPguiy+ys6qZINNNnhKoCgdeEW/yxaW2Xh7UTuZ
zcJ5kq1wKnAdaKFYnHHAR3MuQ7nfs2oeF6MjBNuWX1BM9L9fPubbEh8m6j8nCHJT
ePq8E4RxMt5Zho0riag8JBCd8riMm78te7tYAyU+VvW1CRiXuJmwCxwbs9YDMvB6
b/YoYMEk6ng2qz4QUmOVBsqvvc01TXFBoZCJ2WWEJLF+gJbU0ax6yvf0lOgBS03+
y+UwV6Ak0kqe+Cqu8fBgQ9tITCvG/8/kx/9nvugeOEK8fUtgOw2Mx2fbWbx2oDnM
2tZfkJ5S3+j1/0fCjPjT755qWN/C4Fslpp8kcpTTaWSrJ+Yi/tYv3/wer/ZJt9kT
O58f/Qu8J7R9Kv4tgyazRPxREA65vh9bsWSAkE0T2fdd+QJ7dkPUdcrF7XADQSlw
ngwnnTp/hZS2XKkOFLEvu67JDlTZMHv86RIYs5f5nSI6sqf4E999w3kQTRiNSt6P
Nkq2i0bVADc6dL5VveyY0VbGC1AYHijUkqIxEeWIoKkfXw0iswtOWauIEdpr8izP
nqXjGQ+qboXNDcTtvVXO35X9MJxFQnkLAowhH/CazVpLjegkR5CpkV0gD58SWqIi
bKJ22ACaUuKvSUP/Lu42cw/Q5fxlMS4bd7pBS496ECXLV1JDlb/hJCoCGgaRuvrP
AU2DBLY4BcHndUiX3SVPtrnlvSMT6Bdn+El+3NYwfsUdPHgtD0Zd2qHb9b9LA4fr
dsiVi5GceRwITWXLQdURKrVZKz75rIO4Dil/UzzqS3t1Wa0qyEbLka//RRPLQwPF
aBUJP3NFA8KvF/yXrOBWs3tmKd8l8SpMZmLHx1kf8oEE+UCqqR8KWV/13Ya85p6U
9mcfCNqsGJ24OOeLlMmZ5YPTJG20RqC2yaqCdX1wZx16TkyjIWf8t/Woug/MPmcq
dp6DE1mtdhKzmUH+hq7ySxRfbs4N4pX/QbsaLws233MKdL7enRN/jbPjQxamN6iX
azibQoePWu9UiZ08UnMC7F+ECATcoSy6Y7ch6vtfAHHUzenmktsoNwB8akbjUs81
0JBXjBqIg+I2mXtWaHG/uIcZdQa9hX3xwd0QGDImPoFP2iz97BM6JfH09o/ovwdZ
dK6Oy0XVwISgviLnAMEQQ53h2ukjNtgpc2aLGyFdRgQHYYFwmpAbh9jTAUn2ECAG
zHefnX4ZsPpBRyfG0dLVXPK8eZl64dVSIYFIZpQQNcMNSMToxycTDlSkmi9DEGkJ
7470aOgtMTayxifJ/ViJQxaTlOn4MT2pcqsMTbwbqTQH4TATe/TIQaKnZI3Z7b0r
TLYQkZJzrxaclObVvxgdejP0SKQUtNRU12gGx4xRi2ktrhRJ9N1LPWS4TTtDGAuy
FYfaZ3gVFj1gnp0FkJOtKYuvjgReRKGq/1hYItrr7HWx4cbJwmoUgfO2aomlxVCR
bHF/wCQaSJhI1h+Qvu+X1BsnGO7c2ibkLVBTIM/MnU/DgiI//0jQVLSazac5ur5U
4NaGBYbIfxXeXaOnVTt2cgh9qX68cdi4Hh+NSsn8RtowiK0/xGf5NzUCQ+aNI20+
PiNkzM+4QXiSiyflYsqnSihOPZb7P0ZCyhFEJC0LfvRsAqpyzJhlIOPIwlQ8E6ZB
es26x9ClKpi9fEhlSPGxK1aNoFDJBpxZN18kGpuF/3Kff2DqZentOMxsETt/xcxC
3CVaOrIHr+w0B71j/tEQpkbWLp1FkY1rHyPv8uayop8nbJrLeOxNtI64vsPBSplM
OT/Fuc/hVeUMxeLmzYEC7hJt3WNfT4ZY7l+Z0fijC+f4j2Y3/05fXIxVwnjSG+XO
GE14HH7aANmyotohujAAu4ZGa3qdSudCMzmFunfLktNz9R4tCy+q+gyjwt3M4clQ
foWSnbD2WdFrmF+iNbD1AJZqOfhuctaHJ2haL8GKpFegaw7qijD0rumK/26HNuBA
s6tnxUaiw2V3EYzdhhkccIB8M1zbzCw617RUZfPKaoQuhOUQru3OX6huQ4zKhajm
CZYLvsQ8SInHQEYc2TRYLDmae407rBa/rJO2B/eDif9mMP1JE2d8mvJxnsYAOwc/
7q6MmZoFc+Bd0HFRoN1joKu90b0i3VKJy/rWZOwt2qSLWU93GKjr0wtxBuaJv4dW
kaGjwmimNVON1aP58DKZKx+SX0SiIxvdZyERfrWEX5wuKgvNzHmvlIvS/MjGUsuI
frOfD//KGzRh+U8RzjOP4B7L+WnLR8QnvHqCg0XxKPIQ6FoEA6m+vMun7+AkItDe
QBFKQW0FwdMnSJi6KZ5ATiIL+PTcX71I0FkKkZ6NdM86Hiu60PYxpdcm9F0bhkv8
K6IaRtmdMjz0loZ+o2kxvgbEGdgsHMLyYClQljSOFK+6Bg8AAOCNXLx3Y2pQDMqJ
PI45h06yqQDQZZJvvHjaeCuSSrRxQku0iqmWbL5jG5NmPk1OkUeB8FFQqrHFQUeO
WyxIcRpoVEzHGTkkISiGlShpkAqc8zRB3egJSW9dSJS2SBUMH+3CDQj63dqgrsQM
3LbkLfVIHw1BAUbb0hSJTRE7V6nu6ZjBHS4R1ZeUByGJIg+G8T9/0H+buLajLtGx
h3SoKfmsQYJl+rdcc9ns23Utg8b8kZbQaIp3+6xTzv7K6/BUHrv4el/gq+Wszte+
9wj00y9zML1zuDRbJUU5oISpyD5a3toeSKuqzKi5Te4qj+gL95LvHSgYc6k14WCv
RSFwKjcRhT4vZC0wy51EOfXmGe4lTGgoU64Pc+3eJZBJ8uKs3nLbl5I5GxJjKQWa
VhsXTQy/6pcJPU+mJLe5fSpEvw9P8/USbBwiWHE7HkY8lh8i4wlgLaCJCMBNFvtt
klFip1CMPZWuD63RUiZYF741DPlbOUsAmEkj6Zi+fWTtlXjl5nwiUXpWzydwPgKB
tbOo+SQ7N+P1uNpXPIG2dhmK4dEWAJXEub7I6flzWS7RMQkyAEEBj1/ntg6udTVX
KuKxALmwyjQUcbzK/Wy+AwtwIMRke0DUfTTD92EPK2Kw1gz/qU1KgUW+HArc6HQA
BM67hUW8koj9lD7IxcKys+aqS3w5f8OEJQT9AdbsY6F7xVNAGIxuRNrex3oVWrmu
6Ax37binzN3IVOrbiOVmQBc8e5emwXu8+TuPmB/tdq/lLaqGysxf9tP7Q6driKjI
9xFpZdCrfcZgoRbn0zEAIAmOjrSzwS2SBEyf0hEglkSFWWFddTWB3OPBzBszKn8t
8MovVlF9XaGjZOpWt+yjn7pcTaXF32wPYUOOrbKflBH82U7Tfx+Tf9X4cyYZ6LQ/
ji4R/B7x4pGDHaDLLr3BOlWY4K0/nL5gQtOx3FtIb6TXxDILX5eTu9+mtE7TgIZr
snq0Xaxs6ujYNU0UllXopYIR4DZKznPmwYyTasp86AWNVwBHTaiXtvFEz/WXiB4m
MB694TAqg17zAt4yXQ9OK3crHxKwEhPxpUxqLdSqh2KWO+kuUyhwl9JyCCZ92lsP
QZr6AgPaf8VJ3LCPdefcKJ+ZCzymQq47LQ8ZHheAj2iJCxRuNQvN/YNzF+0t//t2
uHRab/zy6cf6LxE6u3rt19zB/h7hubDKpOzJVkAnrNJTllyWUIUzeVbaBiHdy54c
lvZNkjh7c300LtYu9dg9uPLmYrkHjwrx2Qe4YWR+Y1jxrJjk9/PFnQXvBujLxpG2
RrYXowymxpVeAGyHrUKdIZki9/Cjz2ALY4Foktu7zyfkjKroSrzuwq+7vJYHtv4x
W0h7srihv8Yd23n/mqB+qYdP95ZtcpsAzCjSRnP9BPfVkUd96fkm38JvHcgpIs43
hXFS1yP7s6aTlqBhW8rSoGIp+ZbSc0c5COL8G4xLZp07pFf9HnKt4+uMGFJ69vbK
5Jan20zhowWeH1MOa8qLiCIj7akkmOQMCcwfZQkRrvcL+0pidFl1feHApvoMVuXx
vvtKWexeigKDJX8jmt/sH3WFHv1fBdTsjoa8g8ujmstoLzCMNg2amEr0bduQ6g2r
Qlh0OIhMuzEjGFQpu73/4lzmjkT8W9BCk3ZrW2BTmmDbHNL2zPgqVS0uouRZoTuh
s6MSpYdYdqO7bCuzqOYSA8eUpieiYKDRqr9wpPP75mbJoCS0xiwpvX3Z1IIdrUd9
GuxrAy+ySAe+hu6UPAde3dDh8htlmtcQROyFemFzmUvJ5o4EaPywp0F943/SiarM
xoaUqgHF5j9VNSWNiNFItzIV+h8t6SWA7yS1tqQ494dhiX4PkHLQjoe8sC/RmrgT
8TH5uYqg+pvD7tdv+bY36BdjMBLL9ulXvwpwpv2/M+IxIuKNk8LHaA0BteKk9bxK
FikoRFFxbnsgjCaOr/pVgvoj/LUW32t1IobyQoGO9bCXXXxiwFDMFs7kmfOAKv4X
ybY8v9oO1hYtQoM2m5vKZX/MsiXDfWRyb4rkRrr9yPayWyHk3EXp4f8zhfm/GOtJ
yx8HLhEKBFc4Xe1PhHsVaH8z7b9cwpkOU+caPNm7frO3gwMfUgKTE4wTO6MtI0uT
39Su9cbcNNlQvSGKvetPWiilWVoXiA85X/HvKGSBCEK8MsEC0CZSUukhb0JCOktH
ffTdNQ8Vv8IMt/GzLRXG38BNRwCCalOVhWWDXAlHBi4tcYKh4tmrFxdbMKpvln+2
l/CWkKjYD6aw7d6A4lUIToBaSGCUbuIMnl4rCu5kvRD62aI0g9kcpY2gcVZiYKqy
/hX2B8arC+8Xuugu8hj1C2aHTQXfLavZY6Fs9t+69aqvTdARF09vLbeQxzg30ZVj
uNW8D0gV06BYe8iBeT7NBmIaDIN5Z//+Rhp4xFQVGuF24N3MqvFGthaBYbaXcaqJ
HcoQeAbSrLz9fwuewlCHXf3/qUKA1jwElqlnzZ7VNF4v8vXUCeRRiMwrxrznpR8E
aSkZVw/tnVaX6gTMoiN068RsYVS/La4pwA47+7sUuNo4l5CzqO+I2gHke15NY7o+
qyHOtXszrZeXSIB8i8KL2zyzyn5CWFZnIvx3PH9Xeg9dx0430LCNV3dDEUZRetqr
OgzNqPT7neQFMCl+4UZ5W06RgdVM1Hh8L4bZg6W8GwRY2euiQRdwDn3GM7usuXCA
W4cEzNRe8uDh4iZ7WT9CHE63bWSyxj0XXMPYHZDpTfGdzSlU+R1AcyhUnI0kcvXc
AhTGbxJDxzsygP6YT/nPqZM/OfbEDrnPQ1VhYEvdL9wf3xwpnvZMGpJbQAk16b5G
srjJrYju/SRNNRz17eOT2b28YL002RZj/y2hXnmcA+rGRvlM8IWI8k+RdLgmCpzF
Z0ah/qyj45nCLRXXyfoZsbOpmLChLJcm2C8Dc65/fYVGaAEd0FkxAzc/aukgmy7k
cVnBbga4u3J2/t/+hrY7KFESMq0KpoeiwYO3K4nMs4uqyfbaqd1FllLPGOlmdnrV
c7sBfkaQ6b4L7qv47HzxRHwXFAgTdESrqJwkjTwcsoBLtAxpxln1r66lB+v3beqM
Qe7XdRXdMTglkTpS+hxVwEUgp5Sqa9/7kLZtOfETQNpKlRIW1NuU7Ysd199JAUEl
ZtSGmkojf3PsmITTJjy9vGEDaW/WmeE/myoj91F0a/Eik1xRVR79ygezM3rcKVpk
Q8swXbXvyBTbDbp2Tw+y1AtCs9HZ64QQ8TmYme3ESY8e+l23GEbkIdg+A9+VLVhV
EHLsmKK04Fh+EV1umRjzasJpQ52XRsP8rsekv1LpeQRIyEb/+Rq1axMRw6ifkCge
NDrcHo16rAYRGuzC9muAf+Dh9C2rHyJnjQ29ej5QOLbTYfBlAQiZ0rahX4c4noDr
vlUmnH8cvcKI9tfe8tgKoFWrkJBGZQtkr/Cqf1n3m6P1Sr2lZZcVPwth2hzqcWvF
45qgKknxJo6vYWLgm7PeSoCXPvb4O+uBXkBTURRDU2lXBspHjWv54zGW0Yq9dGRS
lWZKWVkpE1VXMbFd+kudUMcLw1u8vhnJFMziF46zYfydqoQ1fknRY84iTU8gTYlQ
U23OKRnlX07jsjnexRjo5T2kqxyQ5fB0rKsoFSV1I725mkq1dygdJecdZChh4V4B
yzgPPZZ3R8XSNel+JZ5846XdOx5GmLREXbeSSeZ6MCMefMDZqA0IGU3eIT3J1dCJ
Povvvo+3I2AvJ/pmabaop+q+a2s473jOvcOSk2+T0jUp+YjkJtKWWn77diKG+ozi
xl1eLy7KChpbiQRw1iqi3yI3gxJ+uqXZa46/c6V0zaffiINOgnxCxNvpJLKjctUp
0PYvABvLnPcuXlGHXr/W0TZ2ZRm7xr8/lKGilWqaG8X28rmWiZwZJ6mMXdAejFae
pxhJBQZsFd3poopxPkvUX/0AfUloVSoxGnvGCF3Sbxw6N9UY/gdZlaWcIYrK3IW/
bMYMeouEUhk7H3b+ScxyBTKdEKUHT0Qa2020vCGZkP7Rc7UNvIEb4Qr5JVekKgmA
z9qKCsBelC275Kg6nS1FqCRSJuNMUFDLaOFWzi1myH/GZK+rGTztZNCIJhf/BxLk
uQhG9nzaQAm+LEcWP88s2JS1XvFNpxj77BnJtPYp87gxfGQAfo2BJDtlw9wt7pRz
aCcGaXmZF/h6ivXN5+H4iBNsAfD6dS4xVs6mAip9gwK2oCtixhP2LJyuTwx1CW9l
HY49IT0KQ6sQArkzTKryl8P3G4m136R/E6YKYIvIo8lLVqUo+7QMe1nHAjA95nIq
YUIj4l+WebgB2XNnLjaIMFtYkvN5XLnwcmIExoy6z7arwf8Nt2/QjCeIskNKSJcY
JMYVGTOkrdCLVuVMxaD8XKJYBsUn0C+M4qtzogX1HAIGRwoyn9VmawZkVbH+ld49
EoEG/CrauDN1m+QSjJ8cINB2brC1kjBBtJUemL7hhItvx9J8fRDGvbEI2WRfxRiN
9BvvK782sVt07kRUlXPLLFCCjCb3gQpm3lIurdfQZ3obbjY9vaSgm9YVPoD+W4Qo
+bM0qY6mtDFAsexEWwzU9jEOp7kz9AnR6jXdc4e4WoZuOEK7NhdDp6vTxneOoAGx
UoJ2irhMt114sAcxJu3F4d2/RZgWRi81krhVUsE/eo/x52h61yIGL8L+LxEHdEZR
T8qUYrmwWzTGjOhUTFsPNih6B85mkUsGtRchsylriiZDRn4GUWwUnKy+PxRZ1XJe
sBYWTAtIIru/j5sMwRgQEbVbqvPhpgF0crtzwsyF+hfRV6qumluK8gDcA4V1wHZv
uFMeK3k7LdAozmwz+hh+t79CqUaPp0Ufj+hijoipkCuxL/eoC5T6n6xkCWtqYw/G
w20hUuxvmFW+bYRuSbjNOx8oe9ecuGUAdLYduo/79jMOQXTB3MbBtr1y6e91KCay
0IbQseQfoZLzk6ljhKJQ5bapPEjFiOxJqr7lgqhxiCVX3zJOkjvGIu+EfmLkWdcm
nmDOFXZBrMwOrjCEWaZ/UjaYNi8sTr7Hi0m3wLEI5ztzwprafH6anEakfaBpcSGX
GWOmEcuz+5MeW9NpJTGENlneDoRkcVx7CbtnX2uQOoho7I3dELn9PRRy942SbLjU
Vz84v/olq8dpiUdxELH49ikLSD6bfKH35eJz870QoYueXTOw+FCMxJYpqjccEt6/
+f9sgt1XYkWQpV4vZYWkPo5a6OFu450AVBYQdnnh5pEZOLXjfx6JliME86KCW1dk
V1nqcTUPi0SpA5vF28FLHlfVM4ZQ+2+IlwyAKzYa4mxqrF4mfZ8HTwbbPttIj9Ly
RbyyN5gNiUNIlcNBYce3G9uKk+3NNOGjh5hI1av1pMyFmMvKbuh27qmeu6pv7qii
8Gdto6E9aIc1D0G9Q5lV8yabvfrFHGZhqBq9ZmppCgeAXemf+4Ani62qi2caA5kj
vBkcM3uw81ikicL1I9AL62QTLJYAia0yw4P1+MNqMXYRK1k10Y4FQBRjGPkO1ARY
yNo0FS2vij7YR8iaTiorzfM9FJu7/6+ITWG5Fsc7C8kAnTEuodn700/I5xYiKGRf
ujqMOkuqgpNz+2LKhESdglzqPCgrWk/162Xjm/q9URrbSc6aTz9zY5/IpNesKZR0
k0s4YBB7IPJfcpzVOajUVoq28gfZkxeNRbX6tHnHy2pBhBtSPVFHpcpZ8rprdIK2
2MFOFmNTe2rigPhteAKd5uhsghHBrAY35YF5QnJM1Ls++xZkwHhw2MUIDauCMmmK
gdm46A12I04QI/p6aJTTkJsKiCWrjOzxhMv8qx5YhOvbQE9le+c1HY2S6KIw5/DL
HtwLEuPtXFPFLOSXbYiucYENpSETmxcRRQ3qTmaFUBMfaLHPAI9hwGxO1YvhLHw+
oTH2EYq8soYO66DoaahuVttOsNhmOWF241pesImh3RxlWKB8ENDL7ggEiAFEerwQ
UKdYzOaUgNTKYWTHSaqtGJeQ0b46/oVCl8KJNPcnpLhWcq7B1TGGgZXqI6bhs38k
r4atK/MIAjsIHnJTJxxxgk6ElEWJQW5Ir6wcRZZFC//nLsZgnHWHbFJXl/G4Jt1m
j2yHWDPObLu5FLbFTE/ikKPHn66I+EyLv0MpUGXMwGIKbeLtbno3FC3Flzyn8gfD
xwWI9zXTV9VLmww5SweAUBJ6c5HiswH4Dpr05kFDMpm8f6bbqv7ZTY+KnJkCLDKV
HJTtkY9hNpKmPCTHoaE5cszUhTAlhHrsOgg0SivA8GBCir0aEp5yk2bTqsnImHQl
DyJkGwQfEw4wPUXA9zF5l0C28KzCZ41wLlKGF1JVReuYDKatIRx42C1b4qfG84eM
ngH46mWSxVARgkelZl/GSMFYiHqZNqamPInxrJBl2J0NcxJPLM9s+fvFjHpuFqXG
jLhLGoqkSPe4/hsHUpAL10TStWwbrZwN3zVuJCCfL8TDyUjILyNrdZnHPIUw41b7
BFTdq6efBZdbftQL+XExkYJD1hMWmKdDXjdWHWY86zFbCvUFPfuSfSIwsIPbAlLK
bTOM2o6FdBvMIkM5AjuD9c8Oi5wAB8mMMk4QnkwmSWI7rs6ynyzTLQNvCWdrdlg2
JwAb5HZc3tFe1bbQYHGIOwaTKRmhFusMB9gTPKLYlz06wA6b9/ag7JNxXbHPx4mO
NefXNndRqJo1Xr6c1QbEA7sv1f9j7xLK6c3YYDvhn4b+jcXBhfYdbnQli13Zm18O
TVIXHT9FWeqm5wMZSZ8eu8edDB/av/AoOyt5WPLHIytAMWaqJtfSYhNNlWdDnW6l
FNEhFjuKnsnQGEsJKejlPfTWXotVRX619T+vMingtjamxTuliW1azLPCB+JdgAcP
NScZUuEiEh+7snxYfUek10bfNreKXbA7HxYDyesiAs3cIBLbSUSP/Mx1VHmbjiFv
02/L/iBUe141VaepCHdls965Qw1OuusNwH9CSr1fXxgM39sF9K+NTXlbIBGwfBgA
oiIs5JGanIesDkWwbNC4U2dUyrLv8lRC4qeYsf7guPLHo/xNkpWHOVrNcdsfhsAE
U0ROEeAU0XJWL9HVvMbukAOniu89fUkiuk/9aLv6x97l6MFSoNEZRhLF74x10sQ5
HvsrkHhfV3CmE1BZk3YlwH5ZUJQ00OyzzKJSmHm2pWcFJGlAEhOPEq5uXIeMUe3T
NFbhFAkTIjUeo0kbGdHvmtu7+VYheTBtUsmus0lCVlv5Q05/yzY4Xm1dFe6yO/tC
dBQBKvlhmF7uDLqZ8k0F21aLXwSX4BPbKq/AsT10pHbPBuOcoiYpGCMO6w70jqru
2lR+Wfh1a2jLjwSMmw5NGOQ95qRVxtuInaVoqnhq5g/DHwtEBURGp5dOfQxWAkqC
bxY/yt8dgM16RHub6kHJs3n8TwCP3+L5lv78Zd9cOxXV/zXKF7UvSPg0tbnFWzOf
AmXkYqDyT4gZiBYFzyrL2sw0zZJgwCKYHu/MnoxZBlKpDCc9TJVma6RYYcUApCZn
p8xElea+216ObaL3DFXfpKa7fe0JXmw4wTJ8Ii2DYdPSGRiOiYEaOVGbRmE+UXUX
AqdYuXzpo1rTVwnlj4aCkaX/GsKk1H8qw6p0KEUVaLRJc8VhCCJ3N+jdjZHV9CMK
lomggkGnD2fKi7/qD6qiktm1hUj1WpGLgDJG1s4O4N3qz3EMwrSNrXaux0HnEXa2
PpNWBAZKQQF5I0qyssD7OgoCaiwsrQMb35FQa02vxY9GDFndz/Nd4NHiDeYgqwWP
MHLpYb44BttA34cQm1HUlQjlVkamRe5oFzXg4g+RSiqn3BZoCaRSd4HVap/AK7Z7
2rZ/nsqSO/ynuQOSAk6JGroyDrKOBIiRQdN/ZnGtFPlOdAD/QEHVckK4aUvIkquO
7YT/3C8gNYvUPPEXA/y0iB90rQ35Ej0BUL1G5GgdA4WBAUuqSruF/5luY0UFgZxM
h5rkz8s/ToCYfEzMkhS7d3WQkUKtDvV5NEi9QXP2G7ORTlyE8ysL7i5ZK7fCq9B6
+GIUpkFBo0SF8gthBn7SDIoVsQbppCcawls49vHMpIxmifSlO98w4m80hn99kCZ2
BwVMzaY8dFP9SGoqoK5sSIPa25t5AlN1ax/XKuy2q60KUgHFMgs3AprxDhqnIafB
vr3LSAiu6GWdEmxJeJVi0bJj0tpJM9RdehWTDSTVd3olrqy1Y+K6Ak6NqP/hyaoz
H1+8ChsYGEqFYPaueOBj0ZsOh2LFP7KW/VCS3Ilf0k3bJT1FUw4Y53WxNd/HWQuY
yFX4TnJos6CgmanJpJOMTX00LzN/nivwZ6bQWhs7xnDzyzJMw1jvpLc6tV/6SnOo
WR1BrZiSayIELSQe9mgeWla1YE5+19/nH0ejjx/Sps4omEUAxCDdRDF4SHhZTA3W
hpRghHXCPVObjdiqJfQ6/w2dkzx3/9nGT0NSbm0UByh8amuKDmPW6hmY9MSrtOYO
guFgM0y6jCRx8aT6c1m45RKBpVRzT7f2povN2CCIVEN1QnHwvan6ee5PxMvKbrJB
ztWaqEtI+UJve6Ph5NRP15cDkOg1NDLM2UbT/Hg8ztNEafgh5Ff9WEWZhJslgJ7t
kqHOY81fsfueLWyycjZPZRTAppnbG/LAeuVp4RhxaI9jn6DzmvLg5eKsILyEEcqR
JMNA19QgtSlFK9yxogRjtFmhuKe/dEMr4I1tjjdAJIp1iruRla0lyOkGEP/upPHm
ooplBjFpqivTo6OCNjTmZtNtbjZinOQhuFPKJ0yTQcT8ikGkAaWS7df7kfk4BX2D
iLxaMrPb3/GnEaTVV8bB+xpTLUGK+FG0+qoiBPwDPrpym2y3ojpg5ISfbDTmeA3G
L9tlFhkIv+c2FgotUnCUMXgQv1twXiemQbxzH3QmA5jiARcL/S6kBSTZdtZBJ8AC
hN6lA60RkSLNxEN/EK1TZVilFT2DonDRXLCJhoQX5WIyntiAOvXVrd9IKqwfv2ox
54Xe0pLhsx625vEINPTsSzHiSGHzI8MBHqQecLlHnzDBcU5CMBq9YnYqS9wrPQbs
Rm+Fec2cM4qz3t68k8HP/kd8DWfLbWYw2euWAX0x0mrA3BfXOZSr2mR3KDuTv1mh
88gWY+H5C+KrJxNfCW1j1fLBjLruYytBwODJbqSnEyGRLwJo1zAGsKX/iyMOTybG
I/TrJzpWfOTaufW/8gF206hz31BPTqk8fWmE7LKKysJuQoFbqJwijUN8HpFn7Unr
H+TLFnu77AwQusvUZaLatonR64f6hMnTD4Tg0z758OFEbso3hO/0a+OISyeqNqoI
nSVDcqME7MHZTqEBGGkdPiHS87xQA6s4YwEOEcHDP8tdy0w+2pUdJqjiS7ESK/eI
L3UlizqtAF1NRHQp7MJ8OMGOJrtfn/yGANbL9wNdKmFSNSTGvoh19+GeZ1gWAXVa
nOr3TCQYoE6sxz+CGdIW3BurOye1zD7Rl1kOvxlvfw9/1Dfz3wnQ3kGsZNS2cksC
gwsxJau1PdyeDDKgo8Bqz3RZvWY2hbRVbZXOaCXIx4BlMupSKne73XAc/ZgQWb/I
o5wy1+ykJJN/ZXhFGSQRydYggUygEeYm69TP9xtO/MgGj9Tcc946oe1PNk9WJQbW
7pq/wHLHFrZQpBEZtPQbxnEiAcjafkcojtmcAY/qlszyMY2TAovZQuh+aGT4VpTi
Q9W62zA50WrzkAfmgP10fggMy/IvN1/0HMpFBjLuyQv3AGL17mLl2HK7fCGrcK8N
JpnpAyqxADLxsmjCZ6UuNhhajWUa7J7E1S5pV9eJDqYLMVvuAQA1zuKVpEZgwiH/
Kqqlx9w+WJg9NfsL80phakNztpLgStUw0a/yk/G8hF76NoIIAO0cthVQF8BuiHJK
zfflf8A9/gz7fiW2C1rDFfMttdUFpdQHZ/WZujfFJmIAGZ1LajshY84e3gNkulEi
aTOkad6sro+gKSu+zQvtNXfLHMf9Mwty/Rm8Hmb9lm7sfYqFj6jNEn3iNvSn7L1+
SryqLDMM9Prcbv8TPPt3DjapKXLvCdMG6tioA/Qxwxl59OFliKgzrzbc9SeMDKVH
d+F4kRnQS1odxhFO3vEcpVVx1ytJIQbpUKzWP+Aq7OspfHa6X8lN9VORmIF3WoFG
EqcO0jKhzJrMHtDLD4bQ8geGUye5jj9tmYSTDcsTVy29hj2ixFZrBUgzXaMvvn9L
y5sFS3WeTKv561NiQVQcrBmdUCQSykf5CmLhbL5rzGdYkE8zQ6AxryT3ff9ekSmg
Z2nmZ1x+f3qspCYUXI+pS5Jln++2sow0eCAVoify5gr6uvEoIy4J2MR95P1CdDvK
3ubTNULw0XgjItWCfJzuC1ea7mFrK4L5I56GX/tnxRLt+EhqG/mA8Cm2BVil0VVO
KUjd7pJ4iCCx3I+y07YoxyUJryuAdqWgzF7d62EdG5Zno1vzd8AckZRp8kHHA2KE
MzvYSb95GX2jX3tM7OreDzuMG7WQOs1t/yH3EyJ3vUZuDp+l5JcO30gBFB06o63s
kYaHwfm9pgWNPMrslDzOaiF/Tq9w202FX/D/WFMDMWmzhJZC5lQlWrIChv6jAsfB
G2qRuU2J948WjkVQr/aGCeIP9uDRcRIVfKrk2Iqt7Zni+O9aKSgrkHDd9y2Ya4yY
zWRyiuECfLvgGD8UYr/wLPVItNXGd5VC+ignEJUTi1LgKuaBlJpzXeG2Ar0klFeM
oI31aBG5kolyYpFnnAUgaHcrATcLDWjHUqZd85xr6p4NFKBe15hDOy0iiF0ZPO8k
KaNi9cIdEBBa1rk1xadBw3A36ykmF4UcrlsWsHhJLQyNl/S+OMnwH59HGdtr4lSG
BxsY9jQXlcUljIvvR9wQSfDJSgpjAEI6R0/W2eQdKvlayV3RGxtx9qq78BCQFmaj
Hy1zLXfrrgigub8EQPFVMtG+3yvL/ZItIYonyTI+jsTaeQlru8q2jryw5pBwJoPL
DuJCvqJ8tnAkLJbn5T4eF732kT3MjtTUyAm23KvF1HdlXgjopbNgk4NS9nC29ZgC
a+Z3+/baqe8nER33ziYGmZGouazwXYoj3SzsCZJNR7ijHNykljcPMTYgZYgjKjyQ
XzKTQKO9b0wh/VN4ysXK4B/UQ9Yjeh04yOKP0BlyJLilW6DAFQlJp+zoVETinKBY
Wvi/X54u2If2P3NDdaaqJ2esHqSeC8GSUjvaZHKqV5aqRUTHGbeQvddFVHOeNh49
6DOhQqmMrLAe6TmOA8zsEbSHZwwTeycK1qAyNIGzmPVS2OfJmNECnxLviU+Z6/Di
se7hABCZUEqoc/Zvyg73YD8ec+LEv9n9qrqFDbio/7LnTvLzhVd3v63NU3uW5+8w
zuMU83+gAFpQgXWf3PXLGTMfAP+Sizj1ZetuXQueacKTsGoi0u1ZFI7AhZH+4J2e
vVWjemk80j30yskH1j+sVn9OiQwaPaQqfEa/1a4HCvldEX+3E4k7vKZMyPNITM4U
xHp1ReEnXPJDrn5nzM0zA4xhycd+NUL7SBu91JATQeTJtvj8OtWVpLYM58iix+bT
epEcBuJOZOhqSmuyEYoqxf07tbch4izi2N/WNKlsGWs+fv0nmyI5zqEl/UMO2MOR
QOe0xNRmHh+9qYpJjhUsA6QSOZah9zQq5p1JIGg4GQBg8oNh5AQ3o9Zs5/GiraWn
xrG4KYY79NqtrCAcdU4vFXKd7UDC9v5adgT8EzTYL8n4YJKLWix1II+pBZAx7RYq
qJ51PcDUVIfNhjlDHRTPmmPns00XsHb+61xH5ntKvNinhf1nNSKyl+YTuhakail7
+7ebCJ6J2erZ5XnsRzi4srOK8DH+iS/q9kfHCdjHatVJpqfBbh8TXv2/cSFmiaz3
xxr3Cq6W8s30XUIO6wj5McUnkV5VIaeM1hZ9BJf32CB+l5d5V1+kLVaAL6c1nuJC
kb+556OvDuYzvYPCT/t2wt4Sewk2f1mXX4bLrDiJX1AYsGVr1LII9Na8o2K3b4QF
h0kOnNU/mgDkpmgpegJJdb4PcyQmlApAnr47m92gcq9bn/6BUPH/lWUQNAVNgeLj
b2OXTP4QZE+OJD6HVHcw+eVoN5pnVM+z83Vual/WfKrEyIyq4IcgM48Hb5P4Wnh7
IbHqtqCCMPU/L4cglAUdK7YecWADhyqPVD7bXrtHoX4qb1lfdrqc+mEipN7XxLYK
Lfv6D1RxL36jjoALnT11T0JE51L+wwX6tS3O2tMroA03taCvB9gnxnwyVgQK4pwR
CA18gIfY3V1WK1YZQOicAvrtCdvL8H0F3/KSOTbFqocNWXoiwpYk1hENuHudrQE5
UU4WTqZk8aDDRqVd4l+7NUtN56dY9Md5HrPDNExUV1sfEeNBCXNtxVBnicGC89Hh
ZbKgER52k7kfJwIGdIO3AZUSQlhrLvC+7cKcC1p3j7rPvT+UBkkddIROd/D69/ob
Abnb3WRVmrBYZNNmZlYxr4h1/czkYJKyiNxqkZvkMyBwhacOk3ZTXIaYEH2j5MTg
L5IaIYTXJQxarCAO52x/5rw+V2EwC5smFd1kLs3sTtJCFRm5lMDMxZYpIwOA3gru
922nhDF9cVA1jgOyXD8HazD/hbEO3SAU98ssGUq8hz4z02o2enoo1AufZNXku10M
IPMRJNJe0T3qUSiKkj7vviN4tXlUJ1bHd27TUEYzrLJBwJVTZ+RDvTCTR5f56zK7
ni0m+RSuInmALcUhJQ4tWqlqtG1jkopCONZpaAZbfrs0pXxro3xtHrnVEsvRcB1U
j1nK2KSczn0zxX0FHd/pMleC4bLy0JO1Bmf6JOkDYzB7/H/dPCSGWc8mqJrUgE9E
jcXJysCuFa28KCSTSJ6FKLlUKwZIlCGnDqrXxQjF95or009il0eDB1JOpscx9/a0
gmuV8pLTVP0f7RuALy4CZFwMtGFNTBaI4hixm2wU2+JRVS8uTnrR7Dx8m2n9VEXr
MYSMhCiRsJRXn9Y0NHrPe7wWLWiQ5NhIMXsFqKCb5Q0yzvVqslE4cLCEXfLaPTXT
YzVrwf0/RtLpX5o4OktbGuxkAAKdm0L7p6WshP30F1RFYQxMkAdtgiSN14nz3Ycd
rgF1pVmEsPP4+qEARjd1HZCo8xrdwS8hXCWqJVW0NH89jYegF7JSlS4KAogfMeYI
VEqFjEt6rz/rjbGbvFzT1JdUpHdaYgMZpKMez7aSepGhOJbhi9oBBw1u8zAi+fSH
t11HmzVBYM6Y2yjZvFejWl2WQuqpNzm3rvH7cS+ztH/JqmjSBn5TctgZgzDDcyzg
9Crttr+CWLkE3ew/4F3ZhkHio4lhq2jZU6mlgvBGr/BHqXyvP6qlzmyT0KVvzXmx
aGbe9j5GSQ8kbp8OdX1dKuqNkRrURShnc476xBvXe9aOMq3B/mMonO3mBg+RKLfS
j09oqSWqFm7XyQ71HbXqNcBb5nNhLbXTskGHag6cgHcy+BicihqZvlowozSjCRpo
2i0UpvXzcpBb0LN7ig1dPvN3vao630yxLp+vOCXBolgDIBNpBisYyr+PLEN+/fcf
1LCHEkok/AkTxf9tSy+WiwNtysbXdHbYK/VoRlunDgNl5fyQKFLh7FYAZX6gVpav
npyWyktjWVnC2TgbcCtmUv6/RGYaF84faz9kknY+vaRZfvSFsDIhr1B3oTZYEuwQ
eySvzhyybVOFX+n+y5tE182eLzWSrEmEV797rVOZNuinIBDG+y35lz/RY/NPLG/W
8eeXoKZWJ4d0PJWY9DKyoWyTDZWnfFNEMmkWm2CmbK81MfCdROvRfO38ttJNLPTo
QZ6nBeWXLA9gjOr3AQwi8frH869WJv3GN+gmRiqLxElFvePJP0uBXrroylOvb4RT
xl1Oa1kREx4G810DD5KuZoJULFp7hk98wfR6psaPfTwVEYbMBd9V0jJyi5B5cWkM
VCqu2k+DxMtBjLQyme0I7MqqI9Ym3eEf+eSNhkXUqZBlhm8wJtX7Z/1NXzpr8Kk3
GKgpPQOWVSZgBMxXOLX40Ml3LQKg9sKjYyc9C6Bb8bXie2xA1aO7p9ZEeTMRu6+z
UdNHEUV6/D5Z65MPj0Z//RUc3xveB4nXxkFr0ZOLd7xIHqYn88+fBQoNw7YEt3xb
2w/d9JWhFiCgPNowrLgBUJglk9CQ2G66mmQjnpoSFR2jnxKHKBX8s4jdXy3UPeCp
fKHHhYkFn4gaVqjXdPfLD+W6HroTVEyrMjCYVr6WXd6u8rIuGSy5BLa4AC/5S8vb
PsMu/7CrJii0nIb97uHq2d2Q8u3RjP3bR9pH7ShfLVDh/kRoUbPzavFw2Jw96eic
WxTJ+Huv3WddNdiCobZLzAPdTGd8Q0RNgz5eNtLkFIOvFW6N1xaCfX5RLuxU9PQp
EyyBbmcBR6IIA0UOQ+gfdGLGkcbksYbFLhb6ioJiRvgd/bC/Xr/BeNKQyXe/HQWn
zuIYqT17QuCOQ2zxCCe2nHVQYirAfNiwUEs8diQ4Up3c4YGglTQWuoIGqhWeDOaM
1gKrzmAW/R2YhGrAy5e2dgDsqMTPFI4oU4FB9OSuD8Cf2iUxlNNb5vvPyFpIJK+P
4TTSMsF/idQADYj1gknIec7mQotkfVKCeIj6ZLFD5v0O3MmI+uNM1ZzUkwAm/vc3
H6zfcBlYNHk2Py8YhPp9YULbs7vEUcO3/bvQtZt+JK/o+JuxBrZfFZK2uilZOmxd
eFuAVHUGAV4qsGceno24XvdkrgVu76kBYuN//EFgS5Q4rwuzz1yQwRo4OEj8f5VE
6/GPBBt1wDs7uYuJIZXblIYdSeQKemllSYT307h/I2Txkb2lYQ0RPWutCdzUz3Jh
JWZcSfFy2Q5Fl67Ot7+hInboJ+B2q+sOFxF4VUgA21hjz8kCHbJ266YZxKSIYZPZ
eYexicm/a0PGSbRIETdswa8IsQA5c9PHz4Ue6hGGNbyeiPPnWap/VThRuj8xudae
pDFHFkdE1ZBGMPd7nDQ9uFr3a97yqpW6rMt00Gev+YZNp3uAP+PbW73US3uRrL8m
idE/MF/KX6OHeGMImlLq0LZb8biTLYOm1hDgkdoW+FCk+Oh0BgEtkj2v0Q8wDTPu
Msb6Swfy+yXn7Dq2rZhTcA6Ez7oCGxzIx1jpg3g1gLLru52w/HfFB1awuveHcjDU
L7ZvMvdpcahkc5WC5eiUFnnUVvYWok1OtJswwRyVeuqBj97IApqwXCeCU+MJDR94
BwqEB4U6MwHEccO/1y5kwIIZoVhp4DZeV01JueKb3YVEUBLiMA1nLivah0bTDOGI
I5rjnHFKqDxEUVPrK1UkUKsp/thI+EGThJPOy4Il13UUH1GsnwsL2Kcm4Kg3D4Fk
ziQ/dihymUwsZ1tl4oxR1UVPm3zfYjk9nN7Iv/FNA+8q8/ChJD+KTjua7LMpSDoO
TmgvHYwY3y9C5GeDoFWOwfMZ7QDRzvdNyX/AtUcvMnqdICW9xJixwRYGxt96muin
ui2ZmmaT+/PYYe/CTZ4N8kuNjk56lmUS4zTZSD86cSSGhbS+83LI/F+RRZSs5CUk
DHSIVA7bk+E+HSBWE8VjMPOBFl/GhoaVHB27si+SAfZyKUcL0n6oF0hJHxu30J3k
evsLMvRJr9CG2Eua7+/XcH/WvAP8qPrbSbdZqIIr0GrBUX+gewnjMWj8JHMytVsl
vSQK4flAChPKkYSX6I34/BFJumJEdTHNfpxYCtsaOfKe3k7bU0Q8x5FoQg7SJ0qB
UH3hN4P9bDuilbOhDpi8DwEqpSIxHZ6hLigz63sz7W3tucRgwtlRTiYt/d/5xj9Z
vqmx04Hw8O8tCxEbUkf0kmXjA9GQwj5ZZkb4mbIXGrnTMiJp6x0Ct/VFRChIGYfH
JqdyOkVWIHSBwcl8+ADzRMiXLFn5ZFnyXu4PccYeF74VYXz8pwfoFvM5CD+Zvg4W
5mLSwI1KfN5CU/fmxNtHbGj213klh13xY5fsGvxlaSpYTkX8wsF62vuMGzIzQ9/s
lNGk7RaDwaRTuuIW8Zd0sLHV16Tz+CDTLvDTiZZrRtxBfpnRZPb+UKvmktVePEJj
GQE4nlo6pNFK2QtYgVvtx4kT49aVEZZ6Dh61cfGecSBV3gemysCa29kThd6J9+FI
qIfQS455B9gzih3INe6Ww0rao921u0AuEVNhMxe2/iqGpYK5e3bQEjMmx/JYPz6E
GeuEv1THP7fzGOvjU6IpXLntTUrDwRhWlnrFapTjNqC4iX/i7EKDNhoMujEtSjm5
6CWNsh/JfXqRZ8i+htwOd/iJs+qzusL/7CKMsP0N4tZIqjBHcHdD1cqugKmgFc2k
0OM+jl4sUhC7mAp5M2J6H6bxhW37UKAJmTHwuPlDANyj0PKDtUH25bOFSUkXsVTU
pKFwLyQAIghDmO01+X0fi55NaQC/Y9LpzPQ9precpLl81k6omGtElfV6YYddq13k
HXGTFiMZiQEjqvHvsXHDKDFsUnSFI11nCd6pPXmamOL8x4RBTVs87A3wp77UP6XB
hxjjDQz5+QRH6MrcoolaO9Tuid5fcQg73EtN6MgIN9FmjWBvHg7zFrlS14w2pN36
VKmF0T7EOUjsFVXYeZZBSSq3R61/Wx08g+tY0SEuucsMghU2QBnsojgCFTElHFyX
rECGKCf7+Ttv3FcpjNQUP0qeU56gdZ40OD9qXuawiQAFYckK8azHl/TESLVLq6dF
ndNbF155Sc9hpSKfmtfJ34WqhcMXBuM+JsOkm9E0GwAH+GF6LP1CLXS/YdQquzxm
BmFvH7JcfnhQ06DZ1LVsJmM2bg4fNKiW/jPPXOdM5/fMyBbtCTBODVynli4OqLOo
4/SoNJgNu/HzD10ij6IFJt5/gcyXFPbOsC8jUHJfCQRIOeG+Fff8sJ7uuvJIrHt5
4hc8lrGD2Hy3TL8MSQpPzuJ61T3c484SbaqFZ2KSiCyL4rN7a7sxQPFWdpG9S8MY
GvV4Zqy96kTMLzaM5UFnUSBZXKSMKlsVw5yoCxTyGNBe1SRtScdSZ+bwwRKsJzIa
yj5GzPYLsMFFrKhwxJLgeXJIQFyrdJJS6m3ca8rFoyqGdebb+clMUlUuyh3XWJmH
2f3+s3H91KQZS+wR8/NZWzaWZdHtpqdYtF8J9GYr0elGUWqh0j3FM4FE08n9DtMY
Vnau1v3z0YhAJPxf2OzABKjKjddo9Fdbybw6A5NX+lqsPufPJu6u2cBJTZKQuf/k
QiXTG6keOsHz6/pknVlXa8NOFlYsRoNN9TK+LGEAeH/Ko9FjkuzW1BIvQIX66H/N
2FT3YsI4E3rv9Z3a+6gzTVTfwg5/VvRFfUj+5wdIB0mLQ46mVQPnNO2zEw5rLTwu
mjiYvNKiGs5bfX5e9BNtBnfwU3jEiLTgG0LtrgQjQ/eqMZIRZcUgw9Q6F4D3iSHr
TwDRjWUA9FD8Uv0hGnVLrVMSnn91Ki2cQy9ZvO252unPFNVmwYSwuNuz6aHo0k+S
n/tyK5L59ZnRsVNJgLQgxd26/F3esnlyQ5IpFhupu8dfZkh12sZL6aBTd5MK8wus
8UTqF9uHogSdyxqHBi+saf7qGwSxNoAcZ8A5FJoqUhLrpqI9t3WJOWlb9IYhcwun
a/2AxlO/G2CIFArql7VoPjuku9AnWSAQlv63HK7GJuJs7P8CZbBA0GZLI2WrcCUq
zvyOutAGRD5JKu7QkqTJz1B5RocPfm2+zmrLX6ZJyTnlFwlxPhfz2THKpfaDdKo/
wfTnjxXlwtbaTIO8tnlos90/0U1JSrYwPmvJIdJBYCvp4TavA9IX+QE1SJx+LIOB
bRjYB0ebiFwLhtQNdztqq/JY/T2GR1ixrV+dpBBfojsV1wB8LELwfcBS340Qa/uo
hTML1q453REESw1i5BWBc43d9aetdAsHufVRywtHO8YYahon3DDR/WkNlg8h46XH
9vyjua8cW6YM2gUYnCZn4I6ocJrNtyF2ZE05ZOyTRZWEY/fOvEDA0dfAiDiHTGsv
0FsrNLyD2QJTxz8UDrkfwnFaqDjC2yVQoL3PTQDTMqjZ/AXx+RHGXdsy9ZjLndE5
K/w8aSSZNqUmuD+RZxeodRfyVItJf5TUQftwYFpzkAABs2mFd7yuhaIY8fKZJ2Lj
aj84pljGAiAt8azfzW2wk1Fh9VlVpsL8RNewS+MOA2Z6LrZp+iT1CzYNav/1/bjY
UWqilazI0gIKZaEDUlS1GO5WWLDSU6xkdZf+n5xLQUELArd52wJhMEKwQijdeLxw
MXPeFB8sGRZByx2gSNtM9VARdlfZNPs2laPfnJSo+gMuDQtRF11F/WZdyI9lnUjy
3FJqjVvgRaX1QkGD/tz+egwUG09YtmZFeFwgmoBkARgzaFgdNzKEji4axh376NAP
GBxzSwdI4IjuR1FmSAlYlWBU3YS8wjvRMdKg1xBuCy/0DJ1vSlhwNThjVnStpUTa
bckH8b23XBOwt7JvhKo06OWV5rNJ/55BtD0533NxXqKgEeRVn3HBHJAx2s1Zq10d
ZIfuWPS7KRIFOPDXrjPsuHw2RvaTQUB21i5XSwbmk4J6xz0JC3jIYdrIt1M9ohUd
1IwDb9P/lxZoFrAqXll7j746rdw87Tj3XCAwJV5zrmxm1d/fpeoLO2BmqTNJysPr
ufetgzndIrp3msxJNykyXT3rJWtn7pPu9bJkZ9CKQ9qGKFPGQ28/163m7o4QoiMN
g8Hilod5sr7oTc56xCSDyJ1lGzSBLUeWes3IzKii/ai9YfLYjbgc3wZit+rOnWnn
MFd76VAAzhqf8Zl4jxx0q/Wm4lITNNghE/dFgAQA33QEa0e42BvP1b1Bf9qlNs3B
We5reaURGQEDc2yhJ6xQUj0EcBkQMavPumTn8mGHQ0VOoCr9ajbzxXHgsyjALRUX
4GJGxhL3XyExbF62/X+85y+Gw69lyPS/e1tGl6dJ3fFDSNMgJ8fFkhOj+nUbhnj1
dtuR+HiQgAu5R01aUEfrcyYZZ1wgf2LMaTp48JVRu7RItFCem0XyXrXSozbKDA7P
YAu5KDBpeh/i1LKvNDTakKoyL5//YhtKMl1eo2YWmKQ5HctRbInMIkna3KczBjr3
ZdSHdz31fPcxqlRsaYsRDQdtEYViUogPR99LWbWxgACjgZ5mJziEosJEav4zg2Pi
53jvAhmTNgOkKsiRqxURFZii1/gM/iccUt7g+vRez7d9+OVfrReCcYinI8YxdxiZ
gShA2JQl3a/aWo5dWLTuGVH/0KtFbr1iLKABOLvc1xAnMrw4ySzfQs0V5QRLuBzv
TTYsug1DAp8bRXclZ+St8z51yV+nF5TLA4Di69DvAduMnOoHxdjuI3utvH9/0G8Q
FYUrhf6CeBuZsHNUbJ/VmWEteTvtQm5PvHRVfPStKabrkZ95Qeziv2PgekGwOdSU
XYkU+al7zr5ZOd2rDwcPY7pScbq3Ab+GFeW2+GX7kJBX7YgILHF7JZNFX8LNhrH3
LxBZjxTZ75xU2J1+QrSS1cKBfftmXwOWasqR7gjuSJGWSmwCxRGQhVXRVTPIvjK/
zYQIEpHXfD1NtIffzh0wcM9iGnzRNrvH5qtoFeRltqVo98ytqRFy0jR6cKWZR3DW
Oh9UCS9JjL2Us6AuZaCuDcyGB/+r62m482r7HxqerY5Imtwgxp75XLGwioYzKYl3
tHLTgbqrsNGcjgsupZ0M+bx2psf7JKQH94KiM6QHZHbDMCyjLV7+R+yb31ZJsaAu
zgEyYSP97MGz2wm3MnLZ1EyYoIxwY6h8SLBXumCNBrVqhetFZDO73YwAtSE66vpq
hNsKWvQOpKgN3knae68HkrdWqznGgClqmU+yZ+hCyueWCy++FDSyhzbrEVsEjXAq
p5YwyvU2VXkX8Zm0YM6zLca41BATdf/RkIkBXXNa3mSinTzEiZPiVjPqs91c0eiS
83Zl0shWhSF3zNSLR2uyi2qK2jzgJN3+WXx8/OKJA+DnMpAJsWwcBeAB2FspJXXO
z0K+OmvIENF0CoD9eWghElBWSY5MKncU6ADXUPhXhrp925w7K6uyy/2xUzHcUuc5
05kJbMKJVKGvXuYez9tYVo3R3s4MEJVz40dAxT7dzU4I6aV97hCojQeZVlec5KEB
oDeTcl7TmC00CX2xL2otOTO0H7O1fuGYIoTJ7SSTrxfXMW1z2Nqtzq9lh41k6KqW
ctfoCr0Fo4M4pjyI6KXZ+W9fxp93WxWTAGJnRgArNJK/qjShAfbHiYrb/SLZH8Gy
YMYXm2zxeBFbH1d0x35zYX7C1r8kiRCwYGa5xKqjz0YToiiLMah3ruFOtmBrYt0X
iXi2yuBOnkGU7MdF+DO+ccZX6auzjzslCroTOP13jZojSYzKBqdG3gfpMNDqpNnI
BjZCtgmOqKOSAkFjPZnJZkYtVSJPUzCsvrIV1FXmfecVApp4lK66Ost9LPNNYeJf
wC3xZOtUwrBLZOA6lSjVV82KAuZrr8qGRynJVV9qOyY4ayqQ2c9g57ooJADFyfXg
PxYAaMW8Rgu9T4qXCislc6gNx2tgQdJh8q8Az4PdHgEi/e/c4AIZHqcvhxWW0KJh
0B3uuTF27DLtEq+Zcn51mMbxe5EMQamARVptkzSTJwJkVOtWQ9iME2RnJ/Yb4NED
qgbL16syFaZPkP40ZJfR764CiBWFqCUGgWf4g3MOCRCgkFRiCMIGz1qOvS0tOSG9
8SLp1TB6sd3cSRDNeJ3I90fpcZzN1na52WOyqiuh3AJtei4k0Ig8qvOuaWDD0i0U
THD0HuUAH1zJ2QMrAtxTJSAPAgEaKyXUc9DWkzkwG35PK8k9z4fhQ5UeqsVevf+D
+mbGRXTA4/vByQBdYuM61m6shHQf1+tFjcflwLx+zzuclfh0g221I9y+VXDC0xej
378pXPwGANuJpMu7y8T3Eabszdjk0rAHc5MhSXWxWgws9WDqF1H2WRjDm27vR6E3
68LcO7aD+/4W9uFlQ6Brg6KtxxiKnlzE/uLcuCfq1s49pgK/fF/NbXENaBmG/4G2
pphUcJMfkBqnG3N8v7ki9eqKeMkuS7rE6UCrMGX2z3bW559rk+A0k4EmolLWwiEU
Fi3jLYVYNI0lSsEvSOOPqbRkTMp7CGTnu9Vv5aySaAT/U/AWSk+ZZtHtvOh76t26
34BjUtq05VwvSa3ygQ+TGCEnQ7LbCnunSHcO/XVygCKto7yGlk40RUKgF9E8w69Z
TqDLQdkfVIrzR8szr0U+ZqVvvfEIUgVhqoNWWTcwjpy88r8zPtMLvhtV6qr1Qn3J
dGbv9XdBTzGvfo/lIF36EL56TR/pB13jMsbMEZYlEHauKtxung5JsL9vot8pVJIb
cbnE8tidwyvuoZYw9DZbWT9+qk5MCg9zOXPF1yIUWoYWXdi/5/wRaOCIMAd1Ick4
5JH/NQrIm/vWMqEdBXTuGRzkgA1LZ6bcSG6zsKYfP1DEGJigkW7Q/99clWKAKbA1
t+iZVSQzUyaOMYTsgFp4TFAvAlyDiwMo0fepME6ASh5CSg6XCU/drtusop+1UOp4
TNRnZa1vGkV/58dAvtyXXube1I23r7p4X0aA+2J7cn6BNenILQ2MQKkeJaqtAAXP
/25lsAk3FdHgQ5F8r8IVOX9TJAKgLlIcU4072H39SZWAdplAqVxdtQXKIAuxjgep
dqySFBumcqCXrg0rNaK3MAcJI2v3s7G5a8/56St9meWfokhMDSWu+ibZhyiKFCZc
sixG8X69MkTbercv1IAZjzLzarqNXuUv7Kn3D+muHcrhGKoiYUZuqTmSJ/C/Hvio
M8NZmGrXXDVbVwVOtZtQ5vLQAWoaoFT8hcY6H1Fqzn5xjabfPYLJBSrMHvXEGa7q
XU17vENegblGxKW7SeDQ2jOJTO88I2bSgg4JIOx38rScmz+DSaF5tseKMPqh9sM0
9fxFADnu6JBVpxiG18Na6aKgoXalegSGZKjvY3QGm6tiKRzhJxZAoHXxHPxEpmW8
CzbWxYvV/1csxVuc+NoGflMQ0rfElgOOQuPgvLXNeAeTndelEs/ywEGCoAwB7Lv5
V3JnZ/EY24BNc4BS6ZG9D1nlBRb6sPPcc8WzNSWDj+05TRSiJi7+nQiGBZS8VJUv
ERkv9qGmgXeMDqQxm1UzpYo3Y1EwG0Lx8OhOIaMQYBi4r5tHI6DV9qf9PX2ylww6
k5XUzAJqKfzenbCwKr3aSpBI6450yavpUv0+mVYC3D943NV+YfKQ9vE5JW/a4Z7y
GI5LUuN67ki3Ry9j1B6wwDhZJIgEDFhmpOfiTylmydp4wUoZQWSEg9CdBZ7wRTwC
/EUPPvV/lbETy4MCbCernhawzOuGg2uY6QYghmKsWUdrQuEPfB7ShNbWDP8TXzgb
5dQLrWgMWuAC3Kkd5a3J/Qx7YxoK6sVDyNPv9NYlTN0UVvzLWZg3/5pF8s+jyiG4
vUUyNzFdgChzycfAtd2VVrmHvs/bpxE+IkMEKwUc5+Wh1ZG113YM6h2RjSK19kbW
ebnA17HWvkdG2G6h/xfO2+tt9TD9TR9ttw9WzJBdhiRas4fhLXtoGProLKTLy/1X
aRUlh8caS82dwaNaGg0Dd8zjeI6wMvOt90Mh2tita8IDhxjXk09dPFbZs7YG0gYQ
sI3q99RKBc/uMYhDJusLkZ7Nm5qCmfCi8XfneK5xSBrTuSFudj+wNmm9BZ78pAAt
LKCW+j5CZDqAVp3qjSMILqYaLGxyolRg2HjFeQ5VYTq9J2GUITEdSo5tWYLXDu8B
fp9VsmpQBhOOG61ahOjN2adn/8D5xq4U98alUilzK9PRPqgtePJBWalSG/N0wcZI
lTQJJYrDt2DSIUS2UVWkMv8tfJm5mK8tw3O1TxV3gBbFI02/fZV6XJlNZndTvZWB
ueDhH9YJ1dOo1rg1SQ6rQsasHTsWpVPIoS/59KvNZ/7gxsifZ4AamC0LXpoy0bRb
RyjZaiQ/0DRX3dQrngmeIIGU/be2fswW6ymmxeIzn2wgEt7CMJEbFN5yb8fWNqjA
siRQzRhWJYcvMeF2cbQgIveOON0BL6UbGCmu+jqdgPMpCu23XmYQHEb09+uYtKRl
e7kMP4AALIvBNumnSrxGhFVGubLLvEFnIa1YQT2UrAFJvGr779YDjkrMX62XjlBC
RFNEd9D0DLapPJU2t92Btgl+uYvdEqol57iJYjI/jgDU8FYqpa4JI5Xu/C1ju63m
aOqpIXwQAVqgLhN3yerh4IlAwP9aJwJ51VlOPMIAwVjdV3eleoG+xBGWtqS/lwdE
Wa+zU44tLn9/3JCZGXuKhvaYVMqlTw+fTFVMT3eVXeUlq4LYy9D1hcEN+uoWJmHj
/svdG2r78xvkmSq48K2eAO2SUX3eKNIFb4yGpRivDI4x2hZ/QThUh/o3nsJe+2ij
Nu1f33KHKQFry2unHSyTFvzCIKbLyUw1xymbUkLdvPoz02poiXjWm0WyYOn8aYRd
wq9D29LpM6qD6pueFMVxaQ7bn784wkQS/i9zud+0IAmvkBDTJu6qgjXWL1CnJLQP
PiWFgjXMniW/jQBKi4kM1Z2QK56wW3iKpMWHNeKWyLTbmyNiYwGyYqf5xCJvJne8
LHQ7P/CGL68/hXdAgQwwcMfQ5KogZE7rMlInZwdVtNnvYzG9cDt9vRe6wUxnJc9S
deptDImC671YE7O9kXWTy3AoYLSHTZU0BDCUphYN+Uk9DK2+DfgoQBV16F1JUVr/
oCb8vTaxJHUfAt9EwVtvZ+KLMfGSCSmsXil4N9Ks6frem96ffToelJtv30dc/iig
5OBJgKy9AynQlTm+gAjHxvygGODQnXznWLuHDOEUT3GRhwKghGWMIeYuJ8Qkhtvt
6dKD/M5u2zxKGd/TRHdItNrabwvMTHSQGy7na8zQA6f+zdIEwwvSFuFb12rMh3G1
Lnsg8trxIbEWXP+nTxobOhAWnxPBxowYFpcCqxeEzYlaG9+Kh8OY6tsZFtNtpGIO
h6UpZdSvp5cppFGtr0pbu7Nkddf1a0zXT9Gxh/PrHfwsxXyoG1giggLbSM1aj+Wl
mM5JQZiFcusTeNdv2oSumZKTZq2k3e2Y84pPC4ADwyDZMECVWdGGaYxCvShPdWn9
z9Bk/pe6dCRrzK8koTnYVV8Osw+tJ6drEagjMq1O4b6jEkMiKZz8TZ3p4kLkKtcA
c8TZaI7SXKW6K8jfhopyV0LJxLir+sip0ThkxA1LnEmLWSkTe8knTy2lrumTTS9m
X5FZYjy89Dhw2WCWgm0PyC8TwaJXDGq0ByZ7+OMN5/wtIqHLfCWSf/D6AokqygJz
E0NWAUFNb38lKi4nZw18jXlq/0tQvzByGFIiUjNxphVoul+X+9//hripF6eNamTJ
8//PTbEbLoKetUPTdr1xL0iBSAMi3QnDDjZUySo9LP5yTH1pNn2PhN/7kHZ+OnG4
AIoQCFxrrqADxr6EM+gfO1zcchOVHo/ou0KOOo/YKv8EcM/H2EYVtAbKpxfk81Vu
uUic0JEuwM57H+8kQQq0Igf93vmopZEoub5Gxjc3CLSrDKbW4MON2Bgceac49iBX
Bzw2LkVKfEZp3VXJDF7K3IGD7d0Lr0uSAj7Pt/qqzr69oo4babBGy3HC79Khw2RA
4UrfSIzcnqr5Wqbfvw822lPR2Wg7xQBSBEBk3XuuyZXEaHUeEepb54V2vlqflMha
f2UxpVosXxWHsVSeL798iiQoLKam14vj9MHjaAJiBIdlCgQfFV6H1Y3oIHukvRlc
TEm63iUxZ0RVf1pHCapUDCTEfKfVxH27Nyn5n69m7HVRrebJeUstGsh9voYP4Gh3
wjtDomyxbg7Rle9CriqMvUZ9fuxmPeWa4rjd+5DP0wPPOSfolNHUyZR1bUrvZwg7
d5mrC9c+NyKJIO2NBcnDS5eiCT9hWbUeUS+SvBJiP2vnKZMXty/82KILGZ+y+bGE
rWlmefsac/tA6z8BPpH7mgw4HG9uoKqDpn1S3c55Id9IhKTFF8PiTjxD7JsVwyxR
uAXr9KfCuP6bX6MKxVwngpkZwNv67+g+udLblDy/+esZR1atNv0FwwDwDHwTpZRg
yfMtj7bMatUE8EyqAjh7aAXnE2lxqVDyRl1C2OYJfF+syyb6iNrqwRagywLS/YLT
HgaA58t32ADcsRyTZLKku3oVNa2N3X2anmMulyDV9L5go/vlx3yhz+qmq80hHFk0
GA5V06wzErk0DrWMtN0C+nAnrZ6mzaqSeVP89m2A2126UUtfVt80o8HtB6huZnrh
l4pFlOXr34sB03ExkrPhE5P8aIZgI5FDxUZBE4CMfQk+DEdyN6gs5Wm+Nkubj6pJ
UT1xLg0fR2031F2xDfTtwQSQbAGsWjjhqfZUXuUT1yTPhxOvpwWUB/YUf6U1n1/L
aLsr9XtIQd45BGEVfiRwCHlJj43Gx4fCEMfHRXSTw03IM6VFZmlAEwUsRqNHgDG2
gXqfvFnUUSadh0gOkU0Q3TWaAKTrERRHj9P0XvAYytAzPE1KXqOpXHFClGdyryij
SiN62brpZN4yqpav9gI6AixYk0AOi174EicSnTkH6uNlGmXpZqUzlAHdN+Vwose2
MzcvokFLtijk5MHeV+QIUNdejoAyBrarQIlCbqDe+QR7dtfq9idKnfy1p4uoGE/Z
0Vitm/ZE9LJ+qeKkDRRtDWlFwBaG5f0Y1W/BF+I2VbFahozYRKnoMlNMNum5RrJi
4MwphInKDCR5OWpv43SBmrQPMJV1zZkd+nKLfvXfM3HkmQLKo5bOQFDUXM4K8hwd
xnX2k2g6d3nSNHsLFx7+TasrEMOvVMGeePdWoXwcdkgtPIEP9Gah7V7rW2JPNaG8
9NGeSSeStYI6y60/AOHlyB03K6FJRwyAp52ICQzYlywSmZpqzn1rLvl9GqVRypAO
35C5ADtMH65ZsqZvMZEJ9e+B2Zc9fqZcNGN3m2dyCTPte4M+0Jj/tYfGetmEy4mb
0nZcWhoGW4rt1lGcJ5k/b+ltixoMHMD0viGxTifTZo2nZZup3k4gSaWDzIMisHDh
Y08a2pmPEM1ZWRMclaFmbHSmrdCj0G04kerQjriwAZ7ImOv9yw0oW5KmYxVOglSV
LPOjXTSBnYJzfNQOxqK/FRfqyG2pwnVbuAXWz58S5h4nzPWCOhChCA2qOKvAclcR
zqZcm158knmXmpP3th+rqNFSTEjq5zivV9Ku/iGjRnJXyctu7p4W2ASdzK2ETWA2
hW0Wc76r+pZ81T55cAi9oQEYjG2dpcwkxDJHv4UCYr3hpsSa08m97duwVsh8ZClz
vIrzJv4AVok5jXnCnK5w8yClPJx0IpDWpIXnE2ePzgWqGlSOBRdLDYAO2okfCFa1
WMFmhQ0SpBe8IGHABcTKrdlS7vc7tZJVQWg60wUKX5gJmiR2FMBMQVYBN/hCX5fZ
f2lFW1jBGBvkwbCAPKnh4CAUTLPSKwD0BWxCDgOq7G2EBEaEfJ5Utw2aKR6moYN0
m/VFLpFRbSbIpktJ/fvaTfz1o7OPY5afAoKHBCgmU8g0XddxI8ui7RAlM6HAAAfg
4TOm8uzXiJEYD7qwBD71Wwmg1NeWLVX1oOmSQLBL699ynCsHReyXEEB8AN+4Y0gF
jcrFtvub3KI7xvyDX8XSUHd3cztqYUztzNWCpwysnt4jDwFXGtF42rRSFSFYO/d6
KhkBi/eZo8M+3Yoh0d3YPba5NKZ9tAgpqPcfW6hp0KxYKwm0MWTheMr9c8WWa8Ml
ehhsqCNx6TVlq6Re7NpDAFDzFNEd1rpKYl0kDNNuykDUiLfSLXe+f2bpOacdRImS
Zfv4OYS68zrOlkRcg5LIGenNde8aPd/j4+cRQkukluiqWoSV+D982D4XyHQtpP7u
PaNp9c2g3erolY1PnL2eURnnOq/exinmodyQH7C760YFVFqLrl45dxNtRlp/i0pq
b/AP3QXDJo6tmVZ/AfkBaoktAfyvPMN+m4SfNnCMgzpQeVNSnRXjr+67iUdV+DdC
yJ2kONlLWmZCvtib+wiOWE7U/W4+UL4PWFvNvL0ki6/Ym/FhiZGkFMCeyzaNr8Fi
g4ZKnLAPfYnTxQSyhZGaosRD7SGt0DS+z7ioWVy70DELyN4FE4uT+68qEf8KJqzc
TLiaDlo/6WSWJwcVcR/2PiMeobWj7OhDEoWORvh9Yi7scOTKIXhy8iduN1LgKaDB
un+6oORxQ7V30eTqARkV8jcwz2Ud4LVpe7e8oAlVyN1lEHJBc6ZPuFK6/KwPVmro
K4P2+bbelFjkIctL7IZB+A0mJXD8glAMlDNsEtOjaR3ZpK4hfsaGmK+0bfrZ1DjH
gyw5cQeF6M+W++jYGKxXNaP2pEOqvKW06uO5twrIa9WYPGeMHl/knoRtNoet387u
J5muE4ilLYLJ8ccS38+30ZqtBJqK6dQUsBZD9+u6VW7xhLQffasD9fvoc1FmnZaQ
mmwnpabjhty04PqGkfhHNHwti1QQmJ+OvSwmjxjRwMnDiY6mhjMppW3Glhlknl5i
lQDPSi6pqxt3h2eKMkq+eRJc3h2LXx+sTbnITpSInjlMEiLeFwD4KVGznQeQDbk9
JjkuPIch4GtWANULbyfoK8m48XBE10FADjIDY2lV8Wxt32Qp9zGYqYuIsJeDFLOE
G5IEaWYpAZCBjyEohMCAS60ZmmFZkv7gcwzp+SGpPZoeFBu53vhvSOAHvp6S7Iag
evZ7EWQsiYQ2582ahZwNr15WyIG+b/wMc0Ff8P4PShtRIJvQcae5j349qYGFpZZp
IKdoB/upQWgDZpxqIa2WRX+NsnHleX+r/0M5keVjZlznb4ZN+jpZJPxUGlGXnotc
OuZFDBKg0l1WuLkWAP6MyUNBfwhywPdR0U1oqsJHkiRbPlu1sEIvLh0KGFoVZPz/
OaXRxXgEZn0v7n/Ve96RTrWiTJd5pbO5REdTl1S+p30eVoDyQGzvQ51fXn02RsLW
8y4Wrj/2jBTZHFA9xmvwZ1cniTHbDgOiIt6pZdZ0rp/0woAddOEUCd2aG3hr8h9j
aw9tD14OmWPq0m8IJKKaYhIr05IMH/zP7Sc1RtC8cfWTbI+3ho7CUQpm993AjZTv
/BgX4qg2Fel6YVXIvv9nukZ9kcy0XEA8vfvpb6RjSS7dblOf4pgSMW6hFpSMkNID
cxHsRi7CKHlE1Fu8l013tpYS9L3tEJWhHA4skNY6QMaCFH4ER5ScgboZjCUAJzxw
RqDpONvEjy8wof79dtxXn5uURwWH8b2mnAKcvCUmPi0LO/ipuBtDsLhN/NUWhIVz
x+e1X4xaR1ImavPJYtQlHoLEyG+dr5GJ8w4XB3zqF13O/8Lgk354ZXZZHIkwThke
OT7H1t2/ClVrZrhw4DqmMMgS8JPmD/QvXwqk8kNQggZTV8E7RNXVrgrF6kTDUnbK
iaaY0hOi9s4h3H2UR4YVAg5sEURTuI5mZ+5tYYfSVBVLhATtK4qlU1yR5reoSi9F
VHmkCy6AD3TD0tD307HuE1EOsOPrUy4cYje7/Om/ow/iL9vEWIsznjLSbfCQFNCh
vMi/DHEEZ5Jep75lm3kVvV+kVgf8gXdxYk+taJP0/apJp8Zqrve3Cwi8vEmSlhYV
sHwTj/Hi+wpom1bQw26PpNHQa+oSUfBpVRnq+UyvYrURrCYcdWMjyAAtYtpNK2YN
CT41m6j8fnKWaTNAOvEdfLkKzNSA8hfSzziGvdXAspN7cozfUgovSe+6JyeSVDud
9Sgo72fXLU8C0zyTlETiIZcHErumrRTIDQTRW4RMnf+UNAL0iKsMMSZn44ANCXbw
eRaguJHqs6V3tphqJAm+AEgqrhAaKd+6ABFPVo43Tnyxxx1EuBxD/70S9jLiriTH
2ulodKCp4LWWFeVSk3HSdE/YHFp3CeSxvO3LcsOoZl0E3bEHK3rnlrYayp87vg6R
UzT5ZTTe2vA7UrETJRIjZHCrNsKy4x7SZVA5ROZmmYqpTP2MnFi/+GeJm+xOJrG7
mwUD6rggxNft+sLdoO1jJ5bmBs8WRtGKO1QcmY57rCK22I3ER4yC8XF5iD2vh7QE
UzwzTJeq+cQ/wnaG2KDGYIWK3pJ1tPXUSZzftJgsbSIJNrtH/XicuwqEO1gmrS7E
GMinGNQTzTTcf+5H9y3cRttn/JfzA2lQhUO8w0II1HLhPil6pwwW+x8XzMy5qL6k
hvC6rOnTe8zPkSj3mbiUKeJaqxH8/91SFzT/gcB0lZyg2DUQG+EsL7hefdsMBi9Y
zW2JX+wHSElP4vVIUkOsMs45/yOVFfys7hA41uZNVIQ4Hh9wrMhC9+NAv4mhj7D0
sP+i/FdVKsymimRoQ7UqqRnc0g8lL5MDjtCiYu0DrKvR/Okob23YyosPaph0MpZT
D2gzsBR/MSYfi562FjKa+N90NDZQLPaN7TZg2fFFYxtjADyiUQlnjGIA2RhenlqP
uZB1A/TFzfO8y7hsBzqFP7IiarhVs2JsvoPD5rMSGe08HVzAo3LYtB4lvfmVro1U
JnxjWKEzjTQJ6SghNBa4sOK3XpipSPgt9izUy5YvfAw7jtbpu8IAu6fNpyZbgvaf
QfLy+Y9zKIu5s1cP23Evc8DixickRDseQgv5DrTXJ0gFcJa4j8vR8qfunUgk7mi4
fDgu6VCWQJPEqWe+L4JEvf93ONWq4H74iKT4Pwat0hzOjsSjwpolBUJ/Pqo2FdNN
sbPBUOeW46zfmvcMrcBbGwYQmn10GBipTUraZ1ZQxgqWdZg8SJQmps3uULbAMLjf
kl6vuGbqgnDtEGcKWmi5yzvvAaFwaD2t1F332+NMUkCpoTyMwsgRoPSj5xZa+DA+
LuyoWIu1JhMNevx4KEZAOMZNnXjaCDEIdBfptsMxuc6xr/jD0UAgneQfw7/Fz3hx
wQBnGLw6NwaXjWqhr+MzqOI4GeYY58o1tL8Y5TulIKRmoWOU0EDKiEuNj03w6rUN
TnHuM1uRANTf8aEL1h6zeSrUIsVMwzDQV65D9VwgwOUFwisz1ydubo6jtEM3MmAM
bt8CUqUcvqiXWpe0187wMUr5R3GH+tFbgYX/AXktjSgHRDmaTMKjjy8K02f69AH3
vTic+9sgNuICYe4tl2kriUSXbDQCcXPurryu7g3oGSc7oM0XTMgeS9gyFylem0eq
H++Se9xkbzHwnC/rDeJhhZ2DCkvTwPRVr4B71LGCn56dURBxpccLvf12Wt/uE24R
ZE8be2+7YhnnukRpVcJbMT2+pucLmojALekzCgYFhcG6LgHfGRHufO6YIN7SBnC0
7Y2XsoV7oeJn4iR01IcbUm0+KjHhydx2qKB52REzDg09ZP8XJCIFxtwO9lLxfF/P
GVRBdYzh2bZeL2KAz2FkgvKuv3ywFt0fRAnu421xNF40OabuDCCFtG6XtvNvLMv7
XbLJpZhv8SUP+hPa7tckF4oD3hkCD6aYDktc8rxe0/9Esz00ChFB7ba++ZdpSdZE
csGdH2z50ooPW2vg3rj0UDmlgLAOCOxD131o5YL6w5WS6XY9RrX1YwSNT5TH8Ff6
9mhO9pygcxg7+umpsTDxpQmkrO55y/SQ2GneK5iWT6Z9DULZ+vLwMBOpDa9Ega7Z
ifdx3mgNIQ9XGOzonPVmGn1Ex3ciS/YK8KnGuP+vGoY1yeRD1/IprrWCXsmHIbL2
lsQQDtQnOYEPt7BnSkWZWixZB9e3kIEbDAr7+hLI9dOGXyzrSTGEOGXSxDEFHx1C
N6H/Ih6Yigeh7yb/qJOZUa3VTwkImP3OLs+CbX0/pzh0pq+wleq9A8Bni5Gtbws6
qpHG+/7vPqduD0xgV+FMSrMsrbFU8HtqfOIzFpHTHPBSD0WneHVf2L/OapL+7DmU
+LrFWJvcj9CJYa9REHzY2Nl6Kmo5atC2016gYxwOrQ0rhUxJNziO9IHwG+qPDXFU
zRlD/Yorem3d7FwOwbhjEL91J4/GN3m7OxkRZm+7YO7xPtp9xoLkCxTC7WIIvt9l
5W5evtf7vyzl4Ajt8+PkjEz2Wh1kUGQbpryXxtU0HkEDD/OWth6Q9heOTLlzQ3Nd
Bl+zXqnNJsuK2K/nMKEsSjSqAN9UWHEg7VVVcFBvEVG+VKbjWVjWqSVIEbdL/Dp7
Q5/PHf5h12buIFRGNoMCsTeRKWIhVTwTYMNXuaFu5gItKmNP+Z1uvOh+v89dWZaI
PMkWe7cOUfQPPC0Uam5I7T47y7TRhm0UlVsmoxVBrGj/wWTZWQftOjBALDcoHGKv
k/bkBFfpBI065XrhifwNgPsbNEgj7lVNaMqTopPwhe2DPxKM1ePAdDO7kJDwk4rI
LE2GYUZfqi8BuyGUGh1VQXNP0LUSkI0vB0glSS2U+a1jls7n/jOUvEFJv4P/v+U5
Id4TJY6FRUwTIH6Tao437Dp8ucWCbipSIj/rx2rn7mOjIysYlI8g8aQTm5MFqSRI
KedWsQK7ocPiKHrvrZ6VXuU8dN+pDsWQmGJX9us140g+puZFVVwuS4TaSKJwKxtD
0I2x8DGkwWYsdbtYbDv9gRzE1NrV3j9IFtE7m7taL6xCmHr7XpeMYZN+VBRw2YDM
LGUNVCfEzjfmhbh6x6kfjxfoo1bUPmwKuOe+aZR+KY3/gtTe6Nxc0FQMGaq8QZM9
l+VzHtVnINBjROUuPdxnkPrqGRihXNX81P5VpKyl9v85jcYg/Ln0GPEgggrqYg7X
iowZownYCY9IEX05mHscR9gG3F8JEhdHWQH9ZnukswmwQvXUHpIfhksEAy0TS+ig
Msatcmu40OZIbGThF9L6aW2hWIiXRXlDBHL1lwyY8GXI89s1rip+OeGx//rDmKiQ
JW3xQtsRuLEx99e7Fx00HpL4HYKt0KNB06YwT6ifkbNxh4eyH++E5oYEY0p7akv2
W521+KuXiDhOuKdAwGCIgXscKS1EjZ65r0HPrBLU6a6xeqWzd+Ct7p0bVoiEE/ro
OvVwnSc71XjAdkJanTyJjefwQULr47KFvNhn3u+i+7nQqroEMnc78xCUCa2z8qel
NEvvv8dyFV4zhCyItNFwT53cq6EXyoBalIBwSDQex3jPZo1nAlFvzrvBvQWdYggw
UzA6A2v+0Vq1FpKGbqRnUy0ewwNudmF6RVVnd/oHoz3q7gE7HVKmfO36fwgmVs8R
noVsn/kMYFKWIEnpBvig+MQMqrl+1ozFRuC1iaWAOgvdpBfuTkFPgbVhqq2ThbZ3
C1fZz3KVwdGZdpNB9R0X2ZuhQxidBFUsVKnKCGDEGes4AbWYDc/Ir52B3dzdN4q7
VRJ5VUNJ72BANYu78hedeNzaFOVtw3zlyais9p7xJRrTTH4jbf8Q17HNwPrTWY5q
MOqih6o+5B8a798AIug7Mi1tNSkiS9epRyGefVV0i1Csdwpt4VDUiGYCkWWEPsFO
Pnyroe8RTp7ZdZWmNfjA0iTLUBJ8zxah2KHEZlsEzTPSi6PTiwgx4YuAwknaNyos
5NafUrp+L1MNxvtqOzJtPFWn4WfBRlGahrJE0ONkXWiYwagxeBVnAmRoFtbXJ2we
zTmY6DaQWFkUuVzlLFNnPHe7rXYF+XOTglRGcjlxFkZTK799Tp/LyhWfa7FhpK0p
VhvPyNd/pyVkUpbubqzMVvTxHR9vsbQV4/ksNm0qE1xCX+2WZRPxpUkgr9e7KuVm
VQU6iINy4beO6zFad5VkdNLfORcJhNegUNL5I12zjkgZtLR+pzOU8SJCxMqhM466
SsXkAY9dO8pFD73UDnPgXyL+9/ygWYEXduqOgaCzZwF9XXu3SBn9Hg1Dls5qLBBJ
c9EEfxuknhtK+OCuMprh22K5QRc6QQANfJjx/AwDqJ1ybB76KbjokENxBRWZKTnb
xpYytJr/pwHZwluHgxXfTsPmNSjugYnxN3OpMVu7fIi3BirIuINyeHif1T6EiiE0
2V5WQcN2vEGuG7drH3u1QNon/aDiKs1vhxi3te9sTy/8QJTlEh16kYAtR0EcM8SL
q/zNF+oNYUq1KolCCkGH6MEGJd2DF/2n8pzFmc+5tkr+z/8a5/RO9Jku4n1qrCgg
7BXa1FujEHfJbyOhE/VgL8WNxFiw0ukc2+eM1GgTW4UbpfFPj8xwYOOwMWH42xoe
SdRnDA5L7qJdau7G+a32UnUBZuAwataPmjQBoYhoCgoZ53tO59Gpwrn9V7nObS2F
Dbsb7VKLpYWThD/owiS3OqfKfFTG2FuGsVTVHhjx9LDRRmS7X5dtcnJtgMmBQSu9
BCo3CAEEcjkztUZOmMUo58rvKlvcwoYnbwwt+dfb99DiREXq9i7UlXj9vxmsVPst
9R/cPowYIHz9yG67lrhgs0qQjOCmUS7ehVd+iYZk4lu61Kq0760aYMRG98NyAPCl
/XQ/TeDn3FQGx0b9S0iVFOV5ZweSabkFKmxkh8FhK7N76cXnjr2zQTTBQVh+IyRz
04SCyAjYyPo1cB3CSFvIa8UujH0GgcKvP5XKZL6SXx4GEyqM3btJoMeFcpdmdfR0
H7TYDE3od54PrKDTCJnTLNSHme9NK4MAXTsIfyWbNeWvKN/r6u9ThPEZme+zQZsF
qTSmoTqRXTswcrIHWMm0XyC7+oEpXq4NlYiqYRAVTSA3eQpSWzhUxySF7w4fwd1y
naOL2Kb5ET2lUqOWHujq7hHRGBltm4dzBSbJGwyGLknO4NsuUDGmjP0er2puitaB
jYehqkCIcinsSN13KbXgCvfY9HG8weU1rtcGp6Tz1LFeV+0B6a0SMOira6qCMdvq
XfnOl1uicWrVQwKP3uQn9Dlzd8cZWReHHjHNvFTxdz6Oyo/r/M0zaducVfOHtmTq
/YMxmGwD4M8e7QS+/ayzIqOTCfcdIEXb/Pj7FRiz9zF85f0Z0Vj1cOjyFkzvweou
WzPn792ZJT/SdKuqbMWDsvhORQ3XFjIm/x/erQJQ4euCxO5I6tyEZXkcxNe0QE7H
qkjgfyegZDevi8mmUd6c8rOwWryRj59wB++OArt2wZ60HL6+ucwL0E3C+5ZDwEVW
EN8V3Jo4lYucYLBPqzfE9X3QUw72tJb7qX2DJuQwCggvh0n69GItL+t1J9XnFHAi
tWTdoQVoNTreA4K5wnso89B4AmVj1tx2nnTPQY1lk+dpgLBhXcKGiqwpka7FKybx
2fsbO6GXc6o6X3N8vdkA5DVc3RjTftlT5OaEqcl0Q8bIuNDPzPTn+OETmw9lMA16
eFmeOrHjSBqNZ7N4izfeaekGxgISkyUcp8N54HG6I6oxxqzAGbHQEuEAE89pxlKa
gogreoUSjiddWGTQGYPD1Af7hR0d0nj3tjXaKRh6aaatBbmec+J/hFhDve7cuBr/
wIp3LYd6Th6CBsq3ms0WZOqYcL6WwsRQDJmdQhJl94bcbdfDKAemhq2gAkoE+Pp4
j3YD/N8aEkIEDi3P1sqbLRUXcxinaMqSG6NNP7Pydpef2R3HyV+7hS52H93px4oB
tIScgGXNwxX8BZxPv1uABFCRZsccClRVZ2wEnxbyduJO4qZNeXSEU531kuhPaPwm
EB98/o46e7fDRFlF2Iged9lKZcBt+iAOh1heiJv/nBEGrW/tK64CgqdssMYX02qc
HLuOpv5shdh1B4T/WwNgIxy1JqPI5vmKRP7ybGYUxSIKLXYuK+7Fg3k7xxar624Y
ABr30oznz1zcr3nqxkWPqGUE6knzXN2TpQfHr+bb8OadQ375xrw4KgvGNVeUoh+F
V9OMCVjsYxQ8K2aLirX3+/gS5u/yBRmUzLq90U7LQsPaTj7dUsQFJdsetb8k1mfR
k2c2OctdP9wN/H97tDjMWPH+ZEMMrImn470jx97G+WkAvLK1xOMM5/SwT5SrObZ+
0JXqpIzn15IK2N3WeFFUHZTPt/0sqq7zxzZOanWnJcE7LRZaeJKS3sebc03NA70X
I/qJWlEIBf2Bt3VvIM/XzoYEGQK4SEWJBoDzO7G6znICJCqbxvPTW6RBY2SB9FJq
mt99yKsnm/YmRTSBlTaB1i4uboW8haazbjI8cylewXDbU/w4jILIJDxeNNU/u+Pv
vgmJrAj6QwqpthMDWD0CcI/JX23RQceWyouWnoKbXB1b7veEw3yJhph+NqczuYHy
N9sC/njXizXPY99fao6WK9dqOOsaAwJqdksK6Kcdk+9s03HPX2DS+KmId402gFcY
+6cgq1UZzR8f3FLaM2NGixK2kxBNilAaHWcI6i4KOaoQQLk6plPmMJkT90dPST2O
xw/SCNS6BxY07ke+XIb2UAnAziaV3g4TMhK51TENpCr7uO6R3tUBXGJRl2Ji9dj/
w17+0zn1dPvLJTb53QN4wPLdzCkEC+ng31mmhCKY0g5jTZZBHiIHEOeKzgGqrPod
NGAVWB11+ulue//R1xZnxYE9UsaU+DxqH0TSEtqy2XP1ztuCA5ZHB9DbwOPg74GC
5MthTAJRq1uGJjxfzdncDp8ajgsVjOvT/EODvhYJQluDiCQLE/+tj6or61udErLU
Wk7hmQGO+BSonC6alyaesK8HhBDBZheUoHyd7crMoD+lkY2Tu9XLu3YNHkc0hKmg
wken8FRhsySibAB6J7/MfP3OREuKAq3LQh9TGWYD+gaxBhOigP/WzPRUDE0Lgf6X
NV+sIaC6Xx09fZ/GqpBndbyuc13MzaalOgSlznVCCQDjwjbpImyP5Psy0xrzp5hs
w1u9RwVMdpTq9ERJCYRz4wr8QfnWG76fQZKm5bVPiFSAf2QFuY62pUGjdee8cgLj
xWpeeE0v1E9moFvs/UZnzie9lIIxp3ED/rb9zljym1N3c5mPPd2S+lRv5tHVJVJc
m9/siXi2IfdOO5W2bolZ6Gx26z42z9eH9AX8vKvgP/3mD8vyoRbJ92sODg6ZkXFm
uVdqyFBi6zdYrbIfE65aliIIrcPA5LLEWf8lxhx/v40klmRMWCRyM58+x8Boltp4
A6A4RwbrIXVBUN01+7KYvUeS5JPMFvsvuhuUUkPpWX0rWqVfJlf7Q/YcMXwrMoVw
q445R0SzO4uEcCBrmL7k3hHM7Un87ABQmY8DZmAwc+PFs1eWzNNExqZmYULIFVhZ
bWpqEXQfLl+4StaW6+xRQ2RBzNEihYCTG81uuoHM5M1i9qETOk8soPKNKBFd0s38
Jda8LaAw1RpQ13JeEyi0VjkJPNGxrn6qRLaMf6sc5ma+r3XVuEGKm75egCmeJBH4
N1PfI5pSveaYueJ/FoYo6ZI9rApZI36Ueu+beYeOTpZo0E2ZX8tDYWghsBut6nht
L2VrLrX+v3Y+wJ1FwMmaxbT8sECGXGRJK+bHlRl6IGAIodeiFLO+koSbhDndklib
Vi5Xqpq8A+Gsp1O+Pu7ISgA6R9LSqWjkS9j81139/Y9sGB7Uo86nAb8smKvomJj/
dpOEzy6iUHwFfOy2zmrGSkwYBPIshSek1nSo/jTShDfcCANptp1zw8EA53gTroo3
bujeT2OBNYFQEKwGVsh/NWsCp+mhBQpECnNuXsDxLYfcN1ABqS9Jy20BOYjhXRwM
cVPw29NhEZywQsPS0taNzaVfsUNx5y2OH28wvLK9ddtkp057rnTdPooKfnAzwrw3
ZChc0lRaYi+u+G6Y9Z0Egfp1LW+5pTccbK8tLWzY/xWtnPp4CPqsGsfR+TRRb4cj
U0KOJ9289Hn60nIG5pS7ms3xWkw9i5TWMscM+OepMiULhroN41fOEfaCzmD7foOK
IrN2oI4jfU+annUiBTrkS5HhOeNO5PVTg+JCHNwtivMsvWnXA0eABl1WX3uTzadI
DLIwQY0e/uYSc0s+4NTaZ8rJGGWQXz/M9cjmLT+0ag8lCxOK5OgqSsSlwpYKbHnQ
TFmjeyTOUjtVmpPR4jnmtdsXgJgcW3jVdVM0+lV9P07+xsouhioFhjHX1lqpxbNU
cpd/x5TcDE/IdNfLPq4LwD9MwWToOlLkgveCn9gqPRDhxrrjdpRiUGQqLzGkq3Tm
iAQEISKkh6wvb/JFfSoEYUEuxaRAXlDjqdmKcbiQi21nuHtpyASHGqjQSnA/ZqLj
GSUBXIpRuRxnpFp/1FaHU+ICLrYvR1/ZyRT70NWlwvurp9Y7rpVhMGXWVeiAGrgi
aZdzmUwZWDKlolzxcAQUn73c4paWn4HvljiVJWO/en/ycz6WLnwYFOhiIAZYI4s2
bzdKzUgtmCt9I/uA1l7NHopnCr2wcOGgcJcdrgUCKtjQgpIuwiYajqeCXdvoppyc
2w1+J9M7oTXvKnUQ1AlaVAmRgXAqm2j9QblRlxCpRGjtN8nGo//NUQoYnF/dnHb0
srcXSE5gq8w7miwDfpe9yopuDYrFFkGlqqQ6j//3/gGi1GywA7e2lP78j6EZ8raP
67upthgNe3dINEzT7XAUMryIoj1lv+l2rM8Fvotq1EUXkJaIn5cZTbJQFg2uMDxo
rQ+vekFlQvVryC5R2ulNeGDKn13Z1jYTYIn3yLRtoh5guz+yfUQsWsFK7gyRoRWu
jIYU8B+Sg/bvmGZqs8cxtGRr72dcEccRYp6H6wEF20gFeAXSrI2IlSDgmpEudKdh
V3Z+SLtJTClvSX/r/2EUpjZLrookbzHcf+1V++RdKBpYm+TZ4kg+8eJZRV0w1DbI
rlkKcFqp97ACzP1/JDqUJ1dYNCu5+fp6NqfVVKb6Zsb6ULcCvs2TqIKulyD/M+Tx
Y2RUJ2fz7n80nG4ktqjQ1jawQmpwJJTo1DVXf9+qDhaJxZzQlf6a6FRnWj6idxJb
dhimVw7/SEGVI0x47D57jnDki2lJo87UibxuQLRjT0dpAiVl11mRqvB+8jO+MYA2
9HDxI74XA968ai30ZgAkNWE70aRreFdzoodtcw+QiVKIU294eLWx2ZqPs07KX5ez
1TzBCwbaR8RDesUgEYy0x4PUe8XIif2SR+FUqzbok/Z4IaLsltSx83cDFdYgwTcC
Uh/eCDjJal4HJn6VA8bKFdnGiyBzo/A5svl4XPrK2QzKR9dQxI3mNBVJcRohkTQ3
RLrKb4qIZ8cE4sC+zv0uMZQ8Xvs+bdsqSTyjyhswUMmo0AjQnKru5KFVQsMDoBjN
MhcXUc6EToWtTEBprUZPdXyfXeDS/QbwN8zjU62VWsdBOZOrOHz9XI8LzIomhX45
zIGUqJHw0Wpp0/6oGM8AiX3fP3bV+ox0xceNuWpqLRGcDbIEdtZQatGwsjtaX4V5
XsaMVguGLKxpEXXbHLTrMG4kNPkVd5I6keFj6harmHjunH1of3W72a1IZWVYRMyo
+KXM1F96JfOQrXrmKa7hfddsoL0wrBnJaRsslHDwldeDUiBZbSXK7Wg8dC87dkez
3fwzKwB9odt9DgYrzYnSAeMlUn2ENSp1G4MvSfgsmKFxhWDO25GknNPHIgR+8VaL
JILLhGSvsVva+3KHDdcMuGo0dLYHfJtfOpg3Tfip9XoZzWeFPYR1cfFHqZzjV+Nh
lQLVKrY2F6JEPglU/bbfypcHtCErFYvS0W1URw7uydWDn3GWoD7NTTxfwCf/DBqV
M8UOTX4iKD/Cn6CIYsdSE0wwybo3DHa3MaGPKKrxrmcdPR40onaosR/gAAFTEIqn
p/DLw5L+mlETvnKTECvNAuKZS+xVdVMkn8p7UDpkR+jvBjkf4hOaxQeJ7Ts3PjL0
DD6UJ+7JhZu4shGoQPvJiC1O54koq3iSrH8JHad25Soe7bvgPcEQHD5mscsWlmbE
WgQLxHh58EDT6tIwRd1ZrS08dgKQgoHMviEq44xPoFNNxNn8cVbqwrcf3vhJ+xAK
Jn6WTPZmn6tGL+Jgg2PPBZHcZsV+IQoYH+E11octE4Mi+AwG0gZvQwAdXuU3COWj
fJOE+yJWOZr2aPffd9ojx+o8Bo7hBPLnQff6Rn7NRKv47K1SeLALbgCeG5TDkcqi
+JVLQqT7hJi6xSmIr0Ty/Z0eqBaWA6PWZhr5MrdDIuWqLl2te1lvWjNLTIN9UCKI
tl4/5J6QPWCTvUPrg1KkI9fT1Bm+reqpyJGZ9EFZs3VQnMrW/weseDWjaY4Km2YO
n1KRhfdiIvWX3WMVPA9qVh92K1G4Gvhe4QnQ8m4uWGXrbXIIQzC2ADu8sZZ627Aa
B1nSVl1j1uuS06fcWQuZUylDrjjTRUdKy91YQD5Ue80HknlhNLzxUOnmtrYOZOFy
6u+9//kis9thzNscN6rA3TdqlgRuB3kRTYN3KKBrgxWZkshGJ+kOlZIL1rPqrwpp
ddnQvgVDd4ekxcIaHvJIKMfXv8QLawNyQ06dc81DGXiaHAZBoHahZBgzmmJfMZzL
47a0Xtp11YO7o3cV7l3TkRoCGTYpKaeA11MKU2OeIKKMD3iR0i2nsfZ/1krR3YFK
1W2/+iR+ze55+bd4lPUU5dZXZs6a26w/CA7l+Mgeh4eKJN+2r07rU/WLzDq4VAly
OzH6ES3iC1F6QesxjqzLMPdeEANTEtPeceEJZ0ErwHw6Qz4gPyga4AqoUeVlQlxI
80Eo7GYGJ4+Pm0k8u+drj9RWc3TZRUgXCvv4rOFvgBmvoHenBQYxQzzQuuo7NhFl
aDNMf8P/eh5WrOJGqAxeRT7MtTw5OOmAZ+j9W2aPtv2Llr3IbOfgIpD/oS+cgbPE
QQLoaPqa3fJGwR783NVV+ROtkkTG/mdURYHT8CVcz/GRvAGNHkzN5A+8cWXqEInn
jydmDKHpRI2Is5pFLmNJbp27YsckLcqbl/J+x6SZiRvkz0S6SwnbqPJvNgmmPcCJ
d0gDCywO2jclZXwg59A/LaLY0pEAL85snF3ey2Ck9tkHjaCc0BdS+mFY5hTBucnZ
5sVVqxOEne/2FIZgqCJe4JqJp+6es6OzyhIxl3JKKnurO4Sk3/QZnBnnVJo1jszQ
EZ4PJCE+vTeJNfhzBAuwfM5CLG1VB9jb5n5Ns/vKsYwhh+8++KUb/JOcmcZYEmh+
iRPrYN+gSLvgRUQR18ANlxxnGLPGH9eCoxOQxstTNCujPokXMCnTR34Uy4gCBkk0
l1QnvlIGQpMa5ANmz4a+hlGxM6g7yNSlOLEhWMP8BhywvBlV/KZqInRr9jpLb1jf
y/KwbtbF8u0fYYyXtsN9p8EZOEWlU3tl/f9p/9YHfr1t70fpT0ZPkeCuW1juLPFp
xuqI7EYBxcDwazoWTzvF+Xv5Jq2wd3sVhA0Ixe/0nvqM37E8xNGpsqAo+cPQ8giN
QZ+IbIxg47hG3TnSXV9c7xphWiK4z+z164e2ZDFjamOEdP8ZDO1QsiPWYhRDJUzi
8Je2BrIVnsoTGgtHvhg8PXWEwjJ+cXv9z6GwW6Zv+igmzLls5PHrSl0mPchX9JTY
eofqmYeD0IoH9Ff4xSTWrgbIUf7Rkzg3mfgM7fuoUINHFZtKdRweD7aKIhaVldds
87oSsdG57qMum+0PqQboulrIcLbfSrB6GiPQQUYNR4K8nABwCvbGNiy+steskRTu
HUcCAJnTglUiIGhCIdmxcSe2i7EUYkT9KczVPUfw9CadjBVHtLr5ip409WGFtUS2
CHH0LoIJSuBkKgEdBmAxaPVXOfkgDj2Mqb+sHs4aNizM1YpEE67vEYuaAAIIigci
/PkPTtdEwAfK5HFj+Oz85WhQeA2WFw4eGVWAf3dLyt6+j5CDPQrbTitdpyFyq+/F
8EJbrrYwzqo5pbtCGRRMbN5hEA/rYPL1OJ/5BpSCdnSeKwodOCB0J7rnoG+pUfCt
jLACrb7hI9cE5u7VUw85NFuI39Rzmw7lN+sJgkScIKFlRES22bidVZrJM3hckFJO
iyZ/TJw2dP24+UnGdKA9fK2SUyj5fBYbxdn+ArND59f0w1B8LjG5sLnEMHiU+JHm
eZhksVoqgFD1tkTWL+hH2/qKjc0ftFVCXtDAAo4KzSr8kC/LJ002CFwtdWSnAwi/
AHk/BF2qcKFpawnxbo/wM/hQkJfCzbElHuGrxbZ3Y6rng/E7czQ75OhcEP9aPJx0
fk9GqP7oQL36C/fLDV/pOrG0YjNUDUKfvMzdSGZ1xD3NC4niZlwK6RuwJP4Y8ayq
Gt7pd9CCT03WzDICHkYm3DvVUlE47Wq9BsBJF137a54lpUCAaoUVN6jMouDOYV50
EdPT1z8PsmUD4avWeLvU9ywd2TTosm5fpDwEjjJIpXxq0g3Hk6R5xG2iPJxL1Lly
WxYWeB9+v+GpFBppD9dBTKfvv4vf3LOqFjKQuuGWJ4m9Zu7zGpICefRpZX5fK9X4
WBK3PxoLbxjYQmjMEnmog98Zc5F99hRMJ24yAIShKrUzcU6tg7CYD5iL4E8Nj9Xv
msIdJWsRw2oHXP0odTCcEWej4/lUHzXe0eA5gjJSaPwzJVVfTNqEFZBRjlAxQKpT
CdHBSRZA+or9OAJ2YtmSC8s6u3mlrrx+fea6k4/dPq/2m0nlIc3WPZlEFTpiquwD
hX5D7VO3V0jYm98pUpqjIxwOT36HGEghb15kkHXUks8KizaWWE7OIUFhO4Fhw7+l
2r9y8+iO2yWZwGigdpB+kcHi9OYlAvn0pXX8/DCk4e/Nrg0GRJ70bt2lYu9C5qvF
R3/E7eS9ODVETPPsjVvYzxJ4tcOWb5NfiWGSeJj0pqaS2wBf+o0SEfcg3ulvdu6X
u1uedrUrwBm9jHLqIIZkVXrYnzlOKs78H1ZNMmiToYIe6Yu4vCv6OjLcw2GEPlaY
usa8qiMN7pbXzgJf4uwk3B1wU23sapUc2XO3g0+ZUoS4JsB/Z1bAC3YZ71Z4Tf8O
Omg6zoLQBMR2QkRfN2Pkh6CE12q9N0KJvaXuyRCAGV2pqTekPuvkrkHyj24WDkrV
ZlZ1HbpV9kDwKfHmC7DEHhu0FG2bn6NB7RcqF6BpmI1gIfFixwmiAnTCPlDiv8ER
ScJ15EfUGYJ3guZpWqCCfbizUYUh+Y7GQXTY3OxeF3ibcbsK8XHifNqUzOxKgLFR
982NIsfoaJco3eyJnv4a3dGtUSfCBToSXbMd9MbVpYahayI2rKfZpEKQ7v5xIR+L
xTUoEqC5Iyw/ULl9erYhgLTK8/O5zBzH+L3kCnX8ZYwsF6VSFbAS36vKNyQww7RU
zJVAGS8yKajXVXvS7J0CfVyUR0EOifljOWncLGIVjoQcSfZj8NnMsQEkh9eTMEfm
hWXt7liVUyemjIryozC8vGXTJmkkCV0FwdkyW4ugvifytCGasH6WSy99jIG+GVMe
A2L2uze6mStGHrTna6VZyNx14VanttAB/tzs3FwfcPnAtXr/EZGeg8EfNBQX/d5W
7m00OQoVCvME8Fs8MKi+rELGliA5bEELd66VZK65eVrqGANTUPSx9f+x4i/bjRCs
VbcZiQy376sTE9xMcnO/+f+aWVuruXNusNQQcJMAwSMBPB5dUGAkfnF5X+rvFyZt
bnL8i25t4EC09vuXd5OUdY5gFKkg8hWFuxLeOMfuJwJJHUjOpiUTvahHJ/pj50IV
Z0zTvU2xL/xQitvvX0GoMuIgX9HBQZ1aUyuMLvbhKjuWtqgrRtCo6YWXRY+RRwJX
Gh8N0teeCmuFM7poA8j7zcR1AKXfrjG0zTAVRe3yJB73SpsSZXT9fVsVm5UtoPyg
dY7ptMZkfoUngLgYbr/G7vw9z6XlppYe9Df8LxgR+t33AAIpGaMNE6rK5WnlLzU/
W+byBX4xGpmeejhSN+1G5uzYOI8/d1tkMPFp9fua8+Q1pdXeS4XiJRl+k5yOlRan
L4j2vnz9u8thq/oPimlGGhSQQG0OysT1piLPyLgZmaYsYjanQbCcUvEtPozAw7Ac
2aRDqZnUcClBnNfc0dWl0kveuX+bKnrRAS3IPOtnl78OvMZfM0pdSjJ7pRxakIeR
FXNCSHvIIBPDr/CyDzJwXHJSMgl2a8YImFoWaLiGz4ZgEqmSQ2k18MLr/eCN+XcO
cTTxzHUeK5uBN5I4SVZh7tSIudt+BoDl13d63RKI+g8HR3vy+XuRk4cj8dojka2O
JMQjzdEYBbmwz6oAGWMmK4HptIzvEyWx4L9Jq48QNLOgnpsr2iAlvlk9hevuWLKP
pynZ2JR3UHt8jugCXLHDHhhmYw8tnhtAiRZ13lC/8mtfEAOho/0AqubgYRc6kOm1
6KOvZgkjgrHzo5bxtDRFIg==
`protect END_PROTECTED
