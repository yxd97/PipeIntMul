`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AC/0PAcdSfApUHpMxJjG7OZ5zrVpMG2v58G75vpV/28oGQQMAwkMgOGU/xHtydqY
yMPm5EqnlTOSsQPlI49JewPBApRb3Ro3fx3V4g3xygi2nYA3r6fIQq+vrENHw/7O
WqgwgDzrYtH++ISNnXspUcs43xio0/bhhGW0zTgnBXyv/kwbHoS0QXpTASjgQgy6
6hZGAKkzxe3G0mXC2L3MNoPLdvLut024y4rKjp/TkhNbyJ3L4wzwdTpnIQyrhzgy
PkNvaucPoAcBqogwxzVro0AbUhb5T1aVPeVu8v5LE5pVW+H6Rr9DLoR8ey6DDbc+
+xEkS0oe59BB44eaGvvSRen+OT/P4ggmwtW30QNJu6RYGyWsjhlqddyPEMZntoMh
+x5wUIMRoaEnfOC3bsTXSNOvxcKfh9M0l5oO4IApVh5gkmOKgPq4+8M48amhRLd0
uycAIG89l9mH94NCCKg9MmFGhAtCe2OS9mTlemHv88W9gFT+UjPfTqVbCknKmkzq
Ah24EqahUMgLb2O8kMizMiN7CrmEUNL37ZkW5qVbwoziOPIC+mb6WE3D3N+uT6o3
Jj8L/8GA+50vAGsBbQ46i+eAkXxtRGx0HVLFfblyxb0m38yLLMNtxbKSxIrbBPyY
1A4RUNULsq9mNzMFlHw7FXWkfDdxMBut7FY4K/iDNQqR/kPUuhmvWDgAUxJxosw/
iL5ZHS532Vf8s7RkE8KdjArldEG6kgMZagD/+knbW63ldF70eLFsk8foCIESdqgW
qrnD/zi5tKtf80qFEQsags1Y+6KxVLQ5aKCk6qnBBQkEC/XBh8XFaenu3aMk6Jj+
YP7qQIjwJHDPCUxpR5Lpt0BaTmD5ZfmDYHIL8mW8ZQTkIQiVndwfKg0KCepQ5Mb8
GLec5vTDXcIZYjfosqjc/Hcs9/vgALKVBnD96A/u+TsqRIYtAQnKxdxsQFwgLevZ
ezn20p+NFDvpCa+b+txZC7IMN6G5tbdmk4R66KqdJRPIsijp58wJd0Vvb9g6A7U5
gHTtmqeUcE6YE/mZ6HmVNM3Eem/jGxS5pe6qUmk6AHm9n3XH9TSkPnp1/ZdiFT35
0qllwoLNC4WCDYUn3MIrgCLPskll/MbBiMsj7kFzu7FDiDoyydADEvuQw2SZe0zw
Ik0EbCT+PleStYWTVRR6adSdbTgaIrRNbMImBCNq58Hyz9ivQdFaKKNfwQOZUCic
YLVb8prMBdECXrBnz+P0ilcmYns0HCCnc/K9C6zmgxClZE4++64gTtn3XaIN3bdI
Mji2TvI5k6ikHtOMlK2bwAQ8XGRAVqw/XWbhEds+hej9P5jHHdQ2DXTN/YSc2MUa
Z57hz22sOg3dCK/rblIM4O52Ifj/XNoPsjr2b6aoZx7A1e6zUQk52lRUe++gvwy7
yT7OFRiM/UhQ3j6+iRgCBv0H49QXMcjJz/fdKI4zilgfh1uNG0756xK5dVop1tAM
Dj/6SdJd/Cl58Ia/LRPMd9uoX0UMdETk5bPn0g+aQ/EhFeRHIugEm/9qoVlo5OmB
r6buGYCMh5fdvflwb+d4ACURhkTWZk/ZEtFIZk0yji3W4TQOPxOl4mQmom6HBwOG
FzcJp6wcW69A2F1Hm+cVrteevoV6hnAFZGsq+832BWXvpyd7rrIlZ0XFftNLL4kT
F7/YSEQTWS68ztdXmdCQri/+I3XyF4Xzc0nxBhgQM8RJicQAN+KWdjIA7DtMcUu5
ATsyQ4e1G9FnbG5QVPHRfc6+r42OjserK3uTgKAHRLAWcp4a8n503aPosij2RiiF
2FZcQHJ6Gt4S5BebMmSpLIU1IlRK3XYMpQ4IisLzp2FduL+JBjIrSbyEl0N+I6G5
1BM+htNdF51sYUfeCJn9Ir5Gn29KrIHn1lGr2GbcLl7s8LVpQvFAri2o1yc+2Nsg
iO9vK11qQR6vBeyMXlsYsqWvIbo4cpMr0Wg1NY0D31a18wshC4HwWp051yMoYbKM
YcoYeM1/mkAxYyDW1sXbxFJ9vAe93bEea8Pmu+uwg/FCIlZsfUNyjj5Sb3oEcrfC
S4NVg4o106nx0MbeXCzke+yLpHL39xR4y7D4CmkumTC3ytOGSI6Yjkaxwj8BGY92
2P44niMwnCUl9gS+l7LQ7Sfj3ZewTyGF0uVxBBN85s6oRk+il8I9YpL0a52h9S7C
uiDuanUCx1ogs4GwbVR1lmr+n7N2jprckFlnW78BRAZ9oVekxvBSEYgq7i/3oPa8
OyQS0xNBIxq254HpeRaIgje7SQ4FC1v2jhVCTGkRw0vF9e9AoCYgy91N8N1fiHrr
R2R3piM5QyZmaJZYRXYWJgtsx31fU6vibVyWgBAwudU5gaxadXrMqm5W8n28wDnH
b59pDb1Hw02EL9XZIcnexi9XZU0GDGBRQfy+YV5yUN1c04yrhu29pvAZ6HEwsP5R
7MmvAN1ZPJ7qhL+RWel/EX/hOqt82ix0WQeWKVIWsw5jZj/rJMY8YpWtPQl8fS+9
B+ZE77Qf20tGdGcHh6KCufhL5sZDTr+FQ8TQ55vgIgy23s//k9cbgcB6yzKVuo3/
9qBeW6StTE/OmgXqvBo7BApL0pw6t6pJQ6rS2rByIGU2DNAuBltBVCqADCgCN88K
2FbQG2oxglZpuulrqDt6MnYxaUa58nLjyWLV4JSc7iSQ+z4uirGwoX0iE1MTL0IH
+vOKP4a7nuw7SqAsztTBVl6ib/KTyd1p7YM9ph18VKgKVeklvJngK26/FHh9R5M+
3YDlC41VEqS14Q0L5FTCnIK6GSkJGCq2HYlOpRQf03aH79zcVAtLqvIuAivVfy2D
U1CNbuVCPyoFUYW8MnfdsVGe8/y35GK+pVZzv1XuYY9xON1T/IPj46ky4EbyM7ZK
k0TsXrBy9ekGnY5n/caI9YQ/wYVcY8Kf44+2kS6a5z5tZy4Wv9FhfWphxKs1By8R
R8O5IBXKj6h1dRO7F72fEKuk1nHB2LqK/bmDv6hKS7kR71reVBnnCpQIdvRmUd71
E45sUyPAEXod4loJcgTdgXa4CrzNBkSLsozT+bZLyW/3tYWVD8jgHBeNZrl7fdCA
bpGyJx/IlIKeICko6rStTNBgsZ0GGbjsIC3acJfxipizpBl+oITTMiJ/MI7rO3vW
yMgKSYJJVgEZ2UCi198bKXOaG3rqkw7SrwN3UegKRpJAXd3K48mKpUlYhrmN4Ek1
SLXlkA2yqoDIPyVxcO7OZzo0UJacwY4CYqn0WCa0K0WQDfZwIATHegm+FylGn1XR
ZHVSRtA7dkRU6x+5dFN3fKghZpNEusd9K7txzG8Bqds4clwGx10MhY/K+8YbnjN2
sqxGJmg2US0soy+mn6ONgpk8qBBnaG7/WAViO2Qwg+G3D1Pxa3jc9twNnXb9KjCX
4iIlgp5UUrJ+b4D560+UChoMKX3vpkkJP1G4DqCIgTKKDlQQ9uvEI21IzM0xjNFv
VGd06b/FBOkh3ei5hYeSYZpqdb9xrhn7Rn9ESpsEovAuEUrmnbs5WHCfBEHkPz3+
IsVuZZ0b0w4qALiK+dwc9hXCgcvY2QRB7GWYTfYu78/4AwSUHzOe/Rer3qsvluR2
FgRDCSImwwB16ukaxIiaujpMW1dWHmLGHmgK0cVIqcyUQyp3naaLpgZ0i05PWpQw
`protect END_PROTECTED
